magic
tech sky130A
magscale 1 2
timestamp 1634821592
<< error_p >>
rect 170 732 228 738
rect 366 732 424 738
rect 170 698 182 732
rect 366 698 378 732
rect 170 692 228 698
rect 366 692 424 698
<< pwell >>
rect -447 -526 447 526
<< nmos >>
rect -363 -500 -323 500
rect -265 -500 -225 500
rect -167 -500 -127 500
rect -69 -500 -29 500
rect 29 -500 69 500
rect 127 -500 167 500
rect 225 -500 265 500
rect 323 -500 363 500
<< ndiff >>
rect -421 459 -363 500
rect -421 425 -409 459
rect -375 425 -363 459
rect -421 391 -363 425
rect -421 357 -409 391
rect -375 357 -363 391
rect -421 323 -363 357
rect -421 289 -409 323
rect -375 289 -363 323
rect -421 255 -363 289
rect -421 221 -409 255
rect -375 221 -363 255
rect -421 187 -363 221
rect -421 153 -409 187
rect -375 153 -363 187
rect -421 119 -363 153
rect -421 85 -409 119
rect -375 85 -363 119
rect -421 51 -363 85
rect -421 17 -409 51
rect -375 17 -363 51
rect -421 -17 -363 17
rect -421 -51 -409 -17
rect -375 -51 -363 -17
rect -421 -85 -363 -51
rect -421 -119 -409 -85
rect -375 -119 -363 -85
rect -421 -153 -363 -119
rect -421 -187 -409 -153
rect -375 -187 -363 -153
rect -421 -221 -363 -187
rect -421 -255 -409 -221
rect -375 -255 -363 -221
rect -421 -289 -363 -255
rect -421 -323 -409 -289
rect -375 -323 -363 -289
rect -421 -357 -363 -323
rect -421 -391 -409 -357
rect -375 -391 -363 -357
rect -421 -425 -363 -391
rect -421 -459 -409 -425
rect -375 -459 -363 -425
rect -421 -500 -363 -459
rect -323 459 -265 500
rect -323 425 -311 459
rect -277 425 -265 459
rect -323 391 -265 425
rect -323 357 -311 391
rect -277 357 -265 391
rect -323 323 -265 357
rect -323 289 -311 323
rect -277 289 -265 323
rect -323 255 -265 289
rect -323 221 -311 255
rect -277 221 -265 255
rect -323 187 -265 221
rect -323 153 -311 187
rect -277 153 -265 187
rect -323 119 -265 153
rect -323 85 -311 119
rect -277 85 -265 119
rect -323 51 -265 85
rect -323 17 -311 51
rect -277 17 -265 51
rect -323 -17 -265 17
rect -323 -51 -311 -17
rect -277 -51 -265 -17
rect -323 -85 -265 -51
rect -323 -119 -311 -85
rect -277 -119 -265 -85
rect -323 -153 -265 -119
rect -323 -187 -311 -153
rect -277 -187 -265 -153
rect -323 -221 -265 -187
rect -323 -255 -311 -221
rect -277 -255 -265 -221
rect -323 -289 -265 -255
rect -323 -323 -311 -289
rect -277 -323 -265 -289
rect -323 -357 -265 -323
rect -323 -391 -311 -357
rect -277 -391 -265 -357
rect -323 -425 -265 -391
rect -323 -459 -311 -425
rect -277 -459 -265 -425
rect -323 -500 -265 -459
rect -225 459 -167 500
rect -225 425 -213 459
rect -179 425 -167 459
rect -225 391 -167 425
rect -225 357 -213 391
rect -179 357 -167 391
rect -225 323 -167 357
rect -225 289 -213 323
rect -179 289 -167 323
rect -225 255 -167 289
rect -225 221 -213 255
rect -179 221 -167 255
rect -225 187 -167 221
rect -225 153 -213 187
rect -179 153 -167 187
rect -225 119 -167 153
rect -225 85 -213 119
rect -179 85 -167 119
rect -225 51 -167 85
rect -225 17 -213 51
rect -179 17 -167 51
rect -225 -17 -167 17
rect -225 -51 -213 -17
rect -179 -51 -167 -17
rect -225 -85 -167 -51
rect -225 -119 -213 -85
rect -179 -119 -167 -85
rect -225 -153 -167 -119
rect -225 -187 -213 -153
rect -179 -187 -167 -153
rect -225 -221 -167 -187
rect -225 -255 -213 -221
rect -179 -255 -167 -221
rect -225 -289 -167 -255
rect -225 -323 -213 -289
rect -179 -323 -167 -289
rect -225 -357 -167 -323
rect -225 -391 -213 -357
rect -179 -391 -167 -357
rect -225 -425 -167 -391
rect -225 -459 -213 -425
rect -179 -459 -167 -425
rect -225 -500 -167 -459
rect -127 459 -69 500
rect -127 425 -115 459
rect -81 425 -69 459
rect -127 391 -69 425
rect -127 357 -115 391
rect -81 357 -69 391
rect -127 323 -69 357
rect -127 289 -115 323
rect -81 289 -69 323
rect -127 255 -69 289
rect -127 221 -115 255
rect -81 221 -69 255
rect -127 187 -69 221
rect -127 153 -115 187
rect -81 153 -69 187
rect -127 119 -69 153
rect -127 85 -115 119
rect -81 85 -69 119
rect -127 51 -69 85
rect -127 17 -115 51
rect -81 17 -69 51
rect -127 -17 -69 17
rect -127 -51 -115 -17
rect -81 -51 -69 -17
rect -127 -85 -69 -51
rect -127 -119 -115 -85
rect -81 -119 -69 -85
rect -127 -153 -69 -119
rect -127 -187 -115 -153
rect -81 -187 -69 -153
rect -127 -221 -69 -187
rect -127 -255 -115 -221
rect -81 -255 -69 -221
rect -127 -289 -69 -255
rect -127 -323 -115 -289
rect -81 -323 -69 -289
rect -127 -357 -69 -323
rect -127 -391 -115 -357
rect -81 -391 -69 -357
rect -127 -425 -69 -391
rect -127 -459 -115 -425
rect -81 -459 -69 -425
rect -127 -500 -69 -459
rect -29 459 29 500
rect -29 425 -17 459
rect 17 425 29 459
rect -29 391 29 425
rect -29 357 -17 391
rect 17 357 29 391
rect -29 323 29 357
rect -29 289 -17 323
rect 17 289 29 323
rect -29 255 29 289
rect -29 221 -17 255
rect 17 221 29 255
rect -29 187 29 221
rect -29 153 -17 187
rect 17 153 29 187
rect -29 119 29 153
rect -29 85 -17 119
rect 17 85 29 119
rect -29 51 29 85
rect -29 17 -17 51
rect 17 17 29 51
rect -29 -17 29 17
rect -29 -51 -17 -17
rect 17 -51 29 -17
rect -29 -85 29 -51
rect -29 -119 -17 -85
rect 17 -119 29 -85
rect -29 -153 29 -119
rect -29 -187 -17 -153
rect 17 -187 29 -153
rect -29 -221 29 -187
rect -29 -255 -17 -221
rect 17 -255 29 -221
rect -29 -289 29 -255
rect -29 -323 -17 -289
rect 17 -323 29 -289
rect -29 -357 29 -323
rect -29 -391 -17 -357
rect 17 -391 29 -357
rect -29 -425 29 -391
rect -29 -459 -17 -425
rect 17 -459 29 -425
rect -29 -500 29 -459
rect 69 459 127 500
rect 69 425 81 459
rect 115 425 127 459
rect 69 391 127 425
rect 69 357 81 391
rect 115 357 127 391
rect 69 323 127 357
rect 69 289 81 323
rect 115 289 127 323
rect 69 255 127 289
rect 69 221 81 255
rect 115 221 127 255
rect 69 187 127 221
rect 69 153 81 187
rect 115 153 127 187
rect 69 119 127 153
rect 69 85 81 119
rect 115 85 127 119
rect 69 51 127 85
rect 69 17 81 51
rect 115 17 127 51
rect 69 -17 127 17
rect 69 -51 81 -17
rect 115 -51 127 -17
rect 69 -85 127 -51
rect 69 -119 81 -85
rect 115 -119 127 -85
rect 69 -153 127 -119
rect 69 -187 81 -153
rect 115 -187 127 -153
rect 69 -221 127 -187
rect 69 -255 81 -221
rect 115 -255 127 -221
rect 69 -289 127 -255
rect 69 -323 81 -289
rect 115 -323 127 -289
rect 69 -357 127 -323
rect 69 -391 81 -357
rect 115 -391 127 -357
rect 69 -425 127 -391
rect 69 -459 81 -425
rect 115 -459 127 -425
rect 69 -500 127 -459
rect 167 459 225 500
rect 167 425 179 459
rect 213 425 225 459
rect 167 391 225 425
rect 167 357 179 391
rect 213 357 225 391
rect 167 323 225 357
rect 167 289 179 323
rect 213 289 225 323
rect 167 255 225 289
rect 167 221 179 255
rect 213 221 225 255
rect 167 187 225 221
rect 167 153 179 187
rect 213 153 225 187
rect 167 119 225 153
rect 167 85 179 119
rect 213 85 225 119
rect 167 51 225 85
rect 167 17 179 51
rect 213 17 225 51
rect 167 -17 225 17
rect 167 -51 179 -17
rect 213 -51 225 -17
rect 167 -85 225 -51
rect 167 -119 179 -85
rect 213 -119 225 -85
rect 167 -153 225 -119
rect 167 -187 179 -153
rect 213 -187 225 -153
rect 167 -221 225 -187
rect 167 -255 179 -221
rect 213 -255 225 -221
rect 167 -289 225 -255
rect 167 -323 179 -289
rect 213 -323 225 -289
rect 167 -357 225 -323
rect 167 -391 179 -357
rect 213 -391 225 -357
rect 167 -425 225 -391
rect 167 -459 179 -425
rect 213 -459 225 -425
rect 167 -500 225 -459
rect 265 459 323 500
rect 265 425 277 459
rect 311 425 323 459
rect 265 391 323 425
rect 265 357 277 391
rect 311 357 323 391
rect 265 323 323 357
rect 265 289 277 323
rect 311 289 323 323
rect 265 255 323 289
rect 265 221 277 255
rect 311 221 323 255
rect 265 187 323 221
rect 265 153 277 187
rect 311 153 323 187
rect 265 119 323 153
rect 265 85 277 119
rect 311 85 323 119
rect 265 51 323 85
rect 265 17 277 51
rect 311 17 323 51
rect 265 -17 323 17
rect 265 -51 277 -17
rect 311 -51 323 -17
rect 265 -85 323 -51
rect 265 -119 277 -85
rect 311 -119 323 -85
rect 265 -153 323 -119
rect 265 -187 277 -153
rect 311 -187 323 -153
rect 265 -221 323 -187
rect 265 -255 277 -221
rect 311 -255 323 -221
rect 265 -289 323 -255
rect 265 -323 277 -289
rect 311 -323 323 -289
rect 265 -357 323 -323
rect 265 -391 277 -357
rect 311 -391 323 -357
rect 265 -425 323 -391
rect 265 -459 277 -425
rect 311 -459 323 -425
rect 265 -500 323 -459
rect 363 459 421 500
rect 363 425 375 459
rect 409 425 421 459
rect 363 391 421 425
rect 363 357 375 391
rect 409 357 421 391
rect 363 323 421 357
rect 363 289 375 323
rect 409 289 421 323
rect 363 255 421 289
rect 363 221 375 255
rect 409 221 421 255
rect 363 187 421 221
rect 363 153 375 187
rect 409 153 421 187
rect 363 119 421 153
rect 363 85 375 119
rect 409 85 421 119
rect 363 51 421 85
rect 363 17 375 51
rect 409 17 421 51
rect 363 -17 421 17
rect 363 -51 375 -17
rect 409 -51 421 -17
rect 363 -85 421 -51
rect 363 -119 375 -85
rect 409 -119 421 -85
rect 363 -153 421 -119
rect 363 -187 375 -153
rect 409 -187 421 -153
rect 363 -221 421 -187
rect 363 -255 375 -221
rect 409 -255 421 -221
rect 363 -289 421 -255
rect 363 -323 375 -289
rect 409 -323 421 -289
rect 363 -357 421 -323
rect 363 -391 375 -357
rect 409 -391 421 -357
rect 363 -425 421 -391
rect 363 -459 375 -425
rect 409 -459 421 -425
rect 363 -500 421 -459
<< ndiffc >>
rect -409 425 -375 459
rect -409 357 -375 391
rect -409 289 -375 323
rect -409 221 -375 255
rect -409 153 -375 187
rect -409 85 -375 119
rect -409 17 -375 51
rect -409 -51 -375 -17
rect -409 -119 -375 -85
rect -409 -187 -375 -153
rect -409 -255 -375 -221
rect -409 -323 -375 -289
rect -409 -391 -375 -357
rect -409 -459 -375 -425
rect -311 425 -277 459
rect -311 357 -277 391
rect -311 289 -277 323
rect -311 221 -277 255
rect -311 153 -277 187
rect -311 85 -277 119
rect -311 17 -277 51
rect -311 -51 -277 -17
rect -311 -119 -277 -85
rect -311 -187 -277 -153
rect -311 -255 -277 -221
rect -311 -323 -277 -289
rect -311 -391 -277 -357
rect -311 -459 -277 -425
rect -213 425 -179 459
rect -213 357 -179 391
rect -213 289 -179 323
rect -213 221 -179 255
rect -213 153 -179 187
rect -213 85 -179 119
rect -213 17 -179 51
rect -213 -51 -179 -17
rect -213 -119 -179 -85
rect -213 -187 -179 -153
rect -213 -255 -179 -221
rect -213 -323 -179 -289
rect -213 -391 -179 -357
rect -213 -459 -179 -425
rect -115 425 -81 459
rect -115 357 -81 391
rect -115 289 -81 323
rect -115 221 -81 255
rect -115 153 -81 187
rect -115 85 -81 119
rect -115 17 -81 51
rect -115 -51 -81 -17
rect -115 -119 -81 -85
rect -115 -187 -81 -153
rect -115 -255 -81 -221
rect -115 -323 -81 -289
rect -115 -391 -81 -357
rect -115 -459 -81 -425
rect -17 425 17 459
rect -17 357 17 391
rect -17 289 17 323
rect -17 221 17 255
rect -17 153 17 187
rect -17 85 17 119
rect -17 17 17 51
rect -17 -51 17 -17
rect -17 -119 17 -85
rect -17 -187 17 -153
rect -17 -255 17 -221
rect -17 -323 17 -289
rect -17 -391 17 -357
rect -17 -459 17 -425
rect 81 425 115 459
rect 81 357 115 391
rect 81 289 115 323
rect 81 221 115 255
rect 81 153 115 187
rect 81 85 115 119
rect 81 17 115 51
rect 81 -51 115 -17
rect 81 -119 115 -85
rect 81 -187 115 -153
rect 81 -255 115 -221
rect 81 -323 115 -289
rect 81 -391 115 -357
rect 81 -459 115 -425
rect 179 425 213 459
rect 179 357 213 391
rect 179 289 213 323
rect 179 221 213 255
rect 179 153 213 187
rect 179 85 213 119
rect 179 17 213 51
rect 179 -51 213 -17
rect 179 -119 213 -85
rect 179 -187 213 -153
rect 179 -255 213 -221
rect 179 -323 213 -289
rect 179 -391 213 -357
rect 179 -459 213 -425
rect 277 425 311 459
rect 277 357 311 391
rect 277 289 311 323
rect 277 221 311 255
rect 277 153 311 187
rect 277 85 311 119
rect 277 17 311 51
rect 277 -51 311 -17
rect 277 -119 311 -85
rect 277 -187 311 -153
rect 277 -255 311 -221
rect 277 -323 311 -289
rect 277 -391 311 -357
rect 277 -459 311 -425
rect 375 425 409 459
rect 375 357 409 391
rect 375 289 409 323
rect 375 221 409 255
rect 375 153 409 187
rect 375 85 409 119
rect 375 17 409 51
rect 375 -51 409 -17
rect 375 -119 409 -85
rect 375 -187 409 -153
rect 375 -255 409 -221
rect 375 -323 409 -289
rect 375 -391 409 -357
rect 375 -459 409 -425
<< poly >>
rect 166 732 232 748
rect 166 698 182 732
rect 216 698 232 732
rect 166 682 232 698
rect 362 732 428 748
rect 362 698 378 732
rect 412 698 428 732
rect 362 682 428 698
rect 177 614 217 682
rect 373 614 413 682
rect -363 574 419 614
rect -363 500 -323 574
rect -265 500 -225 574
rect -167 500 -127 574
rect -69 500 -29 574
rect 29 500 69 574
rect 127 500 167 574
rect 225 500 265 574
rect 323 500 363 574
rect -363 -526 -323 -500
rect -265 -526 -225 -500
rect -167 -526 -127 -500
rect -69 -526 -29 -500
rect 29 -526 69 -500
rect 127 -526 167 -500
rect 225 -526 265 -500
rect 323 -526 363 -500
<< polycont >>
rect 182 698 216 732
rect 378 698 412 732
<< locali >>
rect 77 698 182 732
rect 216 698 232 732
rect 362 698 378 732
rect 412 698 428 732
rect 77 612 111 698
rect -311 578 311 612
rect -409 485 -375 506
rect -409 413 -375 425
rect -409 341 -375 357
rect -409 269 -375 289
rect -409 197 -375 221
rect -409 125 -375 153
rect -409 53 -375 85
rect -409 -17 -375 17
rect -409 -85 -375 -53
rect -409 -153 -375 -125
rect -409 -221 -375 -197
rect -409 -289 -375 -269
rect -409 -357 -375 -341
rect -409 -425 -375 -413
rect -409 -504 -375 -485
rect -311 485 -277 578
rect -311 413 -277 425
rect -311 341 -277 357
rect -311 269 -277 289
rect -311 197 -277 221
rect -311 125 -277 153
rect -311 53 -277 85
rect -311 -17 -277 17
rect -311 -85 -277 -53
rect -311 -153 -277 -125
rect -311 -221 -277 -197
rect -311 -289 -277 -269
rect -311 -357 -277 -341
rect -311 -425 -277 -413
rect -311 -506 -277 -485
rect -213 485 -179 502
rect -213 413 -179 425
rect -213 341 -179 357
rect -213 269 -179 289
rect -213 197 -179 221
rect -213 125 -179 153
rect -213 53 -179 85
rect -213 -17 -179 17
rect -213 -85 -179 -53
rect -213 -153 -179 -125
rect -213 -221 -179 -197
rect -213 -289 -179 -269
rect -213 -357 -179 -341
rect -213 -425 -179 -413
rect -213 -504 -179 -485
rect -115 485 -81 578
rect -115 413 -81 425
rect -115 341 -81 357
rect -115 269 -81 289
rect -115 197 -81 221
rect -115 125 -81 153
rect -115 53 -81 85
rect -115 -17 -81 17
rect -115 -85 -81 -53
rect -115 -153 -81 -125
rect -115 -221 -81 -197
rect -115 -289 -81 -269
rect -115 -357 -81 -341
rect -115 -425 -81 -413
rect -115 -506 -81 -485
rect -17 485 17 502
rect -17 413 17 425
rect -17 341 17 357
rect -17 269 17 289
rect -17 197 17 221
rect -17 125 17 153
rect -17 53 17 85
rect -17 -17 17 17
rect -17 -85 17 -53
rect -17 -153 17 -125
rect -17 -221 17 -197
rect -17 -289 17 -269
rect -17 -357 17 -341
rect -17 -425 17 -413
rect -17 -504 17 -485
rect 81 485 115 578
rect 81 413 115 425
rect 81 341 115 357
rect 81 269 115 289
rect 81 197 115 221
rect 81 125 115 153
rect 81 53 115 85
rect 81 -17 115 17
rect 81 -85 115 -53
rect 81 -153 115 -125
rect 81 -221 115 -197
rect 81 -289 115 -269
rect 81 -357 115 -341
rect 81 -425 115 -413
rect 81 -506 115 -485
rect 179 485 213 502
rect 179 413 213 425
rect 179 341 213 357
rect 179 269 213 289
rect 179 197 213 221
rect 179 125 213 153
rect 179 53 213 85
rect 179 -17 213 17
rect 179 -85 213 -53
rect 179 -153 213 -125
rect 179 -221 213 -197
rect 179 -289 213 -269
rect 179 -357 213 -341
rect 179 -425 213 -413
rect 179 -504 213 -485
rect 277 485 311 578
rect 277 413 311 425
rect 277 341 311 357
rect 277 269 311 289
rect 277 197 311 221
rect 277 125 311 153
rect 277 53 311 85
rect 277 -17 311 17
rect 277 -85 311 -53
rect 277 -153 311 -125
rect 277 -221 311 -197
rect 277 -289 311 -269
rect 277 -357 311 -341
rect 277 -425 311 -413
rect 277 -506 311 -485
rect 375 485 409 504
rect 375 413 409 425
rect 375 341 409 357
rect 375 269 409 289
rect 375 197 409 221
rect 375 125 409 153
rect 375 53 409 85
rect 375 -17 409 17
rect 375 -85 409 -53
rect 375 -153 409 -125
rect 375 -221 409 -197
rect 375 -289 409 -269
rect 375 -357 409 -341
rect 375 -425 409 -413
rect 375 -504 409 -485
rect -311 -618 313 -584
<< viali >>
rect 182 698 216 732
rect 378 698 412 732
rect -409 459 -375 485
rect -409 451 -375 459
rect -409 391 -375 413
rect -409 379 -375 391
rect -409 323 -375 341
rect -409 307 -375 323
rect -409 255 -375 269
rect -409 235 -375 255
rect -409 187 -375 197
rect -409 163 -375 187
rect -409 119 -375 125
rect -409 91 -375 119
rect -409 51 -375 53
rect -409 19 -375 51
rect -409 -51 -375 -19
rect -409 -53 -375 -51
rect -409 -119 -375 -91
rect -409 -125 -375 -119
rect -409 -187 -375 -163
rect -409 -197 -375 -187
rect -409 -255 -375 -235
rect -409 -269 -375 -255
rect -409 -323 -375 -307
rect -409 -341 -375 -323
rect -409 -391 -375 -379
rect -409 -413 -375 -391
rect -409 -459 -375 -451
rect -409 -485 -375 -459
rect -311 459 -277 485
rect -311 451 -277 459
rect -311 391 -277 413
rect -311 379 -277 391
rect -311 323 -277 341
rect -311 307 -277 323
rect -311 255 -277 269
rect -311 235 -277 255
rect -311 187 -277 197
rect -311 163 -277 187
rect -311 119 -277 125
rect -311 91 -277 119
rect -311 51 -277 53
rect -311 19 -277 51
rect -311 -51 -277 -19
rect -311 -53 -277 -51
rect -311 -119 -277 -91
rect -311 -125 -277 -119
rect -311 -187 -277 -163
rect -311 -197 -277 -187
rect -311 -255 -277 -235
rect -311 -269 -277 -255
rect -311 -323 -277 -307
rect -311 -341 -277 -323
rect -311 -391 -277 -379
rect -311 -413 -277 -391
rect -311 -459 -277 -451
rect -311 -485 -277 -459
rect -213 459 -179 485
rect -213 451 -179 459
rect -213 391 -179 413
rect -213 379 -179 391
rect -213 323 -179 341
rect -213 307 -179 323
rect -213 255 -179 269
rect -213 235 -179 255
rect -213 187 -179 197
rect -213 163 -179 187
rect -213 119 -179 125
rect -213 91 -179 119
rect -213 51 -179 53
rect -213 19 -179 51
rect -213 -51 -179 -19
rect -213 -53 -179 -51
rect -213 -119 -179 -91
rect -213 -125 -179 -119
rect -213 -187 -179 -163
rect -213 -197 -179 -187
rect -213 -255 -179 -235
rect -213 -269 -179 -255
rect -213 -323 -179 -307
rect -213 -341 -179 -323
rect -213 -391 -179 -379
rect -213 -413 -179 -391
rect -213 -459 -179 -451
rect -213 -485 -179 -459
rect -115 459 -81 485
rect -115 451 -81 459
rect -115 391 -81 413
rect -115 379 -81 391
rect -115 323 -81 341
rect -115 307 -81 323
rect -115 255 -81 269
rect -115 235 -81 255
rect -115 187 -81 197
rect -115 163 -81 187
rect -115 119 -81 125
rect -115 91 -81 119
rect -115 51 -81 53
rect -115 19 -81 51
rect -115 -51 -81 -19
rect -115 -53 -81 -51
rect -115 -119 -81 -91
rect -115 -125 -81 -119
rect -115 -187 -81 -163
rect -115 -197 -81 -187
rect -115 -255 -81 -235
rect -115 -269 -81 -255
rect -115 -323 -81 -307
rect -115 -341 -81 -323
rect -115 -391 -81 -379
rect -115 -413 -81 -391
rect -115 -459 -81 -451
rect -115 -485 -81 -459
rect -17 459 17 485
rect -17 451 17 459
rect -17 391 17 413
rect -17 379 17 391
rect -17 323 17 341
rect -17 307 17 323
rect -17 255 17 269
rect -17 235 17 255
rect -17 187 17 197
rect -17 163 17 187
rect -17 119 17 125
rect -17 91 17 119
rect -17 51 17 53
rect -17 19 17 51
rect -17 -51 17 -19
rect -17 -53 17 -51
rect -17 -119 17 -91
rect -17 -125 17 -119
rect -17 -187 17 -163
rect -17 -197 17 -187
rect -17 -255 17 -235
rect -17 -269 17 -255
rect -17 -323 17 -307
rect -17 -341 17 -323
rect -17 -391 17 -379
rect -17 -413 17 -391
rect -17 -459 17 -451
rect -17 -485 17 -459
rect 81 459 115 485
rect 81 451 115 459
rect 81 391 115 413
rect 81 379 115 391
rect 81 323 115 341
rect 81 307 115 323
rect 81 255 115 269
rect 81 235 115 255
rect 81 187 115 197
rect 81 163 115 187
rect 81 119 115 125
rect 81 91 115 119
rect 81 51 115 53
rect 81 19 115 51
rect 81 -51 115 -19
rect 81 -53 115 -51
rect 81 -119 115 -91
rect 81 -125 115 -119
rect 81 -187 115 -163
rect 81 -197 115 -187
rect 81 -255 115 -235
rect 81 -269 115 -255
rect 81 -323 115 -307
rect 81 -341 115 -323
rect 81 -391 115 -379
rect 81 -413 115 -391
rect 81 -459 115 -451
rect 81 -485 115 -459
rect 179 459 213 485
rect 179 451 213 459
rect 179 391 213 413
rect 179 379 213 391
rect 179 323 213 341
rect 179 307 213 323
rect 179 255 213 269
rect 179 235 213 255
rect 179 187 213 197
rect 179 163 213 187
rect 179 119 213 125
rect 179 91 213 119
rect 179 51 213 53
rect 179 19 213 51
rect 179 -51 213 -19
rect 179 -53 213 -51
rect 179 -119 213 -91
rect 179 -125 213 -119
rect 179 -187 213 -163
rect 179 -197 213 -187
rect 179 -255 213 -235
rect 179 -269 213 -255
rect 179 -323 213 -307
rect 179 -341 213 -323
rect 179 -391 213 -379
rect 179 -413 213 -391
rect 179 -459 213 -451
rect 179 -485 213 -459
rect 277 459 311 485
rect 277 451 311 459
rect 277 391 311 413
rect 277 379 311 391
rect 277 323 311 341
rect 277 307 311 323
rect 277 255 311 269
rect 277 235 311 255
rect 277 187 311 197
rect 277 163 311 187
rect 277 119 311 125
rect 277 91 311 119
rect 277 51 311 53
rect 277 19 311 51
rect 277 -51 311 -19
rect 277 -53 311 -51
rect 277 -119 311 -91
rect 277 -125 311 -119
rect 277 -187 311 -163
rect 277 -197 311 -187
rect 277 -255 311 -235
rect 277 -269 311 -255
rect 277 -323 311 -307
rect 277 -341 311 -323
rect 277 -391 311 -379
rect 277 -413 311 -391
rect 277 -459 311 -451
rect 277 -485 311 -459
rect 375 459 409 485
rect 375 451 409 459
rect 375 391 409 413
rect 375 379 409 391
rect 375 323 409 341
rect 375 307 409 323
rect 375 255 409 269
rect 375 235 409 255
rect 375 187 409 197
rect 375 163 409 187
rect 375 119 409 125
rect 375 91 409 119
rect 375 51 409 53
rect 375 19 409 51
rect 375 -51 409 -19
rect 375 -53 409 -51
rect 375 -119 409 -91
rect 375 -125 409 -119
rect 375 -187 409 -163
rect 375 -197 409 -187
rect 375 -255 409 -235
rect 375 -269 409 -255
rect 375 -323 409 -307
rect 375 -341 409 -323
rect 375 -391 409 -379
rect 375 -413 409 -391
rect 375 -459 409 -451
rect 375 -485 409 -459
<< metal1 >>
rect 170 732 228 738
rect 170 698 182 732
rect 216 698 228 732
rect 170 692 228 698
rect 366 732 424 738
rect 366 698 378 732
rect 412 698 424 732
rect 366 692 424 698
rect -415 485 -369 500
rect -415 451 -409 485
rect -375 451 -369 485
rect -415 413 -369 451
rect -415 379 -409 413
rect -375 379 -369 413
rect -415 341 -369 379
rect -415 307 -409 341
rect -375 307 -369 341
rect -415 269 -369 307
rect -415 235 -409 269
rect -375 235 -369 269
rect -415 197 -369 235
rect -415 163 -409 197
rect -375 163 -369 197
rect -415 125 -369 163
rect -415 91 -409 125
rect -375 91 -369 125
rect -415 53 -369 91
rect -415 19 -409 53
rect -375 19 -369 53
rect -415 -19 -369 19
rect -415 -53 -409 -19
rect -375 -53 -369 -19
rect -415 -91 -369 -53
rect -415 -125 -409 -91
rect -375 -125 -369 -91
rect -415 -163 -369 -125
rect -415 -197 -409 -163
rect -375 -197 -369 -163
rect -415 -235 -369 -197
rect -415 -269 -409 -235
rect -375 -269 -369 -235
rect -415 -307 -369 -269
rect -415 -341 -409 -307
rect -375 -341 -369 -307
rect -415 -379 -369 -341
rect -415 -413 -409 -379
rect -375 -413 -369 -379
rect -415 -451 -369 -413
rect -415 -485 -409 -451
rect -375 -485 -369 -451
rect -415 -500 -369 -485
rect -317 485 -271 500
rect -317 451 -311 485
rect -277 451 -271 485
rect -317 413 -271 451
rect -317 379 -311 413
rect -277 379 -271 413
rect -317 341 -271 379
rect -317 307 -311 341
rect -277 307 -271 341
rect -317 269 -271 307
rect -317 235 -311 269
rect -277 235 -271 269
rect -317 197 -271 235
rect -317 163 -311 197
rect -277 163 -271 197
rect -317 125 -271 163
rect -317 91 -311 125
rect -277 91 -271 125
rect -317 53 -271 91
rect -317 19 -311 53
rect -277 19 -271 53
rect -317 -19 -271 19
rect -317 -53 -311 -19
rect -277 -53 -271 -19
rect -317 -91 -271 -53
rect -317 -125 -311 -91
rect -277 -125 -271 -91
rect -317 -163 -271 -125
rect -317 -197 -311 -163
rect -277 -197 -271 -163
rect -317 -235 -271 -197
rect -317 -269 -311 -235
rect -277 -269 -271 -235
rect -317 -307 -271 -269
rect -317 -341 -311 -307
rect -277 -341 -271 -307
rect -317 -379 -271 -341
rect -317 -413 -311 -379
rect -277 -413 -271 -379
rect -317 -451 -271 -413
rect -317 -485 -311 -451
rect -277 -485 -271 -451
rect -317 -500 -271 -485
rect -219 485 -173 500
rect -219 451 -213 485
rect -179 451 -173 485
rect -219 413 -173 451
rect -219 379 -213 413
rect -179 379 -173 413
rect -219 341 -173 379
rect -219 307 -213 341
rect -179 307 -173 341
rect -219 269 -173 307
rect -219 235 -213 269
rect -179 235 -173 269
rect -219 197 -173 235
rect -219 163 -213 197
rect -179 163 -173 197
rect -219 125 -173 163
rect -219 91 -213 125
rect -179 91 -173 125
rect -219 53 -173 91
rect -219 19 -213 53
rect -179 19 -173 53
rect -219 -19 -173 19
rect -219 -53 -213 -19
rect -179 -53 -173 -19
rect -219 -91 -173 -53
rect -219 -125 -213 -91
rect -179 -125 -173 -91
rect -219 -163 -173 -125
rect -219 -197 -213 -163
rect -179 -197 -173 -163
rect -219 -235 -173 -197
rect -219 -269 -213 -235
rect -179 -269 -173 -235
rect -219 -307 -173 -269
rect -219 -341 -213 -307
rect -179 -341 -173 -307
rect -219 -379 -173 -341
rect -219 -413 -213 -379
rect -179 -413 -173 -379
rect -219 -451 -173 -413
rect -219 -485 -213 -451
rect -179 -485 -173 -451
rect -219 -500 -173 -485
rect -121 485 -75 500
rect -121 451 -115 485
rect -81 451 -75 485
rect -121 413 -75 451
rect -121 379 -115 413
rect -81 379 -75 413
rect -121 341 -75 379
rect -121 307 -115 341
rect -81 307 -75 341
rect -121 269 -75 307
rect -121 235 -115 269
rect -81 235 -75 269
rect -121 197 -75 235
rect -121 163 -115 197
rect -81 163 -75 197
rect -121 125 -75 163
rect -121 91 -115 125
rect -81 91 -75 125
rect -121 53 -75 91
rect -121 19 -115 53
rect -81 19 -75 53
rect -121 -19 -75 19
rect -121 -53 -115 -19
rect -81 -53 -75 -19
rect -121 -91 -75 -53
rect -121 -125 -115 -91
rect -81 -125 -75 -91
rect -121 -163 -75 -125
rect -121 -197 -115 -163
rect -81 -197 -75 -163
rect -121 -235 -75 -197
rect -121 -269 -115 -235
rect -81 -269 -75 -235
rect -121 -307 -75 -269
rect -121 -341 -115 -307
rect -81 -341 -75 -307
rect -121 -379 -75 -341
rect -121 -413 -115 -379
rect -81 -413 -75 -379
rect -121 -451 -75 -413
rect -121 -485 -115 -451
rect -81 -485 -75 -451
rect -121 -500 -75 -485
rect -23 485 23 500
rect -23 451 -17 485
rect 17 451 23 485
rect -23 413 23 451
rect -23 379 -17 413
rect 17 379 23 413
rect -23 341 23 379
rect -23 307 -17 341
rect 17 307 23 341
rect -23 269 23 307
rect -23 235 -17 269
rect 17 235 23 269
rect -23 197 23 235
rect -23 163 -17 197
rect 17 163 23 197
rect -23 125 23 163
rect -23 91 -17 125
rect 17 91 23 125
rect -23 53 23 91
rect -23 19 -17 53
rect 17 19 23 53
rect -23 -19 23 19
rect -23 -53 -17 -19
rect 17 -53 23 -19
rect -23 -91 23 -53
rect -23 -125 -17 -91
rect 17 -125 23 -91
rect -23 -163 23 -125
rect -23 -197 -17 -163
rect 17 -197 23 -163
rect -23 -235 23 -197
rect -23 -269 -17 -235
rect 17 -269 23 -235
rect -23 -307 23 -269
rect -23 -341 -17 -307
rect 17 -341 23 -307
rect -23 -379 23 -341
rect -23 -413 -17 -379
rect 17 -413 23 -379
rect -23 -451 23 -413
rect -23 -485 -17 -451
rect 17 -485 23 -451
rect -23 -500 23 -485
rect 75 485 121 500
rect 75 451 81 485
rect 115 451 121 485
rect 75 413 121 451
rect 75 379 81 413
rect 115 379 121 413
rect 75 341 121 379
rect 75 307 81 341
rect 115 307 121 341
rect 75 269 121 307
rect 75 235 81 269
rect 115 235 121 269
rect 75 197 121 235
rect 75 163 81 197
rect 115 163 121 197
rect 75 125 121 163
rect 75 91 81 125
rect 115 91 121 125
rect 75 53 121 91
rect 75 19 81 53
rect 115 19 121 53
rect 75 -19 121 19
rect 75 -53 81 -19
rect 115 -53 121 -19
rect 75 -91 121 -53
rect 75 -125 81 -91
rect 115 -125 121 -91
rect 75 -163 121 -125
rect 75 -197 81 -163
rect 115 -197 121 -163
rect 75 -235 121 -197
rect 75 -269 81 -235
rect 115 -269 121 -235
rect 75 -307 121 -269
rect 75 -341 81 -307
rect 115 -341 121 -307
rect 75 -379 121 -341
rect 75 -413 81 -379
rect 115 -413 121 -379
rect 75 -451 121 -413
rect 75 -485 81 -451
rect 115 -485 121 -451
rect 75 -500 121 -485
rect 173 485 219 500
rect 173 451 179 485
rect 213 451 219 485
rect 173 413 219 451
rect 173 379 179 413
rect 213 379 219 413
rect 173 341 219 379
rect 173 307 179 341
rect 213 307 219 341
rect 173 269 219 307
rect 173 235 179 269
rect 213 235 219 269
rect 173 197 219 235
rect 173 163 179 197
rect 213 163 219 197
rect 173 125 219 163
rect 173 91 179 125
rect 213 91 219 125
rect 173 53 219 91
rect 173 19 179 53
rect 213 19 219 53
rect 173 -19 219 19
rect 173 -53 179 -19
rect 213 -53 219 -19
rect 173 -91 219 -53
rect 173 -125 179 -91
rect 213 -125 219 -91
rect 173 -163 219 -125
rect 173 -197 179 -163
rect 213 -197 219 -163
rect 173 -235 219 -197
rect 173 -269 179 -235
rect 213 -269 219 -235
rect 173 -307 219 -269
rect 173 -341 179 -307
rect 213 -341 219 -307
rect 173 -379 219 -341
rect 173 -413 179 -379
rect 213 -413 219 -379
rect 173 -451 219 -413
rect 173 -485 179 -451
rect 213 -485 219 -451
rect 173 -500 219 -485
rect 271 485 317 500
rect 271 451 277 485
rect 311 451 317 485
rect 271 413 317 451
rect 271 379 277 413
rect 311 379 317 413
rect 271 341 317 379
rect 271 307 277 341
rect 311 307 317 341
rect 271 269 317 307
rect 271 235 277 269
rect 311 235 317 269
rect 271 197 317 235
rect 271 163 277 197
rect 311 163 317 197
rect 271 125 317 163
rect 271 91 277 125
rect 311 91 317 125
rect 271 53 317 91
rect 271 19 277 53
rect 311 19 317 53
rect 271 -19 317 19
rect 271 -53 277 -19
rect 311 -53 317 -19
rect 271 -91 317 -53
rect 271 -125 277 -91
rect 311 -125 317 -91
rect 271 -163 317 -125
rect 271 -197 277 -163
rect 311 -197 317 -163
rect 271 -235 317 -197
rect 271 -269 277 -235
rect 311 -269 317 -235
rect 271 -307 317 -269
rect 271 -341 277 -307
rect 311 -341 317 -307
rect 271 -379 317 -341
rect 271 -413 277 -379
rect 311 -413 317 -379
rect 271 -451 317 -413
rect 271 -485 277 -451
rect 311 -485 317 -451
rect 271 -500 317 -485
rect 369 485 415 500
rect 369 451 375 485
rect 409 451 415 485
rect 369 413 415 451
rect 369 379 375 413
rect 409 379 415 413
rect 369 341 415 379
rect 369 307 375 341
rect 409 307 415 341
rect 369 269 415 307
rect 369 235 375 269
rect 409 235 415 269
rect 369 197 415 235
rect 369 163 375 197
rect 409 163 415 197
rect 369 125 415 163
rect 369 91 375 125
rect 409 91 415 125
rect 369 53 415 91
rect 369 19 375 53
rect 409 19 415 53
rect 369 -19 415 19
rect 369 -53 375 -19
rect 409 -53 415 -19
rect 369 -91 415 -53
rect 369 -125 375 -91
rect 409 -125 415 -91
rect 369 -163 415 -125
rect 369 -197 375 -163
rect 409 -197 415 -163
rect 369 -235 415 -197
rect 369 -269 375 -235
rect 409 -269 415 -235
rect 369 -307 415 -269
rect 369 -341 375 -307
rect 409 -341 415 -307
rect 369 -379 415 -341
rect 369 -413 375 -379
rect 409 -413 415 -379
rect 369 -451 415 -413
rect 369 -485 375 -451
rect 409 -485 415 -451
rect 369 -500 415 -485
<< end >>
