magic
tech sky130A
magscale 1 2
timestamp 1634894729
<< nwell >>
rect -2366 7582 16048 8168
rect -2366 6926 16044 7582
rect -2366 3582 16042 6926
rect -2366 3580 -230 3582
rect 14938 3580 16030 3582
<< pwell >>
rect 15056 3502 15262 3580
rect -2426 -1250 16034 3502
<< nmos >>
rect -1636 2236 -1606 3236
rect -1540 2236 -1510 3236
rect -1444 2236 -1414 3236
rect -1348 2236 -1318 3236
rect -1252 2236 -1222 3236
rect -1156 2236 -1126 3236
rect -1060 2236 -1030 3236
rect -964 2236 -934 3236
rect 1532 1830 1562 2830
rect 1628 1830 1658 2830
rect 1724 1830 1754 2830
rect 1820 1830 1850 2830
rect 2546 2076 2646 2276
rect 4488 1814 4518 2814
rect 4584 1814 4614 2814
rect 4680 1814 4710 2814
rect 4776 1814 4806 2814
rect 5546 2076 5646 2276
rect 7518 1814 7548 2814
rect 7614 1814 7644 2814
rect 7710 1814 7740 2814
rect 7806 1814 7836 2814
rect 8546 2076 8646 2276
rect 10606 1812 10636 2812
rect 10702 1812 10732 2812
rect 10798 1812 10828 2812
rect 10894 1812 10924 2812
rect 11546 2076 11646 2276
rect 13762 1786 13792 2786
rect 13858 1786 13888 2786
rect 13954 1786 13984 2786
rect 14050 1786 14080 2786
rect 14546 2076 14646 2276
rect -1640 66 -1600 1066
rect -1542 66 -1502 1066
rect -1444 66 -1404 1066
rect -1346 66 -1306 1066
rect -1248 66 -1208 1066
rect -1150 66 -1110 1066
rect -1052 66 -1012 1066
rect -954 66 -914 1066
rect 208 268 238 1268
rect 304 268 334 1268
rect 400 268 430 1268
rect 496 268 526 1268
rect 592 268 622 1268
rect 688 268 718 1268
rect 784 268 814 1268
rect 880 268 910 1268
rect 976 268 1006 1268
rect 1072 268 1102 1268
rect 1168 268 1198 1268
rect 1264 268 1294 1268
rect 1976 268 2006 1268
rect 2072 268 2102 1268
rect 2168 268 2198 1268
rect 2264 268 2294 1268
rect 2360 268 2390 1268
rect 2456 268 2486 1268
rect 2552 268 2582 1268
rect 2648 268 2678 1268
rect 2744 268 2774 1268
rect 2840 268 2870 1268
rect 2936 268 2966 1268
rect 3164 252 3194 1252
rect 3260 252 3290 1252
rect 3356 252 3386 1252
rect 3452 252 3482 1252
rect 3548 252 3578 1252
rect 3644 252 3674 1252
rect 3740 252 3770 1252
rect 3836 252 3866 1252
rect 3932 252 3962 1252
rect 4028 252 4058 1252
rect 4124 252 4154 1252
rect 4220 252 4250 1252
rect 4932 252 4962 1252
rect 5028 252 5058 1252
rect 5124 252 5154 1252
rect 5220 252 5250 1252
rect 5316 252 5346 1252
rect 5412 252 5442 1252
rect 5508 252 5538 1252
rect 5604 252 5634 1252
rect 5700 252 5730 1252
rect 5796 252 5826 1252
rect 5892 252 5922 1252
rect 6194 252 6224 1252
rect 6290 252 6320 1252
rect 6386 252 6416 1252
rect 6482 252 6512 1252
rect 6578 252 6608 1252
rect 6674 252 6704 1252
rect 6770 252 6800 1252
rect 6866 252 6896 1252
rect 6962 252 6992 1252
rect 7058 252 7088 1252
rect 7154 252 7184 1252
rect 7250 252 7280 1252
rect 7962 252 7992 1252
rect 8058 252 8088 1252
rect 8154 252 8184 1252
rect 8250 252 8280 1252
rect 8346 252 8376 1252
rect 8442 252 8472 1252
rect 8538 252 8568 1252
rect 8634 252 8664 1252
rect 8730 252 8760 1252
rect 8826 252 8856 1252
rect 8922 252 8952 1252
rect 9282 250 9312 1250
rect 9378 250 9408 1250
rect 9474 250 9504 1250
rect 9570 250 9600 1250
rect 9666 250 9696 1250
rect 9762 250 9792 1250
rect 9858 250 9888 1250
rect 9954 250 9984 1250
rect 10050 250 10080 1250
rect 10146 250 10176 1250
rect 10242 250 10272 1250
rect 10338 250 10368 1250
rect 11050 250 11080 1250
rect 11146 250 11176 1250
rect 11242 250 11272 1250
rect 11338 250 11368 1250
rect 11434 250 11464 1250
rect 11530 250 11560 1250
rect 11626 250 11656 1250
rect 11722 250 11752 1250
rect 11818 250 11848 1250
rect 11914 250 11944 1250
rect 12010 250 12040 1250
rect 12438 224 12468 1224
rect 12534 224 12564 1224
rect 12630 224 12660 1224
rect 12726 224 12756 1224
rect 12822 224 12852 1224
rect 12918 224 12948 1224
rect 13014 224 13044 1224
rect 13110 224 13140 1224
rect 13206 224 13236 1224
rect 13302 224 13332 1224
rect 13398 224 13428 1224
rect 13494 224 13524 1224
rect 14206 224 14236 1224
rect 14302 224 14332 1224
rect 14398 224 14428 1224
rect 14494 224 14524 1224
rect 14590 224 14620 1224
rect 14686 224 14716 1224
rect 14782 224 14812 1224
rect 14878 224 14908 1224
rect 14974 224 15004 1224
rect 15070 224 15100 1224
rect 15166 224 15196 1224
rect 15468 100 15498 1300
<< pmos >>
rect -1606 4936 -1566 5936
rect -1508 4936 -1468 5936
rect -1410 4936 -1370 5936
rect -1312 4936 -1272 5936
rect -1214 4936 -1174 5936
rect -1116 4936 -1076 5936
rect -1018 4936 -978 5936
rect -920 4936 -880 5936
rect 244 5606 274 6606
rect 340 5606 370 6606
rect 436 5606 466 6606
rect 532 5606 562 6606
rect 628 5606 658 6606
rect 724 5606 754 6606
rect 820 5606 850 6606
rect 916 5606 946 6606
rect 1012 5606 1042 6606
rect 1108 5606 1138 6606
rect 1204 5606 1234 6606
rect 1300 5606 1330 6606
rect 2010 5602 2040 6602
rect 2106 5602 2136 6602
rect 2202 5602 2232 6602
rect 2298 5602 2328 6602
rect 2394 5602 2424 6602
rect 2490 5602 2520 6602
rect 2586 5602 2616 6602
rect 2682 5602 2712 6602
rect 3200 5590 3230 6590
rect 3296 5590 3326 6590
rect 3392 5590 3422 6590
rect 3488 5590 3518 6590
rect 3584 5590 3614 6590
rect 3680 5590 3710 6590
rect 3776 5590 3806 6590
rect 3872 5590 3902 6590
rect 3968 5590 3998 6590
rect 4064 5590 4094 6590
rect 4160 5590 4190 6590
rect 4256 5590 4286 6590
rect 4966 5586 4996 6586
rect 5062 5586 5092 6586
rect 5158 5586 5188 6586
rect 5254 5586 5284 6586
rect 5350 5586 5380 6586
rect 5446 5586 5476 6586
rect 5542 5586 5572 6586
rect 5638 5586 5668 6586
rect 6230 5590 6260 6590
rect 6326 5590 6356 6590
rect 6422 5590 6452 6590
rect 6518 5590 6548 6590
rect 6614 5590 6644 6590
rect 6710 5590 6740 6590
rect 6806 5590 6836 6590
rect 6902 5590 6932 6590
rect 6998 5590 7028 6590
rect 7094 5590 7124 6590
rect 7190 5590 7220 6590
rect 7286 5590 7316 6590
rect 7996 5586 8026 6586
rect 8092 5586 8122 6586
rect 8188 5586 8218 6586
rect 8284 5586 8314 6586
rect 8380 5586 8410 6586
rect 8476 5586 8506 6586
rect 8572 5586 8602 6586
rect 8668 5586 8698 6586
rect 9318 5588 9348 6588
rect 9414 5588 9444 6588
rect 9510 5588 9540 6588
rect 9606 5588 9636 6588
rect 9702 5588 9732 6588
rect 9798 5588 9828 6588
rect 9894 5588 9924 6588
rect 9990 5588 10020 6588
rect 10086 5588 10116 6588
rect 10182 5588 10212 6588
rect 10278 5588 10308 6588
rect 10374 5588 10404 6588
rect 11084 5584 11114 6584
rect 11180 5584 11210 6584
rect 11276 5584 11306 6584
rect 11372 5584 11402 6584
rect 11468 5584 11498 6584
rect 11564 5584 11594 6584
rect 11660 5584 11690 6584
rect 11756 5584 11786 6584
rect 12474 5562 12504 6562
rect 12570 5562 12600 6562
rect 12666 5562 12696 6562
rect 12762 5562 12792 6562
rect 12858 5562 12888 6562
rect 12954 5562 12984 6562
rect 13050 5562 13080 6562
rect 13146 5562 13176 6562
rect 13242 5562 13272 6562
rect 13338 5562 13368 6562
rect 13434 5562 13464 6562
rect 13530 5562 13560 6562
rect 14240 5558 14270 6558
rect 14336 5558 14366 6558
rect 14432 5558 14462 6558
rect 14528 5558 14558 6558
rect 14624 5558 14654 6558
rect 14720 5558 14750 6558
rect 14816 5558 14846 6558
rect 14912 5558 14942 6558
rect 1534 3944 1564 4944
rect 1630 3944 1660 4944
rect 1726 3944 1756 4944
rect 1822 3944 1852 4944
rect 4490 3928 4520 4928
rect 4586 3928 4616 4928
rect 4682 3928 4712 4928
rect 4778 3928 4808 4928
rect 7520 3928 7550 4928
rect 7616 3928 7646 4928
rect 7712 3928 7742 4928
rect 7808 3928 7838 4928
rect 10608 3926 10638 4926
rect 10704 3926 10734 4926
rect 10800 3926 10830 4926
rect 10896 3926 10926 4926
rect 13764 3900 13794 4900
rect 13860 3900 13890 4900
rect 13956 3900 13986 4900
rect 14052 3900 14082 4900
rect 15568 3926 15598 5926
rect 15664 3926 15694 5926
<< ndiff >>
rect -1698 3195 -1636 3236
rect -1698 3161 -1686 3195
rect -1652 3161 -1636 3195
rect -1698 3127 -1636 3161
rect -1698 3093 -1686 3127
rect -1652 3093 -1636 3127
rect -1698 3059 -1636 3093
rect -1698 3025 -1686 3059
rect -1652 3025 -1636 3059
rect -1698 2991 -1636 3025
rect -1698 2957 -1686 2991
rect -1652 2957 -1636 2991
rect -1698 2923 -1636 2957
rect -1698 2889 -1686 2923
rect -1652 2889 -1636 2923
rect -1698 2855 -1636 2889
rect -1698 2821 -1686 2855
rect -1652 2821 -1636 2855
rect -1698 2787 -1636 2821
rect -1698 2753 -1686 2787
rect -1652 2753 -1636 2787
rect -1698 2719 -1636 2753
rect -1698 2685 -1686 2719
rect -1652 2685 -1636 2719
rect -1698 2651 -1636 2685
rect -1698 2617 -1686 2651
rect -1652 2617 -1636 2651
rect -1698 2583 -1636 2617
rect -1698 2549 -1686 2583
rect -1652 2549 -1636 2583
rect -1698 2515 -1636 2549
rect -1698 2481 -1686 2515
rect -1652 2481 -1636 2515
rect -1698 2447 -1636 2481
rect -1698 2413 -1686 2447
rect -1652 2413 -1636 2447
rect -1698 2379 -1636 2413
rect -1698 2345 -1686 2379
rect -1652 2345 -1636 2379
rect -1698 2311 -1636 2345
rect -1698 2277 -1686 2311
rect -1652 2277 -1636 2311
rect -1698 2236 -1636 2277
rect -1606 3195 -1540 3236
rect -1606 3161 -1590 3195
rect -1556 3161 -1540 3195
rect -1606 3127 -1540 3161
rect -1606 3093 -1590 3127
rect -1556 3093 -1540 3127
rect -1606 3059 -1540 3093
rect -1606 3025 -1590 3059
rect -1556 3025 -1540 3059
rect -1606 2991 -1540 3025
rect -1606 2957 -1590 2991
rect -1556 2957 -1540 2991
rect -1606 2923 -1540 2957
rect -1606 2889 -1590 2923
rect -1556 2889 -1540 2923
rect -1606 2855 -1540 2889
rect -1606 2821 -1590 2855
rect -1556 2821 -1540 2855
rect -1606 2787 -1540 2821
rect -1606 2753 -1590 2787
rect -1556 2753 -1540 2787
rect -1606 2719 -1540 2753
rect -1606 2685 -1590 2719
rect -1556 2685 -1540 2719
rect -1606 2651 -1540 2685
rect -1606 2617 -1590 2651
rect -1556 2617 -1540 2651
rect -1606 2583 -1540 2617
rect -1606 2549 -1590 2583
rect -1556 2549 -1540 2583
rect -1606 2515 -1540 2549
rect -1606 2481 -1590 2515
rect -1556 2481 -1540 2515
rect -1606 2447 -1540 2481
rect -1606 2413 -1590 2447
rect -1556 2413 -1540 2447
rect -1606 2379 -1540 2413
rect -1606 2345 -1590 2379
rect -1556 2345 -1540 2379
rect -1606 2311 -1540 2345
rect -1606 2277 -1590 2311
rect -1556 2277 -1540 2311
rect -1606 2236 -1540 2277
rect -1510 3195 -1444 3236
rect -1510 3161 -1494 3195
rect -1460 3161 -1444 3195
rect -1510 3127 -1444 3161
rect -1510 3093 -1494 3127
rect -1460 3093 -1444 3127
rect -1510 3059 -1444 3093
rect -1510 3025 -1494 3059
rect -1460 3025 -1444 3059
rect -1510 2991 -1444 3025
rect -1510 2957 -1494 2991
rect -1460 2957 -1444 2991
rect -1510 2923 -1444 2957
rect -1510 2889 -1494 2923
rect -1460 2889 -1444 2923
rect -1510 2855 -1444 2889
rect -1510 2821 -1494 2855
rect -1460 2821 -1444 2855
rect -1510 2787 -1444 2821
rect -1510 2753 -1494 2787
rect -1460 2753 -1444 2787
rect -1510 2719 -1444 2753
rect -1510 2685 -1494 2719
rect -1460 2685 -1444 2719
rect -1510 2651 -1444 2685
rect -1510 2617 -1494 2651
rect -1460 2617 -1444 2651
rect -1510 2583 -1444 2617
rect -1510 2549 -1494 2583
rect -1460 2549 -1444 2583
rect -1510 2515 -1444 2549
rect -1510 2481 -1494 2515
rect -1460 2481 -1444 2515
rect -1510 2447 -1444 2481
rect -1510 2413 -1494 2447
rect -1460 2413 -1444 2447
rect -1510 2379 -1444 2413
rect -1510 2345 -1494 2379
rect -1460 2345 -1444 2379
rect -1510 2311 -1444 2345
rect -1510 2277 -1494 2311
rect -1460 2277 -1444 2311
rect -1510 2236 -1444 2277
rect -1414 3195 -1348 3236
rect -1414 3161 -1398 3195
rect -1364 3161 -1348 3195
rect -1414 3127 -1348 3161
rect -1414 3093 -1398 3127
rect -1364 3093 -1348 3127
rect -1414 3059 -1348 3093
rect -1414 3025 -1398 3059
rect -1364 3025 -1348 3059
rect -1414 2991 -1348 3025
rect -1414 2957 -1398 2991
rect -1364 2957 -1348 2991
rect -1414 2923 -1348 2957
rect -1414 2889 -1398 2923
rect -1364 2889 -1348 2923
rect -1414 2855 -1348 2889
rect -1414 2821 -1398 2855
rect -1364 2821 -1348 2855
rect -1414 2787 -1348 2821
rect -1414 2753 -1398 2787
rect -1364 2753 -1348 2787
rect -1414 2719 -1348 2753
rect -1414 2685 -1398 2719
rect -1364 2685 -1348 2719
rect -1414 2651 -1348 2685
rect -1414 2617 -1398 2651
rect -1364 2617 -1348 2651
rect -1414 2583 -1348 2617
rect -1414 2549 -1398 2583
rect -1364 2549 -1348 2583
rect -1414 2515 -1348 2549
rect -1414 2481 -1398 2515
rect -1364 2481 -1348 2515
rect -1414 2447 -1348 2481
rect -1414 2413 -1398 2447
rect -1364 2413 -1348 2447
rect -1414 2379 -1348 2413
rect -1414 2345 -1398 2379
rect -1364 2345 -1348 2379
rect -1414 2311 -1348 2345
rect -1414 2277 -1398 2311
rect -1364 2277 -1348 2311
rect -1414 2236 -1348 2277
rect -1318 3195 -1252 3236
rect -1318 3161 -1302 3195
rect -1268 3161 -1252 3195
rect -1318 3127 -1252 3161
rect -1318 3093 -1302 3127
rect -1268 3093 -1252 3127
rect -1318 3059 -1252 3093
rect -1318 3025 -1302 3059
rect -1268 3025 -1252 3059
rect -1318 2991 -1252 3025
rect -1318 2957 -1302 2991
rect -1268 2957 -1252 2991
rect -1318 2923 -1252 2957
rect -1318 2889 -1302 2923
rect -1268 2889 -1252 2923
rect -1318 2855 -1252 2889
rect -1318 2821 -1302 2855
rect -1268 2821 -1252 2855
rect -1318 2787 -1252 2821
rect -1318 2753 -1302 2787
rect -1268 2753 -1252 2787
rect -1318 2719 -1252 2753
rect -1318 2685 -1302 2719
rect -1268 2685 -1252 2719
rect -1318 2651 -1252 2685
rect -1318 2617 -1302 2651
rect -1268 2617 -1252 2651
rect -1318 2583 -1252 2617
rect -1318 2549 -1302 2583
rect -1268 2549 -1252 2583
rect -1318 2515 -1252 2549
rect -1318 2481 -1302 2515
rect -1268 2481 -1252 2515
rect -1318 2447 -1252 2481
rect -1318 2413 -1302 2447
rect -1268 2413 -1252 2447
rect -1318 2379 -1252 2413
rect -1318 2345 -1302 2379
rect -1268 2345 -1252 2379
rect -1318 2311 -1252 2345
rect -1318 2277 -1302 2311
rect -1268 2277 -1252 2311
rect -1318 2236 -1252 2277
rect -1222 3195 -1156 3236
rect -1222 3161 -1206 3195
rect -1172 3161 -1156 3195
rect -1222 3127 -1156 3161
rect -1222 3093 -1206 3127
rect -1172 3093 -1156 3127
rect -1222 3059 -1156 3093
rect -1222 3025 -1206 3059
rect -1172 3025 -1156 3059
rect -1222 2991 -1156 3025
rect -1222 2957 -1206 2991
rect -1172 2957 -1156 2991
rect -1222 2923 -1156 2957
rect -1222 2889 -1206 2923
rect -1172 2889 -1156 2923
rect -1222 2855 -1156 2889
rect -1222 2821 -1206 2855
rect -1172 2821 -1156 2855
rect -1222 2787 -1156 2821
rect -1222 2753 -1206 2787
rect -1172 2753 -1156 2787
rect -1222 2719 -1156 2753
rect -1222 2685 -1206 2719
rect -1172 2685 -1156 2719
rect -1222 2651 -1156 2685
rect -1222 2617 -1206 2651
rect -1172 2617 -1156 2651
rect -1222 2583 -1156 2617
rect -1222 2549 -1206 2583
rect -1172 2549 -1156 2583
rect -1222 2515 -1156 2549
rect -1222 2481 -1206 2515
rect -1172 2481 -1156 2515
rect -1222 2447 -1156 2481
rect -1222 2413 -1206 2447
rect -1172 2413 -1156 2447
rect -1222 2379 -1156 2413
rect -1222 2345 -1206 2379
rect -1172 2345 -1156 2379
rect -1222 2311 -1156 2345
rect -1222 2277 -1206 2311
rect -1172 2277 -1156 2311
rect -1222 2236 -1156 2277
rect -1126 3195 -1060 3236
rect -1126 3161 -1110 3195
rect -1076 3161 -1060 3195
rect -1126 3127 -1060 3161
rect -1126 3093 -1110 3127
rect -1076 3093 -1060 3127
rect -1126 3059 -1060 3093
rect -1126 3025 -1110 3059
rect -1076 3025 -1060 3059
rect -1126 2991 -1060 3025
rect -1126 2957 -1110 2991
rect -1076 2957 -1060 2991
rect -1126 2923 -1060 2957
rect -1126 2889 -1110 2923
rect -1076 2889 -1060 2923
rect -1126 2855 -1060 2889
rect -1126 2821 -1110 2855
rect -1076 2821 -1060 2855
rect -1126 2787 -1060 2821
rect -1126 2753 -1110 2787
rect -1076 2753 -1060 2787
rect -1126 2719 -1060 2753
rect -1126 2685 -1110 2719
rect -1076 2685 -1060 2719
rect -1126 2651 -1060 2685
rect -1126 2617 -1110 2651
rect -1076 2617 -1060 2651
rect -1126 2583 -1060 2617
rect -1126 2549 -1110 2583
rect -1076 2549 -1060 2583
rect -1126 2515 -1060 2549
rect -1126 2481 -1110 2515
rect -1076 2481 -1060 2515
rect -1126 2447 -1060 2481
rect -1126 2413 -1110 2447
rect -1076 2413 -1060 2447
rect -1126 2379 -1060 2413
rect -1126 2345 -1110 2379
rect -1076 2345 -1060 2379
rect -1126 2311 -1060 2345
rect -1126 2277 -1110 2311
rect -1076 2277 -1060 2311
rect -1126 2236 -1060 2277
rect -1030 3195 -964 3236
rect -1030 3161 -1014 3195
rect -980 3161 -964 3195
rect -1030 3127 -964 3161
rect -1030 3093 -1014 3127
rect -980 3093 -964 3127
rect -1030 3059 -964 3093
rect -1030 3025 -1014 3059
rect -980 3025 -964 3059
rect -1030 2991 -964 3025
rect -1030 2957 -1014 2991
rect -980 2957 -964 2991
rect -1030 2923 -964 2957
rect -1030 2889 -1014 2923
rect -980 2889 -964 2923
rect -1030 2855 -964 2889
rect -1030 2821 -1014 2855
rect -980 2821 -964 2855
rect -1030 2787 -964 2821
rect -1030 2753 -1014 2787
rect -980 2753 -964 2787
rect -1030 2719 -964 2753
rect -1030 2685 -1014 2719
rect -980 2685 -964 2719
rect -1030 2651 -964 2685
rect -1030 2617 -1014 2651
rect -980 2617 -964 2651
rect -1030 2583 -964 2617
rect -1030 2549 -1014 2583
rect -980 2549 -964 2583
rect -1030 2515 -964 2549
rect -1030 2481 -1014 2515
rect -980 2481 -964 2515
rect -1030 2447 -964 2481
rect -1030 2413 -1014 2447
rect -980 2413 -964 2447
rect -1030 2379 -964 2413
rect -1030 2345 -1014 2379
rect -980 2345 -964 2379
rect -1030 2311 -964 2345
rect -1030 2277 -1014 2311
rect -980 2277 -964 2311
rect -1030 2236 -964 2277
rect -934 3195 -872 3236
rect -934 3161 -918 3195
rect -884 3161 -872 3195
rect -934 3127 -872 3161
rect -934 3093 -918 3127
rect -884 3093 -872 3127
rect -934 3059 -872 3093
rect -934 3025 -918 3059
rect -884 3025 -872 3059
rect -934 2991 -872 3025
rect -934 2957 -918 2991
rect -884 2957 -872 2991
rect -934 2923 -872 2957
rect -934 2889 -918 2923
rect -884 2889 -872 2923
rect -934 2855 -872 2889
rect -934 2821 -918 2855
rect -884 2821 -872 2855
rect -934 2787 -872 2821
rect -934 2753 -918 2787
rect -884 2753 -872 2787
rect -934 2719 -872 2753
rect -934 2685 -918 2719
rect -884 2685 -872 2719
rect -934 2651 -872 2685
rect -934 2617 -918 2651
rect -884 2617 -872 2651
rect -934 2583 -872 2617
rect -934 2549 -918 2583
rect -884 2549 -872 2583
rect -934 2515 -872 2549
rect -934 2481 -918 2515
rect -884 2481 -872 2515
rect -934 2447 -872 2481
rect -934 2413 -918 2447
rect -884 2413 -872 2447
rect -934 2379 -872 2413
rect -934 2345 -918 2379
rect -884 2345 -872 2379
rect -934 2311 -872 2345
rect -934 2277 -918 2311
rect -884 2277 -872 2311
rect -934 2236 -872 2277
rect 1470 2789 1532 2830
rect 1470 2755 1482 2789
rect 1516 2755 1532 2789
rect 1470 2721 1532 2755
rect 1470 2687 1482 2721
rect 1516 2687 1532 2721
rect 1470 2653 1532 2687
rect 1470 2619 1482 2653
rect 1516 2619 1532 2653
rect 1470 2585 1532 2619
rect 1470 2551 1482 2585
rect 1516 2551 1532 2585
rect 1470 2517 1532 2551
rect 1470 2483 1482 2517
rect 1516 2483 1532 2517
rect 1470 2449 1532 2483
rect 1470 2415 1482 2449
rect 1516 2415 1532 2449
rect 1470 2381 1532 2415
rect 1470 2347 1482 2381
rect 1516 2347 1532 2381
rect 1470 2313 1532 2347
rect 1470 2279 1482 2313
rect 1516 2279 1532 2313
rect 1470 2245 1532 2279
rect 1470 2211 1482 2245
rect 1516 2211 1532 2245
rect 1470 2177 1532 2211
rect 1470 2143 1482 2177
rect 1516 2143 1532 2177
rect 1470 2109 1532 2143
rect 1470 2075 1482 2109
rect 1516 2075 1532 2109
rect 1470 2041 1532 2075
rect 1470 2007 1482 2041
rect 1516 2007 1532 2041
rect 1470 1973 1532 2007
rect 1470 1939 1482 1973
rect 1516 1939 1532 1973
rect 1470 1905 1532 1939
rect 1470 1871 1482 1905
rect 1516 1871 1532 1905
rect 1470 1830 1532 1871
rect 1562 2789 1628 2830
rect 1562 2755 1578 2789
rect 1612 2755 1628 2789
rect 1562 2721 1628 2755
rect 1562 2687 1578 2721
rect 1612 2687 1628 2721
rect 1562 2653 1628 2687
rect 1562 2619 1578 2653
rect 1612 2619 1628 2653
rect 1562 2585 1628 2619
rect 1562 2551 1578 2585
rect 1612 2551 1628 2585
rect 1562 2517 1628 2551
rect 1562 2483 1578 2517
rect 1612 2483 1628 2517
rect 1562 2449 1628 2483
rect 1562 2415 1578 2449
rect 1612 2415 1628 2449
rect 1562 2381 1628 2415
rect 1562 2347 1578 2381
rect 1612 2347 1628 2381
rect 1562 2313 1628 2347
rect 1562 2279 1578 2313
rect 1612 2279 1628 2313
rect 1562 2245 1628 2279
rect 1562 2211 1578 2245
rect 1612 2211 1628 2245
rect 1562 2177 1628 2211
rect 1562 2143 1578 2177
rect 1612 2143 1628 2177
rect 1562 2109 1628 2143
rect 1562 2075 1578 2109
rect 1612 2075 1628 2109
rect 1562 2041 1628 2075
rect 1562 2007 1578 2041
rect 1612 2007 1628 2041
rect 1562 1973 1628 2007
rect 1562 1939 1578 1973
rect 1612 1939 1628 1973
rect 1562 1905 1628 1939
rect 1562 1871 1578 1905
rect 1612 1871 1628 1905
rect 1562 1830 1628 1871
rect 1658 2789 1724 2830
rect 1658 2755 1674 2789
rect 1708 2755 1724 2789
rect 1658 2721 1724 2755
rect 1658 2687 1674 2721
rect 1708 2687 1724 2721
rect 1658 2653 1724 2687
rect 1658 2619 1674 2653
rect 1708 2619 1724 2653
rect 1658 2585 1724 2619
rect 1658 2551 1674 2585
rect 1708 2551 1724 2585
rect 1658 2517 1724 2551
rect 1658 2483 1674 2517
rect 1708 2483 1724 2517
rect 1658 2449 1724 2483
rect 1658 2415 1674 2449
rect 1708 2415 1724 2449
rect 1658 2381 1724 2415
rect 1658 2347 1674 2381
rect 1708 2347 1724 2381
rect 1658 2313 1724 2347
rect 1658 2279 1674 2313
rect 1708 2279 1724 2313
rect 1658 2245 1724 2279
rect 1658 2211 1674 2245
rect 1708 2211 1724 2245
rect 1658 2177 1724 2211
rect 1658 2143 1674 2177
rect 1708 2143 1724 2177
rect 1658 2109 1724 2143
rect 1658 2075 1674 2109
rect 1708 2075 1724 2109
rect 1658 2041 1724 2075
rect 1658 2007 1674 2041
rect 1708 2007 1724 2041
rect 1658 1973 1724 2007
rect 1658 1939 1674 1973
rect 1708 1939 1724 1973
rect 1658 1905 1724 1939
rect 1658 1871 1674 1905
rect 1708 1871 1724 1905
rect 1658 1830 1724 1871
rect 1754 2789 1820 2830
rect 1754 2755 1770 2789
rect 1804 2755 1820 2789
rect 1754 2721 1820 2755
rect 1754 2687 1770 2721
rect 1804 2687 1820 2721
rect 1754 2653 1820 2687
rect 1754 2619 1770 2653
rect 1804 2619 1820 2653
rect 1754 2585 1820 2619
rect 1754 2551 1770 2585
rect 1804 2551 1820 2585
rect 1754 2517 1820 2551
rect 1754 2483 1770 2517
rect 1804 2483 1820 2517
rect 1754 2449 1820 2483
rect 1754 2415 1770 2449
rect 1804 2415 1820 2449
rect 1754 2381 1820 2415
rect 1754 2347 1770 2381
rect 1804 2347 1820 2381
rect 1754 2313 1820 2347
rect 1754 2279 1770 2313
rect 1804 2279 1820 2313
rect 1754 2245 1820 2279
rect 1754 2211 1770 2245
rect 1804 2211 1820 2245
rect 1754 2177 1820 2211
rect 1754 2143 1770 2177
rect 1804 2143 1820 2177
rect 1754 2109 1820 2143
rect 1754 2075 1770 2109
rect 1804 2075 1820 2109
rect 1754 2041 1820 2075
rect 1754 2007 1770 2041
rect 1804 2007 1820 2041
rect 1754 1973 1820 2007
rect 1754 1939 1770 1973
rect 1804 1939 1820 1973
rect 1754 1905 1820 1939
rect 1754 1871 1770 1905
rect 1804 1871 1820 1905
rect 1754 1830 1820 1871
rect 1850 2789 1912 2830
rect 1850 2755 1866 2789
rect 1900 2755 1912 2789
rect 1850 2721 1912 2755
rect 1850 2687 1866 2721
rect 1900 2687 1912 2721
rect 1850 2653 1912 2687
rect 1850 2619 1866 2653
rect 1900 2619 1912 2653
rect 1850 2585 1912 2619
rect 1850 2551 1866 2585
rect 1900 2551 1912 2585
rect 1850 2517 1912 2551
rect 1850 2483 1866 2517
rect 1900 2483 1912 2517
rect 1850 2449 1912 2483
rect 1850 2415 1866 2449
rect 1900 2415 1912 2449
rect 4426 2773 4488 2814
rect 4426 2739 4438 2773
rect 4472 2739 4488 2773
rect 4426 2705 4488 2739
rect 4426 2671 4438 2705
rect 4472 2671 4488 2705
rect 4426 2637 4488 2671
rect 4426 2603 4438 2637
rect 4472 2603 4488 2637
rect 4426 2569 4488 2603
rect 4426 2535 4438 2569
rect 4472 2535 4488 2569
rect 4426 2501 4488 2535
rect 4426 2467 4438 2501
rect 4472 2467 4488 2501
rect 1850 2381 1912 2415
rect 1850 2347 1866 2381
rect 1900 2347 1912 2381
rect 1850 2313 1912 2347
rect 1850 2279 1866 2313
rect 1900 2279 1912 2313
rect 1850 2245 1912 2279
rect 4426 2433 4488 2467
rect 4426 2399 4438 2433
rect 4472 2399 4488 2433
rect 4426 2365 4488 2399
rect 4426 2331 4438 2365
rect 4472 2331 4488 2365
rect 4426 2297 4488 2331
rect 1850 2211 1866 2245
rect 1900 2211 1912 2245
rect 1850 2177 1912 2211
rect 1850 2143 1866 2177
rect 1900 2143 1912 2177
rect 1850 2109 1912 2143
rect 1850 2075 1866 2109
rect 1900 2075 1912 2109
rect 2488 2261 2546 2276
rect 2488 2227 2500 2261
rect 2534 2227 2546 2261
rect 2488 2193 2546 2227
rect 2488 2159 2500 2193
rect 2534 2159 2546 2193
rect 2488 2125 2546 2159
rect 2488 2091 2500 2125
rect 2534 2091 2546 2125
rect 2488 2076 2546 2091
rect 2646 2261 2704 2276
rect 2646 2227 2658 2261
rect 2692 2227 2704 2261
rect 2646 2193 2704 2227
rect 2646 2159 2658 2193
rect 2692 2159 2704 2193
rect 2646 2125 2704 2159
rect 2646 2091 2658 2125
rect 2692 2091 2704 2125
rect 2646 2076 2704 2091
rect 4426 2263 4438 2297
rect 4472 2263 4488 2297
rect 4426 2229 4488 2263
rect 4426 2195 4438 2229
rect 4472 2195 4488 2229
rect 4426 2161 4488 2195
rect 4426 2127 4438 2161
rect 4472 2127 4488 2161
rect 4426 2093 4488 2127
rect 1850 2041 1912 2075
rect 4426 2059 4438 2093
rect 4472 2059 4488 2093
rect 1850 2007 1866 2041
rect 1900 2007 1912 2041
rect 1850 1973 1912 2007
rect 1850 1939 1866 1973
rect 1900 1939 1912 1973
rect 1850 1905 1912 1939
rect 1850 1871 1866 1905
rect 1900 1871 1912 1905
rect 1850 1830 1912 1871
rect 4426 2025 4488 2059
rect 4426 1991 4438 2025
rect 4472 1991 4488 2025
rect 4426 1957 4488 1991
rect 4426 1923 4438 1957
rect 4472 1923 4488 1957
rect 4426 1889 4488 1923
rect 4426 1855 4438 1889
rect 4472 1855 4488 1889
rect 4426 1814 4488 1855
rect 4518 2773 4584 2814
rect 4518 2739 4534 2773
rect 4568 2739 4584 2773
rect 4518 2705 4584 2739
rect 4518 2671 4534 2705
rect 4568 2671 4584 2705
rect 4518 2637 4584 2671
rect 4518 2603 4534 2637
rect 4568 2603 4584 2637
rect 4518 2569 4584 2603
rect 4518 2535 4534 2569
rect 4568 2535 4584 2569
rect 4518 2501 4584 2535
rect 4518 2467 4534 2501
rect 4568 2467 4584 2501
rect 4518 2433 4584 2467
rect 4518 2399 4534 2433
rect 4568 2399 4584 2433
rect 4518 2365 4584 2399
rect 4518 2331 4534 2365
rect 4568 2331 4584 2365
rect 4518 2297 4584 2331
rect 4518 2263 4534 2297
rect 4568 2263 4584 2297
rect 4518 2229 4584 2263
rect 4518 2195 4534 2229
rect 4568 2195 4584 2229
rect 4518 2161 4584 2195
rect 4518 2127 4534 2161
rect 4568 2127 4584 2161
rect 4518 2093 4584 2127
rect 4518 2059 4534 2093
rect 4568 2059 4584 2093
rect 4518 2025 4584 2059
rect 4518 1991 4534 2025
rect 4568 1991 4584 2025
rect 4518 1957 4584 1991
rect 4518 1923 4534 1957
rect 4568 1923 4584 1957
rect 4518 1889 4584 1923
rect 4518 1855 4534 1889
rect 4568 1855 4584 1889
rect 4518 1814 4584 1855
rect 4614 2773 4680 2814
rect 4614 2739 4630 2773
rect 4664 2739 4680 2773
rect 4614 2705 4680 2739
rect 4614 2671 4630 2705
rect 4664 2671 4680 2705
rect 4614 2637 4680 2671
rect 4614 2603 4630 2637
rect 4664 2603 4680 2637
rect 4614 2569 4680 2603
rect 4614 2535 4630 2569
rect 4664 2535 4680 2569
rect 4614 2501 4680 2535
rect 4614 2467 4630 2501
rect 4664 2467 4680 2501
rect 4614 2433 4680 2467
rect 4614 2399 4630 2433
rect 4664 2399 4680 2433
rect 4614 2365 4680 2399
rect 4614 2331 4630 2365
rect 4664 2331 4680 2365
rect 4614 2297 4680 2331
rect 4614 2263 4630 2297
rect 4664 2263 4680 2297
rect 4614 2229 4680 2263
rect 4614 2195 4630 2229
rect 4664 2195 4680 2229
rect 4614 2161 4680 2195
rect 4614 2127 4630 2161
rect 4664 2127 4680 2161
rect 4614 2093 4680 2127
rect 4614 2059 4630 2093
rect 4664 2059 4680 2093
rect 4614 2025 4680 2059
rect 4614 1991 4630 2025
rect 4664 1991 4680 2025
rect 4614 1957 4680 1991
rect 4614 1923 4630 1957
rect 4664 1923 4680 1957
rect 4614 1889 4680 1923
rect 4614 1855 4630 1889
rect 4664 1855 4680 1889
rect 4614 1814 4680 1855
rect 4710 2773 4776 2814
rect 4710 2739 4726 2773
rect 4760 2739 4776 2773
rect 4710 2705 4776 2739
rect 4710 2671 4726 2705
rect 4760 2671 4776 2705
rect 4710 2637 4776 2671
rect 4710 2603 4726 2637
rect 4760 2603 4776 2637
rect 4710 2569 4776 2603
rect 4710 2535 4726 2569
rect 4760 2535 4776 2569
rect 4710 2501 4776 2535
rect 4710 2467 4726 2501
rect 4760 2467 4776 2501
rect 4710 2433 4776 2467
rect 4710 2399 4726 2433
rect 4760 2399 4776 2433
rect 4710 2365 4776 2399
rect 4710 2331 4726 2365
rect 4760 2331 4776 2365
rect 4710 2297 4776 2331
rect 4710 2263 4726 2297
rect 4760 2263 4776 2297
rect 4710 2229 4776 2263
rect 4710 2195 4726 2229
rect 4760 2195 4776 2229
rect 4710 2161 4776 2195
rect 4710 2127 4726 2161
rect 4760 2127 4776 2161
rect 4710 2093 4776 2127
rect 4710 2059 4726 2093
rect 4760 2059 4776 2093
rect 4710 2025 4776 2059
rect 4710 1991 4726 2025
rect 4760 1991 4776 2025
rect 4710 1957 4776 1991
rect 4710 1923 4726 1957
rect 4760 1923 4776 1957
rect 4710 1889 4776 1923
rect 4710 1855 4726 1889
rect 4760 1855 4776 1889
rect 4710 1814 4776 1855
rect 4806 2773 4868 2814
rect 4806 2739 4822 2773
rect 4856 2739 4868 2773
rect 4806 2705 4868 2739
rect 4806 2671 4822 2705
rect 4856 2671 4868 2705
rect 4806 2637 4868 2671
rect 4806 2603 4822 2637
rect 4856 2603 4868 2637
rect 4806 2569 4868 2603
rect 4806 2535 4822 2569
rect 4856 2535 4868 2569
rect 4806 2501 4868 2535
rect 4806 2467 4822 2501
rect 4856 2467 4868 2501
rect 4806 2433 4868 2467
rect 7456 2773 7518 2814
rect 7456 2739 7468 2773
rect 7502 2739 7518 2773
rect 7456 2705 7518 2739
rect 7456 2671 7468 2705
rect 7502 2671 7518 2705
rect 7456 2637 7518 2671
rect 7456 2603 7468 2637
rect 7502 2603 7518 2637
rect 7456 2569 7518 2603
rect 7456 2535 7468 2569
rect 7502 2535 7518 2569
rect 7456 2501 7518 2535
rect 7456 2467 7468 2501
rect 7502 2467 7518 2501
rect 4806 2399 4822 2433
rect 4856 2399 4868 2433
rect 4806 2365 4868 2399
rect 4806 2331 4822 2365
rect 4856 2331 4868 2365
rect 4806 2297 4868 2331
rect 4806 2263 4822 2297
rect 4856 2263 4868 2297
rect 7456 2433 7518 2467
rect 7456 2399 7468 2433
rect 7502 2399 7518 2433
rect 7456 2365 7518 2399
rect 7456 2331 7468 2365
rect 7502 2331 7518 2365
rect 7456 2297 7518 2331
rect 4806 2229 4868 2263
rect 4806 2195 4822 2229
rect 4856 2195 4868 2229
rect 4806 2161 4868 2195
rect 4806 2127 4822 2161
rect 4856 2127 4868 2161
rect 4806 2093 4868 2127
rect 4806 2059 4822 2093
rect 4856 2059 4868 2093
rect 5488 2261 5546 2276
rect 5488 2227 5500 2261
rect 5534 2227 5546 2261
rect 5488 2193 5546 2227
rect 5488 2159 5500 2193
rect 5534 2159 5546 2193
rect 5488 2125 5546 2159
rect 5488 2091 5500 2125
rect 5534 2091 5546 2125
rect 5488 2076 5546 2091
rect 5646 2261 5704 2276
rect 5646 2227 5658 2261
rect 5692 2227 5704 2261
rect 5646 2193 5704 2227
rect 5646 2159 5658 2193
rect 5692 2159 5704 2193
rect 5646 2125 5704 2159
rect 5646 2091 5658 2125
rect 5692 2091 5704 2125
rect 5646 2076 5704 2091
rect 7456 2263 7468 2297
rect 7502 2263 7518 2297
rect 7456 2229 7518 2263
rect 7456 2195 7468 2229
rect 7502 2195 7518 2229
rect 7456 2161 7518 2195
rect 7456 2127 7468 2161
rect 7502 2127 7518 2161
rect 7456 2093 7518 2127
rect 4806 2025 4868 2059
rect 7456 2059 7468 2093
rect 7502 2059 7518 2093
rect 4806 1991 4822 2025
rect 4856 1991 4868 2025
rect 4806 1957 4868 1991
rect 4806 1923 4822 1957
rect 4856 1923 4868 1957
rect 4806 1889 4868 1923
rect 4806 1855 4822 1889
rect 4856 1855 4868 1889
rect 4806 1814 4868 1855
rect 7456 2025 7518 2059
rect 7456 1991 7468 2025
rect 7502 1991 7518 2025
rect 7456 1957 7518 1991
rect 7456 1923 7468 1957
rect 7502 1923 7518 1957
rect 7456 1889 7518 1923
rect 7456 1855 7468 1889
rect 7502 1855 7518 1889
rect 7456 1814 7518 1855
rect 7548 2773 7614 2814
rect 7548 2739 7564 2773
rect 7598 2739 7614 2773
rect 7548 2705 7614 2739
rect 7548 2671 7564 2705
rect 7598 2671 7614 2705
rect 7548 2637 7614 2671
rect 7548 2603 7564 2637
rect 7598 2603 7614 2637
rect 7548 2569 7614 2603
rect 7548 2535 7564 2569
rect 7598 2535 7614 2569
rect 7548 2501 7614 2535
rect 7548 2467 7564 2501
rect 7598 2467 7614 2501
rect 7548 2433 7614 2467
rect 7548 2399 7564 2433
rect 7598 2399 7614 2433
rect 7548 2365 7614 2399
rect 7548 2331 7564 2365
rect 7598 2331 7614 2365
rect 7548 2297 7614 2331
rect 7548 2263 7564 2297
rect 7598 2263 7614 2297
rect 7548 2229 7614 2263
rect 7548 2195 7564 2229
rect 7598 2195 7614 2229
rect 7548 2161 7614 2195
rect 7548 2127 7564 2161
rect 7598 2127 7614 2161
rect 7548 2093 7614 2127
rect 7548 2059 7564 2093
rect 7598 2059 7614 2093
rect 7548 2025 7614 2059
rect 7548 1991 7564 2025
rect 7598 1991 7614 2025
rect 7548 1957 7614 1991
rect 7548 1923 7564 1957
rect 7598 1923 7614 1957
rect 7548 1889 7614 1923
rect 7548 1855 7564 1889
rect 7598 1855 7614 1889
rect 7548 1814 7614 1855
rect 7644 2773 7710 2814
rect 7644 2739 7660 2773
rect 7694 2739 7710 2773
rect 7644 2705 7710 2739
rect 7644 2671 7660 2705
rect 7694 2671 7710 2705
rect 7644 2637 7710 2671
rect 7644 2603 7660 2637
rect 7694 2603 7710 2637
rect 7644 2569 7710 2603
rect 7644 2535 7660 2569
rect 7694 2535 7710 2569
rect 7644 2501 7710 2535
rect 7644 2467 7660 2501
rect 7694 2467 7710 2501
rect 7644 2433 7710 2467
rect 7644 2399 7660 2433
rect 7694 2399 7710 2433
rect 7644 2365 7710 2399
rect 7644 2331 7660 2365
rect 7694 2331 7710 2365
rect 7644 2297 7710 2331
rect 7644 2263 7660 2297
rect 7694 2263 7710 2297
rect 7644 2229 7710 2263
rect 7644 2195 7660 2229
rect 7694 2195 7710 2229
rect 7644 2161 7710 2195
rect 7644 2127 7660 2161
rect 7694 2127 7710 2161
rect 7644 2093 7710 2127
rect 7644 2059 7660 2093
rect 7694 2059 7710 2093
rect 7644 2025 7710 2059
rect 7644 1991 7660 2025
rect 7694 1991 7710 2025
rect 7644 1957 7710 1991
rect 7644 1923 7660 1957
rect 7694 1923 7710 1957
rect 7644 1889 7710 1923
rect 7644 1855 7660 1889
rect 7694 1855 7710 1889
rect 7644 1814 7710 1855
rect 7740 2773 7806 2814
rect 7740 2739 7756 2773
rect 7790 2739 7806 2773
rect 7740 2705 7806 2739
rect 7740 2671 7756 2705
rect 7790 2671 7806 2705
rect 7740 2637 7806 2671
rect 7740 2603 7756 2637
rect 7790 2603 7806 2637
rect 7740 2569 7806 2603
rect 7740 2535 7756 2569
rect 7790 2535 7806 2569
rect 7740 2501 7806 2535
rect 7740 2467 7756 2501
rect 7790 2467 7806 2501
rect 7740 2433 7806 2467
rect 7740 2399 7756 2433
rect 7790 2399 7806 2433
rect 7740 2365 7806 2399
rect 7740 2331 7756 2365
rect 7790 2331 7806 2365
rect 7740 2297 7806 2331
rect 7740 2263 7756 2297
rect 7790 2263 7806 2297
rect 7740 2229 7806 2263
rect 7740 2195 7756 2229
rect 7790 2195 7806 2229
rect 7740 2161 7806 2195
rect 7740 2127 7756 2161
rect 7790 2127 7806 2161
rect 7740 2093 7806 2127
rect 7740 2059 7756 2093
rect 7790 2059 7806 2093
rect 7740 2025 7806 2059
rect 7740 1991 7756 2025
rect 7790 1991 7806 2025
rect 7740 1957 7806 1991
rect 7740 1923 7756 1957
rect 7790 1923 7806 1957
rect 7740 1889 7806 1923
rect 7740 1855 7756 1889
rect 7790 1855 7806 1889
rect 7740 1814 7806 1855
rect 7836 2773 7898 2814
rect 7836 2739 7852 2773
rect 7886 2739 7898 2773
rect 7836 2705 7898 2739
rect 7836 2671 7852 2705
rect 7886 2671 7898 2705
rect 7836 2637 7898 2671
rect 7836 2603 7852 2637
rect 7886 2603 7898 2637
rect 7836 2569 7898 2603
rect 7836 2535 7852 2569
rect 7886 2535 7898 2569
rect 7836 2501 7898 2535
rect 7836 2467 7852 2501
rect 7886 2467 7898 2501
rect 7836 2433 7898 2467
rect 10544 2771 10606 2812
rect 10544 2737 10556 2771
rect 10590 2737 10606 2771
rect 10544 2703 10606 2737
rect 10544 2669 10556 2703
rect 10590 2669 10606 2703
rect 10544 2635 10606 2669
rect 10544 2601 10556 2635
rect 10590 2601 10606 2635
rect 10544 2567 10606 2601
rect 10544 2533 10556 2567
rect 10590 2533 10606 2567
rect 10544 2499 10606 2533
rect 10544 2465 10556 2499
rect 10590 2465 10606 2499
rect 7836 2399 7852 2433
rect 7886 2399 7898 2433
rect 7836 2365 7898 2399
rect 7836 2331 7852 2365
rect 7886 2331 7898 2365
rect 7836 2297 7898 2331
rect 7836 2263 7852 2297
rect 7886 2263 7898 2297
rect 10544 2431 10606 2465
rect 10544 2397 10556 2431
rect 10590 2397 10606 2431
rect 10544 2363 10606 2397
rect 10544 2329 10556 2363
rect 10590 2329 10606 2363
rect 10544 2295 10606 2329
rect 7836 2229 7898 2263
rect 7836 2195 7852 2229
rect 7886 2195 7898 2229
rect 7836 2161 7898 2195
rect 7836 2127 7852 2161
rect 7886 2127 7898 2161
rect 7836 2093 7898 2127
rect 7836 2059 7852 2093
rect 7886 2059 7898 2093
rect 8488 2261 8546 2276
rect 8488 2227 8500 2261
rect 8534 2227 8546 2261
rect 8488 2193 8546 2227
rect 8488 2159 8500 2193
rect 8534 2159 8546 2193
rect 8488 2125 8546 2159
rect 8488 2091 8500 2125
rect 8534 2091 8546 2125
rect 8488 2076 8546 2091
rect 8646 2261 8704 2276
rect 8646 2227 8658 2261
rect 8692 2227 8704 2261
rect 8646 2193 8704 2227
rect 8646 2159 8658 2193
rect 8692 2159 8704 2193
rect 8646 2125 8704 2159
rect 8646 2091 8658 2125
rect 8692 2091 8704 2125
rect 8646 2076 8704 2091
rect 10544 2261 10556 2295
rect 10590 2261 10606 2295
rect 10544 2227 10606 2261
rect 10544 2193 10556 2227
rect 10590 2193 10606 2227
rect 10544 2159 10606 2193
rect 10544 2125 10556 2159
rect 10590 2125 10606 2159
rect 10544 2091 10606 2125
rect 7836 2025 7898 2059
rect 10544 2057 10556 2091
rect 10590 2057 10606 2091
rect 7836 1991 7852 2025
rect 7886 1991 7898 2025
rect 7836 1957 7898 1991
rect 7836 1923 7852 1957
rect 7886 1923 7898 1957
rect 7836 1889 7898 1923
rect 7836 1855 7852 1889
rect 7886 1855 7898 1889
rect 7836 1814 7898 1855
rect 10544 2023 10606 2057
rect 10544 1989 10556 2023
rect 10590 1989 10606 2023
rect 10544 1955 10606 1989
rect 10544 1921 10556 1955
rect 10590 1921 10606 1955
rect 10544 1887 10606 1921
rect 10544 1853 10556 1887
rect 10590 1853 10606 1887
rect 10544 1812 10606 1853
rect 10636 2771 10702 2812
rect 10636 2737 10652 2771
rect 10686 2737 10702 2771
rect 10636 2703 10702 2737
rect 10636 2669 10652 2703
rect 10686 2669 10702 2703
rect 10636 2635 10702 2669
rect 10636 2601 10652 2635
rect 10686 2601 10702 2635
rect 10636 2567 10702 2601
rect 10636 2533 10652 2567
rect 10686 2533 10702 2567
rect 10636 2499 10702 2533
rect 10636 2465 10652 2499
rect 10686 2465 10702 2499
rect 10636 2431 10702 2465
rect 10636 2397 10652 2431
rect 10686 2397 10702 2431
rect 10636 2363 10702 2397
rect 10636 2329 10652 2363
rect 10686 2329 10702 2363
rect 10636 2295 10702 2329
rect 10636 2261 10652 2295
rect 10686 2261 10702 2295
rect 10636 2227 10702 2261
rect 10636 2193 10652 2227
rect 10686 2193 10702 2227
rect 10636 2159 10702 2193
rect 10636 2125 10652 2159
rect 10686 2125 10702 2159
rect 10636 2091 10702 2125
rect 10636 2057 10652 2091
rect 10686 2057 10702 2091
rect 10636 2023 10702 2057
rect 10636 1989 10652 2023
rect 10686 1989 10702 2023
rect 10636 1955 10702 1989
rect 10636 1921 10652 1955
rect 10686 1921 10702 1955
rect 10636 1887 10702 1921
rect 10636 1853 10652 1887
rect 10686 1853 10702 1887
rect 10636 1812 10702 1853
rect 10732 2771 10798 2812
rect 10732 2737 10748 2771
rect 10782 2737 10798 2771
rect 10732 2703 10798 2737
rect 10732 2669 10748 2703
rect 10782 2669 10798 2703
rect 10732 2635 10798 2669
rect 10732 2601 10748 2635
rect 10782 2601 10798 2635
rect 10732 2567 10798 2601
rect 10732 2533 10748 2567
rect 10782 2533 10798 2567
rect 10732 2499 10798 2533
rect 10732 2465 10748 2499
rect 10782 2465 10798 2499
rect 10732 2431 10798 2465
rect 10732 2397 10748 2431
rect 10782 2397 10798 2431
rect 10732 2363 10798 2397
rect 10732 2329 10748 2363
rect 10782 2329 10798 2363
rect 10732 2295 10798 2329
rect 10732 2261 10748 2295
rect 10782 2261 10798 2295
rect 10732 2227 10798 2261
rect 10732 2193 10748 2227
rect 10782 2193 10798 2227
rect 10732 2159 10798 2193
rect 10732 2125 10748 2159
rect 10782 2125 10798 2159
rect 10732 2091 10798 2125
rect 10732 2057 10748 2091
rect 10782 2057 10798 2091
rect 10732 2023 10798 2057
rect 10732 1989 10748 2023
rect 10782 1989 10798 2023
rect 10732 1955 10798 1989
rect 10732 1921 10748 1955
rect 10782 1921 10798 1955
rect 10732 1887 10798 1921
rect 10732 1853 10748 1887
rect 10782 1853 10798 1887
rect 10732 1812 10798 1853
rect 10828 2771 10894 2812
rect 10828 2737 10844 2771
rect 10878 2737 10894 2771
rect 10828 2703 10894 2737
rect 10828 2669 10844 2703
rect 10878 2669 10894 2703
rect 10828 2635 10894 2669
rect 10828 2601 10844 2635
rect 10878 2601 10894 2635
rect 10828 2567 10894 2601
rect 10828 2533 10844 2567
rect 10878 2533 10894 2567
rect 10828 2499 10894 2533
rect 10828 2465 10844 2499
rect 10878 2465 10894 2499
rect 10828 2431 10894 2465
rect 10828 2397 10844 2431
rect 10878 2397 10894 2431
rect 10828 2363 10894 2397
rect 10828 2329 10844 2363
rect 10878 2329 10894 2363
rect 10828 2295 10894 2329
rect 10828 2261 10844 2295
rect 10878 2261 10894 2295
rect 10828 2227 10894 2261
rect 10828 2193 10844 2227
rect 10878 2193 10894 2227
rect 10828 2159 10894 2193
rect 10828 2125 10844 2159
rect 10878 2125 10894 2159
rect 10828 2091 10894 2125
rect 10828 2057 10844 2091
rect 10878 2057 10894 2091
rect 10828 2023 10894 2057
rect 10828 1989 10844 2023
rect 10878 1989 10894 2023
rect 10828 1955 10894 1989
rect 10828 1921 10844 1955
rect 10878 1921 10894 1955
rect 10828 1887 10894 1921
rect 10828 1853 10844 1887
rect 10878 1853 10894 1887
rect 10828 1812 10894 1853
rect 10924 2771 10986 2812
rect 10924 2737 10940 2771
rect 10974 2737 10986 2771
rect 10924 2703 10986 2737
rect 10924 2669 10940 2703
rect 10974 2669 10986 2703
rect 10924 2635 10986 2669
rect 10924 2601 10940 2635
rect 10974 2601 10986 2635
rect 10924 2567 10986 2601
rect 10924 2533 10940 2567
rect 10974 2533 10986 2567
rect 10924 2499 10986 2533
rect 10924 2465 10940 2499
rect 10974 2465 10986 2499
rect 10924 2431 10986 2465
rect 13700 2745 13762 2786
rect 13700 2711 13712 2745
rect 13746 2711 13762 2745
rect 13700 2677 13762 2711
rect 13700 2643 13712 2677
rect 13746 2643 13762 2677
rect 13700 2609 13762 2643
rect 13700 2575 13712 2609
rect 13746 2575 13762 2609
rect 13700 2541 13762 2575
rect 13700 2507 13712 2541
rect 13746 2507 13762 2541
rect 13700 2473 13762 2507
rect 10924 2397 10940 2431
rect 10974 2397 10986 2431
rect 10924 2363 10986 2397
rect 10924 2329 10940 2363
rect 10974 2329 10986 2363
rect 10924 2295 10986 2329
rect 10924 2261 10940 2295
rect 10974 2261 10986 2295
rect 13700 2439 13712 2473
rect 13746 2439 13762 2473
rect 13700 2405 13762 2439
rect 13700 2371 13712 2405
rect 13746 2371 13762 2405
rect 13700 2337 13762 2371
rect 13700 2303 13712 2337
rect 13746 2303 13762 2337
rect 10924 2227 10986 2261
rect 10924 2193 10940 2227
rect 10974 2193 10986 2227
rect 10924 2159 10986 2193
rect 10924 2125 10940 2159
rect 10974 2125 10986 2159
rect 10924 2091 10986 2125
rect 10924 2057 10940 2091
rect 10974 2057 10986 2091
rect 11488 2261 11546 2276
rect 11488 2227 11500 2261
rect 11534 2227 11546 2261
rect 11488 2193 11546 2227
rect 11488 2159 11500 2193
rect 11534 2159 11546 2193
rect 11488 2125 11546 2159
rect 11488 2091 11500 2125
rect 11534 2091 11546 2125
rect 11488 2076 11546 2091
rect 11646 2261 11704 2276
rect 11646 2227 11658 2261
rect 11692 2227 11704 2261
rect 11646 2193 11704 2227
rect 11646 2159 11658 2193
rect 11692 2159 11704 2193
rect 11646 2125 11704 2159
rect 11646 2091 11658 2125
rect 11692 2091 11704 2125
rect 11646 2076 11704 2091
rect 13700 2269 13762 2303
rect 13700 2235 13712 2269
rect 13746 2235 13762 2269
rect 13700 2201 13762 2235
rect 13700 2167 13712 2201
rect 13746 2167 13762 2201
rect 13700 2133 13762 2167
rect 13700 2099 13712 2133
rect 13746 2099 13762 2133
rect 10924 2023 10986 2057
rect 13700 2065 13762 2099
rect 10924 1989 10940 2023
rect 10974 1989 10986 2023
rect 10924 1955 10986 1989
rect 10924 1921 10940 1955
rect 10974 1921 10986 1955
rect 10924 1887 10986 1921
rect 10924 1853 10940 1887
rect 10974 1853 10986 1887
rect 10924 1812 10986 1853
rect 13700 2031 13712 2065
rect 13746 2031 13762 2065
rect 13700 1997 13762 2031
rect 13700 1963 13712 1997
rect 13746 1963 13762 1997
rect 13700 1929 13762 1963
rect 13700 1895 13712 1929
rect 13746 1895 13762 1929
rect 13700 1861 13762 1895
rect 13700 1827 13712 1861
rect 13746 1827 13762 1861
rect 13700 1786 13762 1827
rect 13792 2745 13858 2786
rect 13792 2711 13808 2745
rect 13842 2711 13858 2745
rect 13792 2677 13858 2711
rect 13792 2643 13808 2677
rect 13842 2643 13858 2677
rect 13792 2609 13858 2643
rect 13792 2575 13808 2609
rect 13842 2575 13858 2609
rect 13792 2541 13858 2575
rect 13792 2507 13808 2541
rect 13842 2507 13858 2541
rect 13792 2473 13858 2507
rect 13792 2439 13808 2473
rect 13842 2439 13858 2473
rect 13792 2405 13858 2439
rect 13792 2371 13808 2405
rect 13842 2371 13858 2405
rect 13792 2337 13858 2371
rect 13792 2303 13808 2337
rect 13842 2303 13858 2337
rect 13792 2269 13858 2303
rect 13792 2235 13808 2269
rect 13842 2235 13858 2269
rect 13792 2201 13858 2235
rect 13792 2167 13808 2201
rect 13842 2167 13858 2201
rect 13792 2133 13858 2167
rect 13792 2099 13808 2133
rect 13842 2099 13858 2133
rect 13792 2065 13858 2099
rect 13792 2031 13808 2065
rect 13842 2031 13858 2065
rect 13792 1997 13858 2031
rect 13792 1963 13808 1997
rect 13842 1963 13858 1997
rect 13792 1929 13858 1963
rect 13792 1895 13808 1929
rect 13842 1895 13858 1929
rect 13792 1861 13858 1895
rect 13792 1827 13808 1861
rect 13842 1827 13858 1861
rect 13792 1786 13858 1827
rect 13888 2745 13954 2786
rect 13888 2711 13904 2745
rect 13938 2711 13954 2745
rect 13888 2677 13954 2711
rect 13888 2643 13904 2677
rect 13938 2643 13954 2677
rect 13888 2609 13954 2643
rect 13888 2575 13904 2609
rect 13938 2575 13954 2609
rect 13888 2541 13954 2575
rect 13888 2507 13904 2541
rect 13938 2507 13954 2541
rect 13888 2473 13954 2507
rect 13888 2439 13904 2473
rect 13938 2439 13954 2473
rect 13888 2405 13954 2439
rect 13888 2371 13904 2405
rect 13938 2371 13954 2405
rect 13888 2337 13954 2371
rect 13888 2303 13904 2337
rect 13938 2303 13954 2337
rect 13888 2269 13954 2303
rect 13888 2235 13904 2269
rect 13938 2235 13954 2269
rect 13888 2201 13954 2235
rect 13888 2167 13904 2201
rect 13938 2167 13954 2201
rect 13888 2133 13954 2167
rect 13888 2099 13904 2133
rect 13938 2099 13954 2133
rect 13888 2065 13954 2099
rect 13888 2031 13904 2065
rect 13938 2031 13954 2065
rect 13888 1997 13954 2031
rect 13888 1963 13904 1997
rect 13938 1963 13954 1997
rect 13888 1929 13954 1963
rect 13888 1895 13904 1929
rect 13938 1895 13954 1929
rect 13888 1861 13954 1895
rect 13888 1827 13904 1861
rect 13938 1827 13954 1861
rect 13888 1786 13954 1827
rect 13984 2745 14050 2786
rect 13984 2711 14000 2745
rect 14034 2711 14050 2745
rect 13984 2677 14050 2711
rect 13984 2643 14000 2677
rect 14034 2643 14050 2677
rect 13984 2609 14050 2643
rect 13984 2575 14000 2609
rect 14034 2575 14050 2609
rect 13984 2541 14050 2575
rect 13984 2507 14000 2541
rect 14034 2507 14050 2541
rect 13984 2473 14050 2507
rect 13984 2439 14000 2473
rect 14034 2439 14050 2473
rect 13984 2405 14050 2439
rect 13984 2371 14000 2405
rect 14034 2371 14050 2405
rect 13984 2337 14050 2371
rect 13984 2303 14000 2337
rect 14034 2303 14050 2337
rect 13984 2269 14050 2303
rect 13984 2235 14000 2269
rect 14034 2235 14050 2269
rect 13984 2201 14050 2235
rect 13984 2167 14000 2201
rect 14034 2167 14050 2201
rect 13984 2133 14050 2167
rect 13984 2099 14000 2133
rect 14034 2099 14050 2133
rect 13984 2065 14050 2099
rect 13984 2031 14000 2065
rect 14034 2031 14050 2065
rect 13984 1997 14050 2031
rect 13984 1963 14000 1997
rect 14034 1963 14050 1997
rect 13984 1929 14050 1963
rect 13984 1895 14000 1929
rect 14034 1895 14050 1929
rect 13984 1861 14050 1895
rect 13984 1827 14000 1861
rect 14034 1827 14050 1861
rect 13984 1786 14050 1827
rect 14080 2745 14142 2786
rect 14080 2711 14096 2745
rect 14130 2711 14142 2745
rect 14080 2677 14142 2711
rect 14080 2643 14096 2677
rect 14130 2643 14142 2677
rect 14080 2609 14142 2643
rect 14080 2575 14096 2609
rect 14130 2575 14142 2609
rect 14080 2541 14142 2575
rect 14080 2507 14096 2541
rect 14130 2507 14142 2541
rect 14080 2473 14142 2507
rect 14080 2439 14096 2473
rect 14130 2439 14142 2473
rect 14080 2405 14142 2439
rect 14080 2371 14096 2405
rect 14130 2371 14142 2405
rect 14080 2337 14142 2371
rect 14080 2303 14096 2337
rect 14130 2303 14142 2337
rect 14080 2269 14142 2303
rect 14080 2235 14096 2269
rect 14130 2235 14142 2269
rect 14080 2201 14142 2235
rect 14080 2167 14096 2201
rect 14130 2167 14142 2201
rect 14080 2133 14142 2167
rect 14080 2099 14096 2133
rect 14130 2099 14142 2133
rect 14080 2065 14142 2099
rect 14488 2261 14546 2276
rect 14488 2227 14500 2261
rect 14534 2227 14546 2261
rect 14488 2193 14546 2227
rect 14488 2159 14500 2193
rect 14534 2159 14546 2193
rect 14488 2125 14546 2159
rect 14488 2091 14500 2125
rect 14534 2091 14546 2125
rect 14488 2076 14546 2091
rect 14646 2261 14704 2276
rect 14646 2227 14658 2261
rect 14692 2227 14704 2261
rect 14646 2193 14704 2227
rect 14646 2159 14658 2193
rect 14692 2159 14704 2193
rect 14646 2125 14704 2159
rect 14646 2091 14658 2125
rect 14692 2091 14704 2125
rect 14646 2076 14704 2091
rect 14080 2031 14096 2065
rect 14130 2031 14142 2065
rect 14080 1997 14142 2031
rect 14080 1963 14096 1997
rect 14130 1963 14142 1997
rect 14080 1929 14142 1963
rect 14080 1895 14096 1929
rect 14130 1895 14142 1929
rect 14080 1861 14142 1895
rect 14080 1827 14096 1861
rect 14130 1827 14142 1861
rect 14080 1786 14142 1827
rect 146 1227 208 1268
rect 146 1193 158 1227
rect 192 1193 208 1227
rect 146 1159 208 1193
rect 146 1125 158 1159
rect 192 1125 208 1159
rect 146 1091 208 1125
rect -1698 1025 -1640 1066
rect -1698 991 -1686 1025
rect -1652 991 -1640 1025
rect -1698 957 -1640 991
rect -1698 923 -1686 957
rect -1652 923 -1640 957
rect -1698 889 -1640 923
rect -1698 855 -1686 889
rect -1652 855 -1640 889
rect -1698 821 -1640 855
rect -1698 787 -1686 821
rect -1652 787 -1640 821
rect -1698 753 -1640 787
rect -1698 719 -1686 753
rect -1652 719 -1640 753
rect -1698 685 -1640 719
rect -1698 651 -1686 685
rect -1652 651 -1640 685
rect -1698 617 -1640 651
rect -1698 583 -1686 617
rect -1652 583 -1640 617
rect -1698 549 -1640 583
rect -1698 515 -1686 549
rect -1652 515 -1640 549
rect -1698 481 -1640 515
rect -1698 447 -1686 481
rect -1652 447 -1640 481
rect -1698 413 -1640 447
rect -1698 379 -1686 413
rect -1652 379 -1640 413
rect -1698 345 -1640 379
rect -1698 311 -1686 345
rect -1652 311 -1640 345
rect -1698 277 -1640 311
rect -1698 243 -1686 277
rect -1652 243 -1640 277
rect -1698 209 -1640 243
rect -1698 175 -1686 209
rect -1652 175 -1640 209
rect -1698 141 -1640 175
rect -1698 107 -1686 141
rect -1652 107 -1640 141
rect -1698 66 -1640 107
rect -1600 1025 -1542 1066
rect -1600 991 -1588 1025
rect -1554 991 -1542 1025
rect -1600 957 -1542 991
rect -1600 923 -1588 957
rect -1554 923 -1542 957
rect -1600 889 -1542 923
rect -1600 855 -1588 889
rect -1554 855 -1542 889
rect -1600 821 -1542 855
rect -1600 787 -1588 821
rect -1554 787 -1542 821
rect -1600 753 -1542 787
rect -1600 719 -1588 753
rect -1554 719 -1542 753
rect -1600 685 -1542 719
rect -1600 651 -1588 685
rect -1554 651 -1542 685
rect -1600 617 -1542 651
rect -1600 583 -1588 617
rect -1554 583 -1542 617
rect -1600 549 -1542 583
rect -1600 515 -1588 549
rect -1554 515 -1542 549
rect -1600 481 -1542 515
rect -1600 447 -1588 481
rect -1554 447 -1542 481
rect -1600 413 -1542 447
rect -1600 379 -1588 413
rect -1554 379 -1542 413
rect -1600 345 -1542 379
rect -1600 311 -1588 345
rect -1554 311 -1542 345
rect -1600 277 -1542 311
rect -1600 243 -1588 277
rect -1554 243 -1542 277
rect -1600 209 -1542 243
rect -1600 175 -1588 209
rect -1554 175 -1542 209
rect -1600 141 -1542 175
rect -1600 107 -1588 141
rect -1554 107 -1542 141
rect -1600 66 -1542 107
rect -1502 1025 -1444 1066
rect -1502 991 -1490 1025
rect -1456 991 -1444 1025
rect -1502 957 -1444 991
rect -1502 923 -1490 957
rect -1456 923 -1444 957
rect -1502 889 -1444 923
rect -1502 855 -1490 889
rect -1456 855 -1444 889
rect -1502 821 -1444 855
rect -1502 787 -1490 821
rect -1456 787 -1444 821
rect -1502 753 -1444 787
rect -1502 719 -1490 753
rect -1456 719 -1444 753
rect -1502 685 -1444 719
rect -1502 651 -1490 685
rect -1456 651 -1444 685
rect -1502 617 -1444 651
rect -1502 583 -1490 617
rect -1456 583 -1444 617
rect -1502 549 -1444 583
rect -1502 515 -1490 549
rect -1456 515 -1444 549
rect -1502 481 -1444 515
rect -1502 447 -1490 481
rect -1456 447 -1444 481
rect -1502 413 -1444 447
rect -1502 379 -1490 413
rect -1456 379 -1444 413
rect -1502 345 -1444 379
rect -1502 311 -1490 345
rect -1456 311 -1444 345
rect -1502 277 -1444 311
rect -1502 243 -1490 277
rect -1456 243 -1444 277
rect -1502 209 -1444 243
rect -1502 175 -1490 209
rect -1456 175 -1444 209
rect -1502 141 -1444 175
rect -1502 107 -1490 141
rect -1456 107 -1444 141
rect -1502 66 -1444 107
rect -1404 1025 -1346 1066
rect -1404 991 -1392 1025
rect -1358 991 -1346 1025
rect -1404 957 -1346 991
rect -1404 923 -1392 957
rect -1358 923 -1346 957
rect -1404 889 -1346 923
rect -1404 855 -1392 889
rect -1358 855 -1346 889
rect -1404 821 -1346 855
rect -1404 787 -1392 821
rect -1358 787 -1346 821
rect -1404 753 -1346 787
rect -1404 719 -1392 753
rect -1358 719 -1346 753
rect -1404 685 -1346 719
rect -1404 651 -1392 685
rect -1358 651 -1346 685
rect -1404 617 -1346 651
rect -1404 583 -1392 617
rect -1358 583 -1346 617
rect -1404 549 -1346 583
rect -1404 515 -1392 549
rect -1358 515 -1346 549
rect -1404 481 -1346 515
rect -1404 447 -1392 481
rect -1358 447 -1346 481
rect -1404 413 -1346 447
rect -1404 379 -1392 413
rect -1358 379 -1346 413
rect -1404 345 -1346 379
rect -1404 311 -1392 345
rect -1358 311 -1346 345
rect -1404 277 -1346 311
rect -1404 243 -1392 277
rect -1358 243 -1346 277
rect -1404 209 -1346 243
rect -1404 175 -1392 209
rect -1358 175 -1346 209
rect -1404 141 -1346 175
rect -1404 107 -1392 141
rect -1358 107 -1346 141
rect -1404 66 -1346 107
rect -1306 1025 -1248 1066
rect -1306 991 -1294 1025
rect -1260 991 -1248 1025
rect -1306 957 -1248 991
rect -1306 923 -1294 957
rect -1260 923 -1248 957
rect -1306 889 -1248 923
rect -1306 855 -1294 889
rect -1260 855 -1248 889
rect -1306 821 -1248 855
rect -1306 787 -1294 821
rect -1260 787 -1248 821
rect -1306 753 -1248 787
rect -1306 719 -1294 753
rect -1260 719 -1248 753
rect -1306 685 -1248 719
rect -1306 651 -1294 685
rect -1260 651 -1248 685
rect -1306 617 -1248 651
rect -1306 583 -1294 617
rect -1260 583 -1248 617
rect -1306 549 -1248 583
rect -1306 515 -1294 549
rect -1260 515 -1248 549
rect -1306 481 -1248 515
rect -1306 447 -1294 481
rect -1260 447 -1248 481
rect -1306 413 -1248 447
rect -1306 379 -1294 413
rect -1260 379 -1248 413
rect -1306 345 -1248 379
rect -1306 311 -1294 345
rect -1260 311 -1248 345
rect -1306 277 -1248 311
rect -1306 243 -1294 277
rect -1260 243 -1248 277
rect -1306 209 -1248 243
rect -1306 175 -1294 209
rect -1260 175 -1248 209
rect -1306 141 -1248 175
rect -1306 107 -1294 141
rect -1260 107 -1248 141
rect -1306 66 -1248 107
rect -1208 1025 -1150 1066
rect -1208 991 -1196 1025
rect -1162 991 -1150 1025
rect -1208 957 -1150 991
rect -1208 923 -1196 957
rect -1162 923 -1150 957
rect -1208 889 -1150 923
rect -1208 855 -1196 889
rect -1162 855 -1150 889
rect -1208 821 -1150 855
rect -1208 787 -1196 821
rect -1162 787 -1150 821
rect -1208 753 -1150 787
rect -1208 719 -1196 753
rect -1162 719 -1150 753
rect -1208 685 -1150 719
rect -1208 651 -1196 685
rect -1162 651 -1150 685
rect -1208 617 -1150 651
rect -1208 583 -1196 617
rect -1162 583 -1150 617
rect -1208 549 -1150 583
rect -1208 515 -1196 549
rect -1162 515 -1150 549
rect -1208 481 -1150 515
rect -1208 447 -1196 481
rect -1162 447 -1150 481
rect -1208 413 -1150 447
rect -1208 379 -1196 413
rect -1162 379 -1150 413
rect -1208 345 -1150 379
rect -1208 311 -1196 345
rect -1162 311 -1150 345
rect -1208 277 -1150 311
rect -1208 243 -1196 277
rect -1162 243 -1150 277
rect -1208 209 -1150 243
rect -1208 175 -1196 209
rect -1162 175 -1150 209
rect -1208 141 -1150 175
rect -1208 107 -1196 141
rect -1162 107 -1150 141
rect -1208 66 -1150 107
rect -1110 1025 -1052 1066
rect -1110 991 -1098 1025
rect -1064 991 -1052 1025
rect -1110 957 -1052 991
rect -1110 923 -1098 957
rect -1064 923 -1052 957
rect -1110 889 -1052 923
rect -1110 855 -1098 889
rect -1064 855 -1052 889
rect -1110 821 -1052 855
rect -1110 787 -1098 821
rect -1064 787 -1052 821
rect -1110 753 -1052 787
rect -1110 719 -1098 753
rect -1064 719 -1052 753
rect -1110 685 -1052 719
rect -1110 651 -1098 685
rect -1064 651 -1052 685
rect -1110 617 -1052 651
rect -1110 583 -1098 617
rect -1064 583 -1052 617
rect -1110 549 -1052 583
rect -1110 515 -1098 549
rect -1064 515 -1052 549
rect -1110 481 -1052 515
rect -1110 447 -1098 481
rect -1064 447 -1052 481
rect -1110 413 -1052 447
rect -1110 379 -1098 413
rect -1064 379 -1052 413
rect -1110 345 -1052 379
rect -1110 311 -1098 345
rect -1064 311 -1052 345
rect -1110 277 -1052 311
rect -1110 243 -1098 277
rect -1064 243 -1052 277
rect -1110 209 -1052 243
rect -1110 175 -1098 209
rect -1064 175 -1052 209
rect -1110 141 -1052 175
rect -1110 107 -1098 141
rect -1064 107 -1052 141
rect -1110 66 -1052 107
rect -1012 1025 -954 1066
rect -1012 991 -1000 1025
rect -966 991 -954 1025
rect -1012 957 -954 991
rect -1012 923 -1000 957
rect -966 923 -954 957
rect -1012 889 -954 923
rect -1012 855 -1000 889
rect -966 855 -954 889
rect -1012 821 -954 855
rect -1012 787 -1000 821
rect -966 787 -954 821
rect -1012 753 -954 787
rect -1012 719 -1000 753
rect -966 719 -954 753
rect -1012 685 -954 719
rect -1012 651 -1000 685
rect -966 651 -954 685
rect -1012 617 -954 651
rect -1012 583 -1000 617
rect -966 583 -954 617
rect -1012 549 -954 583
rect -1012 515 -1000 549
rect -966 515 -954 549
rect -1012 481 -954 515
rect -1012 447 -1000 481
rect -966 447 -954 481
rect -1012 413 -954 447
rect -1012 379 -1000 413
rect -966 379 -954 413
rect -1012 345 -954 379
rect -1012 311 -1000 345
rect -966 311 -954 345
rect -1012 277 -954 311
rect -1012 243 -1000 277
rect -966 243 -954 277
rect -1012 209 -954 243
rect -1012 175 -1000 209
rect -966 175 -954 209
rect -1012 141 -954 175
rect -1012 107 -1000 141
rect -966 107 -954 141
rect -1012 66 -954 107
rect -914 1025 -856 1066
rect -914 991 -902 1025
rect -868 991 -856 1025
rect -914 957 -856 991
rect -914 923 -902 957
rect -868 923 -856 957
rect -914 889 -856 923
rect -914 855 -902 889
rect -868 855 -856 889
rect -914 821 -856 855
rect -914 787 -902 821
rect -868 787 -856 821
rect -914 753 -856 787
rect -914 719 -902 753
rect -868 719 -856 753
rect -914 685 -856 719
rect -914 651 -902 685
rect -868 651 -856 685
rect -914 617 -856 651
rect -914 583 -902 617
rect -868 583 -856 617
rect -914 549 -856 583
rect -914 515 -902 549
rect -868 515 -856 549
rect -914 481 -856 515
rect -914 447 -902 481
rect -868 447 -856 481
rect -914 413 -856 447
rect -914 379 -902 413
rect -868 379 -856 413
rect -914 345 -856 379
rect -914 311 -902 345
rect -868 311 -856 345
rect -914 277 -856 311
rect -914 243 -902 277
rect -868 243 -856 277
rect 146 1057 158 1091
rect 192 1057 208 1091
rect 146 1023 208 1057
rect 146 989 158 1023
rect 192 989 208 1023
rect 146 955 208 989
rect 146 921 158 955
rect 192 921 208 955
rect 146 887 208 921
rect 146 853 158 887
rect 192 853 208 887
rect 146 819 208 853
rect 146 785 158 819
rect 192 785 208 819
rect 146 751 208 785
rect 146 717 158 751
rect 192 717 208 751
rect 146 683 208 717
rect 146 649 158 683
rect 192 649 208 683
rect 146 615 208 649
rect 146 581 158 615
rect 192 581 208 615
rect 146 547 208 581
rect 146 513 158 547
rect 192 513 208 547
rect 146 479 208 513
rect 146 445 158 479
rect 192 445 208 479
rect 146 411 208 445
rect 146 377 158 411
rect 192 377 208 411
rect 146 343 208 377
rect 146 309 158 343
rect 192 309 208 343
rect 146 268 208 309
rect 238 1227 304 1268
rect 238 1193 254 1227
rect 288 1193 304 1227
rect 238 1159 304 1193
rect 238 1125 254 1159
rect 288 1125 304 1159
rect 238 1091 304 1125
rect 238 1057 254 1091
rect 288 1057 304 1091
rect 238 1023 304 1057
rect 238 989 254 1023
rect 288 989 304 1023
rect 238 955 304 989
rect 238 921 254 955
rect 288 921 304 955
rect 238 887 304 921
rect 238 853 254 887
rect 288 853 304 887
rect 238 819 304 853
rect 238 785 254 819
rect 288 785 304 819
rect 238 751 304 785
rect 238 717 254 751
rect 288 717 304 751
rect 238 683 304 717
rect 238 649 254 683
rect 288 649 304 683
rect 238 615 304 649
rect 238 581 254 615
rect 288 581 304 615
rect 238 547 304 581
rect 238 513 254 547
rect 288 513 304 547
rect 238 479 304 513
rect 238 445 254 479
rect 288 445 304 479
rect 238 411 304 445
rect 238 377 254 411
rect 288 377 304 411
rect 238 343 304 377
rect 238 309 254 343
rect 288 309 304 343
rect 238 268 304 309
rect 334 1227 400 1268
rect 334 1193 350 1227
rect 384 1193 400 1227
rect 334 1159 400 1193
rect 334 1125 350 1159
rect 384 1125 400 1159
rect 334 1091 400 1125
rect 334 1057 350 1091
rect 384 1057 400 1091
rect 334 1023 400 1057
rect 334 989 350 1023
rect 384 989 400 1023
rect 334 955 400 989
rect 334 921 350 955
rect 384 921 400 955
rect 334 887 400 921
rect 334 853 350 887
rect 384 853 400 887
rect 334 819 400 853
rect 334 785 350 819
rect 384 785 400 819
rect 334 751 400 785
rect 334 717 350 751
rect 384 717 400 751
rect 334 683 400 717
rect 334 649 350 683
rect 384 649 400 683
rect 334 615 400 649
rect 334 581 350 615
rect 384 581 400 615
rect 334 547 400 581
rect 334 513 350 547
rect 384 513 400 547
rect 334 479 400 513
rect 334 445 350 479
rect 384 445 400 479
rect 334 411 400 445
rect 334 377 350 411
rect 384 377 400 411
rect 334 343 400 377
rect 334 309 350 343
rect 384 309 400 343
rect 334 268 400 309
rect 430 1227 496 1268
rect 430 1193 446 1227
rect 480 1193 496 1227
rect 430 1159 496 1193
rect 430 1125 446 1159
rect 480 1125 496 1159
rect 430 1091 496 1125
rect 430 1057 446 1091
rect 480 1057 496 1091
rect 430 1023 496 1057
rect 430 989 446 1023
rect 480 989 496 1023
rect 430 955 496 989
rect 430 921 446 955
rect 480 921 496 955
rect 430 887 496 921
rect 430 853 446 887
rect 480 853 496 887
rect 430 819 496 853
rect 430 785 446 819
rect 480 785 496 819
rect 430 751 496 785
rect 430 717 446 751
rect 480 717 496 751
rect 430 683 496 717
rect 430 649 446 683
rect 480 649 496 683
rect 430 615 496 649
rect 430 581 446 615
rect 480 581 496 615
rect 430 547 496 581
rect 430 513 446 547
rect 480 513 496 547
rect 430 479 496 513
rect 430 445 446 479
rect 480 445 496 479
rect 430 411 496 445
rect 430 377 446 411
rect 480 377 496 411
rect 430 343 496 377
rect 430 309 446 343
rect 480 309 496 343
rect 430 268 496 309
rect 526 1227 592 1268
rect 526 1193 542 1227
rect 576 1193 592 1227
rect 526 1159 592 1193
rect 526 1125 542 1159
rect 576 1125 592 1159
rect 526 1091 592 1125
rect 526 1057 542 1091
rect 576 1057 592 1091
rect 526 1023 592 1057
rect 526 989 542 1023
rect 576 989 592 1023
rect 526 955 592 989
rect 526 921 542 955
rect 576 921 592 955
rect 526 887 592 921
rect 526 853 542 887
rect 576 853 592 887
rect 526 819 592 853
rect 526 785 542 819
rect 576 785 592 819
rect 526 751 592 785
rect 526 717 542 751
rect 576 717 592 751
rect 526 683 592 717
rect 526 649 542 683
rect 576 649 592 683
rect 526 615 592 649
rect 526 581 542 615
rect 576 581 592 615
rect 526 547 592 581
rect 526 513 542 547
rect 576 513 592 547
rect 526 479 592 513
rect 526 445 542 479
rect 576 445 592 479
rect 526 411 592 445
rect 526 377 542 411
rect 576 377 592 411
rect 526 343 592 377
rect 526 309 542 343
rect 576 309 592 343
rect 526 268 592 309
rect 622 1227 688 1268
rect 622 1193 638 1227
rect 672 1193 688 1227
rect 622 1159 688 1193
rect 622 1125 638 1159
rect 672 1125 688 1159
rect 622 1091 688 1125
rect 622 1057 638 1091
rect 672 1057 688 1091
rect 622 1023 688 1057
rect 622 989 638 1023
rect 672 989 688 1023
rect 622 955 688 989
rect 622 921 638 955
rect 672 921 688 955
rect 622 887 688 921
rect 622 853 638 887
rect 672 853 688 887
rect 622 819 688 853
rect 622 785 638 819
rect 672 785 688 819
rect 622 751 688 785
rect 622 717 638 751
rect 672 717 688 751
rect 622 683 688 717
rect 622 649 638 683
rect 672 649 688 683
rect 622 615 688 649
rect 622 581 638 615
rect 672 581 688 615
rect 622 547 688 581
rect 622 513 638 547
rect 672 513 688 547
rect 622 479 688 513
rect 622 445 638 479
rect 672 445 688 479
rect 622 411 688 445
rect 622 377 638 411
rect 672 377 688 411
rect 622 343 688 377
rect 622 309 638 343
rect 672 309 688 343
rect 622 268 688 309
rect 718 1227 784 1268
rect 718 1193 734 1227
rect 768 1193 784 1227
rect 718 1159 784 1193
rect 718 1125 734 1159
rect 768 1125 784 1159
rect 718 1091 784 1125
rect 718 1057 734 1091
rect 768 1057 784 1091
rect 718 1023 784 1057
rect 718 989 734 1023
rect 768 989 784 1023
rect 718 955 784 989
rect 718 921 734 955
rect 768 921 784 955
rect 718 887 784 921
rect 718 853 734 887
rect 768 853 784 887
rect 718 819 784 853
rect 718 785 734 819
rect 768 785 784 819
rect 718 751 784 785
rect 718 717 734 751
rect 768 717 784 751
rect 718 683 784 717
rect 718 649 734 683
rect 768 649 784 683
rect 718 615 784 649
rect 718 581 734 615
rect 768 581 784 615
rect 718 547 784 581
rect 718 513 734 547
rect 768 513 784 547
rect 718 479 784 513
rect 718 445 734 479
rect 768 445 784 479
rect 718 411 784 445
rect 718 377 734 411
rect 768 377 784 411
rect 718 343 784 377
rect 718 309 734 343
rect 768 309 784 343
rect 718 268 784 309
rect 814 1227 880 1268
rect 814 1193 830 1227
rect 864 1193 880 1227
rect 814 1159 880 1193
rect 814 1125 830 1159
rect 864 1125 880 1159
rect 814 1091 880 1125
rect 814 1057 830 1091
rect 864 1057 880 1091
rect 814 1023 880 1057
rect 814 989 830 1023
rect 864 989 880 1023
rect 814 955 880 989
rect 814 921 830 955
rect 864 921 880 955
rect 814 887 880 921
rect 814 853 830 887
rect 864 853 880 887
rect 814 819 880 853
rect 814 785 830 819
rect 864 785 880 819
rect 814 751 880 785
rect 814 717 830 751
rect 864 717 880 751
rect 814 683 880 717
rect 814 649 830 683
rect 864 649 880 683
rect 814 615 880 649
rect 814 581 830 615
rect 864 581 880 615
rect 814 547 880 581
rect 814 513 830 547
rect 864 513 880 547
rect 814 479 880 513
rect 814 445 830 479
rect 864 445 880 479
rect 814 411 880 445
rect 814 377 830 411
rect 864 377 880 411
rect 814 343 880 377
rect 814 309 830 343
rect 864 309 880 343
rect 814 268 880 309
rect 910 1227 976 1268
rect 910 1193 926 1227
rect 960 1193 976 1227
rect 910 1159 976 1193
rect 910 1125 926 1159
rect 960 1125 976 1159
rect 910 1091 976 1125
rect 910 1057 926 1091
rect 960 1057 976 1091
rect 910 1023 976 1057
rect 910 989 926 1023
rect 960 989 976 1023
rect 910 955 976 989
rect 910 921 926 955
rect 960 921 976 955
rect 910 887 976 921
rect 910 853 926 887
rect 960 853 976 887
rect 910 819 976 853
rect 910 785 926 819
rect 960 785 976 819
rect 910 751 976 785
rect 910 717 926 751
rect 960 717 976 751
rect 910 683 976 717
rect 910 649 926 683
rect 960 649 976 683
rect 910 615 976 649
rect 910 581 926 615
rect 960 581 976 615
rect 910 547 976 581
rect 910 513 926 547
rect 960 513 976 547
rect 910 479 976 513
rect 910 445 926 479
rect 960 445 976 479
rect 910 411 976 445
rect 910 377 926 411
rect 960 377 976 411
rect 910 343 976 377
rect 910 309 926 343
rect 960 309 976 343
rect 910 268 976 309
rect 1006 1227 1072 1268
rect 1006 1193 1022 1227
rect 1056 1193 1072 1227
rect 1006 1159 1072 1193
rect 1006 1125 1022 1159
rect 1056 1125 1072 1159
rect 1006 1091 1072 1125
rect 1006 1057 1022 1091
rect 1056 1057 1072 1091
rect 1006 1023 1072 1057
rect 1006 989 1022 1023
rect 1056 989 1072 1023
rect 1006 955 1072 989
rect 1006 921 1022 955
rect 1056 921 1072 955
rect 1006 887 1072 921
rect 1006 853 1022 887
rect 1056 853 1072 887
rect 1006 819 1072 853
rect 1006 785 1022 819
rect 1056 785 1072 819
rect 1006 751 1072 785
rect 1006 717 1022 751
rect 1056 717 1072 751
rect 1006 683 1072 717
rect 1006 649 1022 683
rect 1056 649 1072 683
rect 1006 615 1072 649
rect 1006 581 1022 615
rect 1056 581 1072 615
rect 1006 547 1072 581
rect 1006 513 1022 547
rect 1056 513 1072 547
rect 1006 479 1072 513
rect 1006 445 1022 479
rect 1056 445 1072 479
rect 1006 411 1072 445
rect 1006 377 1022 411
rect 1056 377 1072 411
rect 1006 343 1072 377
rect 1006 309 1022 343
rect 1056 309 1072 343
rect 1006 268 1072 309
rect 1102 1227 1168 1268
rect 1102 1193 1118 1227
rect 1152 1193 1168 1227
rect 1102 1159 1168 1193
rect 1102 1125 1118 1159
rect 1152 1125 1168 1159
rect 1102 1091 1168 1125
rect 1102 1057 1118 1091
rect 1152 1057 1168 1091
rect 1102 1023 1168 1057
rect 1102 989 1118 1023
rect 1152 989 1168 1023
rect 1102 955 1168 989
rect 1102 921 1118 955
rect 1152 921 1168 955
rect 1102 887 1168 921
rect 1102 853 1118 887
rect 1152 853 1168 887
rect 1102 819 1168 853
rect 1102 785 1118 819
rect 1152 785 1168 819
rect 1102 751 1168 785
rect 1102 717 1118 751
rect 1152 717 1168 751
rect 1102 683 1168 717
rect 1102 649 1118 683
rect 1152 649 1168 683
rect 1102 615 1168 649
rect 1102 581 1118 615
rect 1152 581 1168 615
rect 1102 547 1168 581
rect 1102 513 1118 547
rect 1152 513 1168 547
rect 1102 479 1168 513
rect 1102 445 1118 479
rect 1152 445 1168 479
rect 1102 411 1168 445
rect 1102 377 1118 411
rect 1152 377 1168 411
rect 1102 343 1168 377
rect 1102 309 1118 343
rect 1152 309 1168 343
rect 1102 268 1168 309
rect 1198 1227 1264 1268
rect 1198 1193 1214 1227
rect 1248 1193 1264 1227
rect 1198 1159 1264 1193
rect 1198 1125 1214 1159
rect 1248 1125 1264 1159
rect 1198 1091 1264 1125
rect 1198 1057 1214 1091
rect 1248 1057 1264 1091
rect 1198 1023 1264 1057
rect 1198 989 1214 1023
rect 1248 989 1264 1023
rect 1198 955 1264 989
rect 1198 921 1214 955
rect 1248 921 1264 955
rect 1198 887 1264 921
rect 1198 853 1214 887
rect 1248 853 1264 887
rect 1198 819 1264 853
rect 1198 785 1214 819
rect 1248 785 1264 819
rect 1198 751 1264 785
rect 1198 717 1214 751
rect 1248 717 1264 751
rect 1198 683 1264 717
rect 1198 649 1214 683
rect 1248 649 1264 683
rect 1198 615 1264 649
rect 1198 581 1214 615
rect 1248 581 1264 615
rect 1198 547 1264 581
rect 1198 513 1214 547
rect 1248 513 1264 547
rect 1198 479 1264 513
rect 1198 445 1214 479
rect 1248 445 1264 479
rect 1198 411 1264 445
rect 1198 377 1214 411
rect 1248 377 1264 411
rect 1198 343 1264 377
rect 1198 309 1214 343
rect 1248 309 1264 343
rect 1198 268 1264 309
rect 1294 1227 1356 1268
rect 1294 1193 1310 1227
rect 1344 1193 1356 1227
rect 1294 1159 1356 1193
rect 1294 1125 1310 1159
rect 1344 1125 1356 1159
rect 1294 1091 1356 1125
rect 1294 1057 1310 1091
rect 1344 1057 1356 1091
rect 1294 1023 1356 1057
rect 1294 989 1310 1023
rect 1344 989 1356 1023
rect 1294 955 1356 989
rect 1294 921 1310 955
rect 1344 921 1356 955
rect 1294 887 1356 921
rect 1294 853 1310 887
rect 1344 853 1356 887
rect 1294 819 1356 853
rect 1294 785 1310 819
rect 1344 785 1356 819
rect 1294 751 1356 785
rect 1294 717 1310 751
rect 1344 717 1356 751
rect 1294 683 1356 717
rect 1294 649 1310 683
rect 1344 649 1356 683
rect 1294 615 1356 649
rect 1294 581 1310 615
rect 1344 581 1356 615
rect 1294 547 1356 581
rect 1294 513 1310 547
rect 1344 513 1356 547
rect 1294 479 1356 513
rect 1294 445 1310 479
rect 1344 445 1356 479
rect 1294 411 1356 445
rect 1294 377 1310 411
rect 1344 377 1356 411
rect 1294 343 1356 377
rect 1294 309 1310 343
rect 1344 309 1356 343
rect 1294 268 1356 309
rect 1914 1227 1976 1268
rect 1914 1193 1926 1227
rect 1960 1193 1976 1227
rect 1914 1159 1976 1193
rect 1914 1125 1926 1159
rect 1960 1125 1976 1159
rect 1914 1091 1976 1125
rect 1914 1057 1926 1091
rect 1960 1057 1976 1091
rect 1914 1023 1976 1057
rect 1914 989 1926 1023
rect 1960 989 1976 1023
rect 1914 955 1976 989
rect 1914 921 1926 955
rect 1960 921 1976 955
rect 1914 887 1976 921
rect 1914 853 1926 887
rect 1960 853 1976 887
rect 1914 819 1976 853
rect 1914 785 1926 819
rect 1960 785 1976 819
rect 1914 751 1976 785
rect 1914 717 1926 751
rect 1960 717 1976 751
rect 1914 683 1976 717
rect 1914 649 1926 683
rect 1960 649 1976 683
rect 1914 615 1976 649
rect 1914 581 1926 615
rect 1960 581 1976 615
rect 1914 547 1976 581
rect 1914 513 1926 547
rect 1960 513 1976 547
rect 1914 479 1976 513
rect 1914 445 1926 479
rect 1960 445 1976 479
rect 1914 411 1976 445
rect 1914 377 1926 411
rect 1960 377 1976 411
rect 1914 343 1976 377
rect 1914 309 1926 343
rect 1960 309 1976 343
rect 1914 268 1976 309
rect 2006 1227 2072 1268
rect 2006 1193 2022 1227
rect 2056 1193 2072 1227
rect 2006 1159 2072 1193
rect 2006 1125 2022 1159
rect 2056 1125 2072 1159
rect 2006 1091 2072 1125
rect 2006 1057 2022 1091
rect 2056 1057 2072 1091
rect 2006 1023 2072 1057
rect 2006 989 2022 1023
rect 2056 989 2072 1023
rect 2006 955 2072 989
rect 2006 921 2022 955
rect 2056 921 2072 955
rect 2006 887 2072 921
rect 2006 853 2022 887
rect 2056 853 2072 887
rect 2006 819 2072 853
rect 2006 785 2022 819
rect 2056 785 2072 819
rect 2006 751 2072 785
rect 2006 717 2022 751
rect 2056 717 2072 751
rect 2006 683 2072 717
rect 2006 649 2022 683
rect 2056 649 2072 683
rect 2006 615 2072 649
rect 2006 581 2022 615
rect 2056 581 2072 615
rect 2006 547 2072 581
rect 2006 513 2022 547
rect 2056 513 2072 547
rect 2006 479 2072 513
rect 2006 445 2022 479
rect 2056 445 2072 479
rect 2006 411 2072 445
rect 2006 377 2022 411
rect 2056 377 2072 411
rect 2006 343 2072 377
rect 2006 309 2022 343
rect 2056 309 2072 343
rect 2006 268 2072 309
rect 2102 1227 2168 1268
rect 2102 1193 2118 1227
rect 2152 1193 2168 1227
rect 2102 1159 2168 1193
rect 2102 1125 2118 1159
rect 2152 1125 2168 1159
rect 2102 1091 2168 1125
rect 2102 1057 2118 1091
rect 2152 1057 2168 1091
rect 2102 1023 2168 1057
rect 2102 989 2118 1023
rect 2152 989 2168 1023
rect 2102 955 2168 989
rect 2102 921 2118 955
rect 2152 921 2168 955
rect 2102 887 2168 921
rect 2102 853 2118 887
rect 2152 853 2168 887
rect 2102 819 2168 853
rect 2102 785 2118 819
rect 2152 785 2168 819
rect 2102 751 2168 785
rect 2102 717 2118 751
rect 2152 717 2168 751
rect 2102 683 2168 717
rect 2102 649 2118 683
rect 2152 649 2168 683
rect 2102 615 2168 649
rect 2102 581 2118 615
rect 2152 581 2168 615
rect 2102 547 2168 581
rect 2102 513 2118 547
rect 2152 513 2168 547
rect 2102 479 2168 513
rect 2102 445 2118 479
rect 2152 445 2168 479
rect 2102 411 2168 445
rect 2102 377 2118 411
rect 2152 377 2168 411
rect 2102 343 2168 377
rect 2102 309 2118 343
rect 2152 309 2168 343
rect 2102 268 2168 309
rect 2198 1227 2264 1268
rect 2198 1193 2214 1227
rect 2248 1193 2264 1227
rect 2198 1159 2264 1193
rect 2198 1125 2214 1159
rect 2248 1125 2264 1159
rect 2198 1091 2264 1125
rect 2198 1057 2214 1091
rect 2248 1057 2264 1091
rect 2198 1023 2264 1057
rect 2198 989 2214 1023
rect 2248 989 2264 1023
rect 2198 955 2264 989
rect 2198 921 2214 955
rect 2248 921 2264 955
rect 2198 887 2264 921
rect 2198 853 2214 887
rect 2248 853 2264 887
rect 2198 819 2264 853
rect 2198 785 2214 819
rect 2248 785 2264 819
rect 2198 751 2264 785
rect 2198 717 2214 751
rect 2248 717 2264 751
rect 2198 683 2264 717
rect 2198 649 2214 683
rect 2248 649 2264 683
rect 2198 615 2264 649
rect 2198 581 2214 615
rect 2248 581 2264 615
rect 2198 547 2264 581
rect 2198 513 2214 547
rect 2248 513 2264 547
rect 2198 479 2264 513
rect 2198 445 2214 479
rect 2248 445 2264 479
rect 2198 411 2264 445
rect 2198 377 2214 411
rect 2248 377 2264 411
rect 2198 343 2264 377
rect 2198 309 2214 343
rect 2248 309 2264 343
rect 2198 268 2264 309
rect 2294 1227 2360 1268
rect 2294 1193 2310 1227
rect 2344 1193 2360 1227
rect 2294 1159 2360 1193
rect 2294 1125 2310 1159
rect 2344 1125 2360 1159
rect 2294 1091 2360 1125
rect 2294 1057 2310 1091
rect 2344 1057 2360 1091
rect 2294 1023 2360 1057
rect 2294 989 2310 1023
rect 2344 989 2360 1023
rect 2294 955 2360 989
rect 2294 921 2310 955
rect 2344 921 2360 955
rect 2294 887 2360 921
rect 2294 853 2310 887
rect 2344 853 2360 887
rect 2294 819 2360 853
rect 2294 785 2310 819
rect 2344 785 2360 819
rect 2294 751 2360 785
rect 2294 717 2310 751
rect 2344 717 2360 751
rect 2294 683 2360 717
rect 2294 649 2310 683
rect 2344 649 2360 683
rect 2294 615 2360 649
rect 2294 581 2310 615
rect 2344 581 2360 615
rect 2294 547 2360 581
rect 2294 513 2310 547
rect 2344 513 2360 547
rect 2294 479 2360 513
rect 2294 445 2310 479
rect 2344 445 2360 479
rect 2294 411 2360 445
rect 2294 377 2310 411
rect 2344 377 2360 411
rect 2294 343 2360 377
rect 2294 309 2310 343
rect 2344 309 2360 343
rect 2294 268 2360 309
rect 2390 1227 2456 1268
rect 2390 1193 2406 1227
rect 2440 1193 2456 1227
rect 2390 1159 2456 1193
rect 2390 1125 2406 1159
rect 2440 1125 2456 1159
rect 2390 1091 2456 1125
rect 2390 1057 2406 1091
rect 2440 1057 2456 1091
rect 2390 1023 2456 1057
rect 2390 989 2406 1023
rect 2440 989 2456 1023
rect 2390 955 2456 989
rect 2390 921 2406 955
rect 2440 921 2456 955
rect 2390 887 2456 921
rect 2390 853 2406 887
rect 2440 853 2456 887
rect 2390 819 2456 853
rect 2390 785 2406 819
rect 2440 785 2456 819
rect 2390 751 2456 785
rect 2390 717 2406 751
rect 2440 717 2456 751
rect 2390 683 2456 717
rect 2390 649 2406 683
rect 2440 649 2456 683
rect 2390 615 2456 649
rect 2390 581 2406 615
rect 2440 581 2456 615
rect 2390 547 2456 581
rect 2390 513 2406 547
rect 2440 513 2456 547
rect 2390 479 2456 513
rect 2390 445 2406 479
rect 2440 445 2456 479
rect 2390 411 2456 445
rect 2390 377 2406 411
rect 2440 377 2456 411
rect 2390 343 2456 377
rect 2390 309 2406 343
rect 2440 309 2456 343
rect 2390 268 2456 309
rect 2486 1227 2552 1268
rect 2486 1193 2502 1227
rect 2536 1193 2552 1227
rect 2486 1159 2552 1193
rect 2486 1125 2502 1159
rect 2536 1125 2552 1159
rect 2486 1091 2552 1125
rect 2486 1057 2502 1091
rect 2536 1057 2552 1091
rect 2486 1023 2552 1057
rect 2486 989 2502 1023
rect 2536 989 2552 1023
rect 2486 955 2552 989
rect 2486 921 2502 955
rect 2536 921 2552 955
rect 2486 887 2552 921
rect 2486 853 2502 887
rect 2536 853 2552 887
rect 2486 819 2552 853
rect 2486 785 2502 819
rect 2536 785 2552 819
rect 2486 751 2552 785
rect 2486 717 2502 751
rect 2536 717 2552 751
rect 2486 683 2552 717
rect 2486 649 2502 683
rect 2536 649 2552 683
rect 2486 615 2552 649
rect 2486 581 2502 615
rect 2536 581 2552 615
rect 2486 547 2552 581
rect 2486 513 2502 547
rect 2536 513 2552 547
rect 2486 479 2552 513
rect 2486 445 2502 479
rect 2536 445 2552 479
rect 2486 411 2552 445
rect 2486 377 2502 411
rect 2536 377 2552 411
rect 2486 343 2552 377
rect 2486 309 2502 343
rect 2536 309 2552 343
rect 2486 268 2552 309
rect 2582 1227 2648 1268
rect 2582 1193 2598 1227
rect 2632 1193 2648 1227
rect 2582 1159 2648 1193
rect 2582 1125 2598 1159
rect 2632 1125 2648 1159
rect 2582 1091 2648 1125
rect 2582 1057 2598 1091
rect 2632 1057 2648 1091
rect 2582 1023 2648 1057
rect 2582 989 2598 1023
rect 2632 989 2648 1023
rect 2582 955 2648 989
rect 2582 921 2598 955
rect 2632 921 2648 955
rect 2582 887 2648 921
rect 2582 853 2598 887
rect 2632 853 2648 887
rect 2582 819 2648 853
rect 2582 785 2598 819
rect 2632 785 2648 819
rect 2582 751 2648 785
rect 2582 717 2598 751
rect 2632 717 2648 751
rect 2582 683 2648 717
rect 2582 649 2598 683
rect 2632 649 2648 683
rect 2582 615 2648 649
rect 2582 581 2598 615
rect 2632 581 2648 615
rect 2582 547 2648 581
rect 2582 513 2598 547
rect 2632 513 2648 547
rect 2582 479 2648 513
rect 2582 445 2598 479
rect 2632 445 2648 479
rect 2582 411 2648 445
rect 2582 377 2598 411
rect 2632 377 2648 411
rect 2582 343 2648 377
rect 2582 309 2598 343
rect 2632 309 2648 343
rect 2582 268 2648 309
rect 2678 1227 2744 1268
rect 2678 1193 2694 1227
rect 2728 1193 2744 1227
rect 2678 1159 2744 1193
rect 2678 1125 2694 1159
rect 2728 1125 2744 1159
rect 2678 1091 2744 1125
rect 2678 1057 2694 1091
rect 2728 1057 2744 1091
rect 2678 1023 2744 1057
rect 2678 989 2694 1023
rect 2728 989 2744 1023
rect 2678 955 2744 989
rect 2678 921 2694 955
rect 2728 921 2744 955
rect 2678 887 2744 921
rect 2678 853 2694 887
rect 2728 853 2744 887
rect 2678 819 2744 853
rect 2678 785 2694 819
rect 2728 785 2744 819
rect 2678 751 2744 785
rect 2678 717 2694 751
rect 2728 717 2744 751
rect 2678 683 2744 717
rect 2678 649 2694 683
rect 2728 649 2744 683
rect 2678 615 2744 649
rect 2678 581 2694 615
rect 2728 581 2744 615
rect 2678 547 2744 581
rect 2678 513 2694 547
rect 2728 513 2744 547
rect 2678 479 2744 513
rect 2678 445 2694 479
rect 2728 445 2744 479
rect 2678 411 2744 445
rect 2678 377 2694 411
rect 2728 377 2744 411
rect 2678 343 2744 377
rect 2678 309 2694 343
rect 2728 309 2744 343
rect 2678 268 2744 309
rect 2774 1227 2840 1268
rect 2774 1193 2790 1227
rect 2824 1193 2840 1227
rect 2774 1159 2840 1193
rect 2774 1125 2790 1159
rect 2824 1125 2840 1159
rect 2774 1091 2840 1125
rect 2774 1057 2790 1091
rect 2824 1057 2840 1091
rect 2774 1023 2840 1057
rect 2774 989 2790 1023
rect 2824 989 2840 1023
rect 2774 955 2840 989
rect 2774 921 2790 955
rect 2824 921 2840 955
rect 2774 887 2840 921
rect 2774 853 2790 887
rect 2824 853 2840 887
rect 2774 819 2840 853
rect 2774 785 2790 819
rect 2824 785 2840 819
rect 2774 751 2840 785
rect 2774 717 2790 751
rect 2824 717 2840 751
rect 2774 683 2840 717
rect 2774 649 2790 683
rect 2824 649 2840 683
rect 2774 615 2840 649
rect 2774 581 2790 615
rect 2824 581 2840 615
rect 2774 547 2840 581
rect 2774 513 2790 547
rect 2824 513 2840 547
rect 2774 479 2840 513
rect 2774 445 2790 479
rect 2824 445 2840 479
rect 2774 411 2840 445
rect 2774 377 2790 411
rect 2824 377 2840 411
rect 2774 343 2840 377
rect 2774 309 2790 343
rect 2824 309 2840 343
rect 2774 268 2840 309
rect 2870 1227 2936 1268
rect 2870 1193 2886 1227
rect 2920 1193 2936 1227
rect 2870 1159 2936 1193
rect 2870 1125 2886 1159
rect 2920 1125 2936 1159
rect 2870 1091 2936 1125
rect 2870 1057 2886 1091
rect 2920 1057 2936 1091
rect 2870 1023 2936 1057
rect 2870 989 2886 1023
rect 2920 989 2936 1023
rect 2870 955 2936 989
rect 2870 921 2886 955
rect 2920 921 2936 955
rect 2870 887 2936 921
rect 2870 853 2886 887
rect 2920 853 2936 887
rect 2870 819 2936 853
rect 2870 785 2886 819
rect 2920 785 2936 819
rect 2870 751 2936 785
rect 2870 717 2886 751
rect 2920 717 2936 751
rect 2870 683 2936 717
rect 2870 649 2886 683
rect 2920 649 2936 683
rect 2870 615 2936 649
rect 2870 581 2886 615
rect 2920 581 2936 615
rect 2870 547 2936 581
rect 2870 513 2886 547
rect 2920 513 2936 547
rect 2870 479 2936 513
rect 2870 445 2886 479
rect 2920 445 2936 479
rect 2870 411 2936 445
rect 2870 377 2886 411
rect 2920 377 2936 411
rect 2870 343 2936 377
rect 2870 309 2886 343
rect 2920 309 2936 343
rect 2870 268 2936 309
rect 2966 1227 3028 1268
rect 2966 1193 2982 1227
rect 3016 1193 3028 1227
rect 2966 1159 3028 1193
rect 2966 1125 2982 1159
rect 3016 1125 3028 1159
rect 2966 1091 3028 1125
rect 2966 1057 2982 1091
rect 3016 1057 3028 1091
rect 2966 1023 3028 1057
rect 2966 989 2982 1023
rect 3016 989 3028 1023
rect 2966 955 3028 989
rect 2966 921 2982 955
rect 3016 921 3028 955
rect 2966 887 3028 921
rect 2966 853 2982 887
rect 3016 853 3028 887
rect 2966 819 3028 853
rect 2966 785 2982 819
rect 3016 785 3028 819
rect 2966 751 3028 785
rect 2966 717 2982 751
rect 3016 717 3028 751
rect 2966 683 3028 717
rect 2966 649 2982 683
rect 3016 649 3028 683
rect 2966 615 3028 649
rect 2966 581 2982 615
rect 3016 581 3028 615
rect 2966 547 3028 581
rect 2966 513 2982 547
rect 3016 513 3028 547
rect 2966 479 3028 513
rect 2966 445 2982 479
rect 3016 445 3028 479
rect 2966 411 3028 445
rect 2966 377 2982 411
rect 3016 377 3028 411
rect 2966 343 3028 377
rect 2966 309 2982 343
rect 3016 309 3028 343
rect 2966 268 3028 309
rect 3102 1211 3164 1252
rect 3102 1177 3114 1211
rect 3148 1177 3164 1211
rect 3102 1143 3164 1177
rect 3102 1109 3114 1143
rect 3148 1109 3164 1143
rect 3102 1075 3164 1109
rect 3102 1041 3114 1075
rect 3148 1041 3164 1075
rect 3102 1007 3164 1041
rect 3102 973 3114 1007
rect 3148 973 3164 1007
rect 3102 939 3164 973
rect 3102 905 3114 939
rect 3148 905 3164 939
rect 3102 871 3164 905
rect 3102 837 3114 871
rect 3148 837 3164 871
rect 3102 803 3164 837
rect 3102 769 3114 803
rect 3148 769 3164 803
rect 3102 735 3164 769
rect 3102 701 3114 735
rect 3148 701 3164 735
rect 3102 667 3164 701
rect 3102 633 3114 667
rect 3148 633 3164 667
rect 3102 599 3164 633
rect 3102 565 3114 599
rect 3148 565 3164 599
rect 3102 531 3164 565
rect 3102 497 3114 531
rect 3148 497 3164 531
rect 3102 463 3164 497
rect 3102 429 3114 463
rect 3148 429 3164 463
rect 3102 395 3164 429
rect 3102 361 3114 395
rect 3148 361 3164 395
rect 3102 327 3164 361
rect 3102 293 3114 327
rect 3148 293 3164 327
rect -914 209 -856 243
rect -914 175 -902 209
rect -868 175 -856 209
rect -914 141 -856 175
rect 3102 252 3164 293
rect 3194 1211 3260 1252
rect 3194 1177 3210 1211
rect 3244 1177 3260 1211
rect 3194 1143 3260 1177
rect 3194 1109 3210 1143
rect 3244 1109 3260 1143
rect 3194 1075 3260 1109
rect 3194 1041 3210 1075
rect 3244 1041 3260 1075
rect 3194 1007 3260 1041
rect 3194 973 3210 1007
rect 3244 973 3260 1007
rect 3194 939 3260 973
rect 3194 905 3210 939
rect 3244 905 3260 939
rect 3194 871 3260 905
rect 3194 837 3210 871
rect 3244 837 3260 871
rect 3194 803 3260 837
rect 3194 769 3210 803
rect 3244 769 3260 803
rect 3194 735 3260 769
rect 3194 701 3210 735
rect 3244 701 3260 735
rect 3194 667 3260 701
rect 3194 633 3210 667
rect 3244 633 3260 667
rect 3194 599 3260 633
rect 3194 565 3210 599
rect 3244 565 3260 599
rect 3194 531 3260 565
rect 3194 497 3210 531
rect 3244 497 3260 531
rect 3194 463 3260 497
rect 3194 429 3210 463
rect 3244 429 3260 463
rect 3194 395 3260 429
rect 3194 361 3210 395
rect 3244 361 3260 395
rect 3194 327 3260 361
rect 3194 293 3210 327
rect 3244 293 3260 327
rect 3194 252 3260 293
rect 3290 1211 3356 1252
rect 3290 1177 3306 1211
rect 3340 1177 3356 1211
rect 3290 1143 3356 1177
rect 3290 1109 3306 1143
rect 3340 1109 3356 1143
rect 3290 1075 3356 1109
rect 3290 1041 3306 1075
rect 3340 1041 3356 1075
rect 3290 1007 3356 1041
rect 3290 973 3306 1007
rect 3340 973 3356 1007
rect 3290 939 3356 973
rect 3290 905 3306 939
rect 3340 905 3356 939
rect 3290 871 3356 905
rect 3290 837 3306 871
rect 3340 837 3356 871
rect 3290 803 3356 837
rect 3290 769 3306 803
rect 3340 769 3356 803
rect 3290 735 3356 769
rect 3290 701 3306 735
rect 3340 701 3356 735
rect 3290 667 3356 701
rect 3290 633 3306 667
rect 3340 633 3356 667
rect 3290 599 3356 633
rect 3290 565 3306 599
rect 3340 565 3356 599
rect 3290 531 3356 565
rect 3290 497 3306 531
rect 3340 497 3356 531
rect 3290 463 3356 497
rect 3290 429 3306 463
rect 3340 429 3356 463
rect 3290 395 3356 429
rect 3290 361 3306 395
rect 3340 361 3356 395
rect 3290 327 3356 361
rect 3290 293 3306 327
rect 3340 293 3356 327
rect 3290 252 3356 293
rect 3386 1211 3452 1252
rect 3386 1177 3402 1211
rect 3436 1177 3452 1211
rect 3386 1143 3452 1177
rect 3386 1109 3402 1143
rect 3436 1109 3452 1143
rect 3386 1075 3452 1109
rect 3386 1041 3402 1075
rect 3436 1041 3452 1075
rect 3386 1007 3452 1041
rect 3386 973 3402 1007
rect 3436 973 3452 1007
rect 3386 939 3452 973
rect 3386 905 3402 939
rect 3436 905 3452 939
rect 3386 871 3452 905
rect 3386 837 3402 871
rect 3436 837 3452 871
rect 3386 803 3452 837
rect 3386 769 3402 803
rect 3436 769 3452 803
rect 3386 735 3452 769
rect 3386 701 3402 735
rect 3436 701 3452 735
rect 3386 667 3452 701
rect 3386 633 3402 667
rect 3436 633 3452 667
rect 3386 599 3452 633
rect 3386 565 3402 599
rect 3436 565 3452 599
rect 3386 531 3452 565
rect 3386 497 3402 531
rect 3436 497 3452 531
rect 3386 463 3452 497
rect 3386 429 3402 463
rect 3436 429 3452 463
rect 3386 395 3452 429
rect 3386 361 3402 395
rect 3436 361 3452 395
rect 3386 327 3452 361
rect 3386 293 3402 327
rect 3436 293 3452 327
rect 3386 252 3452 293
rect 3482 1211 3548 1252
rect 3482 1177 3498 1211
rect 3532 1177 3548 1211
rect 3482 1143 3548 1177
rect 3482 1109 3498 1143
rect 3532 1109 3548 1143
rect 3482 1075 3548 1109
rect 3482 1041 3498 1075
rect 3532 1041 3548 1075
rect 3482 1007 3548 1041
rect 3482 973 3498 1007
rect 3532 973 3548 1007
rect 3482 939 3548 973
rect 3482 905 3498 939
rect 3532 905 3548 939
rect 3482 871 3548 905
rect 3482 837 3498 871
rect 3532 837 3548 871
rect 3482 803 3548 837
rect 3482 769 3498 803
rect 3532 769 3548 803
rect 3482 735 3548 769
rect 3482 701 3498 735
rect 3532 701 3548 735
rect 3482 667 3548 701
rect 3482 633 3498 667
rect 3532 633 3548 667
rect 3482 599 3548 633
rect 3482 565 3498 599
rect 3532 565 3548 599
rect 3482 531 3548 565
rect 3482 497 3498 531
rect 3532 497 3548 531
rect 3482 463 3548 497
rect 3482 429 3498 463
rect 3532 429 3548 463
rect 3482 395 3548 429
rect 3482 361 3498 395
rect 3532 361 3548 395
rect 3482 327 3548 361
rect 3482 293 3498 327
rect 3532 293 3548 327
rect 3482 252 3548 293
rect 3578 1211 3644 1252
rect 3578 1177 3594 1211
rect 3628 1177 3644 1211
rect 3578 1143 3644 1177
rect 3578 1109 3594 1143
rect 3628 1109 3644 1143
rect 3578 1075 3644 1109
rect 3578 1041 3594 1075
rect 3628 1041 3644 1075
rect 3578 1007 3644 1041
rect 3578 973 3594 1007
rect 3628 973 3644 1007
rect 3578 939 3644 973
rect 3578 905 3594 939
rect 3628 905 3644 939
rect 3578 871 3644 905
rect 3578 837 3594 871
rect 3628 837 3644 871
rect 3578 803 3644 837
rect 3578 769 3594 803
rect 3628 769 3644 803
rect 3578 735 3644 769
rect 3578 701 3594 735
rect 3628 701 3644 735
rect 3578 667 3644 701
rect 3578 633 3594 667
rect 3628 633 3644 667
rect 3578 599 3644 633
rect 3578 565 3594 599
rect 3628 565 3644 599
rect 3578 531 3644 565
rect 3578 497 3594 531
rect 3628 497 3644 531
rect 3578 463 3644 497
rect 3578 429 3594 463
rect 3628 429 3644 463
rect 3578 395 3644 429
rect 3578 361 3594 395
rect 3628 361 3644 395
rect 3578 327 3644 361
rect 3578 293 3594 327
rect 3628 293 3644 327
rect 3578 252 3644 293
rect 3674 1211 3740 1252
rect 3674 1177 3690 1211
rect 3724 1177 3740 1211
rect 3674 1143 3740 1177
rect 3674 1109 3690 1143
rect 3724 1109 3740 1143
rect 3674 1075 3740 1109
rect 3674 1041 3690 1075
rect 3724 1041 3740 1075
rect 3674 1007 3740 1041
rect 3674 973 3690 1007
rect 3724 973 3740 1007
rect 3674 939 3740 973
rect 3674 905 3690 939
rect 3724 905 3740 939
rect 3674 871 3740 905
rect 3674 837 3690 871
rect 3724 837 3740 871
rect 3674 803 3740 837
rect 3674 769 3690 803
rect 3724 769 3740 803
rect 3674 735 3740 769
rect 3674 701 3690 735
rect 3724 701 3740 735
rect 3674 667 3740 701
rect 3674 633 3690 667
rect 3724 633 3740 667
rect 3674 599 3740 633
rect 3674 565 3690 599
rect 3724 565 3740 599
rect 3674 531 3740 565
rect 3674 497 3690 531
rect 3724 497 3740 531
rect 3674 463 3740 497
rect 3674 429 3690 463
rect 3724 429 3740 463
rect 3674 395 3740 429
rect 3674 361 3690 395
rect 3724 361 3740 395
rect 3674 327 3740 361
rect 3674 293 3690 327
rect 3724 293 3740 327
rect 3674 252 3740 293
rect 3770 1211 3836 1252
rect 3770 1177 3786 1211
rect 3820 1177 3836 1211
rect 3770 1143 3836 1177
rect 3770 1109 3786 1143
rect 3820 1109 3836 1143
rect 3770 1075 3836 1109
rect 3770 1041 3786 1075
rect 3820 1041 3836 1075
rect 3770 1007 3836 1041
rect 3770 973 3786 1007
rect 3820 973 3836 1007
rect 3770 939 3836 973
rect 3770 905 3786 939
rect 3820 905 3836 939
rect 3770 871 3836 905
rect 3770 837 3786 871
rect 3820 837 3836 871
rect 3770 803 3836 837
rect 3770 769 3786 803
rect 3820 769 3836 803
rect 3770 735 3836 769
rect 3770 701 3786 735
rect 3820 701 3836 735
rect 3770 667 3836 701
rect 3770 633 3786 667
rect 3820 633 3836 667
rect 3770 599 3836 633
rect 3770 565 3786 599
rect 3820 565 3836 599
rect 3770 531 3836 565
rect 3770 497 3786 531
rect 3820 497 3836 531
rect 3770 463 3836 497
rect 3770 429 3786 463
rect 3820 429 3836 463
rect 3770 395 3836 429
rect 3770 361 3786 395
rect 3820 361 3836 395
rect 3770 327 3836 361
rect 3770 293 3786 327
rect 3820 293 3836 327
rect 3770 252 3836 293
rect 3866 1211 3932 1252
rect 3866 1177 3882 1211
rect 3916 1177 3932 1211
rect 3866 1143 3932 1177
rect 3866 1109 3882 1143
rect 3916 1109 3932 1143
rect 3866 1075 3932 1109
rect 3866 1041 3882 1075
rect 3916 1041 3932 1075
rect 3866 1007 3932 1041
rect 3866 973 3882 1007
rect 3916 973 3932 1007
rect 3866 939 3932 973
rect 3866 905 3882 939
rect 3916 905 3932 939
rect 3866 871 3932 905
rect 3866 837 3882 871
rect 3916 837 3932 871
rect 3866 803 3932 837
rect 3866 769 3882 803
rect 3916 769 3932 803
rect 3866 735 3932 769
rect 3866 701 3882 735
rect 3916 701 3932 735
rect 3866 667 3932 701
rect 3866 633 3882 667
rect 3916 633 3932 667
rect 3866 599 3932 633
rect 3866 565 3882 599
rect 3916 565 3932 599
rect 3866 531 3932 565
rect 3866 497 3882 531
rect 3916 497 3932 531
rect 3866 463 3932 497
rect 3866 429 3882 463
rect 3916 429 3932 463
rect 3866 395 3932 429
rect 3866 361 3882 395
rect 3916 361 3932 395
rect 3866 327 3932 361
rect 3866 293 3882 327
rect 3916 293 3932 327
rect 3866 252 3932 293
rect 3962 1211 4028 1252
rect 3962 1177 3978 1211
rect 4012 1177 4028 1211
rect 3962 1143 4028 1177
rect 3962 1109 3978 1143
rect 4012 1109 4028 1143
rect 3962 1075 4028 1109
rect 3962 1041 3978 1075
rect 4012 1041 4028 1075
rect 3962 1007 4028 1041
rect 3962 973 3978 1007
rect 4012 973 4028 1007
rect 3962 939 4028 973
rect 3962 905 3978 939
rect 4012 905 4028 939
rect 3962 871 4028 905
rect 3962 837 3978 871
rect 4012 837 4028 871
rect 3962 803 4028 837
rect 3962 769 3978 803
rect 4012 769 4028 803
rect 3962 735 4028 769
rect 3962 701 3978 735
rect 4012 701 4028 735
rect 3962 667 4028 701
rect 3962 633 3978 667
rect 4012 633 4028 667
rect 3962 599 4028 633
rect 3962 565 3978 599
rect 4012 565 4028 599
rect 3962 531 4028 565
rect 3962 497 3978 531
rect 4012 497 4028 531
rect 3962 463 4028 497
rect 3962 429 3978 463
rect 4012 429 4028 463
rect 3962 395 4028 429
rect 3962 361 3978 395
rect 4012 361 4028 395
rect 3962 327 4028 361
rect 3962 293 3978 327
rect 4012 293 4028 327
rect 3962 252 4028 293
rect 4058 1211 4124 1252
rect 4058 1177 4074 1211
rect 4108 1177 4124 1211
rect 4058 1143 4124 1177
rect 4058 1109 4074 1143
rect 4108 1109 4124 1143
rect 4058 1075 4124 1109
rect 4058 1041 4074 1075
rect 4108 1041 4124 1075
rect 4058 1007 4124 1041
rect 4058 973 4074 1007
rect 4108 973 4124 1007
rect 4058 939 4124 973
rect 4058 905 4074 939
rect 4108 905 4124 939
rect 4058 871 4124 905
rect 4058 837 4074 871
rect 4108 837 4124 871
rect 4058 803 4124 837
rect 4058 769 4074 803
rect 4108 769 4124 803
rect 4058 735 4124 769
rect 4058 701 4074 735
rect 4108 701 4124 735
rect 4058 667 4124 701
rect 4058 633 4074 667
rect 4108 633 4124 667
rect 4058 599 4124 633
rect 4058 565 4074 599
rect 4108 565 4124 599
rect 4058 531 4124 565
rect 4058 497 4074 531
rect 4108 497 4124 531
rect 4058 463 4124 497
rect 4058 429 4074 463
rect 4108 429 4124 463
rect 4058 395 4124 429
rect 4058 361 4074 395
rect 4108 361 4124 395
rect 4058 327 4124 361
rect 4058 293 4074 327
rect 4108 293 4124 327
rect 4058 252 4124 293
rect 4154 1211 4220 1252
rect 4154 1177 4170 1211
rect 4204 1177 4220 1211
rect 4154 1143 4220 1177
rect 4154 1109 4170 1143
rect 4204 1109 4220 1143
rect 4154 1075 4220 1109
rect 4154 1041 4170 1075
rect 4204 1041 4220 1075
rect 4154 1007 4220 1041
rect 4154 973 4170 1007
rect 4204 973 4220 1007
rect 4154 939 4220 973
rect 4154 905 4170 939
rect 4204 905 4220 939
rect 4154 871 4220 905
rect 4154 837 4170 871
rect 4204 837 4220 871
rect 4154 803 4220 837
rect 4154 769 4170 803
rect 4204 769 4220 803
rect 4154 735 4220 769
rect 4154 701 4170 735
rect 4204 701 4220 735
rect 4154 667 4220 701
rect 4154 633 4170 667
rect 4204 633 4220 667
rect 4154 599 4220 633
rect 4154 565 4170 599
rect 4204 565 4220 599
rect 4154 531 4220 565
rect 4154 497 4170 531
rect 4204 497 4220 531
rect 4154 463 4220 497
rect 4154 429 4170 463
rect 4204 429 4220 463
rect 4154 395 4220 429
rect 4154 361 4170 395
rect 4204 361 4220 395
rect 4154 327 4220 361
rect 4154 293 4170 327
rect 4204 293 4220 327
rect 4154 252 4220 293
rect 4250 1211 4312 1252
rect 4250 1177 4266 1211
rect 4300 1177 4312 1211
rect 4250 1143 4312 1177
rect 4250 1109 4266 1143
rect 4300 1109 4312 1143
rect 4250 1075 4312 1109
rect 4250 1041 4266 1075
rect 4300 1041 4312 1075
rect 4250 1007 4312 1041
rect 4250 973 4266 1007
rect 4300 973 4312 1007
rect 4250 939 4312 973
rect 4250 905 4266 939
rect 4300 905 4312 939
rect 4250 871 4312 905
rect 4250 837 4266 871
rect 4300 837 4312 871
rect 4250 803 4312 837
rect 4250 769 4266 803
rect 4300 769 4312 803
rect 4250 735 4312 769
rect 4250 701 4266 735
rect 4300 701 4312 735
rect 4250 667 4312 701
rect 4250 633 4266 667
rect 4300 633 4312 667
rect 4250 599 4312 633
rect 4250 565 4266 599
rect 4300 565 4312 599
rect 4250 531 4312 565
rect 4250 497 4266 531
rect 4300 497 4312 531
rect 4250 463 4312 497
rect 4250 429 4266 463
rect 4300 429 4312 463
rect 4250 395 4312 429
rect 4250 361 4266 395
rect 4300 361 4312 395
rect 4250 327 4312 361
rect 4250 293 4266 327
rect 4300 293 4312 327
rect 4250 252 4312 293
rect 4870 1211 4932 1252
rect 4870 1177 4882 1211
rect 4916 1177 4932 1211
rect 4870 1143 4932 1177
rect 4870 1109 4882 1143
rect 4916 1109 4932 1143
rect 4870 1075 4932 1109
rect 4870 1041 4882 1075
rect 4916 1041 4932 1075
rect 4870 1007 4932 1041
rect 4870 973 4882 1007
rect 4916 973 4932 1007
rect 4870 939 4932 973
rect 4870 905 4882 939
rect 4916 905 4932 939
rect 4870 871 4932 905
rect 4870 837 4882 871
rect 4916 837 4932 871
rect 4870 803 4932 837
rect 4870 769 4882 803
rect 4916 769 4932 803
rect 4870 735 4932 769
rect 4870 701 4882 735
rect 4916 701 4932 735
rect 4870 667 4932 701
rect 4870 633 4882 667
rect 4916 633 4932 667
rect 4870 599 4932 633
rect 4870 565 4882 599
rect 4916 565 4932 599
rect 4870 531 4932 565
rect 4870 497 4882 531
rect 4916 497 4932 531
rect 4870 463 4932 497
rect 4870 429 4882 463
rect 4916 429 4932 463
rect 4870 395 4932 429
rect 4870 361 4882 395
rect 4916 361 4932 395
rect 4870 327 4932 361
rect 4870 293 4882 327
rect 4916 293 4932 327
rect 4870 252 4932 293
rect 4962 1211 5028 1252
rect 4962 1177 4978 1211
rect 5012 1177 5028 1211
rect 4962 1143 5028 1177
rect 4962 1109 4978 1143
rect 5012 1109 5028 1143
rect 4962 1075 5028 1109
rect 4962 1041 4978 1075
rect 5012 1041 5028 1075
rect 4962 1007 5028 1041
rect 4962 973 4978 1007
rect 5012 973 5028 1007
rect 4962 939 5028 973
rect 4962 905 4978 939
rect 5012 905 5028 939
rect 4962 871 5028 905
rect 4962 837 4978 871
rect 5012 837 5028 871
rect 4962 803 5028 837
rect 4962 769 4978 803
rect 5012 769 5028 803
rect 4962 735 5028 769
rect 4962 701 4978 735
rect 5012 701 5028 735
rect 4962 667 5028 701
rect 4962 633 4978 667
rect 5012 633 5028 667
rect 4962 599 5028 633
rect 4962 565 4978 599
rect 5012 565 5028 599
rect 4962 531 5028 565
rect 4962 497 4978 531
rect 5012 497 5028 531
rect 4962 463 5028 497
rect 4962 429 4978 463
rect 5012 429 5028 463
rect 4962 395 5028 429
rect 4962 361 4978 395
rect 5012 361 5028 395
rect 4962 327 5028 361
rect 4962 293 4978 327
rect 5012 293 5028 327
rect 4962 252 5028 293
rect 5058 1211 5124 1252
rect 5058 1177 5074 1211
rect 5108 1177 5124 1211
rect 5058 1143 5124 1177
rect 5058 1109 5074 1143
rect 5108 1109 5124 1143
rect 5058 1075 5124 1109
rect 5058 1041 5074 1075
rect 5108 1041 5124 1075
rect 5058 1007 5124 1041
rect 5058 973 5074 1007
rect 5108 973 5124 1007
rect 5058 939 5124 973
rect 5058 905 5074 939
rect 5108 905 5124 939
rect 5058 871 5124 905
rect 5058 837 5074 871
rect 5108 837 5124 871
rect 5058 803 5124 837
rect 5058 769 5074 803
rect 5108 769 5124 803
rect 5058 735 5124 769
rect 5058 701 5074 735
rect 5108 701 5124 735
rect 5058 667 5124 701
rect 5058 633 5074 667
rect 5108 633 5124 667
rect 5058 599 5124 633
rect 5058 565 5074 599
rect 5108 565 5124 599
rect 5058 531 5124 565
rect 5058 497 5074 531
rect 5108 497 5124 531
rect 5058 463 5124 497
rect 5058 429 5074 463
rect 5108 429 5124 463
rect 5058 395 5124 429
rect 5058 361 5074 395
rect 5108 361 5124 395
rect 5058 327 5124 361
rect 5058 293 5074 327
rect 5108 293 5124 327
rect 5058 252 5124 293
rect 5154 1211 5220 1252
rect 5154 1177 5170 1211
rect 5204 1177 5220 1211
rect 5154 1143 5220 1177
rect 5154 1109 5170 1143
rect 5204 1109 5220 1143
rect 5154 1075 5220 1109
rect 5154 1041 5170 1075
rect 5204 1041 5220 1075
rect 5154 1007 5220 1041
rect 5154 973 5170 1007
rect 5204 973 5220 1007
rect 5154 939 5220 973
rect 5154 905 5170 939
rect 5204 905 5220 939
rect 5154 871 5220 905
rect 5154 837 5170 871
rect 5204 837 5220 871
rect 5154 803 5220 837
rect 5154 769 5170 803
rect 5204 769 5220 803
rect 5154 735 5220 769
rect 5154 701 5170 735
rect 5204 701 5220 735
rect 5154 667 5220 701
rect 5154 633 5170 667
rect 5204 633 5220 667
rect 5154 599 5220 633
rect 5154 565 5170 599
rect 5204 565 5220 599
rect 5154 531 5220 565
rect 5154 497 5170 531
rect 5204 497 5220 531
rect 5154 463 5220 497
rect 5154 429 5170 463
rect 5204 429 5220 463
rect 5154 395 5220 429
rect 5154 361 5170 395
rect 5204 361 5220 395
rect 5154 327 5220 361
rect 5154 293 5170 327
rect 5204 293 5220 327
rect 5154 252 5220 293
rect 5250 1211 5316 1252
rect 5250 1177 5266 1211
rect 5300 1177 5316 1211
rect 5250 1143 5316 1177
rect 5250 1109 5266 1143
rect 5300 1109 5316 1143
rect 5250 1075 5316 1109
rect 5250 1041 5266 1075
rect 5300 1041 5316 1075
rect 5250 1007 5316 1041
rect 5250 973 5266 1007
rect 5300 973 5316 1007
rect 5250 939 5316 973
rect 5250 905 5266 939
rect 5300 905 5316 939
rect 5250 871 5316 905
rect 5250 837 5266 871
rect 5300 837 5316 871
rect 5250 803 5316 837
rect 5250 769 5266 803
rect 5300 769 5316 803
rect 5250 735 5316 769
rect 5250 701 5266 735
rect 5300 701 5316 735
rect 5250 667 5316 701
rect 5250 633 5266 667
rect 5300 633 5316 667
rect 5250 599 5316 633
rect 5250 565 5266 599
rect 5300 565 5316 599
rect 5250 531 5316 565
rect 5250 497 5266 531
rect 5300 497 5316 531
rect 5250 463 5316 497
rect 5250 429 5266 463
rect 5300 429 5316 463
rect 5250 395 5316 429
rect 5250 361 5266 395
rect 5300 361 5316 395
rect 5250 327 5316 361
rect 5250 293 5266 327
rect 5300 293 5316 327
rect 5250 252 5316 293
rect 5346 1211 5412 1252
rect 5346 1177 5362 1211
rect 5396 1177 5412 1211
rect 5346 1143 5412 1177
rect 5346 1109 5362 1143
rect 5396 1109 5412 1143
rect 5346 1075 5412 1109
rect 5346 1041 5362 1075
rect 5396 1041 5412 1075
rect 5346 1007 5412 1041
rect 5346 973 5362 1007
rect 5396 973 5412 1007
rect 5346 939 5412 973
rect 5346 905 5362 939
rect 5396 905 5412 939
rect 5346 871 5412 905
rect 5346 837 5362 871
rect 5396 837 5412 871
rect 5346 803 5412 837
rect 5346 769 5362 803
rect 5396 769 5412 803
rect 5346 735 5412 769
rect 5346 701 5362 735
rect 5396 701 5412 735
rect 5346 667 5412 701
rect 5346 633 5362 667
rect 5396 633 5412 667
rect 5346 599 5412 633
rect 5346 565 5362 599
rect 5396 565 5412 599
rect 5346 531 5412 565
rect 5346 497 5362 531
rect 5396 497 5412 531
rect 5346 463 5412 497
rect 5346 429 5362 463
rect 5396 429 5412 463
rect 5346 395 5412 429
rect 5346 361 5362 395
rect 5396 361 5412 395
rect 5346 327 5412 361
rect 5346 293 5362 327
rect 5396 293 5412 327
rect 5346 252 5412 293
rect 5442 1211 5508 1252
rect 5442 1177 5458 1211
rect 5492 1177 5508 1211
rect 5442 1143 5508 1177
rect 5442 1109 5458 1143
rect 5492 1109 5508 1143
rect 5442 1075 5508 1109
rect 5442 1041 5458 1075
rect 5492 1041 5508 1075
rect 5442 1007 5508 1041
rect 5442 973 5458 1007
rect 5492 973 5508 1007
rect 5442 939 5508 973
rect 5442 905 5458 939
rect 5492 905 5508 939
rect 5442 871 5508 905
rect 5442 837 5458 871
rect 5492 837 5508 871
rect 5442 803 5508 837
rect 5442 769 5458 803
rect 5492 769 5508 803
rect 5442 735 5508 769
rect 5442 701 5458 735
rect 5492 701 5508 735
rect 5442 667 5508 701
rect 5442 633 5458 667
rect 5492 633 5508 667
rect 5442 599 5508 633
rect 5442 565 5458 599
rect 5492 565 5508 599
rect 5442 531 5508 565
rect 5442 497 5458 531
rect 5492 497 5508 531
rect 5442 463 5508 497
rect 5442 429 5458 463
rect 5492 429 5508 463
rect 5442 395 5508 429
rect 5442 361 5458 395
rect 5492 361 5508 395
rect 5442 327 5508 361
rect 5442 293 5458 327
rect 5492 293 5508 327
rect 5442 252 5508 293
rect 5538 1211 5604 1252
rect 5538 1177 5554 1211
rect 5588 1177 5604 1211
rect 5538 1143 5604 1177
rect 5538 1109 5554 1143
rect 5588 1109 5604 1143
rect 5538 1075 5604 1109
rect 5538 1041 5554 1075
rect 5588 1041 5604 1075
rect 5538 1007 5604 1041
rect 5538 973 5554 1007
rect 5588 973 5604 1007
rect 5538 939 5604 973
rect 5538 905 5554 939
rect 5588 905 5604 939
rect 5538 871 5604 905
rect 5538 837 5554 871
rect 5588 837 5604 871
rect 5538 803 5604 837
rect 5538 769 5554 803
rect 5588 769 5604 803
rect 5538 735 5604 769
rect 5538 701 5554 735
rect 5588 701 5604 735
rect 5538 667 5604 701
rect 5538 633 5554 667
rect 5588 633 5604 667
rect 5538 599 5604 633
rect 5538 565 5554 599
rect 5588 565 5604 599
rect 5538 531 5604 565
rect 5538 497 5554 531
rect 5588 497 5604 531
rect 5538 463 5604 497
rect 5538 429 5554 463
rect 5588 429 5604 463
rect 5538 395 5604 429
rect 5538 361 5554 395
rect 5588 361 5604 395
rect 5538 327 5604 361
rect 5538 293 5554 327
rect 5588 293 5604 327
rect 5538 252 5604 293
rect 5634 1211 5700 1252
rect 5634 1177 5650 1211
rect 5684 1177 5700 1211
rect 5634 1143 5700 1177
rect 5634 1109 5650 1143
rect 5684 1109 5700 1143
rect 5634 1075 5700 1109
rect 5634 1041 5650 1075
rect 5684 1041 5700 1075
rect 5634 1007 5700 1041
rect 5634 973 5650 1007
rect 5684 973 5700 1007
rect 5634 939 5700 973
rect 5634 905 5650 939
rect 5684 905 5700 939
rect 5634 871 5700 905
rect 5634 837 5650 871
rect 5684 837 5700 871
rect 5634 803 5700 837
rect 5634 769 5650 803
rect 5684 769 5700 803
rect 5634 735 5700 769
rect 5634 701 5650 735
rect 5684 701 5700 735
rect 5634 667 5700 701
rect 5634 633 5650 667
rect 5684 633 5700 667
rect 5634 599 5700 633
rect 5634 565 5650 599
rect 5684 565 5700 599
rect 5634 531 5700 565
rect 5634 497 5650 531
rect 5684 497 5700 531
rect 5634 463 5700 497
rect 5634 429 5650 463
rect 5684 429 5700 463
rect 5634 395 5700 429
rect 5634 361 5650 395
rect 5684 361 5700 395
rect 5634 327 5700 361
rect 5634 293 5650 327
rect 5684 293 5700 327
rect 5634 252 5700 293
rect 5730 1211 5796 1252
rect 5730 1177 5746 1211
rect 5780 1177 5796 1211
rect 5730 1143 5796 1177
rect 5730 1109 5746 1143
rect 5780 1109 5796 1143
rect 5730 1075 5796 1109
rect 5730 1041 5746 1075
rect 5780 1041 5796 1075
rect 5730 1007 5796 1041
rect 5730 973 5746 1007
rect 5780 973 5796 1007
rect 5730 939 5796 973
rect 5730 905 5746 939
rect 5780 905 5796 939
rect 5730 871 5796 905
rect 5730 837 5746 871
rect 5780 837 5796 871
rect 5730 803 5796 837
rect 5730 769 5746 803
rect 5780 769 5796 803
rect 5730 735 5796 769
rect 5730 701 5746 735
rect 5780 701 5796 735
rect 5730 667 5796 701
rect 5730 633 5746 667
rect 5780 633 5796 667
rect 5730 599 5796 633
rect 5730 565 5746 599
rect 5780 565 5796 599
rect 5730 531 5796 565
rect 5730 497 5746 531
rect 5780 497 5796 531
rect 5730 463 5796 497
rect 5730 429 5746 463
rect 5780 429 5796 463
rect 5730 395 5796 429
rect 5730 361 5746 395
rect 5780 361 5796 395
rect 5730 327 5796 361
rect 5730 293 5746 327
rect 5780 293 5796 327
rect 5730 252 5796 293
rect 5826 1211 5892 1252
rect 5826 1177 5842 1211
rect 5876 1177 5892 1211
rect 5826 1143 5892 1177
rect 5826 1109 5842 1143
rect 5876 1109 5892 1143
rect 5826 1075 5892 1109
rect 5826 1041 5842 1075
rect 5876 1041 5892 1075
rect 5826 1007 5892 1041
rect 5826 973 5842 1007
rect 5876 973 5892 1007
rect 5826 939 5892 973
rect 5826 905 5842 939
rect 5876 905 5892 939
rect 5826 871 5892 905
rect 5826 837 5842 871
rect 5876 837 5892 871
rect 5826 803 5892 837
rect 5826 769 5842 803
rect 5876 769 5892 803
rect 5826 735 5892 769
rect 5826 701 5842 735
rect 5876 701 5892 735
rect 5826 667 5892 701
rect 5826 633 5842 667
rect 5876 633 5892 667
rect 5826 599 5892 633
rect 5826 565 5842 599
rect 5876 565 5892 599
rect 5826 531 5892 565
rect 5826 497 5842 531
rect 5876 497 5892 531
rect 5826 463 5892 497
rect 5826 429 5842 463
rect 5876 429 5892 463
rect 5826 395 5892 429
rect 5826 361 5842 395
rect 5876 361 5892 395
rect 5826 327 5892 361
rect 5826 293 5842 327
rect 5876 293 5892 327
rect 5826 252 5892 293
rect 5922 1211 5984 1252
rect 5922 1177 5938 1211
rect 5972 1177 5984 1211
rect 5922 1143 5984 1177
rect 5922 1109 5938 1143
rect 5972 1109 5984 1143
rect 5922 1075 5984 1109
rect 5922 1041 5938 1075
rect 5972 1041 5984 1075
rect 5922 1007 5984 1041
rect 5922 973 5938 1007
rect 5972 973 5984 1007
rect 5922 939 5984 973
rect 5922 905 5938 939
rect 5972 905 5984 939
rect 5922 871 5984 905
rect 5922 837 5938 871
rect 5972 837 5984 871
rect 5922 803 5984 837
rect 5922 769 5938 803
rect 5972 769 5984 803
rect 5922 735 5984 769
rect 5922 701 5938 735
rect 5972 701 5984 735
rect 5922 667 5984 701
rect 5922 633 5938 667
rect 5972 633 5984 667
rect 5922 599 5984 633
rect 5922 565 5938 599
rect 5972 565 5984 599
rect 5922 531 5984 565
rect 5922 497 5938 531
rect 5972 497 5984 531
rect 5922 463 5984 497
rect 5922 429 5938 463
rect 5972 429 5984 463
rect 5922 395 5984 429
rect 5922 361 5938 395
rect 5972 361 5984 395
rect 5922 327 5984 361
rect 5922 293 5938 327
rect 5972 293 5984 327
rect 5922 252 5984 293
rect 6132 1211 6194 1252
rect 6132 1177 6144 1211
rect 6178 1177 6194 1211
rect 6132 1143 6194 1177
rect 6132 1109 6144 1143
rect 6178 1109 6194 1143
rect 6132 1075 6194 1109
rect 6132 1041 6144 1075
rect 6178 1041 6194 1075
rect 6132 1007 6194 1041
rect 6132 973 6144 1007
rect 6178 973 6194 1007
rect 6132 939 6194 973
rect 6132 905 6144 939
rect 6178 905 6194 939
rect 6132 871 6194 905
rect 6132 837 6144 871
rect 6178 837 6194 871
rect 6132 803 6194 837
rect 6132 769 6144 803
rect 6178 769 6194 803
rect 6132 735 6194 769
rect 6132 701 6144 735
rect 6178 701 6194 735
rect 6132 667 6194 701
rect 6132 633 6144 667
rect 6178 633 6194 667
rect 6132 599 6194 633
rect 6132 565 6144 599
rect 6178 565 6194 599
rect 6132 531 6194 565
rect 6132 497 6144 531
rect 6178 497 6194 531
rect 6132 463 6194 497
rect 6132 429 6144 463
rect 6178 429 6194 463
rect 6132 395 6194 429
rect 6132 361 6144 395
rect 6178 361 6194 395
rect 6132 327 6194 361
rect 6132 293 6144 327
rect 6178 293 6194 327
rect 6132 252 6194 293
rect 6224 1211 6290 1252
rect 6224 1177 6240 1211
rect 6274 1177 6290 1211
rect 6224 1143 6290 1177
rect 6224 1109 6240 1143
rect 6274 1109 6290 1143
rect 6224 1075 6290 1109
rect 6224 1041 6240 1075
rect 6274 1041 6290 1075
rect 6224 1007 6290 1041
rect 6224 973 6240 1007
rect 6274 973 6290 1007
rect 6224 939 6290 973
rect 6224 905 6240 939
rect 6274 905 6290 939
rect 6224 871 6290 905
rect 6224 837 6240 871
rect 6274 837 6290 871
rect 6224 803 6290 837
rect 6224 769 6240 803
rect 6274 769 6290 803
rect 6224 735 6290 769
rect 6224 701 6240 735
rect 6274 701 6290 735
rect 6224 667 6290 701
rect 6224 633 6240 667
rect 6274 633 6290 667
rect 6224 599 6290 633
rect 6224 565 6240 599
rect 6274 565 6290 599
rect 6224 531 6290 565
rect 6224 497 6240 531
rect 6274 497 6290 531
rect 6224 463 6290 497
rect 6224 429 6240 463
rect 6274 429 6290 463
rect 6224 395 6290 429
rect 6224 361 6240 395
rect 6274 361 6290 395
rect 6224 327 6290 361
rect 6224 293 6240 327
rect 6274 293 6290 327
rect 6224 252 6290 293
rect 6320 1211 6386 1252
rect 6320 1177 6336 1211
rect 6370 1177 6386 1211
rect 6320 1143 6386 1177
rect 6320 1109 6336 1143
rect 6370 1109 6386 1143
rect 6320 1075 6386 1109
rect 6320 1041 6336 1075
rect 6370 1041 6386 1075
rect 6320 1007 6386 1041
rect 6320 973 6336 1007
rect 6370 973 6386 1007
rect 6320 939 6386 973
rect 6320 905 6336 939
rect 6370 905 6386 939
rect 6320 871 6386 905
rect 6320 837 6336 871
rect 6370 837 6386 871
rect 6320 803 6386 837
rect 6320 769 6336 803
rect 6370 769 6386 803
rect 6320 735 6386 769
rect 6320 701 6336 735
rect 6370 701 6386 735
rect 6320 667 6386 701
rect 6320 633 6336 667
rect 6370 633 6386 667
rect 6320 599 6386 633
rect 6320 565 6336 599
rect 6370 565 6386 599
rect 6320 531 6386 565
rect 6320 497 6336 531
rect 6370 497 6386 531
rect 6320 463 6386 497
rect 6320 429 6336 463
rect 6370 429 6386 463
rect 6320 395 6386 429
rect 6320 361 6336 395
rect 6370 361 6386 395
rect 6320 327 6386 361
rect 6320 293 6336 327
rect 6370 293 6386 327
rect 6320 252 6386 293
rect 6416 1211 6482 1252
rect 6416 1177 6432 1211
rect 6466 1177 6482 1211
rect 6416 1143 6482 1177
rect 6416 1109 6432 1143
rect 6466 1109 6482 1143
rect 6416 1075 6482 1109
rect 6416 1041 6432 1075
rect 6466 1041 6482 1075
rect 6416 1007 6482 1041
rect 6416 973 6432 1007
rect 6466 973 6482 1007
rect 6416 939 6482 973
rect 6416 905 6432 939
rect 6466 905 6482 939
rect 6416 871 6482 905
rect 6416 837 6432 871
rect 6466 837 6482 871
rect 6416 803 6482 837
rect 6416 769 6432 803
rect 6466 769 6482 803
rect 6416 735 6482 769
rect 6416 701 6432 735
rect 6466 701 6482 735
rect 6416 667 6482 701
rect 6416 633 6432 667
rect 6466 633 6482 667
rect 6416 599 6482 633
rect 6416 565 6432 599
rect 6466 565 6482 599
rect 6416 531 6482 565
rect 6416 497 6432 531
rect 6466 497 6482 531
rect 6416 463 6482 497
rect 6416 429 6432 463
rect 6466 429 6482 463
rect 6416 395 6482 429
rect 6416 361 6432 395
rect 6466 361 6482 395
rect 6416 327 6482 361
rect 6416 293 6432 327
rect 6466 293 6482 327
rect 6416 252 6482 293
rect 6512 1211 6578 1252
rect 6512 1177 6528 1211
rect 6562 1177 6578 1211
rect 6512 1143 6578 1177
rect 6512 1109 6528 1143
rect 6562 1109 6578 1143
rect 6512 1075 6578 1109
rect 6512 1041 6528 1075
rect 6562 1041 6578 1075
rect 6512 1007 6578 1041
rect 6512 973 6528 1007
rect 6562 973 6578 1007
rect 6512 939 6578 973
rect 6512 905 6528 939
rect 6562 905 6578 939
rect 6512 871 6578 905
rect 6512 837 6528 871
rect 6562 837 6578 871
rect 6512 803 6578 837
rect 6512 769 6528 803
rect 6562 769 6578 803
rect 6512 735 6578 769
rect 6512 701 6528 735
rect 6562 701 6578 735
rect 6512 667 6578 701
rect 6512 633 6528 667
rect 6562 633 6578 667
rect 6512 599 6578 633
rect 6512 565 6528 599
rect 6562 565 6578 599
rect 6512 531 6578 565
rect 6512 497 6528 531
rect 6562 497 6578 531
rect 6512 463 6578 497
rect 6512 429 6528 463
rect 6562 429 6578 463
rect 6512 395 6578 429
rect 6512 361 6528 395
rect 6562 361 6578 395
rect 6512 327 6578 361
rect 6512 293 6528 327
rect 6562 293 6578 327
rect 6512 252 6578 293
rect 6608 1211 6674 1252
rect 6608 1177 6624 1211
rect 6658 1177 6674 1211
rect 6608 1143 6674 1177
rect 6608 1109 6624 1143
rect 6658 1109 6674 1143
rect 6608 1075 6674 1109
rect 6608 1041 6624 1075
rect 6658 1041 6674 1075
rect 6608 1007 6674 1041
rect 6608 973 6624 1007
rect 6658 973 6674 1007
rect 6608 939 6674 973
rect 6608 905 6624 939
rect 6658 905 6674 939
rect 6608 871 6674 905
rect 6608 837 6624 871
rect 6658 837 6674 871
rect 6608 803 6674 837
rect 6608 769 6624 803
rect 6658 769 6674 803
rect 6608 735 6674 769
rect 6608 701 6624 735
rect 6658 701 6674 735
rect 6608 667 6674 701
rect 6608 633 6624 667
rect 6658 633 6674 667
rect 6608 599 6674 633
rect 6608 565 6624 599
rect 6658 565 6674 599
rect 6608 531 6674 565
rect 6608 497 6624 531
rect 6658 497 6674 531
rect 6608 463 6674 497
rect 6608 429 6624 463
rect 6658 429 6674 463
rect 6608 395 6674 429
rect 6608 361 6624 395
rect 6658 361 6674 395
rect 6608 327 6674 361
rect 6608 293 6624 327
rect 6658 293 6674 327
rect 6608 252 6674 293
rect 6704 1211 6770 1252
rect 6704 1177 6720 1211
rect 6754 1177 6770 1211
rect 6704 1143 6770 1177
rect 6704 1109 6720 1143
rect 6754 1109 6770 1143
rect 6704 1075 6770 1109
rect 6704 1041 6720 1075
rect 6754 1041 6770 1075
rect 6704 1007 6770 1041
rect 6704 973 6720 1007
rect 6754 973 6770 1007
rect 6704 939 6770 973
rect 6704 905 6720 939
rect 6754 905 6770 939
rect 6704 871 6770 905
rect 6704 837 6720 871
rect 6754 837 6770 871
rect 6704 803 6770 837
rect 6704 769 6720 803
rect 6754 769 6770 803
rect 6704 735 6770 769
rect 6704 701 6720 735
rect 6754 701 6770 735
rect 6704 667 6770 701
rect 6704 633 6720 667
rect 6754 633 6770 667
rect 6704 599 6770 633
rect 6704 565 6720 599
rect 6754 565 6770 599
rect 6704 531 6770 565
rect 6704 497 6720 531
rect 6754 497 6770 531
rect 6704 463 6770 497
rect 6704 429 6720 463
rect 6754 429 6770 463
rect 6704 395 6770 429
rect 6704 361 6720 395
rect 6754 361 6770 395
rect 6704 327 6770 361
rect 6704 293 6720 327
rect 6754 293 6770 327
rect 6704 252 6770 293
rect 6800 1211 6866 1252
rect 6800 1177 6816 1211
rect 6850 1177 6866 1211
rect 6800 1143 6866 1177
rect 6800 1109 6816 1143
rect 6850 1109 6866 1143
rect 6800 1075 6866 1109
rect 6800 1041 6816 1075
rect 6850 1041 6866 1075
rect 6800 1007 6866 1041
rect 6800 973 6816 1007
rect 6850 973 6866 1007
rect 6800 939 6866 973
rect 6800 905 6816 939
rect 6850 905 6866 939
rect 6800 871 6866 905
rect 6800 837 6816 871
rect 6850 837 6866 871
rect 6800 803 6866 837
rect 6800 769 6816 803
rect 6850 769 6866 803
rect 6800 735 6866 769
rect 6800 701 6816 735
rect 6850 701 6866 735
rect 6800 667 6866 701
rect 6800 633 6816 667
rect 6850 633 6866 667
rect 6800 599 6866 633
rect 6800 565 6816 599
rect 6850 565 6866 599
rect 6800 531 6866 565
rect 6800 497 6816 531
rect 6850 497 6866 531
rect 6800 463 6866 497
rect 6800 429 6816 463
rect 6850 429 6866 463
rect 6800 395 6866 429
rect 6800 361 6816 395
rect 6850 361 6866 395
rect 6800 327 6866 361
rect 6800 293 6816 327
rect 6850 293 6866 327
rect 6800 252 6866 293
rect 6896 1211 6962 1252
rect 6896 1177 6912 1211
rect 6946 1177 6962 1211
rect 6896 1143 6962 1177
rect 6896 1109 6912 1143
rect 6946 1109 6962 1143
rect 6896 1075 6962 1109
rect 6896 1041 6912 1075
rect 6946 1041 6962 1075
rect 6896 1007 6962 1041
rect 6896 973 6912 1007
rect 6946 973 6962 1007
rect 6896 939 6962 973
rect 6896 905 6912 939
rect 6946 905 6962 939
rect 6896 871 6962 905
rect 6896 837 6912 871
rect 6946 837 6962 871
rect 6896 803 6962 837
rect 6896 769 6912 803
rect 6946 769 6962 803
rect 6896 735 6962 769
rect 6896 701 6912 735
rect 6946 701 6962 735
rect 6896 667 6962 701
rect 6896 633 6912 667
rect 6946 633 6962 667
rect 6896 599 6962 633
rect 6896 565 6912 599
rect 6946 565 6962 599
rect 6896 531 6962 565
rect 6896 497 6912 531
rect 6946 497 6962 531
rect 6896 463 6962 497
rect 6896 429 6912 463
rect 6946 429 6962 463
rect 6896 395 6962 429
rect 6896 361 6912 395
rect 6946 361 6962 395
rect 6896 327 6962 361
rect 6896 293 6912 327
rect 6946 293 6962 327
rect 6896 252 6962 293
rect 6992 1211 7058 1252
rect 6992 1177 7008 1211
rect 7042 1177 7058 1211
rect 6992 1143 7058 1177
rect 6992 1109 7008 1143
rect 7042 1109 7058 1143
rect 6992 1075 7058 1109
rect 6992 1041 7008 1075
rect 7042 1041 7058 1075
rect 6992 1007 7058 1041
rect 6992 973 7008 1007
rect 7042 973 7058 1007
rect 6992 939 7058 973
rect 6992 905 7008 939
rect 7042 905 7058 939
rect 6992 871 7058 905
rect 6992 837 7008 871
rect 7042 837 7058 871
rect 6992 803 7058 837
rect 6992 769 7008 803
rect 7042 769 7058 803
rect 6992 735 7058 769
rect 6992 701 7008 735
rect 7042 701 7058 735
rect 6992 667 7058 701
rect 6992 633 7008 667
rect 7042 633 7058 667
rect 6992 599 7058 633
rect 6992 565 7008 599
rect 7042 565 7058 599
rect 6992 531 7058 565
rect 6992 497 7008 531
rect 7042 497 7058 531
rect 6992 463 7058 497
rect 6992 429 7008 463
rect 7042 429 7058 463
rect 6992 395 7058 429
rect 6992 361 7008 395
rect 7042 361 7058 395
rect 6992 327 7058 361
rect 6992 293 7008 327
rect 7042 293 7058 327
rect 6992 252 7058 293
rect 7088 1211 7154 1252
rect 7088 1177 7104 1211
rect 7138 1177 7154 1211
rect 7088 1143 7154 1177
rect 7088 1109 7104 1143
rect 7138 1109 7154 1143
rect 7088 1075 7154 1109
rect 7088 1041 7104 1075
rect 7138 1041 7154 1075
rect 7088 1007 7154 1041
rect 7088 973 7104 1007
rect 7138 973 7154 1007
rect 7088 939 7154 973
rect 7088 905 7104 939
rect 7138 905 7154 939
rect 7088 871 7154 905
rect 7088 837 7104 871
rect 7138 837 7154 871
rect 7088 803 7154 837
rect 7088 769 7104 803
rect 7138 769 7154 803
rect 7088 735 7154 769
rect 7088 701 7104 735
rect 7138 701 7154 735
rect 7088 667 7154 701
rect 7088 633 7104 667
rect 7138 633 7154 667
rect 7088 599 7154 633
rect 7088 565 7104 599
rect 7138 565 7154 599
rect 7088 531 7154 565
rect 7088 497 7104 531
rect 7138 497 7154 531
rect 7088 463 7154 497
rect 7088 429 7104 463
rect 7138 429 7154 463
rect 7088 395 7154 429
rect 7088 361 7104 395
rect 7138 361 7154 395
rect 7088 327 7154 361
rect 7088 293 7104 327
rect 7138 293 7154 327
rect 7088 252 7154 293
rect 7184 1211 7250 1252
rect 7184 1177 7200 1211
rect 7234 1177 7250 1211
rect 7184 1143 7250 1177
rect 7184 1109 7200 1143
rect 7234 1109 7250 1143
rect 7184 1075 7250 1109
rect 7184 1041 7200 1075
rect 7234 1041 7250 1075
rect 7184 1007 7250 1041
rect 7184 973 7200 1007
rect 7234 973 7250 1007
rect 7184 939 7250 973
rect 7184 905 7200 939
rect 7234 905 7250 939
rect 7184 871 7250 905
rect 7184 837 7200 871
rect 7234 837 7250 871
rect 7184 803 7250 837
rect 7184 769 7200 803
rect 7234 769 7250 803
rect 7184 735 7250 769
rect 7184 701 7200 735
rect 7234 701 7250 735
rect 7184 667 7250 701
rect 7184 633 7200 667
rect 7234 633 7250 667
rect 7184 599 7250 633
rect 7184 565 7200 599
rect 7234 565 7250 599
rect 7184 531 7250 565
rect 7184 497 7200 531
rect 7234 497 7250 531
rect 7184 463 7250 497
rect 7184 429 7200 463
rect 7234 429 7250 463
rect 7184 395 7250 429
rect 7184 361 7200 395
rect 7234 361 7250 395
rect 7184 327 7250 361
rect 7184 293 7200 327
rect 7234 293 7250 327
rect 7184 252 7250 293
rect 7280 1211 7342 1252
rect 7280 1177 7296 1211
rect 7330 1177 7342 1211
rect 7280 1143 7342 1177
rect 7280 1109 7296 1143
rect 7330 1109 7342 1143
rect 7280 1075 7342 1109
rect 7280 1041 7296 1075
rect 7330 1041 7342 1075
rect 7280 1007 7342 1041
rect 7280 973 7296 1007
rect 7330 973 7342 1007
rect 7280 939 7342 973
rect 7280 905 7296 939
rect 7330 905 7342 939
rect 7280 871 7342 905
rect 7280 837 7296 871
rect 7330 837 7342 871
rect 7280 803 7342 837
rect 7280 769 7296 803
rect 7330 769 7342 803
rect 7280 735 7342 769
rect 7280 701 7296 735
rect 7330 701 7342 735
rect 7280 667 7342 701
rect 7280 633 7296 667
rect 7330 633 7342 667
rect 7280 599 7342 633
rect 7280 565 7296 599
rect 7330 565 7342 599
rect 7280 531 7342 565
rect 7280 497 7296 531
rect 7330 497 7342 531
rect 7280 463 7342 497
rect 7280 429 7296 463
rect 7330 429 7342 463
rect 7280 395 7342 429
rect 7280 361 7296 395
rect 7330 361 7342 395
rect 7280 327 7342 361
rect 7280 293 7296 327
rect 7330 293 7342 327
rect 7280 252 7342 293
rect 7900 1211 7962 1252
rect 7900 1177 7912 1211
rect 7946 1177 7962 1211
rect 7900 1143 7962 1177
rect 7900 1109 7912 1143
rect 7946 1109 7962 1143
rect 7900 1075 7962 1109
rect 7900 1041 7912 1075
rect 7946 1041 7962 1075
rect 7900 1007 7962 1041
rect 7900 973 7912 1007
rect 7946 973 7962 1007
rect 7900 939 7962 973
rect 7900 905 7912 939
rect 7946 905 7962 939
rect 7900 871 7962 905
rect 7900 837 7912 871
rect 7946 837 7962 871
rect 7900 803 7962 837
rect 7900 769 7912 803
rect 7946 769 7962 803
rect 7900 735 7962 769
rect 7900 701 7912 735
rect 7946 701 7962 735
rect 7900 667 7962 701
rect 7900 633 7912 667
rect 7946 633 7962 667
rect 7900 599 7962 633
rect 7900 565 7912 599
rect 7946 565 7962 599
rect 7900 531 7962 565
rect 7900 497 7912 531
rect 7946 497 7962 531
rect 7900 463 7962 497
rect 7900 429 7912 463
rect 7946 429 7962 463
rect 7900 395 7962 429
rect 7900 361 7912 395
rect 7946 361 7962 395
rect 7900 327 7962 361
rect 7900 293 7912 327
rect 7946 293 7962 327
rect 7900 252 7962 293
rect 7992 1211 8058 1252
rect 7992 1177 8008 1211
rect 8042 1177 8058 1211
rect 7992 1143 8058 1177
rect 7992 1109 8008 1143
rect 8042 1109 8058 1143
rect 7992 1075 8058 1109
rect 7992 1041 8008 1075
rect 8042 1041 8058 1075
rect 7992 1007 8058 1041
rect 7992 973 8008 1007
rect 8042 973 8058 1007
rect 7992 939 8058 973
rect 7992 905 8008 939
rect 8042 905 8058 939
rect 7992 871 8058 905
rect 7992 837 8008 871
rect 8042 837 8058 871
rect 7992 803 8058 837
rect 7992 769 8008 803
rect 8042 769 8058 803
rect 7992 735 8058 769
rect 7992 701 8008 735
rect 8042 701 8058 735
rect 7992 667 8058 701
rect 7992 633 8008 667
rect 8042 633 8058 667
rect 7992 599 8058 633
rect 7992 565 8008 599
rect 8042 565 8058 599
rect 7992 531 8058 565
rect 7992 497 8008 531
rect 8042 497 8058 531
rect 7992 463 8058 497
rect 7992 429 8008 463
rect 8042 429 8058 463
rect 7992 395 8058 429
rect 7992 361 8008 395
rect 8042 361 8058 395
rect 7992 327 8058 361
rect 7992 293 8008 327
rect 8042 293 8058 327
rect 7992 252 8058 293
rect 8088 1211 8154 1252
rect 8088 1177 8104 1211
rect 8138 1177 8154 1211
rect 8088 1143 8154 1177
rect 8088 1109 8104 1143
rect 8138 1109 8154 1143
rect 8088 1075 8154 1109
rect 8088 1041 8104 1075
rect 8138 1041 8154 1075
rect 8088 1007 8154 1041
rect 8088 973 8104 1007
rect 8138 973 8154 1007
rect 8088 939 8154 973
rect 8088 905 8104 939
rect 8138 905 8154 939
rect 8088 871 8154 905
rect 8088 837 8104 871
rect 8138 837 8154 871
rect 8088 803 8154 837
rect 8088 769 8104 803
rect 8138 769 8154 803
rect 8088 735 8154 769
rect 8088 701 8104 735
rect 8138 701 8154 735
rect 8088 667 8154 701
rect 8088 633 8104 667
rect 8138 633 8154 667
rect 8088 599 8154 633
rect 8088 565 8104 599
rect 8138 565 8154 599
rect 8088 531 8154 565
rect 8088 497 8104 531
rect 8138 497 8154 531
rect 8088 463 8154 497
rect 8088 429 8104 463
rect 8138 429 8154 463
rect 8088 395 8154 429
rect 8088 361 8104 395
rect 8138 361 8154 395
rect 8088 327 8154 361
rect 8088 293 8104 327
rect 8138 293 8154 327
rect 8088 252 8154 293
rect 8184 1211 8250 1252
rect 8184 1177 8200 1211
rect 8234 1177 8250 1211
rect 8184 1143 8250 1177
rect 8184 1109 8200 1143
rect 8234 1109 8250 1143
rect 8184 1075 8250 1109
rect 8184 1041 8200 1075
rect 8234 1041 8250 1075
rect 8184 1007 8250 1041
rect 8184 973 8200 1007
rect 8234 973 8250 1007
rect 8184 939 8250 973
rect 8184 905 8200 939
rect 8234 905 8250 939
rect 8184 871 8250 905
rect 8184 837 8200 871
rect 8234 837 8250 871
rect 8184 803 8250 837
rect 8184 769 8200 803
rect 8234 769 8250 803
rect 8184 735 8250 769
rect 8184 701 8200 735
rect 8234 701 8250 735
rect 8184 667 8250 701
rect 8184 633 8200 667
rect 8234 633 8250 667
rect 8184 599 8250 633
rect 8184 565 8200 599
rect 8234 565 8250 599
rect 8184 531 8250 565
rect 8184 497 8200 531
rect 8234 497 8250 531
rect 8184 463 8250 497
rect 8184 429 8200 463
rect 8234 429 8250 463
rect 8184 395 8250 429
rect 8184 361 8200 395
rect 8234 361 8250 395
rect 8184 327 8250 361
rect 8184 293 8200 327
rect 8234 293 8250 327
rect 8184 252 8250 293
rect 8280 1211 8346 1252
rect 8280 1177 8296 1211
rect 8330 1177 8346 1211
rect 8280 1143 8346 1177
rect 8280 1109 8296 1143
rect 8330 1109 8346 1143
rect 8280 1075 8346 1109
rect 8280 1041 8296 1075
rect 8330 1041 8346 1075
rect 8280 1007 8346 1041
rect 8280 973 8296 1007
rect 8330 973 8346 1007
rect 8280 939 8346 973
rect 8280 905 8296 939
rect 8330 905 8346 939
rect 8280 871 8346 905
rect 8280 837 8296 871
rect 8330 837 8346 871
rect 8280 803 8346 837
rect 8280 769 8296 803
rect 8330 769 8346 803
rect 8280 735 8346 769
rect 8280 701 8296 735
rect 8330 701 8346 735
rect 8280 667 8346 701
rect 8280 633 8296 667
rect 8330 633 8346 667
rect 8280 599 8346 633
rect 8280 565 8296 599
rect 8330 565 8346 599
rect 8280 531 8346 565
rect 8280 497 8296 531
rect 8330 497 8346 531
rect 8280 463 8346 497
rect 8280 429 8296 463
rect 8330 429 8346 463
rect 8280 395 8346 429
rect 8280 361 8296 395
rect 8330 361 8346 395
rect 8280 327 8346 361
rect 8280 293 8296 327
rect 8330 293 8346 327
rect 8280 252 8346 293
rect 8376 1211 8442 1252
rect 8376 1177 8392 1211
rect 8426 1177 8442 1211
rect 8376 1143 8442 1177
rect 8376 1109 8392 1143
rect 8426 1109 8442 1143
rect 8376 1075 8442 1109
rect 8376 1041 8392 1075
rect 8426 1041 8442 1075
rect 8376 1007 8442 1041
rect 8376 973 8392 1007
rect 8426 973 8442 1007
rect 8376 939 8442 973
rect 8376 905 8392 939
rect 8426 905 8442 939
rect 8376 871 8442 905
rect 8376 837 8392 871
rect 8426 837 8442 871
rect 8376 803 8442 837
rect 8376 769 8392 803
rect 8426 769 8442 803
rect 8376 735 8442 769
rect 8376 701 8392 735
rect 8426 701 8442 735
rect 8376 667 8442 701
rect 8376 633 8392 667
rect 8426 633 8442 667
rect 8376 599 8442 633
rect 8376 565 8392 599
rect 8426 565 8442 599
rect 8376 531 8442 565
rect 8376 497 8392 531
rect 8426 497 8442 531
rect 8376 463 8442 497
rect 8376 429 8392 463
rect 8426 429 8442 463
rect 8376 395 8442 429
rect 8376 361 8392 395
rect 8426 361 8442 395
rect 8376 327 8442 361
rect 8376 293 8392 327
rect 8426 293 8442 327
rect 8376 252 8442 293
rect 8472 1211 8538 1252
rect 8472 1177 8488 1211
rect 8522 1177 8538 1211
rect 8472 1143 8538 1177
rect 8472 1109 8488 1143
rect 8522 1109 8538 1143
rect 8472 1075 8538 1109
rect 8472 1041 8488 1075
rect 8522 1041 8538 1075
rect 8472 1007 8538 1041
rect 8472 973 8488 1007
rect 8522 973 8538 1007
rect 8472 939 8538 973
rect 8472 905 8488 939
rect 8522 905 8538 939
rect 8472 871 8538 905
rect 8472 837 8488 871
rect 8522 837 8538 871
rect 8472 803 8538 837
rect 8472 769 8488 803
rect 8522 769 8538 803
rect 8472 735 8538 769
rect 8472 701 8488 735
rect 8522 701 8538 735
rect 8472 667 8538 701
rect 8472 633 8488 667
rect 8522 633 8538 667
rect 8472 599 8538 633
rect 8472 565 8488 599
rect 8522 565 8538 599
rect 8472 531 8538 565
rect 8472 497 8488 531
rect 8522 497 8538 531
rect 8472 463 8538 497
rect 8472 429 8488 463
rect 8522 429 8538 463
rect 8472 395 8538 429
rect 8472 361 8488 395
rect 8522 361 8538 395
rect 8472 327 8538 361
rect 8472 293 8488 327
rect 8522 293 8538 327
rect 8472 252 8538 293
rect 8568 1211 8634 1252
rect 8568 1177 8584 1211
rect 8618 1177 8634 1211
rect 8568 1143 8634 1177
rect 8568 1109 8584 1143
rect 8618 1109 8634 1143
rect 8568 1075 8634 1109
rect 8568 1041 8584 1075
rect 8618 1041 8634 1075
rect 8568 1007 8634 1041
rect 8568 973 8584 1007
rect 8618 973 8634 1007
rect 8568 939 8634 973
rect 8568 905 8584 939
rect 8618 905 8634 939
rect 8568 871 8634 905
rect 8568 837 8584 871
rect 8618 837 8634 871
rect 8568 803 8634 837
rect 8568 769 8584 803
rect 8618 769 8634 803
rect 8568 735 8634 769
rect 8568 701 8584 735
rect 8618 701 8634 735
rect 8568 667 8634 701
rect 8568 633 8584 667
rect 8618 633 8634 667
rect 8568 599 8634 633
rect 8568 565 8584 599
rect 8618 565 8634 599
rect 8568 531 8634 565
rect 8568 497 8584 531
rect 8618 497 8634 531
rect 8568 463 8634 497
rect 8568 429 8584 463
rect 8618 429 8634 463
rect 8568 395 8634 429
rect 8568 361 8584 395
rect 8618 361 8634 395
rect 8568 327 8634 361
rect 8568 293 8584 327
rect 8618 293 8634 327
rect 8568 252 8634 293
rect 8664 1211 8730 1252
rect 8664 1177 8680 1211
rect 8714 1177 8730 1211
rect 8664 1143 8730 1177
rect 8664 1109 8680 1143
rect 8714 1109 8730 1143
rect 8664 1075 8730 1109
rect 8664 1041 8680 1075
rect 8714 1041 8730 1075
rect 8664 1007 8730 1041
rect 8664 973 8680 1007
rect 8714 973 8730 1007
rect 8664 939 8730 973
rect 8664 905 8680 939
rect 8714 905 8730 939
rect 8664 871 8730 905
rect 8664 837 8680 871
rect 8714 837 8730 871
rect 8664 803 8730 837
rect 8664 769 8680 803
rect 8714 769 8730 803
rect 8664 735 8730 769
rect 8664 701 8680 735
rect 8714 701 8730 735
rect 8664 667 8730 701
rect 8664 633 8680 667
rect 8714 633 8730 667
rect 8664 599 8730 633
rect 8664 565 8680 599
rect 8714 565 8730 599
rect 8664 531 8730 565
rect 8664 497 8680 531
rect 8714 497 8730 531
rect 8664 463 8730 497
rect 8664 429 8680 463
rect 8714 429 8730 463
rect 8664 395 8730 429
rect 8664 361 8680 395
rect 8714 361 8730 395
rect 8664 327 8730 361
rect 8664 293 8680 327
rect 8714 293 8730 327
rect 8664 252 8730 293
rect 8760 1211 8826 1252
rect 8760 1177 8776 1211
rect 8810 1177 8826 1211
rect 8760 1143 8826 1177
rect 8760 1109 8776 1143
rect 8810 1109 8826 1143
rect 8760 1075 8826 1109
rect 8760 1041 8776 1075
rect 8810 1041 8826 1075
rect 8760 1007 8826 1041
rect 8760 973 8776 1007
rect 8810 973 8826 1007
rect 8760 939 8826 973
rect 8760 905 8776 939
rect 8810 905 8826 939
rect 8760 871 8826 905
rect 8760 837 8776 871
rect 8810 837 8826 871
rect 8760 803 8826 837
rect 8760 769 8776 803
rect 8810 769 8826 803
rect 8760 735 8826 769
rect 8760 701 8776 735
rect 8810 701 8826 735
rect 8760 667 8826 701
rect 8760 633 8776 667
rect 8810 633 8826 667
rect 8760 599 8826 633
rect 8760 565 8776 599
rect 8810 565 8826 599
rect 8760 531 8826 565
rect 8760 497 8776 531
rect 8810 497 8826 531
rect 8760 463 8826 497
rect 8760 429 8776 463
rect 8810 429 8826 463
rect 8760 395 8826 429
rect 8760 361 8776 395
rect 8810 361 8826 395
rect 8760 327 8826 361
rect 8760 293 8776 327
rect 8810 293 8826 327
rect 8760 252 8826 293
rect 8856 1211 8922 1252
rect 8856 1177 8872 1211
rect 8906 1177 8922 1211
rect 8856 1143 8922 1177
rect 8856 1109 8872 1143
rect 8906 1109 8922 1143
rect 8856 1075 8922 1109
rect 8856 1041 8872 1075
rect 8906 1041 8922 1075
rect 8856 1007 8922 1041
rect 8856 973 8872 1007
rect 8906 973 8922 1007
rect 8856 939 8922 973
rect 8856 905 8872 939
rect 8906 905 8922 939
rect 8856 871 8922 905
rect 8856 837 8872 871
rect 8906 837 8922 871
rect 8856 803 8922 837
rect 8856 769 8872 803
rect 8906 769 8922 803
rect 8856 735 8922 769
rect 8856 701 8872 735
rect 8906 701 8922 735
rect 8856 667 8922 701
rect 8856 633 8872 667
rect 8906 633 8922 667
rect 8856 599 8922 633
rect 8856 565 8872 599
rect 8906 565 8922 599
rect 8856 531 8922 565
rect 8856 497 8872 531
rect 8906 497 8922 531
rect 8856 463 8922 497
rect 8856 429 8872 463
rect 8906 429 8922 463
rect 8856 395 8922 429
rect 8856 361 8872 395
rect 8906 361 8922 395
rect 8856 327 8922 361
rect 8856 293 8872 327
rect 8906 293 8922 327
rect 8856 252 8922 293
rect 8952 1211 9014 1252
rect 8952 1177 8968 1211
rect 9002 1177 9014 1211
rect 8952 1143 9014 1177
rect 8952 1109 8968 1143
rect 9002 1109 9014 1143
rect 8952 1075 9014 1109
rect 8952 1041 8968 1075
rect 9002 1041 9014 1075
rect 8952 1007 9014 1041
rect 8952 973 8968 1007
rect 9002 973 9014 1007
rect 8952 939 9014 973
rect 8952 905 8968 939
rect 9002 905 9014 939
rect 8952 871 9014 905
rect 8952 837 8968 871
rect 9002 837 9014 871
rect 8952 803 9014 837
rect 8952 769 8968 803
rect 9002 769 9014 803
rect 8952 735 9014 769
rect 8952 701 8968 735
rect 9002 701 9014 735
rect 8952 667 9014 701
rect 8952 633 8968 667
rect 9002 633 9014 667
rect 8952 599 9014 633
rect 8952 565 8968 599
rect 9002 565 9014 599
rect 8952 531 9014 565
rect 8952 497 8968 531
rect 9002 497 9014 531
rect 8952 463 9014 497
rect 8952 429 8968 463
rect 9002 429 9014 463
rect 8952 395 9014 429
rect 8952 361 8968 395
rect 9002 361 9014 395
rect 8952 327 9014 361
rect 8952 293 8968 327
rect 9002 293 9014 327
rect 8952 252 9014 293
rect 9220 1209 9282 1250
rect 9220 1175 9232 1209
rect 9266 1175 9282 1209
rect 9220 1141 9282 1175
rect 9220 1107 9232 1141
rect 9266 1107 9282 1141
rect 9220 1073 9282 1107
rect 9220 1039 9232 1073
rect 9266 1039 9282 1073
rect 9220 1005 9282 1039
rect 9220 971 9232 1005
rect 9266 971 9282 1005
rect 9220 937 9282 971
rect 9220 903 9232 937
rect 9266 903 9282 937
rect 9220 869 9282 903
rect 9220 835 9232 869
rect 9266 835 9282 869
rect 9220 801 9282 835
rect 9220 767 9232 801
rect 9266 767 9282 801
rect 9220 733 9282 767
rect 9220 699 9232 733
rect 9266 699 9282 733
rect 9220 665 9282 699
rect 9220 631 9232 665
rect 9266 631 9282 665
rect 9220 597 9282 631
rect 9220 563 9232 597
rect 9266 563 9282 597
rect 9220 529 9282 563
rect 9220 495 9232 529
rect 9266 495 9282 529
rect 9220 461 9282 495
rect 9220 427 9232 461
rect 9266 427 9282 461
rect 9220 393 9282 427
rect 9220 359 9232 393
rect 9266 359 9282 393
rect 9220 325 9282 359
rect 9220 291 9232 325
rect 9266 291 9282 325
rect -914 107 -902 141
rect -868 107 -856 141
rect -914 66 -856 107
rect 9220 250 9282 291
rect 9312 1209 9378 1250
rect 9312 1175 9328 1209
rect 9362 1175 9378 1209
rect 9312 1141 9378 1175
rect 9312 1107 9328 1141
rect 9362 1107 9378 1141
rect 9312 1073 9378 1107
rect 9312 1039 9328 1073
rect 9362 1039 9378 1073
rect 9312 1005 9378 1039
rect 9312 971 9328 1005
rect 9362 971 9378 1005
rect 9312 937 9378 971
rect 9312 903 9328 937
rect 9362 903 9378 937
rect 9312 869 9378 903
rect 9312 835 9328 869
rect 9362 835 9378 869
rect 9312 801 9378 835
rect 9312 767 9328 801
rect 9362 767 9378 801
rect 9312 733 9378 767
rect 9312 699 9328 733
rect 9362 699 9378 733
rect 9312 665 9378 699
rect 9312 631 9328 665
rect 9362 631 9378 665
rect 9312 597 9378 631
rect 9312 563 9328 597
rect 9362 563 9378 597
rect 9312 529 9378 563
rect 9312 495 9328 529
rect 9362 495 9378 529
rect 9312 461 9378 495
rect 9312 427 9328 461
rect 9362 427 9378 461
rect 9312 393 9378 427
rect 9312 359 9328 393
rect 9362 359 9378 393
rect 9312 325 9378 359
rect 9312 291 9328 325
rect 9362 291 9378 325
rect 9312 250 9378 291
rect 9408 1209 9474 1250
rect 9408 1175 9424 1209
rect 9458 1175 9474 1209
rect 9408 1141 9474 1175
rect 9408 1107 9424 1141
rect 9458 1107 9474 1141
rect 9408 1073 9474 1107
rect 9408 1039 9424 1073
rect 9458 1039 9474 1073
rect 9408 1005 9474 1039
rect 9408 971 9424 1005
rect 9458 971 9474 1005
rect 9408 937 9474 971
rect 9408 903 9424 937
rect 9458 903 9474 937
rect 9408 869 9474 903
rect 9408 835 9424 869
rect 9458 835 9474 869
rect 9408 801 9474 835
rect 9408 767 9424 801
rect 9458 767 9474 801
rect 9408 733 9474 767
rect 9408 699 9424 733
rect 9458 699 9474 733
rect 9408 665 9474 699
rect 9408 631 9424 665
rect 9458 631 9474 665
rect 9408 597 9474 631
rect 9408 563 9424 597
rect 9458 563 9474 597
rect 9408 529 9474 563
rect 9408 495 9424 529
rect 9458 495 9474 529
rect 9408 461 9474 495
rect 9408 427 9424 461
rect 9458 427 9474 461
rect 9408 393 9474 427
rect 9408 359 9424 393
rect 9458 359 9474 393
rect 9408 325 9474 359
rect 9408 291 9424 325
rect 9458 291 9474 325
rect 9408 250 9474 291
rect 9504 1209 9570 1250
rect 9504 1175 9520 1209
rect 9554 1175 9570 1209
rect 9504 1141 9570 1175
rect 9504 1107 9520 1141
rect 9554 1107 9570 1141
rect 9504 1073 9570 1107
rect 9504 1039 9520 1073
rect 9554 1039 9570 1073
rect 9504 1005 9570 1039
rect 9504 971 9520 1005
rect 9554 971 9570 1005
rect 9504 937 9570 971
rect 9504 903 9520 937
rect 9554 903 9570 937
rect 9504 869 9570 903
rect 9504 835 9520 869
rect 9554 835 9570 869
rect 9504 801 9570 835
rect 9504 767 9520 801
rect 9554 767 9570 801
rect 9504 733 9570 767
rect 9504 699 9520 733
rect 9554 699 9570 733
rect 9504 665 9570 699
rect 9504 631 9520 665
rect 9554 631 9570 665
rect 9504 597 9570 631
rect 9504 563 9520 597
rect 9554 563 9570 597
rect 9504 529 9570 563
rect 9504 495 9520 529
rect 9554 495 9570 529
rect 9504 461 9570 495
rect 9504 427 9520 461
rect 9554 427 9570 461
rect 9504 393 9570 427
rect 9504 359 9520 393
rect 9554 359 9570 393
rect 9504 325 9570 359
rect 9504 291 9520 325
rect 9554 291 9570 325
rect 9504 250 9570 291
rect 9600 1209 9666 1250
rect 9600 1175 9616 1209
rect 9650 1175 9666 1209
rect 9600 1141 9666 1175
rect 9600 1107 9616 1141
rect 9650 1107 9666 1141
rect 9600 1073 9666 1107
rect 9600 1039 9616 1073
rect 9650 1039 9666 1073
rect 9600 1005 9666 1039
rect 9600 971 9616 1005
rect 9650 971 9666 1005
rect 9600 937 9666 971
rect 9600 903 9616 937
rect 9650 903 9666 937
rect 9600 869 9666 903
rect 9600 835 9616 869
rect 9650 835 9666 869
rect 9600 801 9666 835
rect 9600 767 9616 801
rect 9650 767 9666 801
rect 9600 733 9666 767
rect 9600 699 9616 733
rect 9650 699 9666 733
rect 9600 665 9666 699
rect 9600 631 9616 665
rect 9650 631 9666 665
rect 9600 597 9666 631
rect 9600 563 9616 597
rect 9650 563 9666 597
rect 9600 529 9666 563
rect 9600 495 9616 529
rect 9650 495 9666 529
rect 9600 461 9666 495
rect 9600 427 9616 461
rect 9650 427 9666 461
rect 9600 393 9666 427
rect 9600 359 9616 393
rect 9650 359 9666 393
rect 9600 325 9666 359
rect 9600 291 9616 325
rect 9650 291 9666 325
rect 9600 250 9666 291
rect 9696 1209 9762 1250
rect 9696 1175 9712 1209
rect 9746 1175 9762 1209
rect 9696 1141 9762 1175
rect 9696 1107 9712 1141
rect 9746 1107 9762 1141
rect 9696 1073 9762 1107
rect 9696 1039 9712 1073
rect 9746 1039 9762 1073
rect 9696 1005 9762 1039
rect 9696 971 9712 1005
rect 9746 971 9762 1005
rect 9696 937 9762 971
rect 9696 903 9712 937
rect 9746 903 9762 937
rect 9696 869 9762 903
rect 9696 835 9712 869
rect 9746 835 9762 869
rect 9696 801 9762 835
rect 9696 767 9712 801
rect 9746 767 9762 801
rect 9696 733 9762 767
rect 9696 699 9712 733
rect 9746 699 9762 733
rect 9696 665 9762 699
rect 9696 631 9712 665
rect 9746 631 9762 665
rect 9696 597 9762 631
rect 9696 563 9712 597
rect 9746 563 9762 597
rect 9696 529 9762 563
rect 9696 495 9712 529
rect 9746 495 9762 529
rect 9696 461 9762 495
rect 9696 427 9712 461
rect 9746 427 9762 461
rect 9696 393 9762 427
rect 9696 359 9712 393
rect 9746 359 9762 393
rect 9696 325 9762 359
rect 9696 291 9712 325
rect 9746 291 9762 325
rect 9696 250 9762 291
rect 9792 1209 9858 1250
rect 9792 1175 9808 1209
rect 9842 1175 9858 1209
rect 9792 1141 9858 1175
rect 9792 1107 9808 1141
rect 9842 1107 9858 1141
rect 9792 1073 9858 1107
rect 9792 1039 9808 1073
rect 9842 1039 9858 1073
rect 9792 1005 9858 1039
rect 9792 971 9808 1005
rect 9842 971 9858 1005
rect 9792 937 9858 971
rect 9792 903 9808 937
rect 9842 903 9858 937
rect 9792 869 9858 903
rect 9792 835 9808 869
rect 9842 835 9858 869
rect 9792 801 9858 835
rect 9792 767 9808 801
rect 9842 767 9858 801
rect 9792 733 9858 767
rect 9792 699 9808 733
rect 9842 699 9858 733
rect 9792 665 9858 699
rect 9792 631 9808 665
rect 9842 631 9858 665
rect 9792 597 9858 631
rect 9792 563 9808 597
rect 9842 563 9858 597
rect 9792 529 9858 563
rect 9792 495 9808 529
rect 9842 495 9858 529
rect 9792 461 9858 495
rect 9792 427 9808 461
rect 9842 427 9858 461
rect 9792 393 9858 427
rect 9792 359 9808 393
rect 9842 359 9858 393
rect 9792 325 9858 359
rect 9792 291 9808 325
rect 9842 291 9858 325
rect 9792 250 9858 291
rect 9888 1209 9954 1250
rect 9888 1175 9904 1209
rect 9938 1175 9954 1209
rect 9888 1141 9954 1175
rect 9888 1107 9904 1141
rect 9938 1107 9954 1141
rect 9888 1073 9954 1107
rect 9888 1039 9904 1073
rect 9938 1039 9954 1073
rect 9888 1005 9954 1039
rect 9888 971 9904 1005
rect 9938 971 9954 1005
rect 9888 937 9954 971
rect 9888 903 9904 937
rect 9938 903 9954 937
rect 9888 869 9954 903
rect 9888 835 9904 869
rect 9938 835 9954 869
rect 9888 801 9954 835
rect 9888 767 9904 801
rect 9938 767 9954 801
rect 9888 733 9954 767
rect 9888 699 9904 733
rect 9938 699 9954 733
rect 9888 665 9954 699
rect 9888 631 9904 665
rect 9938 631 9954 665
rect 9888 597 9954 631
rect 9888 563 9904 597
rect 9938 563 9954 597
rect 9888 529 9954 563
rect 9888 495 9904 529
rect 9938 495 9954 529
rect 9888 461 9954 495
rect 9888 427 9904 461
rect 9938 427 9954 461
rect 9888 393 9954 427
rect 9888 359 9904 393
rect 9938 359 9954 393
rect 9888 325 9954 359
rect 9888 291 9904 325
rect 9938 291 9954 325
rect 9888 250 9954 291
rect 9984 1209 10050 1250
rect 9984 1175 10000 1209
rect 10034 1175 10050 1209
rect 9984 1141 10050 1175
rect 9984 1107 10000 1141
rect 10034 1107 10050 1141
rect 9984 1073 10050 1107
rect 9984 1039 10000 1073
rect 10034 1039 10050 1073
rect 9984 1005 10050 1039
rect 9984 971 10000 1005
rect 10034 971 10050 1005
rect 9984 937 10050 971
rect 9984 903 10000 937
rect 10034 903 10050 937
rect 9984 869 10050 903
rect 9984 835 10000 869
rect 10034 835 10050 869
rect 9984 801 10050 835
rect 9984 767 10000 801
rect 10034 767 10050 801
rect 9984 733 10050 767
rect 9984 699 10000 733
rect 10034 699 10050 733
rect 9984 665 10050 699
rect 9984 631 10000 665
rect 10034 631 10050 665
rect 9984 597 10050 631
rect 9984 563 10000 597
rect 10034 563 10050 597
rect 9984 529 10050 563
rect 9984 495 10000 529
rect 10034 495 10050 529
rect 9984 461 10050 495
rect 9984 427 10000 461
rect 10034 427 10050 461
rect 9984 393 10050 427
rect 9984 359 10000 393
rect 10034 359 10050 393
rect 9984 325 10050 359
rect 9984 291 10000 325
rect 10034 291 10050 325
rect 9984 250 10050 291
rect 10080 1209 10146 1250
rect 10080 1175 10096 1209
rect 10130 1175 10146 1209
rect 10080 1141 10146 1175
rect 10080 1107 10096 1141
rect 10130 1107 10146 1141
rect 10080 1073 10146 1107
rect 10080 1039 10096 1073
rect 10130 1039 10146 1073
rect 10080 1005 10146 1039
rect 10080 971 10096 1005
rect 10130 971 10146 1005
rect 10080 937 10146 971
rect 10080 903 10096 937
rect 10130 903 10146 937
rect 10080 869 10146 903
rect 10080 835 10096 869
rect 10130 835 10146 869
rect 10080 801 10146 835
rect 10080 767 10096 801
rect 10130 767 10146 801
rect 10080 733 10146 767
rect 10080 699 10096 733
rect 10130 699 10146 733
rect 10080 665 10146 699
rect 10080 631 10096 665
rect 10130 631 10146 665
rect 10080 597 10146 631
rect 10080 563 10096 597
rect 10130 563 10146 597
rect 10080 529 10146 563
rect 10080 495 10096 529
rect 10130 495 10146 529
rect 10080 461 10146 495
rect 10080 427 10096 461
rect 10130 427 10146 461
rect 10080 393 10146 427
rect 10080 359 10096 393
rect 10130 359 10146 393
rect 10080 325 10146 359
rect 10080 291 10096 325
rect 10130 291 10146 325
rect 10080 250 10146 291
rect 10176 1209 10242 1250
rect 10176 1175 10192 1209
rect 10226 1175 10242 1209
rect 10176 1141 10242 1175
rect 10176 1107 10192 1141
rect 10226 1107 10242 1141
rect 10176 1073 10242 1107
rect 10176 1039 10192 1073
rect 10226 1039 10242 1073
rect 10176 1005 10242 1039
rect 10176 971 10192 1005
rect 10226 971 10242 1005
rect 10176 937 10242 971
rect 10176 903 10192 937
rect 10226 903 10242 937
rect 10176 869 10242 903
rect 10176 835 10192 869
rect 10226 835 10242 869
rect 10176 801 10242 835
rect 10176 767 10192 801
rect 10226 767 10242 801
rect 10176 733 10242 767
rect 10176 699 10192 733
rect 10226 699 10242 733
rect 10176 665 10242 699
rect 10176 631 10192 665
rect 10226 631 10242 665
rect 10176 597 10242 631
rect 10176 563 10192 597
rect 10226 563 10242 597
rect 10176 529 10242 563
rect 10176 495 10192 529
rect 10226 495 10242 529
rect 10176 461 10242 495
rect 10176 427 10192 461
rect 10226 427 10242 461
rect 10176 393 10242 427
rect 10176 359 10192 393
rect 10226 359 10242 393
rect 10176 325 10242 359
rect 10176 291 10192 325
rect 10226 291 10242 325
rect 10176 250 10242 291
rect 10272 1209 10338 1250
rect 10272 1175 10288 1209
rect 10322 1175 10338 1209
rect 10272 1141 10338 1175
rect 10272 1107 10288 1141
rect 10322 1107 10338 1141
rect 10272 1073 10338 1107
rect 10272 1039 10288 1073
rect 10322 1039 10338 1073
rect 10272 1005 10338 1039
rect 10272 971 10288 1005
rect 10322 971 10338 1005
rect 10272 937 10338 971
rect 10272 903 10288 937
rect 10322 903 10338 937
rect 10272 869 10338 903
rect 10272 835 10288 869
rect 10322 835 10338 869
rect 10272 801 10338 835
rect 10272 767 10288 801
rect 10322 767 10338 801
rect 10272 733 10338 767
rect 10272 699 10288 733
rect 10322 699 10338 733
rect 10272 665 10338 699
rect 10272 631 10288 665
rect 10322 631 10338 665
rect 10272 597 10338 631
rect 10272 563 10288 597
rect 10322 563 10338 597
rect 10272 529 10338 563
rect 10272 495 10288 529
rect 10322 495 10338 529
rect 10272 461 10338 495
rect 10272 427 10288 461
rect 10322 427 10338 461
rect 10272 393 10338 427
rect 10272 359 10288 393
rect 10322 359 10338 393
rect 10272 325 10338 359
rect 10272 291 10288 325
rect 10322 291 10338 325
rect 10272 250 10338 291
rect 10368 1209 10430 1250
rect 10368 1175 10384 1209
rect 10418 1175 10430 1209
rect 10368 1141 10430 1175
rect 10368 1107 10384 1141
rect 10418 1107 10430 1141
rect 10368 1073 10430 1107
rect 10368 1039 10384 1073
rect 10418 1039 10430 1073
rect 10368 1005 10430 1039
rect 10368 971 10384 1005
rect 10418 971 10430 1005
rect 10368 937 10430 971
rect 10368 903 10384 937
rect 10418 903 10430 937
rect 10368 869 10430 903
rect 10368 835 10384 869
rect 10418 835 10430 869
rect 10368 801 10430 835
rect 10368 767 10384 801
rect 10418 767 10430 801
rect 10368 733 10430 767
rect 10368 699 10384 733
rect 10418 699 10430 733
rect 10368 665 10430 699
rect 10368 631 10384 665
rect 10418 631 10430 665
rect 10368 597 10430 631
rect 10368 563 10384 597
rect 10418 563 10430 597
rect 10368 529 10430 563
rect 10368 495 10384 529
rect 10418 495 10430 529
rect 10368 461 10430 495
rect 10368 427 10384 461
rect 10418 427 10430 461
rect 10368 393 10430 427
rect 10368 359 10384 393
rect 10418 359 10430 393
rect 10368 325 10430 359
rect 10368 291 10384 325
rect 10418 291 10430 325
rect 10368 250 10430 291
rect 10988 1209 11050 1250
rect 10988 1175 11000 1209
rect 11034 1175 11050 1209
rect 10988 1141 11050 1175
rect 10988 1107 11000 1141
rect 11034 1107 11050 1141
rect 10988 1073 11050 1107
rect 10988 1039 11000 1073
rect 11034 1039 11050 1073
rect 10988 1005 11050 1039
rect 10988 971 11000 1005
rect 11034 971 11050 1005
rect 10988 937 11050 971
rect 10988 903 11000 937
rect 11034 903 11050 937
rect 10988 869 11050 903
rect 10988 835 11000 869
rect 11034 835 11050 869
rect 10988 801 11050 835
rect 10988 767 11000 801
rect 11034 767 11050 801
rect 10988 733 11050 767
rect 10988 699 11000 733
rect 11034 699 11050 733
rect 10988 665 11050 699
rect 10988 631 11000 665
rect 11034 631 11050 665
rect 10988 597 11050 631
rect 10988 563 11000 597
rect 11034 563 11050 597
rect 10988 529 11050 563
rect 10988 495 11000 529
rect 11034 495 11050 529
rect 10988 461 11050 495
rect 10988 427 11000 461
rect 11034 427 11050 461
rect 10988 393 11050 427
rect 10988 359 11000 393
rect 11034 359 11050 393
rect 10988 325 11050 359
rect 10988 291 11000 325
rect 11034 291 11050 325
rect 10988 250 11050 291
rect 11080 1209 11146 1250
rect 11080 1175 11096 1209
rect 11130 1175 11146 1209
rect 11080 1141 11146 1175
rect 11080 1107 11096 1141
rect 11130 1107 11146 1141
rect 11080 1073 11146 1107
rect 11080 1039 11096 1073
rect 11130 1039 11146 1073
rect 11080 1005 11146 1039
rect 11080 971 11096 1005
rect 11130 971 11146 1005
rect 11080 937 11146 971
rect 11080 903 11096 937
rect 11130 903 11146 937
rect 11080 869 11146 903
rect 11080 835 11096 869
rect 11130 835 11146 869
rect 11080 801 11146 835
rect 11080 767 11096 801
rect 11130 767 11146 801
rect 11080 733 11146 767
rect 11080 699 11096 733
rect 11130 699 11146 733
rect 11080 665 11146 699
rect 11080 631 11096 665
rect 11130 631 11146 665
rect 11080 597 11146 631
rect 11080 563 11096 597
rect 11130 563 11146 597
rect 11080 529 11146 563
rect 11080 495 11096 529
rect 11130 495 11146 529
rect 11080 461 11146 495
rect 11080 427 11096 461
rect 11130 427 11146 461
rect 11080 393 11146 427
rect 11080 359 11096 393
rect 11130 359 11146 393
rect 11080 325 11146 359
rect 11080 291 11096 325
rect 11130 291 11146 325
rect 11080 250 11146 291
rect 11176 1209 11242 1250
rect 11176 1175 11192 1209
rect 11226 1175 11242 1209
rect 11176 1141 11242 1175
rect 11176 1107 11192 1141
rect 11226 1107 11242 1141
rect 11176 1073 11242 1107
rect 11176 1039 11192 1073
rect 11226 1039 11242 1073
rect 11176 1005 11242 1039
rect 11176 971 11192 1005
rect 11226 971 11242 1005
rect 11176 937 11242 971
rect 11176 903 11192 937
rect 11226 903 11242 937
rect 11176 869 11242 903
rect 11176 835 11192 869
rect 11226 835 11242 869
rect 11176 801 11242 835
rect 11176 767 11192 801
rect 11226 767 11242 801
rect 11176 733 11242 767
rect 11176 699 11192 733
rect 11226 699 11242 733
rect 11176 665 11242 699
rect 11176 631 11192 665
rect 11226 631 11242 665
rect 11176 597 11242 631
rect 11176 563 11192 597
rect 11226 563 11242 597
rect 11176 529 11242 563
rect 11176 495 11192 529
rect 11226 495 11242 529
rect 11176 461 11242 495
rect 11176 427 11192 461
rect 11226 427 11242 461
rect 11176 393 11242 427
rect 11176 359 11192 393
rect 11226 359 11242 393
rect 11176 325 11242 359
rect 11176 291 11192 325
rect 11226 291 11242 325
rect 11176 250 11242 291
rect 11272 1209 11338 1250
rect 11272 1175 11288 1209
rect 11322 1175 11338 1209
rect 11272 1141 11338 1175
rect 11272 1107 11288 1141
rect 11322 1107 11338 1141
rect 11272 1073 11338 1107
rect 11272 1039 11288 1073
rect 11322 1039 11338 1073
rect 11272 1005 11338 1039
rect 11272 971 11288 1005
rect 11322 971 11338 1005
rect 11272 937 11338 971
rect 11272 903 11288 937
rect 11322 903 11338 937
rect 11272 869 11338 903
rect 11272 835 11288 869
rect 11322 835 11338 869
rect 11272 801 11338 835
rect 11272 767 11288 801
rect 11322 767 11338 801
rect 11272 733 11338 767
rect 11272 699 11288 733
rect 11322 699 11338 733
rect 11272 665 11338 699
rect 11272 631 11288 665
rect 11322 631 11338 665
rect 11272 597 11338 631
rect 11272 563 11288 597
rect 11322 563 11338 597
rect 11272 529 11338 563
rect 11272 495 11288 529
rect 11322 495 11338 529
rect 11272 461 11338 495
rect 11272 427 11288 461
rect 11322 427 11338 461
rect 11272 393 11338 427
rect 11272 359 11288 393
rect 11322 359 11338 393
rect 11272 325 11338 359
rect 11272 291 11288 325
rect 11322 291 11338 325
rect 11272 250 11338 291
rect 11368 1209 11434 1250
rect 11368 1175 11384 1209
rect 11418 1175 11434 1209
rect 11368 1141 11434 1175
rect 11368 1107 11384 1141
rect 11418 1107 11434 1141
rect 11368 1073 11434 1107
rect 11368 1039 11384 1073
rect 11418 1039 11434 1073
rect 11368 1005 11434 1039
rect 11368 971 11384 1005
rect 11418 971 11434 1005
rect 11368 937 11434 971
rect 11368 903 11384 937
rect 11418 903 11434 937
rect 11368 869 11434 903
rect 11368 835 11384 869
rect 11418 835 11434 869
rect 11368 801 11434 835
rect 11368 767 11384 801
rect 11418 767 11434 801
rect 11368 733 11434 767
rect 11368 699 11384 733
rect 11418 699 11434 733
rect 11368 665 11434 699
rect 11368 631 11384 665
rect 11418 631 11434 665
rect 11368 597 11434 631
rect 11368 563 11384 597
rect 11418 563 11434 597
rect 11368 529 11434 563
rect 11368 495 11384 529
rect 11418 495 11434 529
rect 11368 461 11434 495
rect 11368 427 11384 461
rect 11418 427 11434 461
rect 11368 393 11434 427
rect 11368 359 11384 393
rect 11418 359 11434 393
rect 11368 325 11434 359
rect 11368 291 11384 325
rect 11418 291 11434 325
rect 11368 250 11434 291
rect 11464 1209 11530 1250
rect 11464 1175 11480 1209
rect 11514 1175 11530 1209
rect 11464 1141 11530 1175
rect 11464 1107 11480 1141
rect 11514 1107 11530 1141
rect 11464 1073 11530 1107
rect 11464 1039 11480 1073
rect 11514 1039 11530 1073
rect 11464 1005 11530 1039
rect 11464 971 11480 1005
rect 11514 971 11530 1005
rect 11464 937 11530 971
rect 11464 903 11480 937
rect 11514 903 11530 937
rect 11464 869 11530 903
rect 11464 835 11480 869
rect 11514 835 11530 869
rect 11464 801 11530 835
rect 11464 767 11480 801
rect 11514 767 11530 801
rect 11464 733 11530 767
rect 11464 699 11480 733
rect 11514 699 11530 733
rect 11464 665 11530 699
rect 11464 631 11480 665
rect 11514 631 11530 665
rect 11464 597 11530 631
rect 11464 563 11480 597
rect 11514 563 11530 597
rect 11464 529 11530 563
rect 11464 495 11480 529
rect 11514 495 11530 529
rect 11464 461 11530 495
rect 11464 427 11480 461
rect 11514 427 11530 461
rect 11464 393 11530 427
rect 11464 359 11480 393
rect 11514 359 11530 393
rect 11464 325 11530 359
rect 11464 291 11480 325
rect 11514 291 11530 325
rect 11464 250 11530 291
rect 11560 1209 11626 1250
rect 11560 1175 11576 1209
rect 11610 1175 11626 1209
rect 11560 1141 11626 1175
rect 11560 1107 11576 1141
rect 11610 1107 11626 1141
rect 11560 1073 11626 1107
rect 11560 1039 11576 1073
rect 11610 1039 11626 1073
rect 11560 1005 11626 1039
rect 11560 971 11576 1005
rect 11610 971 11626 1005
rect 11560 937 11626 971
rect 11560 903 11576 937
rect 11610 903 11626 937
rect 11560 869 11626 903
rect 11560 835 11576 869
rect 11610 835 11626 869
rect 11560 801 11626 835
rect 11560 767 11576 801
rect 11610 767 11626 801
rect 11560 733 11626 767
rect 11560 699 11576 733
rect 11610 699 11626 733
rect 11560 665 11626 699
rect 11560 631 11576 665
rect 11610 631 11626 665
rect 11560 597 11626 631
rect 11560 563 11576 597
rect 11610 563 11626 597
rect 11560 529 11626 563
rect 11560 495 11576 529
rect 11610 495 11626 529
rect 11560 461 11626 495
rect 11560 427 11576 461
rect 11610 427 11626 461
rect 11560 393 11626 427
rect 11560 359 11576 393
rect 11610 359 11626 393
rect 11560 325 11626 359
rect 11560 291 11576 325
rect 11610 291 11626 325
rect 11560 250 11626 291
rect 11656 1209 11722 1250
rect 11656 1175 11672 1209
rect 11706 1175 11722 1209
rect 11656 1141 11722 1175
rect 11656 1107 11672 1141
rect 11706 1107 11722 1141
rect 11656 1073 11722 1107
rect 11656 1039 11672 1073
rect 11706 1039 11722 1073
rect 11656 1005 11722 1039
rect 11656 971 11672 1005
rect 11706 971 11722 1005
rect 11656 937 11722 971
rect 11656 903 11672 937
rect 11706 903 11722 937
rect 11656 869 11722 903
rect 11656 835 11672 869
rect 11706 835 11722 869
rect 11656 801 11722 835
rect 11656 767 11672 801
rect 11706 767 11722 801
rect 11656 733 11722 767
rect 11656 699 11672 733
rect 11706 699 11722 733
rect 11656 665 11722 699
rect 11656 631 11672 665
rect 11706 631 11722 665
rect 11656 597 11722 631
rect 11656 563 11672 597
rect 11706 563 11722 597
rect 11656 529 11722 563
rect 11656 495 11672 529
rect 11706 495 11722 529
rect 11656 461 11722 495
rect 11656 427 11672 461
rect 11706 427 11722 461
rect 11656 393 11722 427
rect 11656 359 11672 393
rect 11706 359 11722 393
rect 11656 325 11722 359
rect 11656 291 11672 325
rect 11706 291 11722 325
rect 11656 250 11722 291
rect 11752 1209 11818 1250
rect 11752 1175 11768 1209
rect 11802 1175 11818 1209
rect 11752 1141 11818 1175
rect 11752 1107 11768 1141
rect 11802 1107 11818 1141
rect 11752 1073 11818 1107
rect 11752 1039 11768 1073
rect 11802 1039 11818 1073
rect 11752 1005 11818 1039
rect 11752 971 11768 1005
rect 11802 971 11818 1005
rect 11752 937 11818 971
rect 11752 903 11768 937
rect 11802 903 11818 937
rect 11752 869 11818 903
rect 11752 835 11768 869
rect 11802 835 11818 869
rect 11752 801 11818 835
rect 11752 767 11768 801
rect 11802 767 11818 801
rect 11752 733 11818 767
rect 11752 699 11768 733
rect 11802 699 11818 733
rect 11752 665 11818 699
rect 11752 631 11768 665
rect 11802 631 11818 665
rect 11752 597 11818 631
rect 11752 563 11768 597
rect 11802 563 11818 597
rect 11752 529 11818 563
rect 11752 495 11768 529
rect 11802 495 11818 529
rect 11752 461 11818 495
rect 11752 427 11768 461
rect 11802 427 11818 461
rect 11752 393 11818 427
rect 11752 359 11768 393
rect 11802 359 11818 393
rect 11752 325 11818 359
rect 11752 291 11768 325
rect 11802 291 11818 325
rect 11752 250 11818 291
rect 11848 1209 11914 1250
rect 11848 1175 11864 1209
rect 11898 1175 11914 1209
rect 11848 1141 11914 1175
rect 11848 1107 11864 1141
rect 11898 1107 11914 1141
rect 11848 1073 11914 1107
rect 11848 1039 11864 1073
rect 11898 1039 11914 1073
rect 11848 1005 11914 1039
rect 11848 971 11864 1005
rect 11898 971 11914 1005
rect 11848 937 11914 971
rect 11848 903 11864 937
rect 11898 903 11914 937
rect 11848 869 11914 903
rect 11848 835 11864 869
rect 11898 835 11914 869
rect 11848 801 11914 835
rect 11848 767 11864 801
rect 11898 767 11914 801
rect 11848 733 11914 767
rect 11848 699 11864 733
rect 11898 699 11914 733
rect 11848 665 11914 699
rect 11848 631 11864 665
rect 11898 631 11914 665
rect 11848 597 11914 631
rect 11848 563 11864 597
rect 11898 563 11914 597
rect 11848 529 11914 563
rect 11848 495 11864 529
rect 11898 495 11914 529
rect 11848 461 11914 495
rect 11848 427 11864 461
rect 11898 427 11914 461
rect 11848 393 11914 427
rect 11848 359 11864 393
rect 11898 359 11914 393
rect 11848 325 11914 359
rect 11848 291 11864 325
rect 11898 291 11914 325
rect 11848 250 11914 291
rect 11944 1209 12010 1250
rect 11944 1175 11960 1209
rect 11994 1175 12010 1209
rect 11944 1141 12010 1175
rect 11944 1107 11960 1141
rect 11994 1107 12010 1141
rect 11944 1073 12010 1107
rect 11944 1039 11960 1073
rect 11994 1039 12010 1073
rect 11944 1005 12010 1039
rect 11944 971 11960 1005
rect 11994 971 12010 1005
rect 11944 937 12010 971
rect 11944 903 11960 937
rect 11994 903 12010 937
rect 11944 869 12010 903
rect 11944 835 11960 869
rect 11994 835 12010 869
rect 11944 801 12010 835
rect 11944 767 11960 801
rect 11994 767 12010 801
rect 11944 733 12010 767
rect 11944 699 11960 733
rect 11994 699 12010 733
rect 11944 665 12010 699
rect 11944 631 11960 665
rect 11994 631 12010 665
rect 11944 597 12010 631
rect 11944 563 11960 597
rect 11994 563 12010 597
rect 11944 529 12010 563
rect 11944 495 11960 529
rect 11994 495 12010 529
rect 11944 461 12010 495
rect 11944 427 11960 461
rect 11994 427 12010 461
rect 11944 393 12010 427
rect 11944 359 11960 393
rect 11994 359 12010 393
rect 11944 325 12010 359
rect 11944 291 11960 325
rect 11994 291 12010 325
rect 11944 250 12010 291
rect 12040 1209 12102 1250
rect 15410 1261 15468 1300
rect 15410 1227 15422 1261
rect 15456 1227 15468 1261
rect 12040 1175 12056 1209
rect 12090 1175 12102 1209
rect 12040 1141 12102 1175
rect 12040 1107 12056 1141
rect 12090 1107 12102 1141
rect 12040 1073 12102 1107
rect 12040 1039 12056 1073
rect 12090 1039 12102 1073
rect 12040 1005 12102 1039
rect 12040 971 12056 1005
rect 12090 971 12102 1005
rect 12040 937 12102 971
rect 12040 903 12056 937
rect 12090 903 12102 937
rect 12040 869 12102 903
rect 12040 835 12056 869
rect 12090 835 12102 869
rect 12040 801 12102 835
rect 12040 767 12056 801
rect 12090 767 12102 801
rect 12040 733 12102 767
rect 12040 699 12056 733
rect 12090 699 12102 733
rect 12040 665 12102 699
rect 12040 631 12056 665
rect 12090 631 12102 665
rect 12040 597 12102 631
rect 12040 563 12056 597
rect 12090 563 12102 597
rect 12040 529 12102 563
rect 12040 495 12056 529
rect 12090 495 12102 529
rect 12040 461 12102 495
rect 12040 427 12056 461
rect 12090 427 12102 461
rect 12040 393 12102 427
rect 12040 359 12056 393
rect 12090 359 12102 393
rect 12040 325 12102 359
rect 12040 291 12056 325
rect 12090 291 12102 325
rect 12040 250 12102 291
rect 12376 1183 12438 1224
rect 12376 1149 12388 1183
rect 12422 1149 12438 1183
rect 12376 1115 12438 1149
rect 12376 1081 12388 1115
rect 12422 1081 12438 1115
rect 12376 1047 12438 1081
rect 12376 1013 12388 1047
rect 12422 1013 12438 1047
rect 12376 979 12438 1013
rect 12376 945 12388 979
rect 12422 945 12438 979
rect 12376 911 12438 945
rect 12376 877 12388 911
rect 12422 877 12438 911
rect 12376 843 12438 877
rect 12376 809 12388 843
rect 12422 809 12438 843
rect 12376 775 12438 809
rect 12376 741 12388 775
rect 12422 741 12438 775
rect 12376 707 12438 741
rect 12376 673 12388 707
rect 12422 673 12438 707
rect 12376 639 12438 673
rect 12376 605 12388 639
rect 12422 605 12438 639
rect 12376 571 12438 605
rect 12376 537 12388 571
rect 12422 537 12438 571
rect 12376 503 12438 537
rect 12376 469 12388 503
rect 12422 469 12438 503
rect 12376 435 12438 469
rect 12376 401 12388 435
rect 12422 401 12438 435
rect 12376 367 12438 401
rect 12376 333 12388 367
rect 12422 333 12438 367
rect 12376 299 12438 333
rect 12376 265 12388 299
rect 12422 265 12438 299
rect 12376 224 12438 265
rect 12468 1183 12534 1224
rect 12468 1149 12484 1183
rect 12518 1149 12534 1183
rect 12468 1115 12534 1149
rect 12468 1081 12484 1115
rect 12518 1081 12534 1115
rect 12468 1047 12534 1081
rect 12468 1013 12484 1047
rect 12518 1013 12534 1047
rect 12468 979 12534 1013
rect 12468 945 12484 979
rect 12518 945 12534 979
rect 12468 911 12534 945
rect 12468 877 12484 911
rect 12518 877 12534 911
rect 12468 843 12534 877
rect 12468 809 12484 843
rect 12518 809 12534 843
rect 12468 775 12534 809
rect 12468 741 12484 775
rect 12518 741 12534 775
rect 12468 707 12534 741
rect 12468 673 12484 707
rect 12518 673 12534 707
rect 12468 639 12534 673
rect 12468 605 12484 639
rect 12518 605 12534 639
rect 12468 571 12534 605
rect 12468 537 12484 571
rect 12518 537 12534 571
rect 12468 503 12534 537
rect 12468 469 12484 503
rect 12518 469 12534 503
rect 12468 435 12534 469
rect 12468 401 12484 435
rect 12518 401 12534 435
rect 12468 367 12534 401
rect 12468 333 12484 367
rect 12518 333 12534 367
rect 12468 299 12534 333
rect 12468 265 12484 299
rect 12518 265 12534 299
rect 12468 224 12534 265
rect 12564 1183 12630 1224
rect 12564 1149 12580 1183
rect 12614 1149 12630 1183
rect 12564 1115 12630 1149
rect 12564 1081 12580 1115
rect 12614 1081 12630 1115
rect 12564 1047 12630 1081
rect 12564 1013 12580 1047
rect 12614 1013 12630 1047
rect 12564 979 12630 1013
rect 12564 945 12580 979
rect 12614 945 12630 979
rect 12564 911 12630 945
rect 12564 877 12580 911
rect 12614 877 12630 911
rect 12564 843 12630 877
rect 12564 809 12580 843
rect 12614 809 12630 843
rect 12564 775 12630 809
rect 12564 741 12580 775
rect 12614 741 12630 775
rect 12564 707 12630 741
rect 12564 673 12580 707
rect 12614 673 12630 707
rect 12564 639 12630 673
rect 12564 605 12580 639
rect 12614 605 12630 639
rect 12564 571 12630 605
rect 12564 537 12580 571
rect 12614 537 12630 571
rect 12564 503 12630 537
rect 12564 469 12580 503
rect 12614 469 12630 503
rect 12564 435 12630 469
rect 12564 401 12580 435
rect 12614 401 12630 435
rect 12564 367 12630 401
rect 12564 333 12580 367
rect 12614 333 12630 367
rect 12564 299 12630 333
rect 12564 265 12580 299
rect 12614 265 12630 299
rect 12564 224 12630 265
rect 12660 1183 12726 1224
rect 12660 1149 12676 1183
rect 12710 1149 12726 1183
rect 12660 1115 12726 1149
rect 12660 1081 12676 1115
rect 12710 1081 12726 1115
rect 12660 1047 12726 1081
rect 12660 1013 12676 1047
rect 12710 1013 12726 1047
rect 12660 979 12726 1013
rect 12660 945 12676 979
rect 12710 945 12726 979
rect 12660 911 12726 945
rect 12660 877 12676 911
rect 12710 877 12726 911
rect 12660 843 12726 877
rect 12660 809 12676 843
rect 12710 809 12726 843
rect 12660 775 12726 809
rect 12660 741 12676 775
rect 12710 741 12726 775
rect 12660 707 12726 741
rect 12660 673 12676 707
rect 12710 673 12726 707
rect 12660 639 12726 673
rect 12660 605 12676 639
rect 12710 605 12726 639
rect 12660 571 12726 605
rect 12660 537 12676 571
rect 12710 537 12726 571
rect 12660 503 12726 537
rect 12660 469 12676 503
rect 12710 469 12726 503
rect 12660 435 12726 469
rect 12660 401 12676 435
rect 12710 401 12726 435
rect 12660 367 12726 401
rect 12660 333 12676 367
rect 12710 333 12726 367
rect 12660 299 12726 333
rect 12660 265 12676 299
rect 12710 265 12726 299
rect 12660 224 12726 265
rect 12756 1183 12822 1224
rect 12756 1149 12772 1183
rect 12806 1149 12822 1183
rect 12756 1115 12822 1149
rect 12756 1081 12772 1115
rect 12806 1081 12822 1115
rect 12756 1047 12822 1081
rect 12756 1013 12772 1047
rect 12806 1013 12822 1047
rect 12756 979 12822 1013
rect 12756 945 12772 979
rect 12806 945 12822 979
rect 12756 911 12822 945
rect 12756 877 12772 911
rect 12806 877 12822 911
rect 12756 843 12822 877
rect 12756 809 12772 843
rect 12806 809 12822 843
rect 12756 775 12822 809
rect 12756 741 12772 775
rect 12806 741 12822 775
rect 12756 707 12822 741
rect 12756 673 12772 707
rect 12806 673 12822 707
rect 12756 639 12822 673
rect 12756 605 12772 639
rect 12806 605 12822 639
rect 12756 571 12822 605
rect 12756 537 12772 571
rect 12806 537 12822 571
rect 12756 503 12822 537
rect 12756 469 12772 503
rect 12806 469 12822 503
rect 12756 435 12822 469
rect 12756 401 12772 435
rect 12806 401 12822 435
rect 12756 367 12822 401
rect 12756 333 12772 367
rect 12806 333 12822 367
rect 12756 299 12822 333
rect 12756 265 12772 299
rect 12806 265 12822 299
rect 12756 224 12822 265
rect 12852 1183 12918 1224
rect 12852 1149 12868 1183
rect 12902 1149 12918 1183
rect 12852 1115 12918 1149
rect 12852 1081 12868 1115
rect 12902 1081 12918 1115
rect 12852 1047 12918 1081
rect 12852 1013 12868 1047
rect 12902 1013 12918 1047
rect 12852 979 12918 1013
rect 12852 945 12868 979
rect 12902 945 12918 979
rect 12852 911 12918 945
rect 12852 877 12868 911
rect 12902 877 12918 911
rect 12852 843 12918 877
rect 12852 809 12868 843
rect 12902 809 12918 843
rect 12852 775 12918 809
rect 12852 741 12868 775
rect 12902 741 12918 775
rect 12852 707 12918 741
rect 12852 673 12868 707
rect 12902 673 12918 707
rect 12852 639 12918 673
rect 12852 605 12868 639
rect 12902 605 12918 639
rect 12852 571 12918 605
rect 12852 537 12868 571
rect 12902 537 12918 571
rect 12852 503 12918 537
rect 12852 469 12868 503
rect 12902 469 12918 503
rect 12852 435 12918 469
rect 12852 401 12868 435
rect 12902 401 12918 435
rect 12852 367 12918 401
rect 12852 333 12868 367
rect 12902 333 12918 367
rect 12852 299 12918 333
rect 12852 265 12868 299
rect 12902 265 12918 299
rect 12852 224 12918 265
rect 12948 1183 13014 1224
rect 12948 1149 12964 1183
rect 12998 1149 13014 1183
rect 12948 1115 13014 1149
rect 12948 1081 12964 1115
rect 12998 1081 13014 1115
rect 12948 1047 13014 1081
rect 12948 1013 12964 1047
rect 12998 1013 13014 1047
rect 12948 979 13014 1013
rect 12948 945 12964 979
rect 12998 945 13014 979
rect 12948 911 13014 945
rect 12948 877 12964 911
rect 12998 877 13014 911
rect 12948 843 13014 877
rect 12948 809 12964 843
rect 12998 809 13014 843
rect 12948 775 13014 809
rect 12948 741 12964 775
rect 12998 741 13014 775
rect 12948 707 13014 741
rect 12948 673 12964 707
rect 12998 673 13014 707
rect 12948 639 13014 673
rect 12948 605 12964 639
rect 12998 605 13014 639
rect 12948 571 13014 605
rect 12948 537 12964 571
rect 12998 537 13014 571
rect 12948 503 13014 537
rect 12948 469 12964 503
rect 12998 469 13014 503
rect 12948 435 13014 469
rect 12948 401 12964 435
rect 12998 401 13014 435
rect 12948 367 13014 401
rect 12948 333 12964 367
rect 12998 333 13014 367
rect 12948 299 13014 333
rect 12948 265 12964 299
rect 12998 265 13014 299
rect 12948 224 13014 265
rect 13044 1183 13110 1224
rect 13044 1149 13060 1183
rect 13094 1149 13110 1183
rect 13044 1115 13110 1149
rect 13044 1081 13060 1115
rect 13094 1081 13110 1115
rect 13044 1047 13110 1081
rect 13044 1013 13060 1047
rect 13094 1013 13110 1047
rect 13044 979 13110 1013
rect 13044 945 13060 979
rect 13094 945 13110 979
rect 13044 911 13110 945
rect 13044 877 13060 911
rect 13094 877 13110 911
rect 13044 843 13110 877
rect 13044 809 13060 843
rect 13094 809 13110 843
rect 13044 775 13110 809
rect 13044 741 13060 775
rect 13094 741 13110 775
rect 13044 707 13110 741
rect 13044 673 13060 707
rect 13094 673 13110 707
rect 13044 639 13110 673
rect 13044 605 13060 639
rect 13094 605 13110 639
rect 13044 571 13110 605
rect 13044 537 13060 571
rect 13094 537 13110 571
rect 13044 503 13110 537
rect 13044 469 13060 503
rect 13094 469 13110 503
rect 13044 435 13110 469
rect 13044 401 13060 435
rect 13094 401 13110 435
rect 13044 367 13110 401
rect 13044 333 13060 367
rect 13094 333 13110 367
rect 13044 299 13110 333
rect 13044 265 13060 299
rect 13094 265 13110 299
rect 13044 224 13110 265
rect 13140 1183 13206 1224
rect 13140 1149 13156 1183
rect 13190 1149 13206 1183
rect 13140 1115 13206 1149
rect 13140 1081 13156 1115
rect 13190 1081 13206 1115
rect 13140 1047 13206 1081
rect 13140 1013 13156 1047
rect 13190 1013 13206 1047
rect 13140 979 13206 1013
rect 13140 945 13156 979
rect 13190 945 13206 979
rect 13140 911 13206 945
rect 13140 877 13156 911
rect 13190 877 13206 911
rect 13140 843 13206 877
rect 13140 809 13156 843
rect 13190 809 13206 843
rect 13140 775 13206 809
rect 13140 741 13156 775
rect 13190 741 13206 775
rect 13140 707 13206 741
rect 13140 673 13156 707
rect 13190 673 13206 707
rect 13140 639 13206 673
rect 13140 605 13156 639
rect 13190 605 13206 639
rect 13140 571 13206 605
rect 13140 537 13156 571
rect 13190 537 13206 571
rect 13140 503 13206 537
rect 13140 469 13156 503
rect 13190 469 13206 503
rect 13140 435 13206 469
rect 13140 401 13156 435
rect 13190 401 13206 435
rect 13140 367 13206 401
rect 13140 333 13156 367
rect 13190 333 13206 367
rect 13140 299 13206 333
rect 13140 265 13156 299
rect 13190 265 13206 299
rect 13140 224 13206 265
rect 13236 1183 13302 1224
rect 13236 1149 13252 1183
rect 13286 1149 13302 1183
rect 13236 1115 13302 1149
rect 13236 1081 13252 1115
rect 13286 1081 13302 1115
rect 13236 1047 13302 1081
rect 13236 1013 13252 1047
rect 13286 1013 13302 1047
rect 13236 979 13302 1013
rect 13236 945 13252 979
rect 13286 945 13302 979
rect 13236 911 13302 945
rect 13236 877 13252 911
rect 13286 877 13302 911
rect 13236 843 13302 877
rect 13236 809 13252 843
rect 13286 809 13302 843
rect 13236 775 13302 809
rect 13236 741 13252 775
rect 13286 741 13302 775
rect 13236 707 13302 741
rect 13236 673 13252 707
rect 13286 673 13302 707
rect 13236 639 13302 673
rect 13236 605 13252 639
rect 13286 605 13302 639
rect 13236 571 13302 605
rect 13236 537 13252 571
rect 13286 537 13302 571
rect 13236 503 13302 537
rect 13236 469 13252 503
rect 13286 469 13302 503
rect 13236 435 13302 469
rect 13236 401 13252 435
rect 13286 401 13302 435
rect 13236 367 13302 401
rect 13236 333 13252 367
rect 13286 333 13302 367
rect 13236 299 13302 333
rect 13236 265 13252 299
rect 13286 265 13302 299
rect 13236 224 13302 265
rect 13332 1183 13398 1224
rect 13332 1149 13348 1183
rect 13382 1149 13398 1183
rect 13332 1115 13398 1149
rect 13332 1081 13348 1115
rect 13382 1081 13398 1115
rect 13332 1047 13398 1081
rect 13332 1013 13348 1047
rect 13382 1013 13398 1047
rect 13332 979 13398 1013
rect 13332 945 13348 979
rect 13382 945 13398 979
rect 13332 911 13398 945
rect 13332 877 13348 911
rect 13382 877 13398 911
rect 13332 843 13398 877
rect 13332 809 13348 843
rect 13382 809 13398 843
rect 13332 775 13398 809
rect 13332 741 13348 775
rect 13382 741 13398 775
rect 13332 707 13398 741
rect 13332 673 13348 707
rect 13382 673 13398 707
rect 13332 639 13398 673
rect 13332 605 13348 639
rect 13382 605 13398 639
rect 13332 571 13398 605
rect 13332 537 13348 571
rect 13382 537 13398 571
rect 13332 503 13398 537
rect 13332 469 13348 503
rect 13382 469 13398 503
rect 13332 435 13398 469
rect 13332 401 13348 435
rect 13382 401 13398 435
rect 13332 367 13398 401
rect 13332 333 13348 367
rect 13382 333 13398 367
rect 13332 299 13398 333
rect 13332 265 13348 299
rect 13382 265 13398 299
rect 13332 224 13398 265
rect 13428 1183 13494 1224
rect 13428 1149 13444 1183
rect 13478 1149 13494 1183
rect 13428 1115 13494 1149
rect 13428 1081 13444 1115
rect 13478 1081 13494 1115
rect 13428 1047 13494 1081
rect 13428 1013 13444 1047
rect 13478 1013 13494 1047
rect 13428 979 13494 1013
rect 13428 945 13444 979
rect 13478 945 13494 979
rect 13428 911 13494 945
rect 13428 877 13444 911
rect 13478 877 13494 911
rect 13428 843 13494 877
rect 13428 809 13444 843
rect 13478 809 13494 843
rect 13428 775 13494 809
rect 13428 741 13444 775
rect 13478 741 13494 775
rect 13428 707 13494 741
rect 13428 673 13444 707
rect 13478 673 13494 707
rect 13428 639 13494 673
rect 13428 605 13444 639
rect 13478 605 13494 639
rect 13428 571 13494 605
rect 13428 537 13444 571
rect 13478 537 13494 571
rect 13428 503 13494 537
rect 13428 469 13444 503
rect 13478 469 13494 503
rect 13428 435 13494 469
rect 13428 401 13444 435
rect 13478 401 13494 435
rect 13428 367 13494 401
rect 13428 333 13444 367
rect 13478 333 13494 367
rect 13428 299 13494 333
rect 13428 265 13444 299
rect 13478 265 13494 299
rect 13428 224 13494 265
rect 13524 1183 13586 1224
rect 13524 1149 13540 1183
rect 13574 1149 13586 1183
rect 13524 1115 13586 1149
rect 13524 1081 13540 1115
rect 13574 1081 13586 1115
rect 13524 1047 13586 1081
rect 13524 1013 13540 1047
rect 13574 1013 13586 1047
rect 13524 979 13586 1013
rect 13524 945 13540 979
rect 13574 945 13586 979
rect 13524 911 13586 945
rect 13524 877 13540 911
rect 13574 877 13586 911
rect 13524 843 13586 877
rect 13524 809 13540 843
rect 13574 809 13586 843
rect 13524 775 13586 809
rect 13524 741 13540 775
rect 13574 741 13586 775
rect 13524 707 13586 741
rect 13524 673 13540 707
rect 13574 673 13586 707
rect 13524 639 13586 673
rect 13524 605 13540 639
rect 13574 605 13586 639
rect 13524 571 13586 605
rect 13524 537 13540 571
rect 13574 537 13586 571
rect 13524 503 13586 537
rect 13524 469 13540 503
rect 13574 469 13586 503
rect 13524 435 13586 469
rect 13524 401 13540 435
rect 13574 401 13586 435
rect 13524 367 13586 401
rect 13524 333 13540 367
rect 13574 333 13586 367
rect 13524 299 13586 333
rect 13524 265 13540 299
rect 13574 265 13586 299
rect 13524 224 13586 265
rect 14144 1183 14206 1224
rect 14144 1149 14156 1183
rect 14190 1149 14206 1183
rect 14144 1115 14206 1149
rect 14144 1081 14156 1115
rect 14190 1081 14206 1115
rect 14144 1047 14206 1081
rect 14144 1013 14156 1047
rect 14190 1013 14206 1047
rect 14144 979 14206 1013
rect 14144 945 14156 979
rect 14190 945 14206 979
rect 14144 911 14206 945
rect 14144 877 14156 911
rect 14190 877 14206 911
rect 14144 843 14206 877
rect 14144 809 14156 843
rect 14190 809 14206 843
rect 14144 775 14206 809
rect 14144 741 14156 775
rect 14190 741 14206 775
rect 14144 707 14206 741
rect 14144 673 14156 707
rect 14190 673 14206 707
rect 14144 639 14206 673
rect 14144 605 14156 639
rect 14190 605 14206 639
rect 14144 571 14206 605
rect 14144 537 14156 571
rect 14190 537 14206 571
rect 14144 503 14206 537
rect 14144 469 14156 503
rect 14190 469 14206 503
rect 14144 435 14206 469
rect 14144 401 14156 435
rect 14190 401 14206 435
rect 14144 367 14206 401
rect 14144 333 14156 367
rect 14190 333 14206 367
rect 14144 299 14206 333
rect 14144 265 14156 299
rect 14190 265 14206 299
rect 14144 224 14206 265
rect 14236 1183 14302 1224
rect 14236 1149 14252 1183
rect 14286 1149 14302 1183
rect 14236 1115 14302 1149
rect 14236 1081 14252 1115
rect 14286 1081 14302 1115
rect 14236 1047 14302 1081
rect 14236 1013 14252 1047
rect 14286 1013 14302 1047
rect 14236 979 14302 1013
rect 14236 945 14252 979
rect 14286 945 14302 979
rect 14236 911 14302 945
rect 14236 877 14252 911
rect 14286 877 14302 911
rect 14236 843 14302 877
rect 14236 809 14252 843
rect 14286 809 14302 843
rect 14236 775 14302 809
rect 14236 741 14252 775
rect 14286 741 14302 775
rect 14236 707 14302 741
rect 14236 673 14252 707
rect 14286 673 14302 707
rect 14236 639 14302 673
rect 14236 605 14252 639
rect 14286 605 14302 639
rect 14236 571 14302 605
rect 14236 537 14252 571
rect 14286 537 14302 571
rect 14236 503 14302 537
rect 14236 469 14252 503
rect 14286 469 14302 503
rect 14236 435 14302 469
rect 14236 401 14252 435
rect 14286 401 14302 435
rect 14236 367 14302 401
rect 14236 333 14252 367
rect 14286 333 14302 367
rect 14236 299 14302 333
rect 14236 265 14252 299
rect 14286 265 14302 299
rect 14236 224 14302 265
rect 14332 1183 14398 1224
rect 14332 1149 14348 1183
rect 14382 1149 14398 1183
rect 14332 1115 14398 1149
rect 14332 1081 14348 1115
rect 14382 1081 14398 1115
rect 14332 1047 14398 1081
rect 14332 1013 14348 1047
rect 14382 1013 14398 1047
rect 14332 979 14398 1013
rect 14332 945 14348 979
rect 14382 945 14398 979
rect 14332 911 14398 945
rect 14332 877 14348 911
rect 14382 877 14398 911
rect 14332 843 14398 877
rect 14332 809 14348 843
rect 14382 809 14398 843
rect 14332 775 14398 809
rect 14332 741 14348 775
rect 14382 741 14398 775
rect 14332 707 14398 741
rect 14332 673 14348 707
rect 14382 673 14398 707
rect 14332 639 14398 673
rect 14332 605 14348 639
rect 14382 605 14398 639
rect 14332 571 14398 605
rect 14332 537 14348 571
rect 14382 537 14398 571
rect 14332 503 14398 537
rect 14332 469 14348 503
rect 14382 469 14398 503
rect 14332 435 14398 469
rect 14332 401 14348 435
rect 14382 401 14398 435
rect 14332 367 14398 401
rect 14332 333 14348 367
rect 14382 333 14398 367
rect 14332 299 14398 333
rect 14332 265 14348 299
rect 14382 265 14398 299
rect 14332 224 14398 265
rect 14428 1183 14494 1224
rect 14428 1149 14444 1183
rect 14478 1149 14494 1183
rect 14428 1115 14494 1149
rect 14428 1081 14444 1115
rect 14478 1081 14494 1115
rect 14428 1047 14494 1081
rect 14428 1013 14444 1047
rect 14478 1013 14494 1047
rect 14428 979 14494 1013
rect 14428 945 14444 979
rect 14478 945 14494 979
rect 14428 911 14494 945
rect 14428 877 14444 911
rect 14478 877 14494 911
rect 14428 843 14494 877
rect 14428 809 14444 843
rect 14478 809 14494 843
rect 14428 775 14494 809
rect 14428 741 14444 775
rect 14478 741 14494 775
rect 14428 707 14494 741
rect 14428 673 14444 707
rect 14478 673 14494 707
rect 14428 639 14494 673
rect 14428 605 14444 639
rect 14478 605 14494 639
rect 14428 571 14494 605
rect 14428 537 14444 571
rect 14478 537 14494 571
rect 14428 503 14494 537
rect 14428 469 14444 503
rect 14478 469 14494 503
rect 14428 435 14494 469
rect 14428 401 14444 435
rect 14478 401 14494 435
rect 14428 367 14494 401
rect 14428 333 14444 367
rect 14478 333 14494 367
rect 14428 299 14494 333
rect 14428 265 14444 299
rect 14478 265 14494 299
rect 14428 224 14494 265
rect 14524 1183 14590 1224
rect 14524 1149 14540 1183
rect 14574 1149 14590 1183
rect 14524 1115 14590 1149
rect 14524 1081 14540 1115
rect 14574 1081 14590 1115
rect 14524 1047 14590 1081
rect 14524 1013 14540 1047
rect 14574 1013 14590 1047
rect 14524 979 14590 1013
rect 14524 945 14540 979
rect 14574 945 14590 979
rect 14524 911 14590 945
rect 14524 877 14540 911
rect 14574 877 14590 911
rect 14524 843 14590 877
rect 14524 809 14540 843
rect 14574 809 14590 843
rect 14524 775 14590 809
rect 14524 741 14540 775
rect 14574 741 14590 775
rect 14524 707 14590 741
rect 14524 673 14540 707
rect 14574 673 14590 707
rect 14524 639 14590 673
rect 14524 605 14540 639
rect 14574 605 14590 639
rect 14524 571 14590 605
rect 14524 537 14540 571
rect 14574 537 14590 571
rect 14524 503 14590 537
rect 14524 469 14540 503
rect 14574 469 14590 503
rect 14524 435 14590 469
rect 14524 401 14540 435
rect 14574 401 14590 435
rect 14524 367 14590 401
rect 14524 333 14540 367
rect 14574 333 14590 367
rect 14524 299 14590 333
rect 14524 265 14540 299
rect 14574 265 14590 299
rect 14524 224 14590 265
rect 14620 1183 14686 1224
rect 14620 1149 14636 1183
rect 14670 1149 14686 1183
rect 14620 1115 14686 1149
rect 14620 1081 14636 1115
rect 14670 1081 14686 1115
rect 14620 1047 14686 1081
rect 14620 1013 14636 1047
rect 14670 1013 14686 1047
rect 14620 979 14686 1013
rect 14620 945 14636 979
rect 14670 945 14686 979
rect 14620 911 14686 945
rect 14620 877 14636 911
rect 14670 877 14686 911
rect 14620 843 14686 877
rect 14620 809 14636 843
rect 14670 809 14686 843
rect 14620 775 14686 809
rect 14620 741 14636 775
rect 14670 741 14686 775
rect 14620 707 14686 741
rect 14620 673 14636 707
rect 14670 673 14686 707
rect 14620 639 14686 673
rect 14620 605 14636 639
rect 14670 605 14686 639
rect 14620 571 14686 605
rect 14620 537 14636 571
rect 14670 537 14686 571
rect 14620 503 14686 537
rect 14620 469 14636 503
rect 14670 469 14686 503
rect 14620 435 14686 469
rect 14620 401 14636 435
rect 14670 401 14686 435
rect 14620 367 14686 401
rect 14620 333 14636 367
rect 14670 333 14686 367
rect 14620 299 14686 333
rect 14620 265 14636 299
rect 14670 265 14686 299
rect 14620 224 14686 265
rect 14716 1183 14782 1224
rect 14716 1149 14732 1183
rect 14766 1149 14782 1183
rect 14716 1115 14782 1149
rect 14716 1081 14732 1115
rect 14766 1081 14782 1115
rect 14716 1047 14782 1081
rect 14716 1013 14732 1047
rect 14766 1013 14782 1047
rect 14716 979 14782 1013
rect 14716 945 14732 979
rect 14766 945 14782 979
rect 14716 911 14782 945
rect 14716 877 14732 911
rect 14766 877 14782 911
rect 14716 843 14782 877
rect 14716 809 14732 843
rect 14766 809 14782 843
rect 14716 775 14782 809
rect 14716 741 14732 775
rect 14766 741 14782 775
rect 14716 707 14782 741
rect 14716 673 14732 707
rect 14766 673 14782 707
rect 14716 639 14782 673
rect 14716 605 14732 639
rect 14766 605 14782 639
rect 14716 571 14782 605
rect 14716 537 14732 571
rect 14766 537 14782 571
rect 14716 503 14782 537
rect 14716 469 14732 503
rect 14766 469 14782 503
rect 14716 435 14782 469
rect 14716 401 14732 435
rect 14766 401 14782 435
rect 14716 367 14782 401
rect 14716 333 14732 367
rect 14766 333 14782 367
rect 14716 299 14782 333
rect 14716 265 14732 299
rect 14766 265 14782 299
rect 14716 224 14782 265
rect 14812 1183 14878 1224
rect 14812 1149 14828 1183
rect 14862 1149 14878 1183
rect 14812 1115 14878 1149
rect 14812 1081 14828 1115
rect 14862 1081 14878 1115
rect 14812 1047 14878 1081
rect 14812 1013 14828 1047
rect 14862 1013 14878 1047
rect 14812 979 14878 1013
rect 14812 945 14828 979
rect 14862 945 14878 979
rect 14812 911 14878 945
rect 14812 877 14828 911
rect 14862 877 14878 911
rect 14812 843 14878 877
rect 14812 809 14828 843
rect 14862 809 14878 843
rect 14812 775 14878 809
rect 14812 741 14828 775
rect 14862 741 14878 775
rect 14812 707 14878 741
rect 14812 673 14828 707
rect 14862 673 14878 707
rect 14812 639 14878 673
rect 14812 605 14828 639
rect 14862 605 14878 639
rect 14812 571 14878 605
rect 14812 537 14828 571
rect 14862 537 14878 571
rect 14812 503 14878 537
rect 14812 469 14828 503
rect 14862 469 14878 503
rect 14812 435 14878 469
rect 14812 401 14828 435
rect 14862 401 14878 435
rect 14812 367 14878 401
rect 14812 333 14828 367
rect 14862 333 14878 367
rect 14812 299 14878 333
rect 14812 265 14828 299
rect 14862 265 14878 299
rect 14812 224 14878 265
rect 14908 1183 14974 1224
rect 14908 1149 14924 1183
rect 14958 1149 14974 1183
rect 14908 1115 14974 1149
rect 14908 1081 14924 1115
rect 14958 1081 14974 1115
rect 14908 1047 14974 1081
rect 14908 1013 14924 1047
rect 14958 1013 14974 1047
rect 14908 979 14974 1013
rect 14908 945 14924 979
rect 14958 945 14974 979
rect 14908 911 14974 945
rect 14908 877 14924 911
rect 14958 877 14974 911
rect 14908 843 14974 877
rect 14908 809 14924 843
rect 14958 809 14974 843
rect 14908 775 14974 809
rect 14908 741 14924 775
rect 14958 741 14974 775
rect 14908 707 14974 741
rect 14908 673 14924 707
rect 14958 673 14974 707
rect 14908 639 14974 673
rect 14908 605 14924 639
rect 14958 605 14974 639
rect 14908 571 14974 605
rect 14908 537 14924 571
rect 14958 537 14974 571
rect 14908 503 14974 537
rect 14908 469 14924 503
rect 14958 469 14974 503
rect 14908 435 14974 469
rect 14908 401 14924 435
rect 14958 401 14974 435
rect 14908 367 14974 401
rect 14908 333 14924 367
rect 14958 333 14974 367
rect 14908 299 14974 333
rect 14908 265 14924 299
rect 14958 265 14974 299
rect 14908 224 14974 265
rect 15004 1183 15070 1224
rect 15004 1149 15020 1183
rect 15054 1149 15070 1183
rect 15004 1115 15070 1149
rect 15004 1081 15020 1115
rect 15054 1081 15070 1115
rect 15004 1047 15070 1081
rect 15004 1013 15020 1047
rect 15054 1013 15070 1047
rect 15004 979 15070 1013
rect 15004 945 15020 979
rect 15054 945 15070 979
rect 15004 911 15070 945
rect 15004 877 15020 911
rect 15054 877 15070 911
rect 15004 843 15070 877
rect 15004 809 15020 843
rect 15054 809 15070 843
rect 15004 775 15070 809
rect 15004 741 15020 775
rect 15054 741 15070 775
rect 15004 707 15070 741
rect 15004 673 15020 707
rect 15054 673 15070 707
rect 15004 639 15070 673
rect 15004 605 15020 639
rect 15054 605 15070 639
rect 15004 571 15070 605
rect 15004 537 15020 571
rect 15054 537 15070 571
rect 15004 503 15070 537
rect 15004 469 15020 503
rect 15054 469 15070 503
rect 15004 435 15070 469
rect 15004 401 15020 435
rect 15054 401 15070 435
rect 15004 367 15070 401
rect 15004 333 15020 367
rect 15054 333 15070 367
rect 15004 299 15070 333
rect 15004 265 15020 299
rect 15054 265 15070 299
rect 15004 224 15070 265
rect 15100 1183 15166 1224
rect 15100 1149 15116 1183
rect 15150 1149 15166 1183
rect 15100 1115 15166 1149
rect 15100 1081 15116 1115
rect 15150 1081 15166 1115
rect 15100 1047 15166 1081
rect 15100 1013 15116 1047
rect 15150 1013 15166 1047
rect 15100 979 15166 1013
rect 15100 945 15116 979
rect 15150 945 15166 979
rect 15100 911 15166 945
rect 15100 877 15116 911
rect 15150 877 15166 911
rect 15100 843 15166 877
rect 15100 809 15116 843
rect 15150 809 15166 843
rect 15100 775 15166 809
rect 15100 741 15116 775
rect 15150 741 15166 775
rect 15100 707 15166 741
rect 15100 673 15116 707
rect 15150 673 15166 707
rect 15100 639 15166 673
rect 15100 605 15116 639
rect 15150 605 15166 639
rect 15100 571 15166 605
rect 15100 537 15116 571
rect 15150 537 15166 571
rect 15100 503 15166 537
rect 15100 469 15116 503
rect 15150 469 15166 503
rect 15100 435 15166 469
rect 15100 401 15116 435
rect 15150 401 15166 435
rect 15100 367 15166 401
rect 15100 333 15116 367
rect 15150 333 15166 367
rect 15100 299 15166 333
rect 15100 265 15116 299
rect 15150 265 15166 299
rect 15100 224 15166 265
rect 15196 1183 15258 1224
rect 15196 1149 15212 1183
rect 15246 1149 15258 1183
rect 15196 1115 15258 1149
rect 15196 1081 15212 1115
rect 15246 1081 15258 1115
rect 15196 1047 15258 1081
rect 15196 1013 15212 1047
rect 15246 1013 15258 1047
rect 15196 979 15258 1013
rect 15196 945 15212 979
rect 15246 945 15258 979
rect 15196 911 15258 945
rect 15196 877 15212 911
rect 15246 877 15258 911
rect 15196 843 15258 877
rect 15196 809 15212 843
rect 15246 809 15258 843
rect 15196 775 15258 809
rect 15196 741 15212 775
rect 15246 741 15258 775
rect 15196 707 15258 741
rect 15196 673 15212 707
rect 15246 673 15258 707
rect 15196 639 15258 673
rect 15196 605 15212 639
rect 15246 605 15258 639
rect 15196 571 15258 605
rect 15196 537 15212 571
rect 15246 537 15258 571
rect 15196 503 15258 537
rect 15196 469 15212 503
rect 15246 469 15258 503
rect 15196 435 15258 469
rect 15196 401 15212 435
rect 15246 401 15258 435
rect 15196 367 15258 401
rect 15196 333 15212 367
rect 15246 333 15258 367
rect 15196 299 15258 333
rect 15196 265 15212 299
rect 15246 265 15258 299
rect 15196 224 15258 265
rect 15410 1193 15468 1227
rect 15410 1159 15422 1193
rect 15456 1159 15468 1193
rect 15410 1125 15468 1159
rect 15410 1091 15422 1125
rect 15456 1091 15468 1125
rect 15410 1057 15468 1091
rect 15410 1023 15422 1057
rect 15456 1023 15468 1057
rect 15410 989 15468 1023
rect 15410 955 15422 989
rect 15456 955 15468 989
rect 15410 921 15468 955
rect 15410 887 15422 921
rect 15456 887 15468 921
rect 15410 853 15468 887
rect 15410 819 15422 853
rect 15456 819 15468 853
rect 15410 785 15468 819
rect 15410 751 15422 785
rect 15456 751 15468 785
rect 15410 717 15468 751
rect 15410 683 15422 717
rect 15456 683 15468 717
rect 15410 649 15468 683
rect 15410 615 15422 649
rect 15456 615 15468 649
rect 15410 581 15468 615
rect 15410 547 15422 581
rect 15456 547 15468 581
rect 15410 513 15468 547
rect 15410 479 15422 513
rect 15456 479 15468 513
rect 15410 445 15468 479
rect 15410 411 15422 445
rect 15456 411 15468 445
rect 15410 377 15468 411
rect 15410 343 15422 377
rect 15456 343 15468 377
rect 15410 309 15468 343
rect 15410 275 15422 309
rect 15456 275 15468 309
rect 15410 241 15468 275
rect 15410 207 15422 241
rect 15456 207 15468 241
rect 15410 173 15468 207
rect 15410 139 15422 173
rect 15456 139 15468 173
rect 15410 100 15468 139
rect 15498 1261 15556 1300
rect 15498 1227 15510 1261
rect 15544 1227 15556 1261
rect 15498 1193 15556 1227
rect 15498 1159 15510 1193
rect 15544 1159 15556 1193
rect 15498 1125 15556 1159
rect 15498 1091 15510 1125
rect 15544 1091 15556 1125
rect 15498 1057 15556 1091
rect 15498 1023 15510 1057
rect 15544 1023 15556 1057
rect 15498 989 15556 1023
rect 15498 955 15510 989
rect 15544 955 15556 989
rect 15498 921 15556 955
rect 15498 887 15510 921
rect 15544 887 15556 921
rect 15498 853 15556 887
rect 15498 819 15510 853
rect 15544 819 15556 853
rect 15498 785 15556 819
rect 15498 751 15510 785
rect 15544 751 15556 785
rect 15498 717 15556 751
rect 15498 683 15510 717
rect 15544 683 15556 717
rect 15498 649 15556 683
rect 15498 615 15510 649
rect 15544 615 15556 649
rect 15498 581 15556 615
rect 15498 547 15510 581
rect 15544 547 15556 581
rect 15498 513 15556 547
rect 15498 479 15510 513
rect 15544 479 15556 513
rect 15498 445 15556 479
rect 15498 411 15510 445
rect 15544 411 15556 445
rect 15498 377 15556 411
rect 15498 343 15510 377
rect 15544 343 15556 377
rect 15498 309 15556 343
rect 15498 275 15510 309
rect 15544 275 15556 309
rect 15498 241 15556 275
rect 15498 207 15510 241
rect 15544 207 15556 241
rect 15498 173 15556 207
rect 15498 139 15510 173
rect 15544 139 15556 173
rect 15498 100 15556 139
<< pdiff >>
rect 182 6565 244 6606
rect 182 6531 194 6565
rect 228 6531 244 6565
rect 182 6497 244 6531
rect 182 6463 194 6497
rect 228 6463 244 6497
rect 182 6429 244 6463
rect 182 6395 194 6429
rect 228 6395 244 6429
rect 182 6361 244 6395
rect 182 6327 194 6361
rect 228 6327 244 6361
rect 182 6293 244 6327
rect 182 6259 194 6293
rect 228 6259 244 6293
rect 182 6225 244 6259
rect 182 6191 194 6225
rect 228 6191 244 6225
rect 182 6157 244 6191
rect 182 6123 194 6157
rect 228 6123 244 6157
rect 182 6089 244 6123
rect 182 6055 194 6089
rect 228 6055 244 6089
rect 182 6021 244 6055
rect 182 5987 194 6021
rect 228 5987 244 6021
rect 182 5953 244 5987
rect -1664 5895 -1606 5936
rect -1664 5861 -1652 5895
rect -1618 5861 -1606 5895
rect -1664 5827 -1606 5861
rect -1664 5793 -1652 5827
rect -1618 5793 -1606 5827
rect -1664 5759 -1606 5793
rect -1664 5725 -1652 5759
rect -1618 5725 -1606 5759
rect -1664 5691 -1606 5725
rect -1664 5657 -1652 5691
rect -1618 5657 -1606 5691
rect -1664 5623 -1606 5657
rect -1664 5589 -1652 5623
rect -1618 5589 -1606 5623
rect -1664 5555 -1606 5589
rect -1664 5521 -1652 5555
rect -1618 5521 -1606 5555
rect -1664 5487 -1606 5521
rect -1664 5453 -1652 5487
rect -1618 5453 -1606 5487
rect -1664 5419 -1606 5453
rect -1664 5385 -1652 5419
rect -1618 5385 -1606 5419
rect -1664 5351 -1606 5385
rect -1664 5317 -1652 5351
rect -1618 5317 -1606 5351
rect -1664 5283 -1606 5317
rect -1664 5249 -1652 5283
rect -1618 5249 -1606 5283
rect -1664 5215 -1606 5249
rect -1664 5181 -1652 5215
rect -1618 5181 -1606 5215
rect -1664 5147 -1606 5181
rect -1664 5113 -1652 5147
rect -1618 5113 -1606 5147
rect -1664 5079 -1606 5113
rect -1664 5045 -1652 5079
rect -1618 5045 -1606 5079
rect -1664 5011 -1606 5045
rect -1664 4977 -1652 5011
rect -1618 4977 -1606 5011
rect -1664 4936 -1606 4977
rect -1566 5895 -1508 5936
rect -1566 5861 -1554 5895
rect -1520 5861 -1508 5895
rect -1566 5827 -1508 5861
rect -1566 5793 -1554 5827
rect -1520 5793 -1508 5827
rect -1566 5759 -1508 5793
rect -1566 5725 -1554 5759
rect -1520 5725 -1508 5759
rect -1566 5691 -1508 5725
rect -1566 5657 -1554 5691
rect -1520 5657 -1508 5691
rect -1566 5623 -1508 5657
rect -1566 5589 -1554 5623
rect -1520 5589 -1508 5623
rect -1566 5555 -1508 5589
rect -1566 5521 -1554 5555
rect -1520 5521 -1508 5555
rect -1566 5487 -1508 5521
rect -1566 5453 -1554 5487
rect -1520 5453 -1508 5487
rect -1566 5419 -1508 5453
rect -1566 5385 -1554 5419
rect -1520 5385 -1508 5419
rect -1566 5351 -1508 5385
rect -1566 5317 -1554 5351
rect -1520 5317 -1508 5351
rect -1566 5283 -1508 5317
rect -1566 5249 -1554 5283
rect -1520 5249 -1508 5283
rect -1566 5215 -1508 5249
rect -1566 5181 -1554 5215
rect -1520 5181 -1508 5215
rect -1566 5147 -1508 5181
rect -1566 5113 -1554 5147
rect -1520 5113 -1508 5147
rect -1566 5079 -1508 5113
rect -1566 5045 -1554 5079
rect -1520 5045 -1508 5079
rect -1566 5011 -1508 5045
rect -1566 4977 -1554 5011
rect -1520 4977 -1508 5011
rect -1566 4936 -1508 4977
rect -1468 5895 -1410 5936
rect -1468 5861 -1456 5895
rect -1422 5861 -1410 5895
rect -1468 5827 -1410 5861
rect -1468 5793 -1456 5827
rect -1422 5793 -1410 5827
rect -1468 5759 -1410 5793
rect -1468 5725 -1456 5759
rect -1422 5725 -1410 5759
rect -1468 5691 -1410 5725
rect -1468 5657 -1456 5691
rect -1422 5657 -1410 5691
rect -1468 5623 -1410 5657
rect -1468 5589 -1456 5623
rect -1422 5589 -1410 5623
rect -1468 5555 -1410 5589
rect -1468 5521 -1456 5555
rect -1422 5521 -1410 5555
rect -1468 5487 -1410 5521
rect -1468 5453 -1456 5487
rect -1422 5453 -1410 5487
rect -1468 5419 -1410 5453
rect -1468 5385 -1456 5419
rect -1422 5385 -1410 5419
rect -1468 5351 -1410 5385
rect -1468 5317 -1456 5351
rect -1422 5317 -1410 5351
rect -1468 5283 -1410 5317
rect -1468 5249 -1456 5283
rect -1422 5249 -1410 5283
rect -1468 5215 -1410 5249
rect -1468 5181 -1456 5215
rect -1422 5181 -1410 5215
rect -1468 5147 -1410 5181
rect -1468 5113 -1456 5147
rect -1422 5113 -1410 5147
rect -1468 5079 -1410 5113
rect -1468 5045 -1456 5079
rect -1422 5045 -1410 5079
rect -1468 5011 -1410 5045
rect -1468 4977 -1456 5011
rect -1422 4977 -1410 5011
rect -1468 4936 -1410 4977
rect -1370 5895 -1312 5936
rect -1370 5861 -1358 5895
rect -1324 5861 -1312 5895
rect -1370 5827 -1312 5861
rect -1370 5793 -1358 5827
rect -1324 5793 -1312 5827
rect -1370 5759 -1312 5793
rect -1370 5725 -1358 5759
rect -1324 5725 -1312 5759
rect -1370 5691 -1312 5725
rect -1370 5657 -1358 5691
rect -1324 5657 -1312 5691
rect -1370 5623 -1312 5657
rect -1370 5589 -1358 5623
rect -1324 5589 -1312 5623
rect -1370 5555 -1312 5589
rect -1370 5521 -1358 5555
rect -1324 5521 -1312 5555
rect -1370 5487 -1312 5521
rect -1370 5453 -1358 5487
rect -1324 5453 -1312 5487
rect -1370 5419 -1312 5453
rect -1370 5385 -1358 5419
rect -1324 5385 -1312 5419
rect -1370 5351 -1312 5385
rect -1370 5317 -1358 5351
rect -1324 5317 -1312 5351
rect -1370 5283 -1312 5317
rect -1370 5249 -1358 5283
rect -1324 5249 -1312 5283
rect -1370 5215 -1312 5249
rect -1370 5181 -1358 5215
rect -1324 5181 -1312 5215
rect -1370 5147 -1312 5181
rect -1370 5113 -1358 5147
rect -1324 5113 -1312 5147
rect -1370 5079 -1312 5113
rect -1370 5045 -1358 5079
rect -1324 5045 -1312 5079
rect -1370 5011 -1312 5045
rect -1370 4977 -1358 5011
rect -1324 4977 -1312 5011
rect -1370 4936 -1312 4977
rect -1272 5895 -1214 5936
rect -1272 5861 -1260 5895
rect -1226 5861 -1214 5895
rect -1272 5827 -1214 5861
rect -1272 5793 -1260 5827
rect -1226 5793 -1214 5827
rect -1272 5759 -1214 5793
rect -1272 5725 -1260 5759
rect -1226 5725 -1214 5759
rect -1272 5691 -1214 5725
rect -1272 5657 -1260 5691
rect -1226 5657 -1214 5691
rect -1272 5623 -1214 5657
rect -1272 5589 -1260 5623
rect -1226 5589 -1214 5623
rect -1272 5555 -1214 5589
rect -1272 5521 -1260 5555
rect -1226 5521 -1214 5555
rect -1272 5487 -1214 5521
rect -1272 5453 -1260 5487
rect -1226 5453 -1214 5487
rect -1272 5419 -1214 5453
rect -1272 5385 -1260 5419
rect -1226 5385 -1214 5419
rect -1272 5351 -1214 5385
rect -1272 5317 -1260 5351
rect -1226 5317 -1214 5351
rect -1272 5283 -1214 5317
rect -1272 5249 -1260 5283
rect -1226 5249 -1214 5283
rect -1272 5215 -1214 5249
rect -1272 5181 -1260 5215
rect -1226 5181 -1214 5215
rect -1272 5147 -1214 5181
rect -1272 5113 -1260 5147
rect -1226 5113 -1214 5147
rect -1272 5079 -1214 5113
rect -1272 5045 -1260 5079
rect -1226 5045 -1214 5079
rect -1272 5011 -1214 5045
rect -1272 4977 -1260 5011
rect -1226 4977 -1214 5011
rect -1272 4936 -1214 4977
rect -1174 5895 -1116 5936
rect -1174 5861 -1162 5895
rect -1128 5861 -1116 5895
rect -1174 5827 -1116 5861
rect -1174 5793 -1162 5827
rect -1128 5793 -1116 5827
rect -1174 5759 -1116 5793
rect -1174 5725 -1162 5759
rect -1128 5725 -1116 5759
rect -1174 5691 -1116 5725
rect -1174 5657 -1162 5691
rect -1128 5657 -1116 5691
rect -1174 5623 -1116 5657
rect -1174 5589 -1162 5623
rect -1128 5589 -1116 5623
rect -1174 5555 -1116 5589
rect -1174 5521 -1162 5555
rect -1128 5521 -1116 5555
rect -1174 5487 -1116 5521
rect -1174 5453 -1162 5487
rect -1128 5453 -1116 5487
rect -1174 5419 -1116 5453
rect -1174 5385 -1162 5419
rect -1128 5385 -1116 5419
rect -1174 5351 -1116 5385
rect -1174 5317 -1162 5351
rect -1128 5317 -1116 5351
rect -1174 5283 -1116 5317
rect -1174 5249 -1162 5283
rect -1128 5249 -1116 5283
rect -1174 5215 -1116 5249
rect -1174 5181 -1162 5215
rect -1128 5181 -1116 5215
rect -1174 5147 -1116 5181
rect -1174 5113 -1162 5147
rect -1128 5113 -1116 5147
rect -1174 5079 -1116 5113
rect -1174 5045 -1162 5079
rect -1128 5045 -1116 5079
rect -1174 5011 -1116 5045
rect -1174 4977 -1162 5011
rect -1128 4977 -1116 5011
rect -1174 4936 -1116 4977
rect -1076 5895 -1018 5936
rect -1076 5861 -1064 5895
rect -1030 5861 -1018 5895
rect -1076 5827 -1018 5861
rect -1076 5793 -1064 5827
rect -1030 5793 -1018 5827
rect -1076 5759 -1018 5793
rect -1076 5725 -1064 5759
rect -1030 5725 -1018 5759
rect -1076 5691 -1018 5725
rect -1076 5657 -1064 5691
rect -1030 5657 -1018 5691
rect -1076 5623 -1018 5657
rect -1076 5589 -1064 5623
rect -1030 5589 -1018 5623
rect -1076 5555 -1018 5589
rect -1076 5521 -1064 5555
rect -1030 5521 -1018 5555
rect -1076 5487 -1018 5521
rect -1076 5453 -1064 5487
rect -1030 5453 -1018 5487
rect -1076 5419 -1018 5453
rect -1076 5385 -1064 5419
rect -1030 5385 -1018 5419
rect -1076 5351 -1018 5385
rect -1076 5317 -1064 5351
rect -1030 5317 -1018 5351
rect -1076 5283 -1018 5317
rect -1076 5249 -1064 5283
rect -1030 5249 -1018 5283
rect -1076 5215 -1018 5249
rect -1076 5181 -1064 5215
rect -1030 5181 -1018 5215
rect -1076 5147 -1018 5181
rect -1076 5113 -1064 5147
rect -1030 5113 -1018 5147
rect -1076 5079 -1018 5113
rect -1076 5045 -1064 5079
rect -1030 5045 -1018 5079
rect -1076 5011 -1018 5045
rect -1076 4977 -1064 5011
rect -1030 4977 -1018 5011
rect -1076 4936 -1018 4977
rect -978 5895 -920 5936
rect -978 5861 -966 5895
rect -932 5861 -920 5895
rect -978 5827 -920 5861
rect -978 5793 -966 5827
rect -932 5793 -920 5827
rect -978 5759 -920 5793
rect -978 5725 -966 5759
rect -932 5725 -920 5759
rect -978 5691 -920 5725
rect -978 5657 -966 5691
rect -932 5657 -920 5691
rect -978 5623 -920 5657
rect -978 5589 -966 5623
rect -932 5589 -920 5623
rect -978 5555 -920 5589
rect -978 5521 -966 5555
rect -932 5521 -920 5555
rect -978 5487 -920 5521
rect -978 5453 -966 5487
rect -932 5453 -920 5487
rect -978 5419 -920 5453
rect -978 5385 -966 5419
rect -932 5385 -920 5419
rect -978 5351 -920 5385
rect -978 5317 -966 5351
rect -932 5317 -920 5351
rect -978 5283 -920 5317
rect -978 5249 -966 5283
rect -932 5249 -920 5283
rect -978 5215 -920 5249
rect -978 5181 -966 5215
rect -932 5181 -920 5215
rect -978 5147 -920 5181
rect -978 5113 -966 5147
rect -932 5113 -920 5147
rect -978 5079 -920 5113
rect -978 5045 -966 5079
rect -932 5045 -920 5079
rect -978 5011 -920 5045
rect -978 4977 -966 5011
rect -932 4977 -920 5011
rect -978 4936 -920 4977
rect -880 5895 -822 5936
rect -880 5861 -868 5895
rect -834 5861 -822 5895
rect -880 5827 -822 5861
rect -880 5793 -868 5827
rect -834 5793 -822 5827
rect -880 5759 -822 5793
rect -880 5725 -868 5759
rect -834 5725 -822 5759
rect -880 5691 -822 5725
rect -880 5657 -868 5691
rect -834 5657 -822 5691
rect -880 5623 -822 5657
rect -880 5589 -868 5623
rect -834 5589 -822 5623
rect 182 5919 194 5953
rect 228 5919 244 5953
rect 182 5885 244 5919
rect 182 5851 194 5885
rect 228 5851 244 5885
rect 182 5817 244 5851
rect 182 5783 194 5817
rect 228 5783 244 5817
rect 182 5749 244 5783
rect 182 5715 194 5749
rect 228 5715 244 5749
rect 182 5681 244 5715
rect 182 5647 194 5681
rect 228 5647 244 5681
rect 182 5606 244 5647
rect 274 6565 340 6606
rect 274 6531 290 6565
rect 324 6531 340 6565
rect 274 6497 340 6531
rect 274 6463 290 6497
rect 324 6463 340 6497
rect 274 6429 340 6463
rect 274 6395 290 6429
rect 324 6395 340 6429
rect 274 6361 340 6395
rect 274 6327 290 6361
rect 324 6327 340 6361
rect 274 6293 340 6327
rect 274 6259 290 6293
rect 324 6259 340 6293
rect 274 6225 340 6259
rect 274 6191 290 6225
rect 324 6191 340 6225
rect 274 6157 340 6191
rect 274 6123 290 6157
rect 324 6123 340 6157
rect 274 6089 340 6123
rect 274 6055 290 6089
rect 324 6055 340 6089
rect 274 6021 340 6055
rect 274 5987 290 6021
rect 324 5987 340 6021
rect 274 5953 340 5987
rect 274 5919 290 5953
rect 324 5919 340 5953
rect 274 5885 340 5919
rect 274 5851 290 5885
rect 324 5851 340 5885
rect 274 5817 340 5851
rect 274 5783 290 5817
rect 324 5783 340 5817
rect 274 5749 340 5783
rect 274 5715 290 5749
rect 324 5715 340 5749
rect 274 5681 340 5715
rect 274 5647 290 5681
rect 324 5647 340 5681
rect 274 5606 340 5647
rect 370 6565 436 6606
rect 370 6531 386 6565
rect 420 6531 436 6565
rect 370 6497 436 6531
rect 370 6463 386 6497
rect 420 6463 436 6497
rect 370 6429 436 6463
rect 370 6395 386 6429
rect 420 6395 436 6429
rect 370 6361 436 6395
rect 370 6327 386 6361
rect 420 6327 436 6361
rect 370 6293 436 6327
rect 370 6259 386 6293
rect 420 6259 436 6293
rect 370 6225 436 6259
rect 370 6191 386 6225
rect 420 6191 436 6225
rect 370 6157 436 6191
rect 370 6123 386 6157
rect 420 6123 436 6157
rect 370 6089 436 6123
rect 370 6055 386 6089
rect 420 6055 436 6089
rect 370 6021 436 6055
rect 370 5987 386 6021
rect 420 5987 436 6021
rect 370 5953 436 5987
rect 370 5919 386 5953
rect 420 5919 436 5953
rect 370 5885 436 5919
rect 370 5851 386 5885
rect 420 5851 436 5885
rect 370 5817 436 5851
rect 370 5783 386 5817
rect 420 5783 436 5817
rect 370 5749 436 5783
rect 370 5715 386 5749
rect 420 5715 436 5749
rect 370 5681 436 5715
rect 370 5647 386 5681
rect 420 5647 436 5681
rect 370 5606 436 5647
rect 466 6565 532 6606
rect 466 6531 482 6565
rect 516 6531 532 6565
rect 466 6497 532 6531
rect 466 6463 482 6497
rect 516 6463 532 6497
rect 466 6429 532 6463
rect 466 6395 482 6429
rect 516 6395 532 6429
rect 466 6361 532 6395
rect 466 6327 482 6361
rect 516 6327 532 6361
rect 466 6293 532 6327
rect 466 6259 482 6293
rect 516 6259 532 6293
rect 466 6225 532 6259
rect 466 6191 482 6225
rect 516 6191 532 6225
rect 466 6157 532 6191
rect 466 6123 482 6157
rect 516 6123 532 6157
rect 466 6089 532 6123
rect 466 6055 482 6089
rect 516 6055 532 6089
rect 466 6021 532 6055
rect 466 5987 482 6021
rect 516 5987 532 6021
rect 466 5953 532 5987
rect 466 5919 482 5953
rect 516 5919 532 5953
rect 466 5885 532 5919
rect 466 5851 482 5885
rect 516 5851 532 5885
rect 466 5817 532 5851
rect 466 5783 482 5817
rect 516 5783 532 5817
rect 466 5749 532 5783
rect 466 5715 482 5749
rect 516 5715 532 5749
rect 466 5681 532 5715
rect 466 5647 482 5681
rect 516 5647 532 5681
rect 466 5606 532 5647
rect 562 6565 628 6606
rect 562 6531 578 6565
rect 612 6531 628 6565
rect 562 6497 628 6531
rect 562 6463 578 6497
rect 612 6463 628 6497
rect 562 6429 628 6463
rect 562 6395 578 6429
rect 612 6395 628 6429
rect 562 6361 628 6395
rect 562 6327 578 6361
rect 612 6327 628 6361
rect 562 6293 628 6327
rect 562 6259 578 6293
rect 612 6259 628 6293
rect 562 6225 628 6259
rect 562 6191 578 6225
rect 612 6191 628 6225
rect 562 6157 628 6191
rect 562 6123 578 6157
rect 612 6123 628 6157
rect 562 6089 628 6123
rect 562 6055 578 6089
rect 612 6055 628 6089
rect 562 6021 628 6055
rect 562 5987 578 6021
rect 612 5987 628 6021
rect 562 5953 628 5987
rect 562 5919 578 5953
rect 612 5919 628 5953
rect 562 5885 628 5919
rect 562 5851 578 5885
rect 612 5851 628 5885
rect 562 5817 628 5851
rect 562 5783 578 5817
rect 612 5783 628 5817
rect 562 5749 628 5783
rect 562 5715 578 5749
rect 612 5715 628 5749
rect 562 5681 628 5715
rect 562 5647 578 5681
rect 612 5647 628 5681
rect 562 5606 628 5647
rect 658 6565 724 6606
rect 658 6531 674 6565
rect 708 6531 724 6565
rect 658 6497 724 6531
rect 658 6463 674 6497
rect 708 6463 724 6497
rect 658 6429 724 6463
rect 658 6395 674 6429
rect 708 6395 724 6429
rect 658 6361 724 6395
rect 658 6327 674 6361
rect 708 6327 724 6361
rect 658 6293 724 6327
rect 658 6259 674 6293
rect 708 6259 724 6293
rect 658 6225 724 6259
rect 658 6191 674 6225
rect 708 6191 724 6225
rect 658 6157 724 6191
rect 658 6123 674 6157
rect 708 6123 724 6157
rect 658 6089 724 6123
rect 658 6055 674 6089
rect 708 6055 724 6089
rect 658 6021 724 6055
rect 658 5987 674 6021
rect 708 5987 724 6021
rect 658 5953 724 5987
rect 658 5919 674 5953
rect 708 5919 724 5953
rect 658 5885 724 5919
rect 658 5851 674 5885
rect 708 5851 724 5885
rect 658 5817 724 5851
rect 658 5783 674 5817
rect 708 5783 724 5817
rect 658 5749 724 5783
rect 658 5715 674 5749
rect 708 5715 724 5749
rect 658 5681 724 5715
rect 658 5647 674 5681
rect 708 5647 724 5681
rect 658 5606 724 5647
rect 754 6565 820 6606
rect 754 6531 770 6565
rect 804 6531 820 6565
rect 754 6497 820 6531
rect 754 6463 770 6497
rect 804 6463 820 6497
rect 754 6429 820 6463
rect 754 6395 770 6429
rect 804 6395 820 6429
rect 754 6361 820 6395
rect 754 6327 770 6361
rect 804 6327 820 6361
rect 754 6293 820 6327
rect 754 6259 770 6293
rect 804 6259 820 6293
rect 754 6225 820 6259
rect 754 6191 770 6225
rect 804 6191 820 6225
rect 754 6157 820 6191
rect 754 6123 770 6157
rect 804 6123 820 6157
rect 754 6089 820 6123
rect 754 6055 770 6089
rect 804 6055 820 6089
rect 754 6021 820 6055
rect 754 5987 770 6021
rect 804 5987 820 6021
rect 754 5953 820 5987
rect 754 5919 770 5953
rect 804 5919 820 5953
rect 754 5885 820 5919
rect 754 5851 770 5885
rect 804 5851 820 5885
rect 754 5817 820 5851
rect 754 5783 770 5817
rect 804 5783 820 5817
rect 754 5749 820 5783
rect 754 5715 770 5749
rect 804 5715 820 5749
rect 754 5681 820 5715
rect 754 5647 770 5681
rect 804 5647 820 5681
rect 754 5606 820 5647
rect 850 6565 916 6606
rect 850 6531 866 6565
rect 900 6531 916 6565
rect 850 6497 916 6531
rect 850 6463 866 6497
rect 900 6463 916 6497
rect 850 6429 916 6463
rect 850 6395 866 6429
rect 900 6395 916 6429
rect 850 6361 916 6395
rect 850 6327 866 6361
rect 900 6327 916 6361
rect 850 6293 916 6327
rect 850 6259 866 6293
rect 900 6259 916 6293
rect 850 6225 916 6259
rect 850 6191 866 6225
rect 900 6191 916 6225
rect 850 6157 916 6191
rect 850 6123 866 6157
rect 900 6123 916 6157
rect 850 6089 916 6123
rect 850 6055 866 6089
rect 900 6055 916 6089
rect 850 6021 916 6055
rect 850 5987 866 6021
rect 900 5987 916 6021
rect 850 5953 916 5987
rect 850 5919 866 5953
rect 900 5919 916 5953
rect 850 5885 916 5919
rect 850 5851 866 5885
rect 900 5851 916 5885
rect 850 5817 916 5851
rect 850 5783 866 5817
rect 900 5783 916 5817
rect 850 5749 916 5783
rect 850 5715 866 5749
rect 900 5715 916 5749
rect 850 5681 916 5715
rect 850 5647 866 5681
rect 900 5647 916 5681
rect 850 5606 916 5647
rect 946 6565 1012 6606
rect 946 6531 962 6565
rect 996 6531 1012 6565
rect 946 6497 1012 6531
rect 946 6463 962 6497
rect 996 6463 1012 6497
rect 946 6429 1012 6463
rect 946 6395 962 6429
rect 996 6395 1012 6429
rect 946 6361 1012 6395
rect 946 6327 962 6361
rect 996 6327 1012 6361
rect 946 6293 1012 6327
rect 946 6259 962 6293
rect 996 6259 1012 6293
rect 946 6225 1012 6259
rect 946 6191 962 6225
rect 996 6191 1012 6225
rect 946 6157 1012 6191
rect 946 6123 962 6157
rect 996 6123 1012 6157
rect 946 6089 1012 6123
rect 946 6055 962 6089
rect 996 6055 1012 6089
rect 946 6021 1012 6055
rect 946 5987 962 6021
rect 996 5987 1012 6021
rect 946 5953 1012 5987
rect 946 5919 962 5953
rect 996 5919 1012 5953
rect 946 5885 1012 5919
rect 946 5851 962 5885
rect 996 5851 1012 5885
rect 946 5817 1012 5851
rect 946 5783 962 5817
rect 996 5783 1012 5817
rect 946 5749 1012 5783
rect 946 5715 962 5749
rect 996 5715 1012 5749
rect 946 5681 1012 5715
rect 946 5647 962 5681
rect 996 5647 1012 5681
rect 946 5606 1012 5647
rect 1042 6565 1108 6606
rect 1042 6531 1058 6565
rect 1092 6531 1108 6565
rect 1042 6497 1108 6531
rect 1042 6463 1058 6497
rect 1092 6463 1108 6497
rect 1042 6429 1108 6463
rect 1042 6395 1058 6429
rect 1092 6395 1108 6429
rect 1042 6361 1108 6395
rect 1042 6327 1058 6361
rect 1092 6327 1108 6361
rect 1042 6293 1108 6327
rect 1042 6259 1058 6293
rect 1092 6259 1108 6293
rect 1042 6225 1108 6259
rect 1042 6191 1058 6225
rect 1092 6191 1108 6225
rect 1042 6157 1108 6191
rect 1042 6123 1058 6157
rect 1092 6123 1108 6157
rect 1042 6089 1108 6123
rect 1042 6055 1058 6089
rect 1092 6055 1108 6089
rect 1042 6021 1108 6055
rect 1042 5987 1058 6021
rect 1092 5987 1108 6021
rect 1042 5953 1108 5987
rect 1042 5919 1058 5953
rect 1092 5919 1108 5953
rect 1042 5885 1108 5919
rect 1042 5851 1058 5885
rect 1092 5851 1108 5885
rect 1042 5817 1108 5851
rect 1042 5783 1058 5817
rect 1092 5783 1108 5817
rect 1042 5749 1108 5783
rect 1042 5715 1058 5749
rect 1092 5715 1108 5749
rect 1042 5681 1108 5715
rect 1042 5647 1058 5681
rect 1092 5647 1108 5681
rect 1042 5606 1108 5647
rect 1138 6565 1204 6606
rect 1138 6531 1154 6565
rect 1188 6531 1204 6565
rect 1138 6497 1204 6531
rect 1138 6463 1154 6497
rect 1188 6463 1204 6497
rect 1138 6429 1204 6463
rect 1138 6395 1154 6429
rect 1188 6395 1204 6429
rect 1138 6361 1204 6395
rect 1138 6327 1154 6361
rect 1188 6327 1204 6361
rect 1138 6293 1204 6327
rect 1138 6259 1154 6293
rect 1188 6259 1204 6293
rect 1138 6225 1204 6259
rect 1138 6191 1154 6225
rect 1188 6191 1204 6225
rect 1138 6157 1204 6191
rect 1138 6123 1154 6157
rect 1188 6123 1204 6157
rect 1138 6089 1204 6123
rect 1138 6055 1154 6089
rect 1188 6055 1204 6089
rect 1138 6021 1204 6055
rect 1138 5987 1154 6021
rect 1188 5987 1204 6021
rect 1138 5953 1204 5987
rect 1138 5919 1154 5953
rect 1188 5919 1204 5953
rect 1138 5885 1204 5919
rect 1138 5851 1154 5885
rect 1188 5851 1204 5885
rect 1138 5817 1204 5851
rect 1138 5783 1154 5817
rect 1188 5783 1204 5817
rect 1138 5749 1204 5783
rect 1138 5715 1154 5749
rect 1188 5715 1204 5749
rect 1138 5681 1204 5715
rect 1138 5647 1154 5681
rect 1188 5647 1204 5681
rect 1138 5606 1204 5647
rect 1234 6565 1300 6606
rect 1234 6531 1250 6565
rect 1284 6531 1300 6565
rect 1234 6497 1300 6531
rect 1234 6463 1250 6497
rect 1284 6463 1300 6497
rect 1234 6429 1300 6463
rect 1234 6395 1250 6429
rect 1284 6395 1300 6429
rect 1234 6361 1300 6395
rect 1234 6327 1250 6361
rect 1284 6327 1300 6361
rect 1234 6293 1300 6327
rect 1234 6259 1250 6293
rect 1284 6259 1300 6293
rect 1234 6225 1300 6259
rect 1234 6191 1250 6225
rect 1284 6191 1300 6225
rect 1234 6157 1300 6191
rect 1234 6123 1250 6157
rect 1284 6123 1300 6157
rect 1234 6089 1300 6123
rect 1234 6055 1250 6089
rect 1284 6055 1300 6089
rect 1234 6021 1300 6055
rect 1234 5987 1250 6021
rect 1284 5987 1300 6021
rect 1234 5953 1300 5987
rect 1234 5919 1250 5953
rect 1284 5919 1300 5953
rect 1234 5885 1300 5919
rect 1234 5851 1250 5885
rect 1284 5851 1300 5885
rect 1234 5817 1300 5851
rect 1234 5783 1250 5817
rect 1284 5783 1300 5817
rect 1234 5749 1300 5783
rect 1234 5715 1250 5749
rect 1284 5715 1300 5749
rect 1234 5681 1300 5715
rect 1234 5647 1250 5681
rect 1284 5647 1300 5681
rect 1234 5606 1300 5647
rect 1330 6565 1392 6606
rect 1330 6531 1346 6565
rect 1380 6531 1392 6565
rect 1330 6497 1392 6531
rect 1330 6463 1346 6497
rect 1380 6463 1392 6497
rect 1330 6429 1392 6463
rect 1330 6395 1346 6429
rect 1380 6395 1392 6429
rect 1330 6361 1392 6395
rect 1330 6327 1346 6361
rect 1380 6327 1392 6361
rect 1330 6293 1392 6327
rect 1330 6259 1346 6293
rect 1380 6259 1392 6293
rect 1330 6225 1392 6259
rect 1330 6191 1346 6225
rect 1380 6191 1392 6225
rect 1330 6157 1392 6191
rect 1330 6123 1346 6157
rect 1380 6123 1392 6157
rect 1330 6089 1392 6123
rect 1330 6055 1346 6089
rect 1380 6055 1392 6089
rect 1330 6021 1392 6055
rect 1330 5987 1346 6021
rect 1380 5987 1392 6021
rect 1330 5953 1392 5987
rect 1330 5919 1346 5953
rect 1380 5919 1392 5953
rect 1330 5885 1392 5919
rect 1330 5851 1346 5885
rect 1380 5851 1392 5885
rect 1330 5817 1392 5851
rect 1330 5783 1346 5817
rect 1380 5783 1392 5817
rect 1330 5749 1392 5783
rect 1330 5715 1346 5749
rect 1380 5715 1392 5749
rect 1330 5681 1392 5715
rect 1330 5647 1346 5681
rect 1380 5647 1392 5681
rect 1330 5606 1392 5647
rect 1948 6561 2010 6602
rect 1948 6527 1960 6561
rect 1994 6527 2010 6561
rect 1948 6493 2010 6527
rect 1948 6459 1960 6493
rect 1994 6459 2010 6493
rect 1948 6425 2010 6459
rect 1948 6391 1960 6425
rect 1994 6391 2010 6425
rect 1948 6357 2010 6391
rect 1948 6323 1960 6357
rect 1994 6323 2010 6357
rect 1948 6289 2010 6323
rect 1948 6255 1960 6289
rect 1994 6255 2010 6289
rect 1948 6221 2010 6255
rect 1948 6187 1960 6221
rect 1994 6187 2010 6221
rect 1948 6153 2010 6187
rect 1948 6119 1960 6153
rect 1994 6119 2010 6153
rect 1948 6085 2010 6119
rect 1948 6051 1960 6085
rect 1994 6051 2010 6085
rect 1948 6017 2010 6051
rect 1948 5983 1960 6017
rect 1994 5983 2010 6017
rect 1948 5949 2010 5983
rect 1948 5915 1960 5949
rect 1994 5915 2010 5949
rect 1948 5881 2010 5915
rect 1948 5847 1960 5881
rect 1994 5847 2010 5881
rect 1948 5813 2010 5847
rect 1948 5779 1960 5813
rect 1994 5779 2010 5813
rect 1948 5745 2010 5779
rect 1948 5711 1960 5745
rect 1994 5711 2010 5745
rect 1948 5677 2010 5711
rect 1948 5643 1960 5677
rect 1994 5643 2010 5677
rect -880 5555 -822 5589
rect 1948 5602 2010 5643
rect 2040 6561 2106 6602
rect 2040 6527 2056 6561
rect 2090 6527 2106 6561
rect 2040 6493 2106 6527
rect 2040 6459 2056 6493
rect 2090 6459 2106 6493
rect 2040 6425 2106 6459
rect 2040 6391 2056 6425
rect 2090 6391 2106 6425
rect 2040 6357 2106 6391
rect 2040 6323 2056 6357
rect 2090 6323 2106 6357
rect 2040 6289 2106 6323
rect 2040 6255 2056 6289
rect 2090 6255 2106 6289
rect 2040 6221 2106 6255
rect 2040 6187 2056 6221
rect 2090 6187 2106 6221
rect 2040 6153 2106 6187
rect 2040 6119 2056 6153
rect 2090 6119 2106 6153
rect 2040 6085 2106 6119
rect 2040 6051 2056 6085
rect 2090 6051 2106 6085
rect 2040 6017 2106 6051
rect 2040 5983 2056 6017
rect 2090 5983 2106 6017
rect 2040 5949 2106 5983
rect 2040 5915 2056 5949
rect 2090 5915 2106 5949
rect 2040 5881 2106 5915
rect 2040 5847 2056 5881
rect 2090 5847 2106 5881
rect 2040 5813 2106 5847
rect 2040 5779 2056 5813
rect 2090 5779 2106 5813
rect 2040 5745 2106 5779
rect 2040 5711 2056 5745
rect 2090 5711 2106 5745
rect 2040 5677 2106 5711
rect 2040 5643 2056 5677
rect 2090 5643 2106 5677
rect 2040 5602 2106 5643
rect 2136 6561 2202 6602
rect 2136 6527 2152 6561
rect 2186 6527 2202 6561
rect 2136 6493 2202 6527
rect 2136 6459 2152 6493
rect 2186 6459 2202 6493
rect 2136 6425 2202 6459
rect 2136 6391 2152 6425
rect 2186 6391 2202 6425
rect 2136 6357 2202 6391
rect 2136 6323 2152 6357
rect 2186 6323 2202 6357
rect 2136 6289 2202 6323
rect 2136 6255 2152 6289
rect 2186 6255 2202 6289
rect 2136 6221 2202 6255
rect 2136 6187 2152 6221
rect 2186 6187 2202 6221
rect 2136 6153 2202 6187
rect 2136 6119 2152 6153
rect 2186 6119 2202 6153
rect 2136 6085 2202 6119
rect 2136 6051 2152 6085
rect 2186 6051 2202 6085
rect 2136 6017 2202 6051
rect 2136 5983 2152 6017
rect 2186 5983 2202 6017
rect 2136 5949 2202 5983
rect 2136 5915 2152 5949
rect 2186 5915 2202 5949
rect 2136 5881 2202 5915
rect 2136 5847 2152 5881
rect 2186 5847 2202 5881
rect 2136 5813 2202 5847
rect 2136 5779 2152 5813
rect 2186 5779 2202 5813
rect 2136 5745 2202 5779
rect 2136 5711 2152 5745
rect 2186 5711 2202 5745
rect 2136 5677 2202 5711
rect 2136 5643 2152 5677
rect 2186 5643 2202 5677
rect 2136 5602 2202 5643
rect 2232 6561 2298 6602
rect 2232 6527 2248 6561
rect 2282 6527 2298 6561
rect 2232 6493 2298 6527
rect 2232 6459 2248 6493
rect 2282 6459 2298 6493
rect 2232 6425 2298 6459
rect 2232 6391 2248 6425
rect 2282 6391 2298 6425
rect 2232 6357 2298 6391
rect 2232 6323 2248 6357
rect 2282 6323 2298 6357
rect 2232 6289 2298 6323
rect 2232 6255 2248 6289
rect 2282 6255 2298 6289
rect 2232 6221 2298 6255
rect 2232 6187 2248 6221
rect 2282 6187 2298 6221
rect 2232 6153 2298 6187
rect 2232 6119 2248 6153
rect 2282 6119 2298 6153
rect 2232 6085 2298 6119
rect 2232 6051 2248 6085
rect 2282 6051 2298 6085
rect 2232 6017 2298 6051
rect 2232 5983 2248 6017
rect 2282 5983 2298 6017
rect 2232 5949 2298 5983
rect 2232 5915 2248 5949
rect 2282 5915 2298 5949
rect 2232 5881 2298 5915
rect 2232 5847 2248 5881
rect 2282 5847 2298 5881
rect 2232 5813 2298 5847
rect 2232 5779 2248 5813
rect 2282 5779 2298 5813
rect 2232 5745 2298 5779
rect 2232 5711 2248 5745
rect 2282 5711 2298 5745
rect 2232 5677 2298 5711
rect 2232 5643 2248 5677
rect 2282 5643 2298 5677
rect 2232 5602 2298 5643
rect 2328 6561 2394 6602
rect 2328 6527 2344 6561
rect 2378 6527 2394 6561
rect 2328 6493 2394 6527
rect 2328 6459 2344 6493
rect 2378 6459 2394 6493
rect 2328 6425 2394 6459
rect 2328 6391 2344 6425
rect 2378 6391 2394 6425
rect 2328 6357 2394 6391
rect 2328 6323 2344 6357
rect 2378 6323 2394 6357
rect 2328 6289 2394 6323
rect 2328 6255 2344 6289
rect 2378 6255 2394 6289
rect 2328 6221 2394 6255
rect 2328 6187 2344 6221
rect 2378 6187 2394 6221
rect 2328 6153 2394 6187
rect 2328 6119 2344 6153
rect 2378 6119 2394 6153
rect 2328 6085 2394 6119
rect 2328 6051 2344 6085
rect 2378 6051 2394 6085
rect 2328 6017 2394 6051
rect 2328 5983 2344 6017
rect 2378 5983 2394 6017
rect 2328 5949 2394 5983
rect 2328 5915 2344 5949
rect 2378 5915 2394 5949
rect 2328 5881 2394 5915
rect 2328 5847 2344 5881
rect 2378 5847 2394 5881
rect 2328 5813 2394 5847
rect 2328 5779 2344 5813
rect 2378 5779 2394 5813
rect 2328 5745 2394 5779
rect 2328 5711 2344 5745
rect 2378 5711 2394 5745
rect 2328 5677 2394 5711
rect 2328 5643 2344 5677
rect 2378 5643 2394 5677
rect 2328 5602 2394 5643
rect 2424 6561 2490 6602
rect 2424 6527 2440 6561
rect 2474 6527 2490 6561
rect 2424 6493 2490 6527
rect 2424 6459 2440 6493
rect 2474 6459 2490 6493
rect 2424 6425 2490 6459
rect 2424 6391 2440 6425
rect 2474 6391 2490 6425
rect 2424 6357 2490 6391
rect 2424 6323 2440 6357
rect 2474 6323 2490 6357
rect 2424 6289 2490 6323
rect 2424 6255 2440 6289
rect 2474 6255 2490 6289
rect 2424 6221 2490 6255
rect 2424 6187 2440 6221
rect 2474 6187 2490 6221
rect 2424 6153 2490 6187
rect 2424 6119 2440 6153
rect 2474 6119 2490 6153
rect 2424 6085 2490 6119
rect 2424 6051 2440 6085
rect 2474 6051 2490 6085
rect 2424 6017 2490 6051
rect 2424 5983 2440 6017
rect 2474 5983 2490 6017
rect 2424 5949 2490 5983
rect 2424 5915 2440 5949
rect 2474 5915 2490 5949
rect 2424 5881 2490 5915
rect 2424 5847 2440 5881
rect 2474 5847 2490 5881
rect 2424 5813 2490 5847
rect 2424 5779 2440 5813
rect 2474 5779 2490 5813
rect 2424 5745 2490 5779
rect 2424 5711 2440 5745
rect 2474 5711 2490 5745
rect 2424 5677 2490 5711
rect 2424 5643 2440 5677
rect 2474 5643 2490 5677
rect 2424 5602 2490 5643
rect 2520 6561 2586 6602
rect 2520 6527 2536 6561
rect 2570 6527 2586 6561
rect 2520 6493 2586 6527
rect 2520 6459 2536 6493
rect 2570 6459 2586 6493
rect 2520 6425 2586 6459
rect 2520 6391 2536 6425
rect 2570 6391 2586 6425
rect 2520 6357 2586 6391
rect 2520 6323 2536 6357
rect 2570 6323 2586 6357
rect 2520 6289 2586 6323
rect 2520 6255 2536 6289
rect 2570 6255 2586 6289
rect 2520 6221 2586 6255
rect 2520 6187 2536 6221
rect 2570 6187 2586 6221
rect 2520 6153 2586 6187
rect 2520 6119 2536 6153
rect 2570 6119 2586 6153
rect 2520 6085 2586 6119
rect 2520 6051 2536 6085
rect 2570 6051 2586 6085
rect 2520 6017 2586 6051
rect 2520 5983 2536 6017
rect 2570 5983 2586 6017
rect 2520 5949 2586 5983
rect 2520 5915 2536 5949
rect 2570 5915 2586 5949
rect 2520 5881 2586 5915
rect 2520 5847 2536 5881
rect 2570 5847 2586 5881
rect 2520 5813 2586 5847
rect 2520 5779 2536 5813
rect 2570 5779 2586 5813
rect 2520 5745 2586 5779
rect 2520 5711 2536 5745
rect 2570 5711 2586 5745
rect 2520 5677 2586 5711
rect 2520 5643 2536 5677
rect 2570 5643 2586 5677
rect 2520 5602 2586 5643
rect 2616 6561 2682 6602
rect 2616 6527 2632 6561
rect 2666 6527 2682 6561
rect 2616 6493 2682 6527
rect 2616 6459 2632 6493
rect 2666 6459 2682 6493
rect 2616 6425 2682 6459
rect 2616 6391 2632 6425
rect 2666 6391 2682 6425
rect 2616 6357 2682 6391
rect 2616 6323 2632 6357
rect 2666 6323 2682 6357
rect 2616 6289 2682 6323
rect 2616 6255 2632 6289
rect 2666 6255 2682 6289
rect 2616 6221 2682 6255
rect 2616 6187 2632 6221
rect 2666 6187 2682 6221
rect 2616 6153 2682 6187
rect 2616 6119 2632 6153
rect 2666 6119 2682 6153
rect 2616 6085 2682 6119
rect 2616 6051 2632 6085
rect 2666 6051 2682 6085
rect 2616 6017 2682 6051
rect 2616 5983 2632 6017
rect 2666 5983 2682 6017
rect 2616 5949 2682 5983
rect 2616 5915 2632 5949
rect 2666 5915 2682 5949
rect 2616 5881 2682 5915
rect 2616 5847 2632 5881
rect 2666 5847 2682 5881
rect 2616 5813 2682 5847
rect 2616 5779 2632 5813
rect 2666 5779 2682 5813
rect 2616 5745 2682 5779
rect 2616 5711 2632 5745
rect 2666 5711 2682 5745
rect 2616 5677 2682 5711
rect 2616 5643 2632 5677
rect 2666 5643 2682 5677
rect 2616 5602 2682 5643
rect 2712 6561 2774 6602
rect 2712 6527 2728 6561
rect 2762 6527 2774 6561
rect 2712 6493 2774 6527
rect 2712 6459 2728 6493
rect 2762 6459 2774 6493
rect 2712 6425 2774 6459
rect 2712 6391 2728 6425
rect 2762 6391 2774 6425
rect 2712 6357 2774 6391
rect 2712 6323 2728 6357
rect 2762 6323 2774 6357
rect 2712 6289 2774 6323
rect 2712 6255 2728 6289
rect 2762 6255 2774 6289
rect 2712 6221 2774 6255
rect 2712 6187 2728 6221
rect 2762 6187 2774 6221
rect 2712 6153 2774 6187
rect 2712 6119 2728 6153
rect 2762 6119 2774 6153
rect 2712 6085 2774 6119
rect 2712 6051 2728 6085
rect 2762 6051 2774 6085
rect 2712 6017 2774 6051
rect 2712 5983 2728 6017
rect 2762 5983 2774 6017
rect 2712 5949 2774 5983
rect 2712 5915 2728 5949
rect 2762 5915 2774 5949
rect 2712 5881 2774 5915
rect 2712 5847 2728 5881
rect 2762 5847 2774 5881
rect 2712 5813 2774 5847
rect 2712 5779 2728 5813
rect 2762 5779 2774 5813
rect 2712 5745 2774 5779
rect 2712 5711 2728 5745
rect 2762 5711 2774 5745
rect 2712 5677 2774 5711
rect 2712 5643 2728 5677
rect 2762 5643 2774 5677
rect 2712 5602 2774 5643
rect 3138 6549 3200 6590
rect 3138 6515 3150 6549
rect 3184 6515 3200 6549
rect 3138 6481 3200 6515
rect 3138 6447 3150 6481
rect 3184 6447 3200 6481
rect 3138 6413 3200 6447
rect 3138 6379 3150 6413
rect 3184 6379 3200 6413
rect 3138 6345 3200 6379
rect 3138 6311 3150 6345
rect 3184 6311 3200 6345
rect 3138 6277 3200 6311
rect 3138 6243 3150 6277
rect 3184 6243 3200 6277
rect 3138 6209 3200 6243
rect 3138 6175 3150 6209
rect 3184 6175 3200 6209
rect 3138 6141 3200 6175
rect 3138 6107 3150 6141
rect 3184 6107 3200 6141
rect 3138 6073 3200 6107
rect 3138 6039 3150 6073
rect 3184 6039 3200 6073
rect 3138 6005 3200 6039
rect 3138 5971 3150 6005
rect 3184 5971 3200 6005
rect 3138 5937 3200 5971
rect 3138 5903 3150 5937
rect 3184 5903 3200 5937
rect 3138 5869 3200 5903
rect 3138 5835 3150 5869
rect 3184 5835 3200 5869
rect 3138 5801 3200 5835
rect 3138 5767 3150 5801
rect 3184 5767 3200 5801
rect 3138 5733 3200 5767
rect 3138 5699 3150 5733
rect 3184 5699 3200 5733
rect 3138 5665 3200 5699
rect 3138 5631 3150 5665
rect 3184 5631 3200 5665
rect 3138 5590 3200 5631
rect 3230 6549 3296 6590
rect 3230 6515 3246 6549
rect 3280 6515 3296 6549
rect 3230 6481 3296 6515
rect 3230 6447 3246 6481
rect 3280 6447 3296 6481
rect 3230 6413 3296 6447
rect 3230 6379 3246 6413
rect 3280 6379 3296 6413
rect 3230 6345 3296 6379
rect 3230 6311 3246 6345
rect 3280 6311 3296 6345
rect 3230 6277 3296 6311
rect 3230 6243 3246 6277
rect 3280 6243 3296 6277
rect 3230 6209 3296 6243
rect 3230 6175 3246 6209
rect 3280 6175 3296 6209
rect 3230 6141 3296 6175
rect 3230 6107 3246 6141
rect 3280 6107 3296 6141
rect 3230 6073 3296 6107
rect 3230 6039 3246 6073
rect 3280 6039 3296 6073
rect 3230 6005 3296 6039
rect 3230 5971 3246 6005
rect 3280 5971 3296 6005
rect 3230 5937 3296 5971
rect 3230 5903 3246 5937
rect 3280 5903 3296 5937
rect 3230 5869 3296 5903
rect 3230 5835 3246 5869
rect 3280 5835 3296 5869
rect 3230 5801 3296 5835
rect 3230 5767 3246 5801
rect 3280 5767 3296 5801
rect 3230 5733 3296 5767
rect 3230 5699 3246 5733
rect 3280 5699 3296 5733
rect 3230 5665 3296 5699
rect 3230 5631 3246 5665
rect 3280 5631 3296 5665
rect 3230 5590 3296 5631
rect 3326 6549 3392 6590
rect 3326 6515 3342 6549
rect 3376 6515 3392 6549
rect 3326 6481 3392 6515
rect 3326 6447 3342 6481
rect 3376 6447 3392 6481
rect 3326 6413 3392 6447
rect 3326 6379 3342 6413
rect 3376 6379 3392 6413
rect 3326 6345 3392 6379
rect 3326 6311 3342 6345
rect 3376 6311 3392 6345
rect 3326 6277 3392 6311
rect 3326 6243 3342 6277
rect 3376 6243 3392 6277
rect 3326 6209 3392 6243
rect 3326 6175 3342 6209
rect 3376 6175 3392 6209
rect 3326 6141 3392 6175
rect 3326 6107 3342 6141
rect 3376 6107 3392 6141
rect 3326 6073 3392 6107
rect 3326 6039 3342 6073
rect 3376 6039 3392 6073
rect 3326 6005 3392 6039
rect 3326 5971 3342 6005
rect 3376 5971 3392 6005
rect 3326 5937 3392 5971
rect 3326 5903 3342 5937
rect 3376 5903 3392 5937
rect 3326 5869 3392 5903
rect 3326 5835 3342 5869
rect 3376 5835 3392 5869
rect 3326 5801 3392 5835
rect 3326 5767 3342 5801
rect 3376 5767 3392 5801
rect 3326 5733 3392 5767
rect 3326 5699 3342 5733
rect 3376 5699 3392 5733
rect 3326 5665 3392 5699
rect 3326 5631 3342 5665
rect 3376 5631 3392 5665
rect 3326 5590 3392 5631
rect 3422 6549 3488 6590
rect 3422 6515 3438 6549
rect 3472 6515 3488 6549
rect 3422 6481 3488 6515
rect 3422 6447 3438 6481
rect 3472 6447 3488 6481
rect 3422 6413 3488 6447
rect 3422 6379 3438 6413
rect 3472 6379 3488 6413
rect 3422 6345 3488 6379
rect 3422 6311 3438 6345
rect 3472 6311 3488 6345
rect 3422 6277 3488 6311
rect 3422 6243 3438 6277
rect 3472 6243 3488 6277
rect 3422 6209 3488 6243
rect 3422 6175 3438 6209
rect 3472 6175 3488 6209
rect 3422 6141 3488 6175
rect 3422 6107 3438 6141
rect 3472 6107 3488 6141
rect 3422 6073 3488 6107
rect 3422 6039 3438 6073
rect 3472 6039 3488 6073
rect 3422 6005 3488 6039
rect 3422 5971 3438 6005
rect 3472 5971 3488 6005
rect 3422 5937 3488 5971
rect 3422 5903 3438 5937
rect 3472 5903 3488 5937
rect 3422 5869 3488 5903
rect 3422 5835 3438 5869
rect 3472 5835 3488 5869
rect 3422 5801 3488 5835
rect 3422 5767 3438 5801
rect 3472 5767 3488 5801
rect 3422 5733 3488 5767
rect 3422 5699 3438 5733
rect 3472 5699 3488 5733
rect 3422 5665 3488 5699
rect 3422 5631 3438 5665
rect 3472 5631 3488 5665
rect 3422 5590 3488 5631
rect 3518 6549 3584 6590
rect 3518 6515 3534 6549
rect 3568 6515 3584 6549
rect 3518 6481 3584 6515
rect 3518 6447 3534 6481
rect 3568 6447 3584 6481
rect 3518 6413 3584 6447
rect 3518 6379 3534 6413
rect 3568 6379 3584 6413
rect 3518 6345 3584 6379
rect 3518 6311 3534 6345
rect 3568 6311 3584 6345
rect 3518 6277 3584 6311
rect 3518 6243 3534 6277
rect 3568 6243 3584 6277
rect 3518 6209 3584 6243
rect 3518 6175 3534 6209
rect 3568 6175 3584 6209
rect 3518 6141 3584 6175
rect 3518 6107 3534 6141
rect 3568 6107 3584 6141
rect 3518 6073 3584 6107
rect 3518 6039 3534 6073
rect 3568 6039 3584 6073
rect 3518 6005 3584 6039
rect 3518 5971 3534 6005
rect 3568 5971 3584 6005
rect 3518 5937 3584 5971
rect 3518 5903 3534 5937
rect 3568 5903 3584 5937
rect 3518 5869 3584 5903
rect 3518 5835 3534 5869
rect 3568 5835 3584 5869
rect 3518 5801 3584 5835
rect 3518 5767 3534 5801
rect 3568 5767 3584 5801
rect 3518 5733 3584 5767
rect 3518 5699 3534 5733
rect 3568 5699 3584 5733
rect 3518 5665 3584 5699
rect 3518 5631 3534 5665
rect 3568 5631 3584 5665
rect 3518 5590 3584 5631
rect 3614 6549 3680 6590
rect 3614 6515 3630 6549
rect 3664 6515 3680 6549
rect 3614 6481 3680 6515
rect 3614 6447 3630 6481
rect 3664 6447 3680 6481
rect 3614 6413 3680 6447
rect 3614 6379 3630 6413
rect 3664 6379 3680 6413
rect 3614 6345 3680 6379
rect 3614 6311 3630 6345
rect 3664 6311 3680 6345
rect 3614 6277 3680 6311
rect 3614 6243 3630 6277
rect 3664 6243 3680 6277
rect 3614 6209 3680 6243
rect 3614 6175 3630 6209
rect 3664 6175 3680 6209
rect 3614 6141 3680 6175
rect 3614 6107 3630 6141
rect 3664 6107 3680 6141
rect 3614 6073 3680 6107
rect 3614 6039 3630 6073
rect 3664 6039 3680 6073
rect 3614 6005 3680 6039
rect 3614 5971 3630 6005
rect 3664 5971 3680 6005
rect 3614 5937 3680 5971
rect 3614 5903 3630 5937
rect 3664 5903 3680 5937
rect 3614 5869 3680 5903
rect 3614 5835 3630 5869
rect 3664 5835 3680 5869
rect 3614 5801 3680 5835
rect 3614 5767 3630 5801
rect 3664 5767 3680 5801
rect 3614 5733 3680 5767
rect 3614 5699 3630 5733
rect 3664 5699 3680 5733
rect 3614 5665 3680 5699
rect 3614 5631 3630 5665
rect 3664 5631 3680 5665
rect 3614 5590 3680 5631
rect 3710 6549 3776 6590
rect 3710 6515 3726 6549
rect 3760 6515 3776 6549
rect 3710 6481 3776 6515
rect 3710 6447 3726 6481
rect 3760 6447 3776 6481
rect 3710 6413 3776 6447
rect 3710 6379 3726 6413
rect 3760 6379 3776 6413
rect 3710 6345 3776 6379
rect 3710 6311 3726 6345
rect 3760 6311 3776 6345
rect 3710 6277 3776 6311
rect 3710 6243 3726 6277
rect 3760 6243 3776 6277
rect 3710 6209 3776 6243
rect 3710 6175 3726 6209
rect 3760 6175 3776 6209
rect 3710 6141 3776 6175
rect 3710 6107 3726 6141
rect 3760 6107 3776 6141
rect 3710 6073 3776 6107
rect 3710 6039 3726 6073
rect 3760 6039 3776 6073
rect 3710 6005 3776 6039
rect 3710 5971 3726 6005
rect 3760 5971 3776 6005
rect 3710 5937 3776 5971
rect 3710 5903 3726 5937
rect 3760 5903 3776 5937
rect 3710 5869 3776 5903
rect 3710 5835 3726 5869
rect 3760 5835 3776 5869
rect 3710 5801 3776 5835
rect 3710 5767 3726 5801
rect 3760 5767 3776 5801
rect 3710 5733 3776 5767
rect 3710 5699 3726 5733
rect 3760 5699 3776 5733
rect 3710 5665 3776 5699
rect 3710 5631 3726 5665
rect 3760 5631 3776 5665
rect 3710 5590 3776 5631
rect 3806 6549 3872 6590
rect 3806 6515 3822 6549
rect 3856 6515 3872 6549
rect 3806 6481 3872 6515
rect 3806 6447 3822 6481
rect 3856 6447 3872 6481
rect 3806 6413 3872 6447
rect 3806 6379 3822 6413
rect 3856 6379 3872 6413
rect 3806 6345 3872 6379
rect 3806 6311 3822 6345
rect 3856 6311 3872 6345
rect 3806 6277 3872 6311
rect 3806 6243 3822 6277
rect 3856 6243 3872 6277
rect 3806 6209 3872 6243
rect 3806 6175 3822 6209
rect 3856 6175 3872 6209
rect 3806 6141 3872 6175
rect 3806 6107 3822 6141
rect 3856 6107 3872 6141
rect 3806 6073 3872 6107
rect 3806 6039 3822 6073
rect 3856 6039 3872 6073
rect 3806 6005 3872 6039
rect 3806 5971 3822 6005
rect 3856 5971 3872 6005
rect 3806 5937 3872 5971
rect 3806 5903 3822 5937
rect 3856 5903 3872 5937
rect 3806 5869 3872 5903
rect 3806 5835 3822 5869
rect 3856 5835 3872 5869
rect 3806 5801 3872 5835
rect 3806 5767 3822 5801
rect 3856 5767 3872 5801
rect 3806 5733 3872 5767
rect 3806 5699 3822 5733
rect 3856 5699 3872 5733
rect 3806 5665 3872 5699
rect 3806 5631 3822 5665
rect 3856 5631 3872 5665
rect 3806 5590 3872 5631
rect 3902 6549 3968 6590
rect 3902 6515 3918 6549
rect 3952 6515 3968 6549
rect 3902 6481 3968 6515
rect 3902 6447 3918 6481
rect 3952 6447 3968 6481
rect 3902 6413 3968 6447
rect 3902 6379 3918 6413
rect 3952 6379 3968 6413
rect 3902 6345 3968 6379
rect 3902 6311 3918 6345
rect 3952 6311 3968 6345
rect 3902 6277 3968 6311
rect 3902 6243 3918 6277
rect 3952 6243 3968 6277
rect 3902 6209 3968 6243
rect 3902 6175 3918 6209
rect 3952 6175 3968 6209
rect 3902 6141 3968 6175
rect 3902 6107 3918 6141
rect 3952 6107 3968 6141
rect 3902 6073 3968 6107
rect 3902 6039 3918 6073
rect 3952 6039 3968 6073
rect 3902 6005 3968 6039
rect 3902 5971 3918 6005
rect 3952 5971 3968 6005
rect 3902 5937 3968 5971
rect 3902 5903 3918 5937
rect 3952 5903 3968 5937
rect 3902 5869 3968 5903
rect 3902 5835 3918 5869
rect 3952 5835 3968 5869
rect 3902 5801 3968 5835
rect 3902 5767 3918 5801
rect 3952 5767 3968 5801
rect 3902 5733 3968 5767
rect 3902 5699 3918 5733
rect 3952 5699 3968 5733
rect 3902 5665 3968 5699
rect 3902 5631 3918 5665
rect 3952 5631 3968 5665
rect 3902 5590 3968 5631
rect 3998 6549 4064 6590
rect 3998 6515 4014 6549
rect 4048 6515 4064 6549
rect 3998 6481 4064 6515
rect 3998 6447 4014 6481
rect 4048 6447 4064 6481
rect 3998 6413 4064 6447
rect 3998 6379 4014 6413
rect 4048 6379 4064 6413
rect 3998 6345 4064 6379
rect 3998 6311 4014 6345
rect 4048 6311 4064 6345
rect 3998 6277 4064 6311
rect 3998 6243 4014 6277
rect 4048 6243 4064 6277
rect 3998 6209 4064 6243
rect 3998 6175 4014 6209
rect 4048 6175 4064 6209
rect 3998 6141 4064 6175
rect 3998 6107 4014 6141
rect 4048 6107 4064 6141
rect 3998 6073 4064 6107
rect 3998 6039 4014 6073
rect 4048 6039 4064 6073
rect 3998 6005 4064 6039
rect 3998 5971 4014 6005
rect 4048 5971 4064 6005
rect 3998 5937 4064 5971
rect 3998 5903 4014 5937
rect 4048 5903 4064 5937
rect 3998 5869 4064 5903
rect 3998 5835 4014 5869
rect 4048 5835 4064 5869
rect 3998 5801 4064 5835
rect 3998 5767 4014 5801
rect 4048 5767 4064 5801
rect 3998 5733 4064 5767
rect 3998 5699 4014 5733
rect 4048 5699 4064 5733
rect 3998 5665 4064 5699
rect 3998 5631 4014 5665
rect 4048 5631 4064 5665
rect 3998 5590 4064 5631
rect 4094 6549 4160 6590
rect 4094 6515 4110 6549
rect 4144 6515 4160 6549
rect 4094 6481 4160 6515
rect 4094 6447 4110 6481
rect 4144 6447 4160 6481
rect 4094 6413 4160 6447
rect 4094 6379 4110 6413
rect 4144 6379 4160 6413
rect 4094 6345 4160 6379
rect 4094 6311 4110 6345
rect 4144 6311 4160 6345
rect 4094 6277 4160 6311
rect 4094 6243 4110 6277
rect 4144 6243 4160 6277
rect 4094 6209 4160 6243
rect 4094 6175 4110 6209
rect 4144 6175 4160 6209
rect 4094 6141 4160 6175
rect 4094 6107 4110 6141
rect 4144 6107 4160 6141
rect 4094 6073 4160 6107
rect 4094 6039 4110 6073
rect 4144 6039 4160 6073
rect 4094 6005 4160 6039
rect 4094 5971 4110 6005
rect 4144 5971 4160 6005
rect 4094 5937 4160 5971
rect 4094 5903 4110 5937
rect 4144 5903 4160 5937
rect 4094 5869 4160 5903
rect 4094 5835 4110 5869
rect 4144 5835 4160 5869
rect 4094 5801 4160 5835
rect 4094 5767 4110 5801
rect 4144 5767 4160 5801
rect 4094 5733 4160 5767
rect 4094 5699 4110 5733
rect 4144 5699 4160 5733
rect 4094 5665 4160 5699
rect 4094 5631 4110 5665
rect 4144 5631 4160 5665
rect 4094 5590 4160 5631
rect 4190 6549 4256 6590
rect 4190 6515 4206 6549
rect 4240 6515 4256 6549
rect 4190 6481 4256 6515
rect 4190 6447 4206 6481
rect 4240 6447 4256 6481
rect 4190 6413 4256 6447
rect 4190 6379 4206 6413
rect 4240 6379 4256 6413
rect 4190 6345 4256 6379
rect 4190 6311 4206 6345
rect 4240 6311 4256 6345
rect 4190 6277 4256 6311
rect 4190 6243 4206 6277
rect 4240 6243 4256 6277
rect 4190 6209 4256 6243
rect 4190 6175 4206 6209
rect 4240 6175 4256 6209
rect 4190 6141 4256 6175
rect 4190 6107 4206 6141
rect 4240 6107 4256 6141
rect 4190 6073 4256 6107
rect 4190 6039 4206 6073
rect 4240 6039 4256 6073
rect 4190 6005 4256 6039
rect 4190 5971 4206 6005
rect 4240 5971 4256 6005
rect 4190 5937 4256 5971
rect 4190 5903 4206 5937
rect 4240 5903 4256 5937
rect 4190 5869 4256 5903
rect 4190 5835 4206 5869
rect 4240 5835 4256 5869
rect 4190 5801 4256 5835
rect 4190 5767 4206 5801
rect 4240 5767 4256 5801
rect 4190 5733 4256 5767
rect 4190 5699 4206 5733
rect 4240 5699 4256 5733
rect 4190 5665 4256 5699
rect 4190 5631 4206 5665
rect 4240 5631 4256 5665
rect 4190 5590 4256 5631
rect 4286 6549 4348 6590
rect 4286 6515 4302 6549
rect 4336 6515 4348 6549
rect 4286 6481 4348 6515
rect 4286 6447 4302 6481
rect 4336 6447 4348 6481
rect 4286 6413 4348 6447
rect 4286 6379 4302 6413
rect 4336 6379 4348 6413
rect 4286 6345 4348 6379
rect 4286 6311 4302 6345
rect 4336 6311 4348 6345
rect 4286 6277 4348 6311
rect 4286 6243 4302 6277
rect 4336 6243 4348 6277
rect 4286 6209 4348 6243
rect 4286 6175 4302 6209
rect 4336 6175 4348 6209
rect 4286 6141 4348 6175
rect 4286 6107 4302 6141
rect 4336 6107 4348 6141
rect 4286 6073 4348 6107
rect 4286 6039 4302 6073
rect 4336 6039 4348 6073
rect 4286 6005 4348 6039
rect 4286 5971 4302 6005
rect 4336 5971 4348 6005
rect 4286 5937 4348 5971
rect 4286 5903 4302 5937
rect 4336 5903 4348 5937
rect 4286 5869 4348 5903
rect 4286 5835 4302 5869
rect 4336 5835 4348 5869
rect 4286 5801 4348 5835
rect 4286 5767 4302 5801
rect 4336 5767 4348 5801
rect 4286 5733 4348 5767
rect 4286 5699 4302 5733
rect 4336 5699 4348 5733
rect 4286 5665 4348 5699
rect 4286 5631 4302 5665
rect 4336 5631 4348 5665
rect 4286 5590 4348 5631
rect 4904 6545 4966 6586
rect 4904 6511 4916 6545
rect 4950 6511 4966 6545
rect 4904 6477 4966 6511
rect 4904 6443 4916 6477
rect 4950 6443 4966 6477
rect 4904 6409 4966 6443
rect 4904 6375 4916 6409
rect 4950 6375 4966 6409
rect 4904 6341 4966 6375
rect 4904 6307 4916 6341
rect 4950 6307 4966 6341
rect 4904 6273 4966 6307
rect 4904 6239 4916 6273
rect 4950 6239 4966 6273
rect 4904 6205 4966 6239
rect 4904 6171 4916 6205
rect 4950 6171 4966 6205
rect 4904 6137 4966 6171
rect 4904 6103 4916 6137
rect 4950 6103 4966 6137
rect 4904 6069 4966 6103
rect 4904 6035 4916 6069
rect 4950 6035 4966 6069
rect 4904 6001 4966 6035
rect 4904 5967 4916 6001
rect 4950 5967 4966 6001
rect 4904 5933 4966 5967
rect 4904 5899 4916 5933
rect 4950 5899 4966 5933
rect 4904 5865 4966 5899
rect 4904 5831 4916 5865
rect 4950 5831 4966 5865
rect 4904 5797 4966 5831
rect 4904 5763 4916 5797
rect 4950 5763 4966 5797
rect 4904 5729 4966 5763
rect 4904 5695 4916 5729
rect 4950 5695 4966 5729
rect 4904 5661 4966 5695
rect 4904 5627 4916 5661
rect 4950 5627 4966 5661
rect 4904 5586 4966 5627
rect 4996 6545 5062 6586
rect 4996 6511 5012 6545
rect 5046 6511 5062 6545
rect 4996 6477 5062 6511
rect 4996 6443 5012 6477
rect 5046 6443 5062 6477
rect 4996 6409 5062 6443
rect 4996 6375 5012 6409
rect 5046 6375 5062 6409
rect 4996 6341 5062 6375
rect 4996 6307 5012 6341
rect 5046 6307 5062 6341
rect 4996 6273 5062 6307
rect 4996 6239 5012 6273
rect 5046 6239 5062 6273
rect 4996 6205 5062 6239
rect 4996 6171 5012 6205
rect 5046 6171 5062 6205
rect 4996 6137 5062 6171
rect 4996 6103 5012 6137
rect 5046 6103 5062 6137
rect 4996 6069 5062 6103
rect 4996 6035 5012 6069
rect 5046 6035 5062 6069
rect 4996 6001 5062 6035
rect 4996 5967 5012 6001
rect 5046 5967 5062 6001
rect 4996 5933 5062 5967
rect 4996 5899 5012 5933
rect 5046 5899 5062 5933
rect 4996 5865 5062 5899
rect 4996 5831 5012 5865
rect 5046 5831 5062 5865
rect 4996 5797 5062 5831
rect 4996 5763 5012 5797
rect 5046 5763 5062 5797
rect 4996 5729 5062 5763
rect 4996 5695 5012 5729
rect 5046 5695 5062 5729
rect 4996 5661 5062 5695
rect 4996 5627 5012 5661
rect 5046 5627 5062 5661
rect 4996 5586 5062 5627
rect 5092 6545 5158 6586
rect 5092 6511 5108 6545
rect 5142 6511 5158 6545
rect 5092 6477 5158 6511
rect 5092 6443 5108 6477
rect 5142 6443 5158 6477
rect 5092 6409 5158 6443
rect 5092 6375 5108 6409
rect 5142 6375 5158 6409
rect 5092 6341 5158 6375
rect 5092 6307 5108 6341
rect 5142 6307 5158 6341
rect 5092 6273 5158 6307
rect 5092 6239 5108 6273
rect 5142 6239 5158 6273
rect 5092 6205 5158 6239
rect 5092 6171 5108 6205
rect 5142 6171 5158 6205
rect 5092 6137 5158 6171
rect 5092 6103 5108 6137
rect 5142 6103 5158 6137
rect 5092 6069 5158 6103
rect 5092 6035 5108 6069
rect 5142 6035 5158 6069
rect 5092 6001 5158 6035
rect 5092 5967 5108 6001
rect 5142 5967 5158 6001
rect 5092 5933 5158 5967
rect 5092 5899 5108 5933
rect 5142 5899 5158 5933
rect 5092 5865 5158 5899
rect 5092 5831 5108 5865
rect 5142 5831 5158 5865
rect 5092 5797 5158 5831
rect 5092 5763 5108 5797
rect 5142 5763 5158 5797
rect 5092 5729 5158 5763
rect 5092 5695 5108 5729
rect 5142 5695 5158 5729
rect 5092 5661 5158 5695
rect 5092 5627 5108 5661
rect 5142 5627 5158 5661
rect 5092 5586 5158 5627
rect 5188 6545 5254 6586
rect 5188 6511 5204 6545
rect 5238 6511 5254 6545
rect 5188 6477 5254 6511
rect 5188 6443 5204 6477
rect 5238 6443 5254 6477
rect 5188 6409 5254 6443
rect 5188 6375 5204 6409
rect 5238 6375 5254 6409
rect 5188 6341 5254 6375
rect 5188 6307 5204 6341
rect 5238 6307 5254 6341
rect 5188 6273 5254 6307
rect 5188 6239 5204 6273
rect 5238 6239 5254 6273
rect 5188 6205 5254 6239
rect 5188 6171 5204 6205
rect 5238 6171 5254 6205
rect 5188 6137 5254 6171
rect 5188 6103 5204 6137
rect 5238 6103 5254 6137
rect 5188 6069 5254 6103
rect 5188 6035 5204 6069
rect 5238 6035 5254 6069
rect 5188 6001 5254 6035
rect 5188 5967 5204 6001
rect 5238 5967 5254 6001
rect 5188 5933 5254 5967
rect 5188 5899 5204 5933
rect 5238 5899 5254 5933
rect 5188 5865 5254 5899
rect 5188 5831 5204 5865
rect 5238 5831 5254 5865
rect 5188 5797 5254 5831
rect 5188 5763 5204 5797
rect 5238 5763 5254 5797
rect 5188 5729 5254 5763
rect 5188 5695 5204 5729
rect 5238 5695 5254 5729
rect 5188 5661 5254 5695
rect 5188 5627 5204 5661
rect 5238 5627 5254 5661
rect 5188 5586 5254 5627
rect 5284 6545 5350 6586
rect 5284 6511 5300 6545
rect 5334 6511 5350 6545
rect 5284 6477 5350 6511
rect 5284 6443 5300 6477
rect 5334 6443 5350 6477
rect 5284 6409 5350 6443
rect 5284 6375 5300 6409
rect 5334 6375 5350 6409
rect 5284 6341 5350 6375
rect 5284 6307 5300 6341
rect 5334 6307 5350 6341
rect 5284 6273 5350 6307
rect 5284 6239 5300 6273
rect 5334 6239 5350 6273
rect 5284 6205 5350 6239
rect 5284 6171 5300 6205
rect 5334 6171 5350 6205
rect 5284 6137 5350 6171
rect 5284 6103 5300 6137
rect 5334 6103 5350 6137
rect 5284 6069 5350 6103
rect 5284 6035 5300 6069
rect 5334 6035 5350 6069
rect 5284 6001 5350 6035
rect 5284 5967 5300 6001
rect 5334 5967 5350 6001
rect 5284 5933 5350 5967
rect 5284 5899 5300 5933
rect 5334 5899 5350 5933
rect 5284 5865 5350 5899
rect 5284 5831 5300 5865
rect 5334 5831 5350 5865
rect 5284 5797 5350 5831
rect 5284 5763 5300 5797
rect 5334 5763 5350 5797
rect 5284 5729 5350 5763
rect 5284 5695 5300 5729
rect 5334 5695 5350 5729
rect 5284 5661 5350 5695
rect 5284 5627 5300 5661
rect 5334 5627 5350 5661
rect 5284 5586 5350 5627
rect 5380 6545 5446 6586
rect 5380 6511 5396 6545
rect 5430 6511 5446 6545
rect 5380 6477 5446 6511
rect 5380 6443 5396 6477
rect 5430 6443 5446 6477
rect 5380 6409 5446 6443
rect 5380 6375 5396 6409
rect 5430 6375 5446 6409
rect 5380 6341 5446 6375
rect 5380 6307 5396 6341
rect 5430 6307 5446 6341
rect 5380 6273 5446 6307
rect 5380 6239 5396 6273
rect 5430 6239 5446 6273
rect 5380 6205 5446 6239
rect 5380 6171 5396 6205
rect 5430 6171 5446 6205
rect 5380 6137 5446 6171
rect 5380 6103 5396 6137
rect 5430 6103 5446 6137
rect 5380 6069 5446 6103
rect 5380 6035 5396 6069
rect 5430 6035 5446 6069
rect 5380 6001 5446 6035
rect 5380 5967 5396 6001
rect 5430 5967 5446 6001
rect 5380 5933 5446 5967
rect 5380 5899 5396 5933
rect 5430 5899 5446 5933
rect 5380 5865 5446 5899
rect 5380 5831 5396 5865
rect 5430 5831 5446 5865
rect 5380 5797 5446 5831
rect 5380 5763 5396 5797
rect 5430 5763 5446 5797
rect 5380 5729 5446 5763
rect 5380 5695 5396 5729
rect 5430 5695 5446 5729
rect 5380 5661 5446 5695
rect 5380 5627 5396 5661
rect 5430 5627 5446 5661
rect 5380 5586 5446 5627
rect 5476 6545 5542 6586
rect 5476 6511 5492 6545
rect 5526 6511 5542 6545
rect 5476 6477 5542 6511
rect 5476 6443 5492 6477
rect 5526 6443 5542 6477
rect 5476 6409 5542 6443
rect 5476 6375 5492 6409
rect 5526 6375 5542 6409
rect 5476 6341 5542 6375
rect 5476 6307 5492 6341
rect 5526 6307 5542 6341
rect 5476 6273 5542 6307
rect 5476 6239 5492 6273
rect 5526 6239 5542 6273
rect 5476 6205 5542 6239
rect 5476 6171 5492 6205
rect 5526 6171 5542 6205
rect 5476 6137 5542 6171
rect 5476 6103 5492 6137
rect 5526 6103 5542 6137
rect 5476 6069 5542 6103
rect 5476 6035 5492 6069
rect 5526 6035 5542 6069
rect 5476 6001 5542 6035
rect 5476 5967 5492 6001
rect 5526 5967 5542 6001
rect 5476 5933 5542 5967
rect 5476 5899 5492 5933
rect 5526 5899 5542 5933
rect 5476 5865 5542 5899
rect 5476 5831 5492 5865
rect 5526 5831 5542 5865
rect 5476 5797 5542 5831
rect 5476 5763 5492 5797
rect 5526 5763 5542 5797
rect 5476 5729 5542 5763
rect 5476 5695 5492 5729
rect 5526 5695 5542 5729
rect 5476 5661 5542 5695
rect 5476 5627 5492 5661
rect 5526 5627 5542 5661
rect 5476 5586 5542 5627
rect 5572 6545 5638 6586
rect 5572 6511 5588 6545
rect 5622 6511 5638 6545
rect 5572 6477 5638 6511
rect 5572 6443 5588 6477
rect 5622 6443 5638 6477
rect 5572 6409 5638 6443
rect 5572 6375 5588 6409
rect 5622 6375 5638 6409
rect 5572 6341 5638 6375
rect 5572 6307 5588 6341
rect 5622 6307 5638 6341
rect 5572 6273 5638 6307
rect 5572 6239 5588 6273
rect 5622 6239 5638 6273
rect 5572 6205 5638 6239
rect 5572 6171 5588 6205
rect 5622 6171 5638 6205
rect 5572 6137 5638 6171
rect 5572 6103 5588 6137
rect 5622 6103 5638 6137
rect 5572 6069 5638 6103
rect 5572 6035 5588 6069
rect 5622 6035 5638 6069
rect 5572 6001 5638 6035
rect 5572 5967 5588 6001
rect 5622 5967 5638 6001
rect 5572 5933 5638 5967
rect 5572 5899 5588 5933
rect 5622 5899 5638 5933
rect 5572 5865 5638 5899
rect 5572 5831 5588 5865
rect 5622 5831 5638 5865
rect 5572 5797 5638 5831
rect 5572 5763 5588 5797
rect 5622 5763 5638 5797
rect 5572 5729 5638 5763
rect 5572 5695 5588 5729
rect 5622 5695 5638 5729
rect 5572 5661 5638 5695
rect 5572 5627 5588 5661
rect 5622 5627 5638 5661
rect 5572 5586 5638 5627
rect 5668 6545 5730 6586
rect 5668 6511 5684 6545
rect 5718 6511 5730 6545
rect 5668 6477 5730 6511
rect 5668 6443 5684 6477
rect 5718 6443 5730 6477
rect 5668 6409 5730 6443
rect 5668 6375 5684 6409
rect 5718 6375 5730 6409
rect 5668 6341 5730 6375
rect 5668 6307 5684 6341
rect 5718 6307 5730 6341
rect 5668 6273 5730 6307
rect 5668 6239 5684 6273
rect 5718 6239 5730 6273
rect 5668 6205 5730 6239
rect 5668 6171 5684 6205
rect 5718 6171 5730 6205
rect 5668 6137 5730 6171
rect 5668 6103 5684 6137
rect 5718 6103 5730 6137
rect 5668 6069 5730 6103
rect 5668 6035 5684 6069
rect 5718 6035 5730 6069
rect 5668 6001 5730 6035
rect 5668 5967 5684 6001
rect 5718 5967 5730 6001
rect 5668 5933 5730 5967
rect 5668 5899 5684 5933
rect 5718 5899 5730 5933
rect 5668 5865 5730 5899
rect 5668 5831 5684 5865
rect 5718 5831 5730 5865
rect 5668 5797 5730 5831
rect 5668 5763 5684 5797
rect 5718 5763 5730 5797
rect 5668 5729 5730 5763
rect 5668 5695 5684 5729
rect 5718 5695 5730 5729
rect 5668 5661 5730 5695
rect 5668 5627 5684 5661
rect 5718 5627 5730 5661
rect 5668 5586 5730 5627
rect 6168 6549 6230 6590
rect 6168 6515 6180 6549
rect 6214 6515 6230 6549
rect 6168 6481 6230 6515
rect 6168 6447 6180 6481
rect 6214 6447 6230 6481
rect 6168 6413 6230 6447
rect 6168 6379 6180 6413
rect 6214 6379 6230 6413
rect 6168 6345 6230 6379
rect 6168 6311 6180 6345
rect 6214 6311 6230 6345
rect 6168 6277 6230 6311
rect 6168 6243 6180 6277
rect 6214 6243 6230 6277
rect 6168 6209 6230 6243
rect 6168 6175 6180 6209
rect 6214 6175 6230 6209
rect 6168 6141 6230 6175
rect 6168 6107 6180 6141
rect 6214 6107 6230 6141
rect 6168 6073 6230 6107
rect 6168 6039 6180 6073
rect 6214 6039 6230 6073
rect 6168 6005 6230 6039
rect 6168 5971 6180 6005
rect 6214 5971 6230 6005
rect 6168 5937 6230 5971
rect 6168 5903 6180 5937
rect 6214 5903 6230 5937
rect 6168 5869 6230 5903
rect 6168 5835 6180 5869
rect 6214 5835 6230 5869
rect 6168 5801 6230 5835
rect 6168 5767 6180 5801
rect 6214 5767 6230 5801
rect 6168 5733 6230 5767
rect 6168 5699 6180 5733
rect 6214 5699 6230 5733
rect 6168 5665 6230 5699
rect 6168 5631 6180 5665
rect 6214 5631 6230 5665
rect 6168 5590 6230 5631
rect 6260 6549 6326 6590
rect 6260 6515 6276 6549
rect 6310 6515 6326 6549
rect 6260 6481 6326 6515
rect 6260 6447 6276 6481
rect 6310 6447 6326 6481
rect 6260 6413 6326 6447
rect 6260 6379 6276 6413
rect 6310 6379 6326 6413
rect 6260 6345 6326 6379
rect 6260 6311 6276 6345
rect 6310 6311 6326 6345
rect 6260 6277 6326 6311
rect 6260 6243 6276 6277
rect 6310 6243 6326 6277
rect 6260 6209 6326 6243
rect 6260 6175 6276 6209
rect 6310 6175 6326 6209
rect 6260 6141 6326 6175
rect 6260 6107 6276 6141
rect 6310 6107 6326 6141
rect 6260 6073 6326 6107
rect 6260 6039 6276 6073
rect 6310 6039 6326 6073
rect 6260 6005 6326 6039
rect 6260 5971 6276 6005
rect 6310 5971 6326 6005
rect 6260 5937 6326 5971
rect 6260 5903 6276 5937
rect 6310 5903 6326 5937
rect 6260 5869 6326 5903
rect 6260 5835 6276 5869
rect 6310 5835 6326 5869
rect 6260 5801 6326 5835
rect 6260 5767 6276 5801
rect 6310 5767 6326 5801
rect 6260 5733 6326 5767
rect 6260 5699 6276 5733
rect 6310 5699 6326 5733
rect 6260 5665 6326 5699
rect 6260 5631 6276 5665
rect 6310 5631 6326 5665
rect 6260 5590 6326 5631
rect 6356 6549 6422 6590
rect 6356 6515 6372 6549
rect 6406 6515 6422 6549
rect 6356 6481 6422 6515
rect 6356 6447 6372 6481
rect 6406 6447 6422 6481
rect 6356 6413 6422 6447
rect 6356 6379 6372 6413
rect 6406 6379 6422 6413
rect 6356 6345 6422 6379
rect 6356 6311 6372 6345
rect 6406 6311 6422 6345
rect 6356 6277 6422 6311
rect 6356 6243 6372 6277
rect 6406 6243 6422 6277
rect 6356 6209 6422 6243
rect 6356 6175 6372 6209
rect 6406 6175 6422 6209
rect 6356 6141 6422 6175
rect 6356 6107 6372 6141
rect 6406 6107 6422 6141
rect 6356 6073 6422 6107
rect 6356 6039 6372 6073
rect 6406 6039 6422 6073
rect 6356 6005 6422 6039
rect 6356 5971 6372 6005
rect 6406 5971 6422 6005
rect 6356 5937 6422 5971
rect 6356 5903 6372 5937
rect 6406 5903 6422 5937
rect 6356 5869 6422 5903
rect 6356 5835 6372 5869
rect 6406 5835 6422 5869
rect 6356 5801 6422 5835
rect 6356 5767 6372 5801
rect 6406 5767 6422 5801
rect 6356 5733 6422 5767
rect 6356 5699 6372 5733
rect 6406 5699 6422 5733
rect 6356 5665 6422 5699
rect 6356 5631 6372 5665
rect 6406 5631 6422 5665
rect 6356 5590 6422 5631
rect 6452 6549 6518 6590
rect 6452 6515 6468 6549
rect 6502 6515 6518 6549
rect 6452 6481 6518 6515
rect 6452 6447 6468 6481
rect 6502 6447 6518 6481
rect 6452 6413 6518 6447
rect 6452 6379 6468 6413
rect 6502 6379 6518 6413
rect 6452 6345 6518 6379
rect 6452 6311 6468 6345
rect 6502 6311 6518 6345
rect 6452 6277 6518 6311
rect 6452 6243 6468 6277
rect 6502 6243 6518 6277
rect 6452 6209 6518 6243
rect 6452 6175 6468 6209
rect 6502 6175 6518 6209
rect 6452 6141 6518 6175
rect 6452 6107 6468 6141
rect 6502 6107 6518 6141
rect 6452 6073 6518 6107
rect 6452 6039 6468 6073
rect 6502 6039 6518 6073
rect 6452 6005 6518 6039
rect 6452 5971 6468 6005
rect 6502 5971 6518 6005
rect 6452 5937 6518 5971
rect 6452 5903 6468 5937
rect 6502 5903 6518 5937
rect 6452 5869 6518 5903
rect 6452 5835 6468 5869
rect 6502 5835 6518 5869
rect 6452 5801 6518 5835
rect 6452 5767 6468 5801
rect 6502 5767 6518 5801
rect 6452 5733 6518 5767
rect 6452 5699 6468 5733
rect 6502 5699 6518 5733
rect 6452 5665 6518 5699
rect 6452 5631 6468 5665
rect 6502 5631 6518 5665
rect 6452 5590 6518 5631
rect 6548 6549 6614 6590
rect 6548 6515 6564 6549
rect 6598 6515 6614 6549
rect 6548 6481 6614 6515
rect 6548 6447 6564 6481
rect 6598 6447 6614 6481
rect 6548 6413 6614 6447
rect 6548 6379 6564 6413
rect 6598 6379 6614 6413
rect 6548 6345 6614 6379
rect 6548 6311 6564 6345
rect 6598 6311 6614 6345
rect 6548 6277 6614 6311
rect 6548 6243 6564 6277
rect 6598 6243 6614 6277
rect 6548 6209 6614 6243
rect 6548 6175 6564 6209
rect 6598 6175 6614 6209
rect 6548 6141 6614 6175
rect 6548 6107 6564 6141
rect 6598 6107 6614 6141
rect 6548 6073 6614 6107
rect 6548 6039 6564 6073
rect 6598 6039 6614 6073
rect 6548 6005 6614 6039
rect 6548 5971 6564 6005
rect 6598 5971 6614 6005
rect 6548 5937 6614 5971
rect 6548 5903 6564 5937
rect 6598 5903 6614 5937
rect 6548 5869 6614 5903
rect 6548 5835 6564 5869
rect 6598 5835 6614 5869
rect 6548 5801 6614 5835
rect 6548 5767 6564 5801
rect 6598 5767 6614 5801
rect 6548 5733 6614 5767
rect 6548 5699 6564 5733
rect 6598 5699 6614 5733
rect 6548 5665 6614 5699
rect 6548 5631 6564 5665
rect 6598 5631 6614 5665
rect 6548 5590 6614 5631
rect 6644 6549 6710 6590
rect 6644 6515 6660 6549
rect 6694 6515 6710 6549
rect 6644 6481 6710 6515
rect 6644 6447 6660 6481
rect 6694 6447 6710 6481
rect 6644 6413 6710 6447
rect 6644 6379 6660 6413
rect 6694 6379 6710 6413
rect 6644 6345 6710 6379
rect 6644 6311 6660 6345
rect 6694 6311 6710 6345
rect 6644 6277 6710 6311
rect 6644 6243 6660 6277
rect 6694 6243 6710 6277
rect 6644 6209 6710 6243
rect 6644 6175 6660 6209
rect 6694 6175 6710 6209
rect 6644 6141 6710 6175
rect 6644 6107 6660 6141
rect 6694 6107 6710 6141
rect 6644 6073 6710 6107
rect 6644 6039 6660 6073
rect 6694 6039 6710 6073
rect 6644 6005 6710 6039
rect 6644 5971 6660 6005
rect 6694 5971 6710 6005
rect 6644 5937 6710 5971
rect 6644 5903 6660 5937
rect 6694 5903 6710 5937
rect 6644 5869 6710 5903
rect 6644 5835 6660 5869
rect 6694 5835 6710 5869
rect 6644 5801 6710 5835
rect 6644 5767 6660 5801
rect 6694 5767 6710 5801
rect 6644 5733 6710 5767
rect 6644 5699 6660 5733
rect 6694 5699 6710 5733
rect 6644 5665 6710 5699
rect 6644 5631 6660 5665
rect 6694 5631 6710 5665
rect 6644 5590 6710 5631
rect 6740 6549 6806 6590
rect 6740 6515 6756 6549
rect 6790 6515 6806 6549
rect 6740 6481 6806 6515
rect 6740 6447 6756 6481
rect 6790 6447 6806 6481
rect 6740 6413 6806 6447
rect 6740 6379 6756 6413
rect 6790 6379 6806 6413
rect 6740 6345 6806 6379
rect 6740 6311 6756 6345
rect 6790 6311 6806 6345
rect 6740 6277 6806 6311
rect 6740 6243 6756 6277
rect 6790 6243 6806 6277
rect 6740 6209 6806 6243
rect 6740 6175 6756 6209
rect 6790 6175 6806 6209
rect 6740 6141 6806 6175
rect 6740 6107 6756 6141
rect 6790 6107 6806 6141
rect 6740 6073 6806 6107
rect 6740 6039 6756 6073
rect 6790 6039 6806 6073
rect 6740 6005 6806 6039
rect 6740 5971 6756 6005
rect 6790 5971 6806 6005
rect 6740 5937 6806 5971
rect 6740 5903 6756 5937
rect 6790 5903 6806 5937
rect 6740 5869 6806 5903
rect 6740 5835 6756 5869
rect 6790 5835 6806 5869
rect 6740 5801 6806 5835
rect 6740 5767 6756 5801
rect 6790 5767 6806 5801
rect 6740 5733 6806 5767
rect 6740 5699 6756 5733
rect 6790 5699 6806 5733
rect 6740 5665 6806 5699
rect 6740 5631 6756 5665
rect 6790 5631 6806 5665
rect 6740 5590 6806 5631
rect 6836 6549 6902 6590
rect 6836 6515 6852 6549
rect 6886 6515 6902 6549
rect 6836 6481 6902 6515
rect 6836 6447 6852 6481
rect 6886 6447 6902 6481
rect 6836 6413 6902 6447
rect 6836 6379 6852 6413
rect 6886 6379 6902 6413
rect 6836 6345 6902 6379
rect 6836 6311 6852 6345
rect 6886 6311 6902 6345
rect 6836 6277 6902 6311
rect 6836 6243 6852 6277
rect 6886 6243 6902 6277
rect 6836 6209 6902 6243
rect 6836 6175 6852 6209
rect 6886 6175 6902 6209
rect 6836 6141 6902 6175
rect 6836 6107 6852 6141
rect 6886 6107 6902 6141
rect 6836 6073 6902 6107
rect 6836 6039 6852 6073
rect 6886 6039 6902 6073
rect 6836 6005 6902 6039
rect 6836 5971 6852 6005
rect 6886 5971 6902 6005
rect 6836 5937 6902 5971
rect 6836 5903 6852 5937
rect 6886 5903 6902 5937
rect 6836 5869 6902 5903
rect 6836 5835 6852 5869
rect 6886 5835 6902 5869
rect 6836 5801 6902 5835
rect 6836 5767 6852 5801
rect 6886 5767 6902 5801
rect 6836 5733 6902 5767
rect 6836 5699 6852 5733
rect 6886 5699 6902 5733
rect 6836 5665 6902 5699
rect 6836 5631 6852 5665
rect 6886 5631 6902 5665
rect 6836 5590 6902 5631
rect 6932 6549 6998 6590
rect 6932 6515 6948 6549
rect 6982 6515 6998 6549
rect 6932 6481 6998 6515
rect 6932 6447 6948 6481
rect 6982 6447 6998 6481
rect 6932 6413 6998 6447
rect 6932 6379 6948 6413
rect 6982 6379 6998 6413
rect 6932 6345 6998 6379
rect 6932 6311 6948 6345
rect 6982 6311 6998 6345
rect 6932 6277 6998 6311
rect 6932 6243 6948 6277
rect 6982 6243 6998 6277
rect 6932 6209 6998 6243
rect 6932 6175 6948 6209
rect 6982 6175 6998 6209
rect 6932 6141 6998 6175
rect 6932 6107 6948 6141
rect 6982 6107 6998 6141
rect 6932 6073 6998 6107
rect 6932 6039 6948 6073
rect 6982 6039 6998 6073
rect 6932 6005 6998 6039
rect 6932 5971 6948 6005
rect 6982 5971 6998 6005
rect 6932 5937 6998 5971
rect 6932 5903 6948 5937
rect 6982 5903 6998 5937
rect 6932 5869 6998 5903
rect 6932 5835 6948 5869
rect 6982 5835 6998 5869
rect 6932 5801 6998 5835
rect 6932 5767 6948 5801
rect 6982 5767 6998 5801
rect 6932 5733 6998 5767
rect 6932 5699 6948 5733
rect 6982 5699 6998 5733
rect 6932 5665 6998 5699
rect 6932 5631 6948 5665
rect 6982 5631 6998 5665
rect 6932 5590 6998 5631
rect 7028 6549 7094 6590
rect 7028 6515 7044 6549
rect 7078 6515 7094 6549
rect 7028 6481 7094 6515
rect 7028 6447 7044 6481
rect 7078 6447 7094 6481
rect 7028 6413 7094 6447
rect 7028 6379 7044 6413
rect 7078 6379 7094 6413
rect 7028 6345 7094 6379
rect 7028 6311 7044 6345
rect 7078 6311 7094 6345
rect 7028 6277 7094 6311
rect 7028 6243 7044 6277
rect 7078 6243 7094 6277
rect 7028 6209 7094 6243
rect 7028 6175 7044 6209
rect 7078 6175 7094 6209
rect 7028 6141 7094 6175
rect 7028 6107 7044 6141
rect 7078 6107 7094 6141
rect 7028 6073 7094 6107
rect 7028 6039 7044 6073
rect 7078 6039 7094 6073
rect 7028 6005 7094 6039
rect 7028 5971 7044 6005
rect 7078 5971 7094 6005
rect 7028 5937 7094 5971
rect 7028 5903 7044 5937
rect 7078 5903 7094 5937
rect 7028 5869 7094 5903
rect 7028 5835 7044 5869
rect 7078 5835 7094 5869
rect 7028 5801 7094 5835
rect 7028 5767 7044 5801
rect 7078 5767 7094 5801
rect 7028 5733 7094 5767
rect 7028 5699 7044 5733
rect 7078 5699 7094 5733
rect 7028 5665 7094 5699
rect 7028 5631 7044 5665
rect 7078 5631 7094 5665
rect 7028 5590 7094 5631
rect 7124 6549 7190 6590
rect 7124 6515 7140 6549
rect 7174 6515 7190 6549
rect 7124 6481 7190 6515
rect 7124 6447 7140 6481
rect 7174 6447 7190 6481
rect 7124 6413 7190 6447
rect 7124 6379 7140 6413
rect 7174 6379 7190 6413
rect 7124 6345 7190 6379
rect 7124 6311 7140 6345
rect 7174 6311 7190 6345
rect 7124 6277 7190 6311
rect 7124 6243 7140 6277
rect 7174 6243 7190 6277
rect 7124 6209 7190 6243
rect 7124 6175 7140 6209
rect 7174 6175 7190 6209
rect 7124 6141 7190 6175
rect 7124 6107 7140 6141
rect 7174 6107 7190 6141
rect 7124 6073 7190 6107
rect 7124 6039 7140 6073
rect 7174 6039 7190 6073
rect 7124 6005 7190 6039
rect 7124 5971 7140 6005
rect 7174 5971 7190 6005
rect 7124 5937 7190 5971
rect 7124 5903 7140 5937
rect 7174 5903 7190 5937
rect 7124 5869 7190 5903
rect 7124 5835 7140 5869
rect 7174 5835 7190 5869
rect 7124 5801 7190 5835
rect 7124 5767 7140 5801
rect 7174 5767 7190 5801
rect 7124 5733 7190 5767
rect 7124 5699 7140 5733
rect 7174 5699 7190 5733
rect 7124 5665 7190 5699
rect 7124 5631 7140 5665
rect 7174 5631 7190 5665
rect 7124 5590 7190 5631
rect 7220 6549 7286 6590
rect 7220 6515 7236 6549
rect 7270 6515 7286 6549
rect 7220 6481 7286 6515
rect 7220 6447 7236 6481
rect 7270 6447 7286 6481
rect 7220 6413 7286 6447
rect 7220 6379 7236 6413
rect 7270 6379 7286 6413
rect 7220 6345 7286 6379
rect 7220 6311 7236 6345
rect 7270 6311 7286 6345
rect 7220 6277 7286 6311
rect 7220 6243 7236 6277
rect 7270 6243 7286 6277
rect 7220 6209 7286 6243
rect 7220 6175 7236 6209
rect 7270 6175 7286 6209
rect 7220 6141 7286 6175
rect 7220 6107 7236 6141
rect 7270 6107 7286 6141
rect 7220 6073 7286 6107
rect 7220 6039 7236 6073
rect 7270 6039 7286 6073
rect 7220 6005 7286 6039
rect 7220 5971 7236 6005
rect 7270 5971 7286 6005
rect 7220 5937 7286 5971
rect 7220 5903 7236 5937
rect 7270 5903 7286 5937
rect 7220 5869 7286 5903
rect 7220 5835 7236 5869
rect 7270 5835 7286 5869
rect 7220 5801 7286 5835
rect 7220 5767 7236 5801
rect 7270 5767 7286 5801
rect 7220 5733 7286 5767
rect 7220 5699 7236 5733
rect 7270 5699 7286 5733
rect 7220 5665 7286 5699
rect 7220 5631 7236 5665
rect 7270 5631 7286 5665
rect 7220 5590 7286 5631
rect 7316 6549 7378 6590
rect 7316 6515 7332 6549
rect 7366 6515 7378 6549
rect 7316 6481 7378 6515
rect 7316 6447 7332 6481
rect 7366 6447 7378 6481
rect 7316 6413 7378 6447
rect 7316 6379 7332 6413
rect 7366 6379 7378 6413
rect 7316 6345 7378 6379
rect 7316 6311 7332 6345
rect 7366 6311 7378 6345
rect 7316 6277 7378 6311
rect 7316 6243 7332 6277
rect 7366 6243 7378 6277
rect 7316 6209 7378 6243
rect 7316 6175 7332 6209
rect 7366 6175 7378 6209
rect 7316 6141 7378 6175
rect 7316 6107 7332 6141
rect 7366 6107 7378 6141
rect 7316 6073 7378 6107
rect 7316 6039 7332 6073
rect 7366 6039 7378 6073
rect 7316 6005 7378 6039
rect 7316 5971 7332 6005
rect 7366 5971 7378 6005
rect 7316 5937 7378 5971
rect 7316 5903 7332 5937
rect 7366 5903 7378 5937
rect 7316 5869 7378 5903
rect 7316 5835 7332 5869
rect 7366 5835 7378 5869
rect 7316 5801 7378 5835
rect 7316 5767 7332 5801
rect 7366 5767 7378 5801
rect 7316 5733 7378 5767
rect 7316 5699 7332 5733
rect 7366 5699 7378 5733
rect 7316 5665 7378 5699
rect 7316 5631 7332 5665
rect 7366 5631 7378 5665
rect 7316 5590 7378 5631
rect 7934 6545 7996 6586
rect 7934 6511 7946 6545
rect 7980 6511 7996 6545
rect 7934 6477 7996 6511
rect 7934 6443 7946 6477
rect 7980 6443 7996 6477
rect 7934 6409 7996 6443
rect 7934 6375 7946 6409
rect 7980 6375 7996 6409
rect 7934 6341 7996 6375
rect 7934 6307 7946 6341
rect 7980 6307 7996 6341
rect 7934 6273 7996 6307
rect 7934 6239 7946 6273
rect 7980 6239 7996 6273
rect 7934 6205 7996 6239
rect 7934 6171 7946 6205
rect 7980 6171 7996 6205
rect 7934 6137 7996 6171
rect 7934 6103 7946 6137
rect 7980 6103 7996 6137
rect 7934 6069 7996 6103
rect 7934 6035 7946 6069
rect 7980 6035 7996 6069
rect 7934 6001 7996 6035
rect 7934 5967 7946 6001
rect 7980 5967 7996 6001
rect 7934 5933 7996 5967
rect 7934 5899 7946 5933
rect 7980 5899 7996 5933
rect 7934 5865 7996 5899
rect 7934 5831 7946 5865
rect 7980 5831 7996 5865
rect 7934 5797 7996 5831
rect 7934 5763 7946 5797
rect 7980 5763 7996 5797
rect 7934 5729 7996 5763
rect 7934 5695 7946 5729
rect 7980 5695 7996 5729
rect 7934 5661 7996 5695
rect 7934 5627 7946 5661
rect 7980 5627 7996 5661
rect 7934 5586 7996 5627
rect 8026 6545 8092 6586
rect 8026 6511 8042 6545
rect 8076 6511 8092 6545
rect 8026 6477 8092 6511
rect 8026 6443 8042 6477
rect 8076 6443 8092 6477
rect 8026 6409 8092 6443
rect 8026 6375 8042 6409
rect 8076 6375 8092 6409
rect 8026 6341 8092 6375
rect 8026 6307 8042 6341
rect 8076 6307 8092 6341
rect 8026 6273 8092 6307
rect 8026 6239 8042 6273
rect 8076 6239 8092 6273
rect 8026 6205 8092 6239
rect 8026 6171 8042 6205
rect 8076 6171 8092 6205
rect 8026 6137 8092 6171
rect 8026 6103 8042 6137
rect 8076 6103 8092 6137
rect 8026 6069 8092 6103
rect 8026 6035 8042 6069
rect 8076 6035 8092 6069
rect 8026 6001 8092 6035
rect 8026 5967 8042 6001
rect 8076 5967 8092 6001
rect 8026 5933 8092 5967
rect 8026 5899 8042 5933
rect 8076 5899 8092 5933
rect 8026 5865 8092 5899
rect 8026 5831 8042 5865
rect 8076 5831 8092 5865
rect 8026 5797 8092 5831
rect 8026 5763 8042 5797
rect 8076 5763 8092 5797
rect 8026 5729 8092 5763
rect 8026 5695 8042 5729
rect 8076 5695 8092 5729
rect 8026 5661 8092 5695
rect 8026 5627 8042 5661
rect 8076 5627 8092 5661
rect 8026 5586 8092 5627
rect 8122 6545 8188 6586
rect 8122 6511 8138 6545
rect 8172 6511 8188 6545
rect 8122 6477 8188 6511
rect 8122 6443 8138 6477
rect 8172 6443 8188 6477
rect 8122 6409 8188 6443
rect 8122 6375 8138 6409
rect 8172 6375 8188 6409
rect 8122 6341 8188 6375
rect 8122 6307 8138 6341
rect 8172 6307 8188 6341
rect 8122 6273 8188 6307
rect 8122 6239 8138 6273
rect 8172 6239 8188 6273
rect 8122 6205 8188 6239
rect 8122 6171 8138 6205
rect 8172 6171 8188 6205
rect 8122 6137 8188 6171
rect 8122 6103 8138 6137
rect 8172 6103 8188 6137
rect 8122 6069 8188 6103
rect 8122 6035 8138 6069
rect 8172 6035 8188 6069
rect 8122 6001 8188 6035
rect 8122 5967 8138 6001
rect 8172 5967 8188 6001
rect 8122 5933 8188 5967
rect 8122 5899 8138 5933
rect 8172 5899 8188 5933
rect 8122 5865 8188 5899
rect 8122 5831 8138 5865
rect 8172 5831 8188 5865
rect 8122 5797 8188 5831
rect 8122 5763 8138 5797
rect 8172 5763 8188 5797
rect 8122 5729 8188 5763
rect 8122 5695 8138 5729
rect 8172 5695 8188 5729
rect 8122 5661 8188 5695
rect 8122 5627 8138 5661
rect 8172 5627 8188 5661
rect 8122 5586 8188 5627
rect 8218 6545 8284 6586
rect 8218 6511 8234 6545
rect 8268 6511 8284 6545
rect 8218 6477 8284 6511
rect 8218 6443 8234 6477
rect 8268 6443 8284 6477
rect 8218 6409 8284 6443
rect 8218 6375 8234 6409
rect 8268 6375 8284 6409
rect 8218 6341 8284 6375
rect 8218 6307 8234 6341
rect 8268 6307 8284 6341
rect 8218 6273 8284 6307
rect 8218 6239 8234 6273
rect 8268 6239 8284 6273
rect 8218 6205 8284 6239
rect 8218 6171 8234 6205
rect 8268 6171 8284 6205
rect 8218 6137 8284 6171
rect 8218 6103 8234 6137
rect 8268 6103 8284 6137
rect 8218 6069 8284 6103
rect 8218 6035 8234 6069
rect 8268 6035 8284 6069
rect 8218 6001 8284 6035
rect 8218 5967 8234 6001
rect 8268 5967 8284 6001
rect 8218 5933 8284 5967
rect 8218 5899 8234 5933
rect 8268 5899 8284 5933
rect 8218 5865 8284 5899
rect 8218 5831 8234 5865
rect 8268 5831 8284 5865
rect 8218 5797 8284 5831
rect 8218 5763 8234 5797
rect 8268 5763 8284 5797
rect 8218 5729 8284 5763
rect 8218 5695 8234 5729
rect 8268 5695 8284 5729
rect 8218 5661 8284 5695
rect 8218 5627 8234 5661
rect 8268 5627 8284 5661
rect 8218 5586 8284 5627
rect 8314 6545 8380 6586
rect 8314 6511 8330 6545
rect 8364 6511 8380 6545
rect 8314 6477 8380 6511
rect 8314 6443 8330 6477
rect 8364 6443 8380 6477
rect 8314 6409 8380 6443
rect 8314 6375 8330 6409
rect 8364 6375 8380 6409
rect 8314 6341 8380 6375
rect 8314 6307 8330 6341
rect 8364 6307 8380 6341
rect 8314 6273 8380 6307
rect 8314 6239 8330 6273
rect 8364 6239 8380 6273
rect 8314 6205 8380 6239
rect 8314 6171 8330 6205
rect 8364 6171 8380 6205
rect 8314 6137 8380 6171
rect 8314 6103 8330 6137
rect 8364 6103 8380 6137
rect 8314 6069 8380 6103
rect 8314 6035 8330 6069
rect 8364 6035 8380 6069
rect 8314 6001 8380 6035
rect 8314 5967 8330 6001
rect 8364 5967 8380 6001
rect 8314 5933 8380 5967
rect 8314 5899 8330 5933
rect 8364 5899 8380 5933
rect 8314 5865 8380 5899
rect 8314 5831 8330 5865
rect 8364 5831 8380 5865
rect 8314 5797 8380 5831
rect 8314 5763 8330 5797
rect 8364 5763 8380 5797
rect 8314 5729 8380 5763
rect 8314 5695 8330 5729
rect 8364 5695 8380 5729
rect 8314 5661 8380 5695
rect 8314 5627 8330 5661
rect 8364 5627 8380 5661
rect 8314 5586 8380 5627
rect 8410 6545 8476 6586
rect 8410 6511 8426 6545
rect 8460 6511 8476 6545
rect 8410 6477 8476 6511
rect 8410 6443 8426 6477
rect 8460 6443 8476 6477
rect 8410 6409 8476 6443
rect 8410 6375 8426 6409
rect 8460 6375 8476 6409
rect 8410 6341 8476 6375
rect 8410 6307 8426 6341
rect 8460 6307 8476 6341
rect 8410 6273 8476 6307
rect 8410 6239 8426 6273
rect 8460 6239 8476 6273
rect 8410 6205 8476 6239
rect 8410 6171 8426 6205
rect 8460 6171 8476 6205
rect 8410 6137 8476 6171
rect 8410 6103 8426 6137
rect 8460 6103 8476 6137
rect 8410 6069 8476 6103
rect 8410 6035 8426 6069
rect 8460 6035 8476 6069
rect 8410 6001 8476 6035
rect 8410 5967 8426 6001
rect 8460 5967 8476 6001
rect 8410 5933 8476 5967
rect 8410 5899 8426 5933
rect 8460 5899 8476 5933
rect 8410 5865 8476 5899
rect 8410 5831 8426 5865
rect 8460 5831 8476 5865
rect 8410 5797 8476 5831
rect 8410 5763 8426 5797
rect 8460 5763 8476 5797
rect 8410 5729 8476 5763
rect 8410 5695 8426 5729
rect 8460 5695 8476 5729
rect 8410 5661 8476 5695
rect 8410 5627 8426 5661
rect 8460 5627 8476 5661
rect 8410 5586 8476 5627
rect 8506 6545 8572 6586
rect 8506 6511 8522 6545
rect 8556 6511 8572 6545
rect 8506 6477 8572 6511
rect 8506 6443 8522 6477
rect 8556 6443 8572 6477
rect 8506 6409 8572 6443
rect 8506 6375 8522 6409
rect 8556 6375 8572 6409
rect 8506 6341 8572 6375
rect 8506 6307 8522 6341
rect 8556 6307 8572 6341
rect 8506 6273 8572 6307
rect 8506 6239 8522 6273
rect 8556 6239 8572 6273
rect 8506 6205 8572 6239
rect 8506 6171 8522 6205
rect 8556 6171 8572 6205
rect 8506 6137 8572 6171
rect 8506 6103 8522 6137
rect 8556 6103 8572 6137
rect 8506 6069 8572 6103
rect 8506 6035 8522 6069
rect 8556 6035 8572 6069
rect 8506 6001 8572 6035
rect 8506 5967 8522 6001
rect 8556 5967 8572 6001
rect 8506 5933 8572 5967
rect 8506 5899 8522 5933
rect 8556 5899 8572 5933
rect 8506 5865 8572 5899
rect 8506 5831 8522 5865
rect 8556 5831 8572 5865
rect 8506 5797 8572 5831
rect 8506 5763 8522 5797
rect 8556 5763 8572 5797
rect 8506 5729 8572 5763
rect 8506 5695 8522 5729
rect 8556 5695 8572 5729
rect 8506 5661 8572 5695
rect 8506 5627 8522 5661
rect 8556 5627 8572 5661
rect 8506 5586 8572 5627
rect 8602 6545 8668 6586
rect 8602 6511 8618 6545
rect 8652 6511 8668 6545
rect 8602 6477 8668 6511
rect 8602 6443 8618 6477
rect 8652 6443 8668 6477
rect 8602 6409 8668 6443
rect 8602 6375 8618 6409
rect 8652 6375 8668 6409
rect 8602 6341 8668 6375
rect 8602 6307 8618 6341
rect 8652 6307 8668 6341
rect 8602 6273 8668 6307
rect 8602 6239 8618 6273
rect 8652 6239 8668 6273
rect 8602 6205 8668 6239
rect 8602 6171 8618 6205
rect 8652 6171 8668 6205
rect 8602 6137 8668 6171
rect 8602 6103 8618 6137
rect 8652 6103 8668 6137
rect 8602 6069 8668 6103
rect 8602 6035 8618 6069
rect 8652 6035 8668 6069
rect 8602 6001 8668 6035
rect 8602 5967 8618 6001
rect 8652 5967 8668 6001
rect 8602 5933 8668 5967
rect 8602 5899 8618 5933
rect 8652 5899 8668 5933
rect 8602 5865 8668 5899
rect 8602 5831 8618 5865
rect 8652 5831 8668 5865
rect 8602 5797 8668 5831
rect 8602 5763 8618 5797
rect 8652 5763 8668 5797
rect 8602 5729 8668 5763
rect 8602 5695 8618 5729
rect 8652 5695 8668 5729
rect 8602 5661 8668 5695
rect 8602 5627 8618 5661
rect 8652 5627 8668 5661
rect 8602 5586 8668 5627
rect 8698 6545 8760 6586
rect 8698 6511 8714 6545
rect 8748 6511 8760 6545
rect 8698 6477 8760 6511
rect 8698 6443 8714 6477
rect 8748 6443 8760 6477
rect 8698 6409 8760 6443
rect 8698 6375 8714 6409
rect 8748 6375 8760 6409
rect 8698 6341 8760 6375
rect 8698 6307 8714 6341
rect 8748 6307 8760 6341
rect 8698 6273 8760 6307
rect 8698 6239 8714 6273
rect 8748 6239 8760 6273
rect 8698 6205 8760 6239
rect 8698 6171 8714 6205
rect 8748 6171 8760 6205
rect 8698 6137 8760 6171
rect 8698 6103 8714 6137
rect 8748 6103 8760 6137
rect 8698 6069 8760 6103
rect 8698 6035 8714 6069
rect 8748 6035 8760 6069
rect 8698 6001 8760 6035
rect 8698 5967 8714 6001
rect 8748 5967 8760 6001
rect 8698 5933 8760 5967
rect 8698 5899 8714 5933
rect 8748 5899 8760 5933
rect 8698 5865 8760 5899
rect 8698 5831 8714 5865
rect 8748 5831 8760 5865
rect 8698 5797 8760 5831
rect 8698 5763 8714 5797
rect 8748 5763 8760 5797
rect 8698 5729 8760 5763
rect 8698 5695 8714 5729
rect 8748 5695 8760 5729
rect 8698 5661 8760 5695
rect 8698 5627 8714 5661
rect 8748 5627 8760 5661
rect 8698 5586 8760 5627
rect 9256 6547 9318 6588
rect 9256 6513 9268 6547
rect 9302 6513 9318 6547
rect 9256 6479 9318 6513
rect 9256 6445 9268 6479
rect 9302 6445 9318 6479
rect 9256 6411 9318 6445
rect 9256 6377 9268 6411
rect 9302 6377 9318 6411
rect 9256 6343 9318 6377
rect 9256 6309 9268 6343
rect 9302 6309 9318 6343
rect 9256 6275 9318 6309
rect 9256 6241 9268 6275
rect 9302 6241 9318 6275
rect 9256 6207 9318 6241
rect 9256 6173 9268 6207
rect 9302 6173 9318 6207
rect 9256 6139 9318 6173
rect 9256 6105 9268 6139
rect 9302 6105 9318 6139
rect 9256 6071 9318 6105
rect 9256 6037 9268 6071
rect 9302 6037 9318 6071
rect 9256 6003 9318 6037
rect 9256 5969 9268 6003
rect 9302 5969 9318 6003
rect 9256 5935 9318 5969
rect 9256 5901 9268 5935
rect 9302 5901 9318 5935
rect 9256 5867 9318 5901
rect 9256 5833 9268 5867
rect 9302 5833 9318 5867
rect 9256 5799 9318 5833
rect 9256 5765 9268 5799
rect 9302 5765 9318 5799
rect 9256 5731 9318 5765
rect 9256 5697 9268 5731
rect 9302 5697 9318 5731
rect 9256 5663 9318 5697
rect 9256 5629 9268 5663
rect 9302 5629 9318 5663
rect 9256 5588 9318 5629
rect 9348 6547 9414 6588
rect 9348 6513 9364 6547
rect 9398 6513 9414 6547
rect 9348 6479 9414 6513
rect 9348 6445 9364 6479
rect 9398 6445 9414 6479
rect 9348 6411 9414 6445
rect 9348 6377 9364 6411
rect 9398 6377 9414 6411
rect 9348 6343 9414 6377
rect 9348 6309 9364 6343
rect 9398 6309 9414 6343
rect 9348 6275 9414 6309
rect 9348 6241 9364 6275
rect 9398 6241 9414 6275
rect 9348 6207 9414 6241
rect 9348 6173 9364 6207
rect 9398 6173 9414 6207
rect 9348 6139 9414 6173
rect 9348 6105 9364 6139
rect 9398 6105 9414 6139
rect 9348 6071 9414 6105
rect 9348 6037 9364 6071
rect 9398 6037 9414 6071
rect 9348 6003 9414 6037
rect 9348 5969 9364 6003
rect 9398 5969 9414 6003
rect 9348 5935 9414 5969
rect 9348 5901 9364 5935
rect 9398 5901 9414 5935
rect 9348 5867 9414 5901
rect 9348 5833 9364 5867
rect 9398 5833 9414 5867
rect 9348 5799 9414 5833
rect 9348 5765 9364 5799
rect 9398 5765 9414 5799
rect 9348 5731 9414 5765
rect 9348 5697 9364 5731
rect 9398 5697 9414 5731
rect 9348 5663 9414 5697
rect 9348 5629 9364 5663
rect 9398 5629 9414 5663
rect 9348 5588 9414 5629
rect 9444 6547 9510 6588
rect 9444 6513 9460 6547
rect 9494 6513 9510 6547
rect 9444 6479 9510 6513
rect 9444 6445 9460 6479
rect 9494 6445 9510 6479
rect 9444 6411 9510 6445
rect 9444 6377 9460 6411
rect 9494 6377 9510 6411
rect 9444 6343 9510 6377
rect 9444 6309 9460 6343
rect 9494 6309 9510 6343
rect 9444 6275 9510 6309
rect 9444 6241 9460 6275
rect 9494 6241 9510 6275
rect 9444 6207 9510 6241
rect 9444 6173 9460 6207
rect 9494 6173 9510 6207
rect 9444 6139 9510 6173
rect 9444 6105 9460 6139
rect 9494 6105 9510 6139
rect 9444 6071 9510 6105
rect 9444 6037 9460 6071
rect 9494 6037 9510 6071
rect 9444 6003 9510 6037
rect 9444 5969 9460 6003
rect 9494 5969 9510 6003
rect 9444 5935 9510 5969
rect 9444 5901 9460 5935
rect 9494 5901 9510 5935
rect 9444 5867 9510 5901
rect 9444 5833 9460 5867
rect 9494 5833 9510 5867
rect 9444 5799 9510 5833
rect 9444 5765 9460 5799
rect 9494 5765 9510 5799
rect 9444 5731 9510 5765
rect 9444 5697 9460 5731
rect 9494 5697 9510 5731
rect 9444 5663 9510 5697
rect 9444 5629 9460 5663
rect 9494 5629 9510 5663
rect 9444 5588 9510 5629
rect 9540 6547 9606 6588
rect 9540 6513 9556 6547
rect 9590 6513 9606 6547
rect 9540 6479 9606 6513
rect 9540 6445 9556 6479
rect 9590 6445 9606 6479
rect 9540 6411 9606 6445
rect 9540 6377 9556 6411
rect 9590 6377 9606 6411
rect 9540 6343 9606 6377
rect 9540 6309 9556 6343
rect 9590 6309 9606 6343
rect 9540 6275 9606 6309
rect 9540 6241 9556 6275
rect 9590 6241 9606 6275
rect 9540 6207 9606 6241
rect 9540 6173 9556 6207
rect 9590 6173 9606 6207
rect 9540 6139 9606 6173
rect 9540 6105 9556 6139
rect 9590 6105 9606 6139
rect 9540 6071 9606 6105
rect 9540 6037 9556 6071
rect 9590 6037 9606 6071
rect 9540 6003 9606 6037
rect 9540 5969 9556 6003
rect 9590 5969 9606 6003
rect 9540 5935 9606 5969
rect 9540 5901 9556 5935
rect 9590 5901 9606 5935
rect 9540 5867 9606 5901
rect 9540 5833 9556 5867
rect 9590 5833 9606 5867
rect 9540 5799 9606 5833
rect 9540 5765 9556 5799
rect 9590 5765 9606 5799
rect 9540 5731 9606 5765
rect 9540 5697 9556 5731
rect 9590 5697 9606 5731
rect 9540 5663 9606 5697
rect 9540 5629 9556 5663
rect 9590 5629 9606 5663
rect 9540 5588 9606 5629
rect 9636 6547 9702 6588
rect 9636 6513 9652 6547
rect 9686 6513 9702 6547
rect 9636 6479 9702 6513
rect 9636 6445 9652 6479
rect 9686 6445 9702 6479
rect 9636 6411 9702 6445
rect 9636 6377 9652 6411
rect 9686 6377 9702 6411
rect 9636 6343 9702 6377
rect 9636 6309 9652 6343
rect 9686 6309 9702 6343
rect 9636 6275 9702 6309
rect 9636 6241 9652 6275
rect 9686 6241 9702 6275
rect 9636 6207 9702 6241
rect 9636 6173 9652 6207
rect 9686 6173 9702 6207
rect 9636 6139 9702 6173
rect 9636 6105 9652 6139
rect 9686 6105 9702 6139
rect 9636 6071 9702 6105
rect 9636 6037 9652 6071
rect 9686 6037 9702 6071
rect 9636 6003 9702 6037
rect 9636 5969 9652 6003
rect 9686 5969 9702 6003
rect 9636 5935 9702 5969
rect 9636 5901 9652 5935
rect 9686 5901 9702 5935
rect 9636 5867 9702 5901
rect 9636 5833 9652 5867
rect 9686 5833 9702 5867
rect 9636 5799 9702 5833
rect 9636 5765 9652 5799
rect 9686 5765 9702 5799
rect 9636 5731 9702 5765
rect 9636 5697 9652 5731
rect 9686 5697 9702 5731
rect 9636 5663 9702 5697
rect 9636 5629 9652 5663
rect 9686 5629 9702 5663
rect 9636 5588 9702 5629
rect 9732 6547 9798 6588
rect 9732 6513 9748 6547
rect 9782 6513 9798 6547
rect 9732 6479 9798 6513
rect 9732 6445 9748 6479
rect 9782 6445 9798 6479
rect 9732 6411 9798 6445
rect 9732 6377 9748 6411
rect 9782 6377 9798 6411
rect 9732 6343 9798 6377
rect 9732 6309 9748 6343
rect 9782 6309 9798 6343
rect 9732 6275 9798 6309
rect 9732 6241 9748 6275
rect 9782 6241 9798 6275
rect 9732 6207 9798 6241
rect 9732 6173 9748 6207
rect 9782 6173 9798 6207
rect 9732 6139 9798 6173
rect 9732 6105 9748 6139
rect 9782 6105 9798 6139
rect 9732 6071 9798 6105
rect 9732 6037 9748 6071
rect 9782 6037 9798 6071
rect 9732 6003 9798 6037
rect 9732 5969 9748 6003
rect 9782 5969 9798 6003
rect 9732 5935 9798 5969
rect 9732 5901 9748 5935
rect 9782 5901 9798 5935
rect 9732 5867 9798 5901
rect 9732 5833 9748 5867
rect 9782 5833 9798 5867
rect 9732 5799 9798 5833
rect 9732 5765 9748 5799
rect 9782 5765 9798 5799
rect 9732 5731 9798 5765
rect 9732 5697 9748 5731
rect 9782 5697 9798 5731
rect 9732 5663 9798 5697
rect 9732 5629 9748 5663
rect 9782 5629 9798 5663
rect 9732 5588 9798 5629
rect 9828 6547 9894 6588
rect 9828 6513 9844 6547
rect 9878 6513 9894 6547
rect 9828 6479 9894 6513
rect 9828 6445 9844 6479
rect 9878 6445 9894 6479
rect 9828 6411 9894 6445
rect 9828 6377 9844 6411
rect 9878 6377 9894 6411
rect 9828 6343 9894 6377
rect 9828 6309 9844 6343
rect 9878 6309 9894 6343
rect 9828 6275 9894 6309
rect 9828 6241 9844 6275
rect 9878 6241 9894 6275
rect 9828 6207 9894 6241
rect 9828 6173 9844 6207
rect 9878 6173 9894 6207
rect 9828 6139 9894 6173
rect 9828 6105 9844 6139
rect 9878 6105 9894 6139
rect 9828 6071 9894 6105
rect 9828 6037 9844 6071
rect 9878 6037 9894 6071
rect 9828 6003 9894 6037
rect 9828 5969 9844 6003
rect 9878 5969 9894 6003
rect 9828 5935 9894 5969
rect 9828 5901 9844 5935
rect 9878 5901 9894 5935
rect 9828 5867 9894 5901
rect 9828 5833 9844 5867
rect 9878 5833 9894 5867
rect 9828 5799 9894 5833
rect 9828 5765 9844 5799
rect 9878 5765 9894 5799
rect 9828 5731 9894 5765
rect 9828 5697 9844 5731
rect 9878 5697 9894 5731
rect 9828 5663 9894 5697
rect 9828 5629 9844 5663
rect 9878 5629 9894 5663
rect 9828 5588 9894 5629
rect 9924 6547 9990 6588
rect 9924 6513 9940 6547
rect 9974 6513 9990 6547
rect 9924 6479 9990 6513
rect 9924 6445 9940 6479
rect 9974 6445 9990 6479
rect 9924 6411 9990 6445
rect 9924 6377 9940 6411
rect 9974 6377 9990 6411
rect 9924 6343 9990 6377
rect 9924 6309 9940 6343
rect 9974 6309 9990 6343
rect 9924 6275 9990 6309
rect 9924 6241 9940 6275
rect 9974 6241 9990 6275
rect 9924 6207 9990 6241
rect 9924 6173 9940 6207
rect 9974 6173 9990 6207
rect 9924 6139 9990 6173
rect 9924 6105 9940 6139
rect 9974 6105 9990 6139
rect 9924 6071 9990 6105
rect 9924 6037 9940 6071
rect 9974 6037 9990 6071
rect 9924 6003 9990 6037
rect 9924 5969 9940 6003
rect 9974 5969 9990 6003
rect 9924 5935 9990 5969
rect 9924 5901 9940 5935
rect 9974 5901 9990 5935
rect 9924 5867 9990 5901
rect 9924 5833 9940 5867
rect 9974 5833 9990 5867
rect 9924 5799 9990 5833
rect 9924 5765 9940 5799
rect 9974 5765 9990 5799
rect 9924 5731 9990 5765
rect 9924 5697 9940 5731
rect 9974 5697 9990 5731
rect 9924 5663 9990 5697
rect 9924 5629 9940 5663
rect 9974 5629 9990 5663
rect 9924 5588 9990 5629
rect 10020 6547 10086 6588
rect 10020 6513 10036 6547
rect 10070 6513 10086 6547
rect 10020 6479 10086 6513
rect 10020 6445 10036 6479
rect 10070 6445 10086 6479
rect 10020 6411 10086 6445
rect 10020 6377 10036 6411
rect 10070 6377 10086 6411
rect 10020 6343 10086 6377
rect 10020 6309 10036 6343
rect 10070 6309 10086 6343
rect 10020 6275 10086 6309
rect 10020 6241 10036 6275
rect 10070 6241 10086 6275
rect 10020 6207 10086 6241
rect 10020 6173 10036 6207
rect 10070 6173 10086 6207
rect 10020 6139 10086 6173
rect 10020 6105 10036 6139
rect 10070 6105 10086 6139
rect 10020 6071 10086 6105
rect 10020 6037 10036 6071
rect 10070 6037 10086 6071
rect 10020 6003 10086 6037
rect 10020 5969 10036 6003
rect 10070 5969 10086 6003
rect 10020 5935 10086 5969
rect 10020 5901 10036 5935
rect 10070 5901 10086 5935
rect 10020 5867 10086 5901
rect 10020 5833 10036 5867
rect 10070 5833 10086 5867
rect 10020 5799 10086 5833
rect 10020 5765 10036 5799
rect 10070 5765 10086 5799
rect 10020 5731 10086 5765
rect 10020 5697 10036 5731
rect 10070 5697 10086 5731
rect 10020 5663 10086 5697
rect 10020 5629 10036 5663
rect 10070 5629 10086 5663
rect 10020 5588 10086 5629
rect 10116 6547 10182 6588
rect 10116 6513 10132 6547
rect 10166 6513 10182 6547
rect 10116 6479 10182 6513
rect 10116 6445 10132 6479
rect 10166 6445 10182 6479
rect 10116 6411 10182 6445
rect 10116 6377 10132 6411
rect 10166 6377 10182 6411
rect 10116 6343 10182 6377
rect 10116 6309 10132 6343
rect 10166 6309 10182 6343
rect 10116 6275 10182 6309
rect 10116 6241 10132 6275
rect 10166 6241 10182 6275
rect 10116 6207 10182 6241
rect 10116 6173 10132 6207
rect 10166 6173 10182 6207
rect 10116 6139 10182 6173
rect 10116 6105 10132 6139
rect 10166 6105 10182 6139
rect 10116 6071 10182 6105
rect 10116 6037 10132 6071
rect 10166 6037 10182 6071
rect 10116 6003 10182 6037
rect 10116 5969 10132 6003
rect 10166 5969 10182 6003
rect 10116 5935 10182 5969
rect 10116 5901 10132 5935
rect 10166 5901 10182 5935
rect 10116 5867 10182 5901
rect 10116 5833 10132 5867
rect 10166 5833 10182 5867
rect 10116 5799 10182 5833
rect 10116 5765 10132 5799
rect 10166 5765 10182 5799
rect 10116 5731 10182 5765
rect 10116 5697 10132 5731
rect 10166 5697 10182 5731
rect 10116 5663 10182 5697
rect 10116 5629 10132 5663
rect 10166 5629 10182 5663
rect 10116 5588 10182 5629
rect 10212 6547 10278 6588
rect 10212 6513 10228 6547
rect 10262 6513 10278 6547
rect 10212 6479 10278 6513
rect 10212 6445 10228 6479
rect 10262 6445 10278 6479
rect 10212 6411 10278 6445
rect 10212 6377 10228 6411
rect 10262 6377 10278 6411
rect 10212 6343 10278 6377
rect 10212 6309 10228 6343
rect 10262 6309 10278 6343
rect 10212 6275 10278 6309
rect 10212 6241 10228 6275
rect 10262 6241 10278 6275
rect 10212 6207 10278 6241
rect 10212 6173 10228 6207
rect 10262 6173 10278 6207
rect 10212 6139 10278 6173
rect 10212 6105 10228 6139
rect 10262 6105 10278 6139
rect 10212 6071 10278 6105
rect 10212 6037 10228 6071
rect 10262 6037 10278 6071
rect 10212 6003 10278 6037
rect 10212 5969 10228 6003
rect 10262 5969 10278 6003
rect 10212 5935 10278 5969
rect 10212 5901 10228 5935
rect 10262 5901 10278 5935
rect 10212 5867 10278 5901
rect 10212 5833 10228 5867
rect 10262 5833 10278 5867
rect 10212 5799 10278 5833
rect 10212 5765 10228 5799
rect 10262 5765 10278 5799
rect 10212 5731 10278 5765
rect 10212 5697 10228 5731
rect 10262 5697 10278 5731
rect 10212 5663 10278 5697
rect 10212 5629 10228 5663
rect 10262 5629 10278 5663
rect 10212 5588 10278 5629
rect 10308 6547 10374 6588
rect 10308 6513 10324 6547
rect 10358 6513 10374 6547
rect 10308 6479 10374 6513
rect 10308 6445 10324 6479
rect 10358 6445 10374 6479
rect 10308 6411 10374 6445
rect 10308 6377 10324 6411
rect 10358 6377 10374 6411
rect 10308 6343 10374 6377
rect 10308 6309 10324 6343
rect 10358 6309 10374 6343
rect 10308 6275 10374 6309
rect 10308 6241 10324 6275
rect 10358 6241 10374 6275
rect 10308 6207 10374 6241
rect 10308 6173 10324 6207
rect 10358 6173 10374 6207
rect 10308 6139 10374 6173
rect 10308 6105 10324 6139
rect 10358 6105 10374 6139
rect 10308 6071 10374 6105
rect 10308 6037 10324 6071
rect 10358 6037 10374 6071
rect 10308 6003 10374 6037
rect 10308 5969 10324 6003
rect 10358 5969 10374 6003
rect 10308 5935 10374 5969
rect 10308 5901 10324 5935
rect 10358 5901 10374 5935
rect 10308 5867 10374 5901
rect 10308 5833 10324 5867
rect 10358 5833 10374 5867
rect 10308 5799 10374 5833
rect 10308 5765 10324 5799
rect 10358 5765 10374 5799
rect 10308 5731 10374 5765
rect 10308 5697 10324 5731
rect 10358 5697 10374 5731
rect 10308 5663 10374 5697
rect 10308 5629 10324 5663
rect 10358 5629 10374 5663
rect 10308 5588 10374 5629
rect 10404 6547 10466 6588
rect 10404 6513 10420 6547
rect 10454 6513 10466 6547
rect 10404 6479 10466 6513
rect 10404 6445 10420 6479
rect 10454 6445 10466 6479
rect 10404 6411 10466 6445
rect 10404 6377 10420 6411
rect 10454 6377 10466 6411
rect 10404 6343 10466 6377
rect 10404 6309 10420 6343
rect 10454 6309 10466 6343
rect 10404 6275 10466 6309
rect 10404 6241 10420 6275
rect 10454 6241 10466 6275
rect 10404 6207 10466 6241
rect 10404 6173 10420 6207
rect 10454 6173 10466 6207
rect 10404 6139 10466 6173
rect 10404 6105 10420 6139
rect 10454 6105 10466 6139
rect 10404 6071 10466 6105
rect 10404 6037 10420 6071
rect 10454 6037 10466 6071
rect 10404 6003 10466 6037
rect 10404 5969 10420 6003
rect 10454 5969 10466 6003
rect 10404 5935 10466 5969
rect 10404 5901 10420 5935
rect 10454 5901 10466 5935
rect 10404 5867 10466 5901
rect 10404 5833 10420 5867
rect 10454 5833 10466 5867
rect 10404 5799 10466 5833
rect 10404 5765 10420 5799
rect 10454 5765 10466 5799
rect 10404 5731 10466 5765
rect 10404 5697 10420 5731
rect 10454 5697 10466 5731
rect 10404 5663 10466 5697
rect 10404 5629 10420 5663
rect 10454 5629 10466 5663
rect 10404 5588 10466 5629
rect 11022 6543 11084 6584
rect 11022 6509 11034 6543
rect 11068 6509 11084 6543
rect 11022 6475 11084 6509
rect 11022 6441 11034 6475
rect 11068 6441 11084 6475
rect 11022 6407 11084 6441
rect 11022 6373 11034 6407
rect 11068 6373 11084 6407
rect 11022 6339 11084 6373
rect 11022 6305 11034 6339
rect 11068 6305 11084 6339
rect 11022 6271 11084 6305
rect 11022 6237 11034 6271
rect 11068 6237 11084 6271
rect 11022 6203 11084 6237
rect 11022 6169 11034 6203
rect 11068 6169 11084 6203
rect 11022 6135 11084 6169
rect 11022 6101 11034 6135
rect 11068 6101 11084 6135
rect 11022 6067 11084 6101
rect 11022 6033 11034 6067
rect 11068 6033 11084 6067
rect 11022 5999 11084 6033
rect 11022 5965 11034 5999
rect 11068 5965 11084 5999
rect 11022 5931 11084 5965
rect 11022 5897 11034 5931
rect 11068 5897 11084 5931
rect 11022 5863 11084 5897
rect 11022 5829 11034 5863
rect 11068 5829 11084 5863
rect 11022 5795 11084 5829
rect 11022 5761 11034 5795
rect 11068 5761 11084 5795
rect 11022 5727 11084 5761
rect 11022 5693 11034 5727
rect 11068 5693 11084 5727
rect 11022 5659 11084 5693
rect 11022 5625 11034 5659
rect 11068 5625 11084 5659
rect 11022 5584 11084 5625
rect 11114 6543 11180 6584
rect 11114 6509 11130 6543
rect 11164 6509 11180 6543
rect 11114 6475 11180 6509
rect 11114 6441 11130 6475
rect 11164 6441 11180 6475
rect 11114 6407 11180 6441
rect 11114 6373 11130 6407
rect 11164 6373 11180 6407
rect 11114 6339 11180 6373
rect 11114 6305 11130 6339
rect 11164 6305 11180 6339
rect 11114 6271 11180 6305
rect 11114 6237 11130 6271
rect 11164 6237 11180 6271
rect 11114 6203 11180 6237
rect 11114 6169 11130 6203
rect 11164 6169 11180 6203
rect 11114 6135 11180 6169
rect 11114 6101 11130 6135
rect 11164 6101 11180 6135
rect 11114 6067 11180 6101
rect 11114 6033 11130 6067
rect 11164 6033 11180 6067
rect 11114 5999 11180 6033
rect 11114 5965 11130 5999
rect 11164 5965 11180 5999
rect 11114 5931 11180 5965
rect 11114 5897 11130 5931
rect 11164 5897 11180 5931
rect 11114 5863 11180 5897
rect 11114 5829 11130 5863
rect 11164 5829 11180 5863
rect 11114 5795 11180 5829
rect 11114 5761 11130 5795
rect 11164 5761 11180 5795
rect 11114 5727 11180 5761
rect 11114 5693 11130 5727
rect 11164 5693 11180 5727
rect 11114 5659 11180 5693
rect 11114 5625 11130 5659
rect 11164 5625 11180 5659
rect 11114 5584 11180 5625
rect 11210 6543 11276 6584
rect 11210 6509 11226 6543
rect 11260 6509 11276 6543
rect 11210 6475 11276 6509
rect 11210 6441 11226 6475
rect 11260 6441 11276 6475
rect 11210 6407 11276 6441
rect 11210 6373 11226 6407
rect 11260 6373 11276 6407
rect 11210 6339 11276 6373
rect 11210 6305 11226 6339
rect 11260 6305 11276 6339
rect 11210 6271 11276 6305
rect 11210 6237 11226 6271
rect 11260 6237 11276 6271
rect 11210 6203 11276 6237
rect 11210 6169 11226 6203
rect 11260 6169 11276 6203
rect 11210 6135 11276 6169
rect 11210 6101 11226 6135
rect 11260 6101 11276 6135
rect 11210 6067 11276 6101
rect 11210 6033 11226 6067
rect 11260 6033 11276 6067
rect 11210 5999 11276 6033
rect 11210 5965 11226 5999
rect 11260 5965 11276 5999
rect 11210 5931 11276 5965
rect 11210 5897 11226 5931
rect 11260 5897 11276 5931
rect 11210 5863 11276 5897
rect 11210 5829 11226 5863
rect 11260 5829 11276 5863
rect 11210 5795 11276 5829
rect 11210 5761 11226 5795
rect 11260 5761 11276 5795
rect 11210 5727 11276 5761
rect 11210 5693 11226 5727
rect 11260 5693 11276 5727
rect 11210 5659 11276 5693
rect 11210 5625 11226 5659
rect 11260 5625 11276 5659
rect 11210 5584 11276 5625
rect 11306 6543 11372 6584
rect 11306 6509 11322 6543
rect 11356 6509 11372 6543
rect 11306 6475 11372 6509
rect 11306 6441 11322 6475
rect 11356 6441 11372 6475
rect 11306 6407 11372 6441
rect 11306 6373 11322 6407
rect 11356 6373 11372 6407
rect 11306 6339 11372 6373
rect 11306 6305 11322 6339
rect 11356 6305 11372 6339
rect 11306 6271 11372 6305
rect 11306 6237 11322 6271
rect 11356 6237 11372 6271
rect 11306 6203 11372 6237
rect 11306 6169 11322 6203
rect 11356 6169 11372 6203
rect 11306 6135 11372 6169
rect 11306 6101 11322 6135
rect 11356 6101 11372 6135
rect 11306 6067 11372 6101
rect 11306 6033 11322 6067
rect 11356 6033 11372 6067
rect 11306 5999 11372 6033
rect 11306 5965 11322 5999
rect 11356 5965 11372 5999
rect 11306 5931 11372 5965
rect 11306 5897 11322 5931
rect 11356 5897 11372 5931
rect 11306 5863 11372 5897
rect 11306 5829 11322 5863
rect 11356 5829 11372 5863
rect 11306 5795 11372 5829
rect 11306 5761 11322 5795
rect 11356 5761 11372 5795
rect 11306 5727 11372 5761
rect 11306 5693 11322 5727
rect 11356 5693 11372 5727
rect 11306 5659 11372 5693
rect 11306 5625 11322 5659
rect 11356 5625 11372 5659
rect 11306 5584 11372 5625
rect 11402 6543 11468 6584
rect 11402 6509 11418 6543
rect 11452 6509 11468 6543
rect 11402 6475 11468 6509
rect 11402 6441 11418 6475
rect 11452 6441 11468 6475
rect 11402 6407 11468 6441
rect 11402 6373 11418 6407
rect 11452 6373 11468 6407
rect 11402 6339 11468 6373
rect 11402 6305 11418 6339
rect 11452 6305 11468 6339
rect 11402 6271 11468 6305
rect 11402 6237 11418 6271
rect 11452 6237 11468 6271
rect 11402 6203 11468 6237
rect 11402 6169 11418 6203
rect 11452 6169 11468 6203
rect 11402 6135 11468 6169
rect 11402 6101 11418 6135
rect 11452 6101 11468 6135
rect 11402 6067 11468 6101
rect 11402 6033 11418 6067
rect 11452 6033 11468 6067
rect 11402 5999 11468 6033
rect 11402 5965 11418 5999
rect 11452 5965 11468 5999
rect 11402 5931 11468 5965
rect 11402 5897 11418 5931
rect 11452 5897 11468 5931
rect 11402 5863 11468 5897
rect 11402 5829 11418 5863
rect 11452 5829 11468 5863
rect 11402 5795 11468 5829
rect 11402 5761 11418 5795
rect 11452 5761 11468 5795
rect 11402 5727 11468 5761
rect 11402 5693 11418 5727
rect 11452 5693 11468 5727
rect 11402 5659 11468 5693
rect 11402 5625 11418 5659
rect 11452 5625 11468 5659
rect 11402 5584 11468 5625
rect 11498 6543 11564 6584
rect 11498 6509 11514 6543
rect 11548 6509 11564 6543
rect 11498 6475 11564 6509
rect 11498 6441 11514 6475
rect 11548 6441 11564 6475
rect 11498 6407 11564 6441
rect 11498 6373 11514 6407
rect 11548 6373 11564 6407
rect 11498 6339 11564 6373
rect 11498 6305 11514 6339
rect 11548 6305 11564 6339
rect 11498 6271 11564 6305
rect 11498 6237 11514 6271
rect 11548 6237 11564 6271
rect 11498 6203 11564 6237
rect 11498 6169 11514 6203
rect 11548 6169 11564 6203
rect 11498 6135 11564 6169
rect 11498 6101 11514 6135
rect 11548 6101 11564 6135
rect 11498 6067 11564 6101
rect 11498 6033 11514 6067
rect 11548 6033 11564 6067
rect 11498 5999 11564 6033
rect 11498 5965 11514 5999
rect 11548 5965 11564 5999
rect 11498 5931 11564 5965
rect 11498 5897 11514 5931
rect 11548 5897 11564 5931
rect 11498 5863 11564 5897
rect 11498 5829 11514 5863
rect 11548 5829 11564 5863
rect 11498 5795 11564 5829
rect 11498 5761 11514 5795
rect 11548 5761 11564 5795
rect 11498 5727 11564 5761
rect 11498 5693 11514 5727
rect 11548 5693 11564 5727
rect 11498 5659 11564 5693
rect 11498 5625 11514 5659
rect 11548 5625 11564 5659
rect 11498 5584 11564 5625
rect 11594 6543 11660 6584
rect 11594 6509 11610 6543
rect 11644 6509 11660 6543
rect 11594 6475 11660 6509
rect 11594 6441 11610 6475
rect 11644 6441 11660 6475
rect 11594 6407 11660 6441
rect 11594 6373 11610 6407
rect 11644 6373 11660 6407
rect 11594 6339 11660 6373
rect 11594 6305 11610 6339
rect 11644 6305 11660 6339
rect 11594 6271 11660 6305
rect 11594 6237 11610 6271
rect 11644 6237 11660 6271
rect 11594 6203 11660 6237
rect 11594 6169 11610 6203
rect 11644 6169 11660 6203
rect 11594 6135 11660 6169
rect 11594 6101 11610 6135
rect 11644 6101 11660 6135
rect 11594 6067 11660 6101
rect 11594 6033 11610 6067
rect 11644 6033 11660 6067
rect 11594 5999 11660 6033
rect 11594 5965 11610 5999
rect 11644 5965 11660 5999
rect 11594 5931 11660 5965
rect 11594 5897 11610 5931
rect 11644 5897 11660 5931
rect 11594 5863 11660 5897
rect 11594 5829 11610 5863
rect 11644 5829 11660 5863
rect 11594 5795 11660 5829
rect 11594 5761 11610 5795
rect 11644 5761 11660 5795
rect 11594 5727 11660 5761
rect 11594 5693 11610 5727
rect 11644 5693 11660 5727
rect 11594 5659 11660 5693
rect 11594 5625 11610 5659
rect 11644 5625 11660 5659
rect 11594 5584 11660 5625
rect 11690 6543 11756 6584
rect 11690 6509 11706 6543
rect 11740 6509 11756 6543
rect 11690 6475 11756 6509
rect 11690 6441 11706 6475
rect 11740 6441 11756 6475
rect 11690 6407 11756 6441
rect 11690 6373 11706 6407
rect 11740 6373 11756 6407
rect 11690 6339 11756 6373
rect 11690 6305 11706 6339
rect 11740 6305 11756 6339
rect 11690 6271 11756 6305
rect 11690 6237 11706 6271
rect 11740 6237 11756 6271
rect 11690 6203 11756 6237
rect 11690 6169 11706 6203
rect 11740 6169 11756 6203
rect 11690 6135 11756 6169
rect 11690 6101 11706 6135
rect 11740 6101 11756 6135
rect 11690 6067 11756 6101
rect 11690 6033 11706 6067
rect 11740 6033 11756 6067
rect 11690 5999 11756 6033
rect 11690 5965 11706 5999
rect 11740 5965 11756 5999
rect 11690 5931 11756 5965
rect 11690 5897 11706 5931
rect 11740 5897 11756 5931
rect 11690 5863 11756 5897
rect 11690 5829 11706 5863
rect 11740 5829 11756 5863
rect 11690 5795 11756 5829
rect 11690 5761 11706 5795
rect 11740 5761 11756 5795
rect 11690 5727 11756 5761
rect 11690 5693 11706 5727
rect 11740 5693 11756 5727
rect 11690 5659 11756 5693
rect 11690 5625 11706 5659
rect 11740 5625 11756 5659
rect 11690 5584 11756 5625
rect 11786 6543 11848 6584
rect 11786 6509 11802 6543
rect 11836 6509 11848 6543
rect 11786 6475 11848 6509
rect 11786 6441 11802 6475
rect 11836 6441 11848 6475
rect 11786 6407 11848 6441
rect 11786 6373 11802 6407
rect 11836 6373 11848 6407
rect 11786 6339 11848 6373
rect 11786 6305 11802 6339
rect 11836 6305 11848 6339
rect 11786 6271 11848 6305
rect 11786 6237 11802 6271
rect 11836 6237 11848 6271
rect 11786 6203 11848 6237
rect 11786 6169 11802 6203
rect 11836 6169 11848 6203
rect 11786 6135 11848 6169
rect 11786 6101 11802 6135
rect 11836 6101 11848 6135
rect 11786 6067 11848 6101
rect 11786 6033 11802 6067
rect 11836 6033 11848 6067
rect 11786 5999 11848 6033
rect 11786 5965 11802 5999
rect 11836 5965 11848 5999
rect 11786 5931 11848 5965
rect 11786 5897 11802 5931
rect 11836 5897 11848 5931
rect 11786 5863 11848 5897
rect 11786 5829 11802 5863
rect 11836 5829 11848 5863
rect 11786 5795 11848 5829
rect 11786 5761 11802 5795
rect 11836 5761 11848 5795
rect 11786 5727 11848 5761
rect 11786 5693 11802 5727
rect 11836 5693 11848 5727
rect 11786 5659 11848 5693
rect 11786 5625 11802 5659
rect 11836 5625 11848 5659
rect 11786 5584 11848 5625
rect 12412 6521 12474 6562
rect 12412 6487 12424 6521
rect 12458 6487 12474 6521
rect 12412 6453 12474 6487
rect 12412 6419 12424 6453
rect 12458 6419 12474 6453
rect 12412 6385 12474 6419
rect 12412 6351 12424 6385
rect 12458 6351 12474 6385
rect 12412 6317 12474 6351
rect 12412 6283 12424 6317
rect 12458 6283 12474 6317
rect 12412 6249 12474 6283
rect 12412 6215 12424 6249
rect 12458 6215 12474 6249
rect 12412 6181 12474 6215
rect 12412 6147 12424 6181
rect 12458 6147 12474 6181
rect 12412 6113 12474 6147
rect 12412 6079 12424 6113
rect 12458 6079 12474 6113
rect 12412 6045 12474 6079
rect 12412 6011 12424 6045
rect 12458 6011 12474 6045
rect 12412 5977 12474 6011
rect 12412 5943 12424 5977
rect 12458 5943 12474 5977
rect 12412 5909 12474 5943
rect 12412 5875 12424 5909
rect 12458 5875 12474 5909
rect 12412 5841 12474 5875
rect 12412 5807 12424 5841
rect 12458 5807 12474 5841
rect 12412 5773 12474 5807
rect 12412 5739 12424 5773
rect 12458 5739 12474 5773
rect 12412 5705 12474 5739
rect 12412 5671 12424 5705
rect 12458 5671 12474 5705
rect 12412 5637 12474 5671
rect 12412 5603 12424 5637
rect 12458 5603 12474 5637
rect 12412 5562 12474 5603
rect 12504 6521 12570 6562
rect 12504 6487 12520 6521
rect 12554 6487 12570 6521
rect 12504 6453 12570 6487
rect 12504 6419 12520 6453
rect 12554 6419 12570 6453
rect 12504 6385 12570 6419
rect 12504 6351 12520 6385
rect 12554 6351 12570 6385
rect 12504 6317 12570 6351
rect 12504 6283 12520 6317
rect 12554 6283 12570 6317
rect 12504 6249 12570 6283
rect 12504 6215 12520 6249
rect 12554 6215 12570 6249
rect 12504 6181 12570 6215
rect 12504 6147 12520 6181
rect 12554 6147 12570 6181
rect 12504 6113 12570 6147
rect 12504 6079 12520 6113
rect 12554 6079 12570 6113
rect 12504 6045 12570 6079
rect 12504 6011 12520 6045
rect 12554 6011 12570 6045
rect 12504 5977 12570 6011
rect 12504 5943 12520 5977
rect 12554 5943 12570 5977
rect 12504 5909 12570 5943
rect 12504 5875 12520 5909
rect 12554 5875 12570 5909
rect 12504 5841 12570 5875
rect 12504 5807 12520 5841
rect 12554 5807 12570 5841
rect 12504 5773 12570 5807
rect 12504 5739 12520 5773
rect 12554 5739 12570 5773
rect 12504 5705 12570 5739
rect 12504 5671 12520 5705
rect 12554 5671 12570 5705
rect 12504 5637 12570 5671
rect 12504 5603 12520 5637
rect 12554 5603 12570 5637
rect 12504 5562 12570 5603
rect 12600 6521 12666 6562
rect 12600 6487 12616 6521
rect 12650 6487 12666 6521
rect 12600 6453 12666 6487
rect 12600 6419 12616 6453
rect 12650 6419 12666 6453
rect 12600 6385 12666 6419
rect 12600 6351 12616 6385
rect 12650 6351 12666 6385
rect 12600 6317 12666 6351
rect 12600 6283 12616 6317
rect 12650 6283 12666 6317
rect 12600 6249 12666 6283
rect 12600 6215 12616 6249
rect 12650 6215 12666 6249
rect 12600 6181 12666 6215
rect 12600 6147 12616 6181
rect 12650 6147 12666 6181
rect 12600 6113 12666 6147
rect 12600 6079 12616 6113
rect 12650 6079 12666 6113
rect 12600 6045 12666 6079
rect 12600 6011 12616 6045
rect 12650 6011 12666 6045
rect 12600 5977 12666 6011
rect 12600 5943 12616 5977
rect 12650 5943 12666 5977
rect 12600 5909 12666 5943
rect 12600 5875 12616 5909
rect 12650 5875 12666 5909
rect 12600 5841 12666 5875
rect 12600 5807 12616 5841
rect 12650 5807 12666 5841
rect 12600 5773 12666 5807
rect 12600 5739 12616 5773
rect 12650 5739 12666 5773
rect 12600 5705 12666 5739
rect 12600 5671 12616 5705
rect 12650 5671 12666 5705
rect 12600 5637 12666 5671
rect 12600 5603 12616 5637
rect 12650 5603 12666 5637
rect 12600 5562 12666 5603
rect 12696 6521 12762 6562
rect 12696 6487 12712 6521
rect 12746 6487 12762 6521
rect 12696 6453 12762 6487
rect 12696 6419 12712 6453
rect 12746 6419 12762 6453
rect 12696 6385 12762 6419
rect 12696 6351 12712 6385
rect 12746 6351 12762 6385
rect 12696 6317 12762 6351
rect 12696 6283 12712 6317
rect 12746 6283 12762 6317
rect 12696 6249 12762 6283
rect 12696 6215 12712 6249
rect 12746 6215 12762 6249
rect 12696 6181 12762 6215
rect 12696 6147 12712 6181
rect 12746 6147 12762 6181
rect 12696 6113 12762 6147
rect 12696 6079 12712 6113
rect 12746 6079 12762 6113
rect 12696 6045 12762 6079
rect 12696 6011 12712 6045
rect 12746 6011 12762 6045
rect 12696 5977 12762 6011
rect 12696 5943 12712 5977
rect 12746 5943 12762 5977
rect 12696 5909 12762 5943
rect 12696 5875 12712 5909
rect 12746 5875 12762 5909
rect 12696 5841 12762 5875
rect 12696 5807 12712 5841
rect 12746 5807 12762 5841
rect 12696 5773 12762 5807
rect 12696 5739 12712 5773
rect 12746 5739 12762 5773
rect 12696 5705 12762 5739
rect 12696 5671 12712 5705
rect 12746 5671 12762 5705
rect 12696 5637 12762 5671
rect 12696 5603 12712 5637
rect 12746 5603 12762 5637
rect 12696 5562 12762 5603
rect 12792 6521 12858 6562
rect 12792 6487 12808 6521
rect 12842 6487 12858 6521
rect 12792 6453 12858 6487
rect 12792 6419 12808 6453
rect 12842 6419 12858 6453
rect 12792 6385 12858 6419
rect 12792 6351 12808 6385
rect 12842 6351 12858 6385
rect 12792 6317 12858 6351
rect 12792 6283 12808 6317
rect 12842 6283 12858 6317
rect 12792 6249 12858 6283
rect 12792 6215 12808 6249
rect 12842 6215 12858 6249
rect 12792 6181 12858 6215
rect 12792 6147 12808 6181
rect 12842 6147 12858 6181
rect 12792 6113 12858 6147
rect 12792 6079 12808 6113
rect 12842 6079 12858 6113
rect 12792 6045 12858 6079
rect 12792 6011 12808 6045
rect 12842 6011 12858 6045
rect 12792 5977 12858 6011
rect 12792 5943 12808 5977
rect 12842 5943 12858 5977
rect 12792 5909 12858 5943
rect 12792 5875 12808 5909
rect 12842 5875 12858 5909
rect 12792 5841 12858 5875
rect 12792 5807 12808 5841
rect 12842 5807 12858 5841
rect 12792 5773 12858 5807
rect 12792 5739 12808 5773
rect 12842 5739 12858 5773
rect 12792 5705 12858 5739
rect 12792 5671 12808 5705
rect 12842 5671 12858 5705
rect 12792 5637 12858 5671
rect 12792 5603 12808 5637
rect 12842 5603 12858 5637
rect 12792 5562 12858 5603
rect 12888 6521 12954 6562
rect 12888 6487 12904 6521
rect 12938 6487 12954 6521
rect 12888 6453 12954 6487
rect 12888 6419 12904 6453
rect 12938 6419 12954 6453
rect 12888 6385 12954 6419
rect 12888 6351 12904 6385
rect 12938 6351 12954 6385
rect 12888 6317 12954 6351
rect 12888 6283 12904 6317
rect 12938 6283 12954 6317
rect 12888 6249 12954 6283
rect 12888 6215 12904 6249
rect 12938 6215 12954 6249
rect 12888 6181 12954 6215
rect 12888 6147 12904 6181
rect 12938 6147 12954 6181
rect 12888 6113 12954 6147
rect 12888 6079 12904 6113
rect 12938 6079 12954 6113
rect 12888 6045 12954 6079
rect 12888 6011 12904 6045
rect 12938 6011 12954 6045
rect 12888 5977 12954 6011
rect 12888 5943 12904 5977
rect 12938 5943 12954 5977
rect 12888 5909 12954 5943
rect 12888 5875 12904 5909
rect 12938 5875 12954 5909
rect 12888 5841 12954 5875
rect 12888 5807 12904 5841
rect 12938 5807 12954 5841
rect 12888 5773 12954 5807
rect 12888 5739 12904 5773
rect 12938 5739 12954 5773
rect 12888 5705 12954 5739
rect 12888 5671 12904 5705
rect 12938 5671 12954 5705
rect 12888 5637 12954 5671
rect 12888 5603 12904 5637
rect 12938 5603 12954 5637
rect 12888 5562 12954 5603
rect 12984 6521 13050 6562
rect 12984 6487 13000 6521
rect 13034 6487 13050 6521
rect 12984 6453 13050 6487
rect 12984 6419 13000 6453
rect 13034 6419 13050 6453
rect 12984 6385 13050 6419
rect 12984 6351 13000 6385
rect 13034 6351 13050 6385
rect 12984 6317 13050 6351
rect 12984 6283 13000 6317
rect 13034 6283 13050 6317
rect 12984 6249 13050 6283
rect 12984 6215 13000 6249
rect 13034 6215 13050 6249
rect 12984 6181 13050 6215
rect 12984 6147 13000 6181
rect 13034 6147 13050 6181
rect 12984 6113 13050 6147
rect 12984 6079 13000 6113
rect 13034 6079 13050 6113
rect 12984 6045 13050 6079
rect 12984 6011 13000 6045
rect 13034 6011 13050 6045
rect 12984 5977 13050 6011
rect 12984 5943 13000 5977
rect 13034 5943 13050 5977
rect 12984 5909 13050 5943
rect 12984 5875 13000 5909
rect 13034 5875 13050 5909
rect 12984 5841 13050 5875
rect 12984 5807 13000 5841
rect 13034 5807 13050 5841
rect 12984 5773 13050 5807
rect 12984 5739 13000 5773
rect 13034 5739 13050 5773
rect 12984 5705 13050 5739
rect 12984 5671 13000 5705
rect 13034 5671 13050 5705
rect 12984 5637 13050 5671
rect 12984 5603 13000 5637
rect 13034 5603 13050 5637
rect 12984 5562 13050 5603
rect 13080 6521 13146 6562
rect 13080 6487 13096 6521
rect 13130 6487 13146 6521
rect 13080 6453 13146 6487
rect 13080 6419 13096 6453
rect 13130 6419 13146 6453
rect 13080 6385 13146 6419
rect 13080 6351 13096 6385
rect 13130 6351 13146 6385
rect 13080 6317 13146 6351
rect 13080 6283 13096 6317
rect 13130 6283 13146 6317
rect 13080 6249 13146 6283
rect 13080 6215 13096 6249
rect 13130 6215 13146 6249
rect 13080 6181 13146 6215
rect 13080 6147 13096 6181
rect 13130 6147 13146 6181
rect 13080 6113 13146 6147
rect 13080 6079 13096 6113
rect 13130 6079 13146 6113
rect 13080 6045 13146 6079
rect 13080 6011 13096 6045
rect 13130 6011 13146 6045
rect 13080 5977 13146 6011
rect 13080 5943 13096 5977
rect 13130 5943 13146 5977
rect 13080 5909 13146 5943
rect 13080 5875 13096 5909
rect 13130 5875 13146 5909
rect 13080 5841 13146 5875
rect 13080 5807 13096 5841
rect 13130 5807 13146 5841
rect 13080 5773 13146 5807
rect 13080 5739 13096 5773
rect 13130 5739 13146 5773
rect 13080 5705 13146 5739
rect 13080 5671 13096 5705
rect 13130 5671 13146 5705
rect 13080 5637 13146 5671
rect 13080 5603 13096 5637
rect 13130 5603 13146 5637
rect 13080 5562 13146 5603
rect 13176 6521 13242 6562
rect 13176 6487 13192 6521
rect 13226 6487 13242 6521
rect 13176 6453 13242 6487
rect 13176 6419 13192 6453
rect 13226 6419 13242 6453
rect 13176 6385 13242 6419
rect 13176 6351 13192 6385
rect 13226 6351 13242 6385
rect 13176 6317 13242 6351
rect 13176 6283 13192 6317
rect 13226 6283 13242 6317
rect 13176 6249 13242 6283
rect 13176 6215 13192 6249
rect 13226 6215 13242 6249
rect 13176 6181 13242 6215
rect 13176 6147 13192 6181
rect 13226 6147 13242 6181
rect 13176 6113 13242 6147
rect 13176 6079 13192 6113
rect 13226 6079 13242 6113
rect 13176 6045 13242 6079
rect 13176 6011 13192 6045
rect 13226 6011 13242 6045
rect 13176 5977 13242 6011
rect 13176 5943 13192 5977
rect 13226 5943 13242 5977
rect 13176 5909 13242 5943
rect 13176 5875 13192 5909
rect 13226 5875 13242 5909
rect 13176 5841 13242 5875
rect 13176 5807 13192 5841
rect 13226 5807 13242 5841
rect 13176 5773 13242 5807
rect 13176 5739 13192 5773
rect 13226 5739 13242 5773
rect 13176 5705 13242 5739
rect 13176 5671 13192 5705
rect 13226 5671 13242 5705
rect 13176 5637 13242 5671
rect 13176 5603 13192 5637
rect 13226 5603 13242 5637
rect 13176 5562 13242 5603
rect 13272 6521 13338 6562
rect 13272 6487 13288 6521
rect 13322 6487 13338 6521
rect 13272 6453 13338 6487
rect 13272 6419 13288 6453
rect 13322 6419 13338 6453
rect 13272 6385 13338 6419
rect 13272 6351 13288 6385
rect 13322 6351 13338 6385
rect 13272 6317 13338 6351
rect 13272 6283 13288 6317
rect 13322 6283 13338 6317
rect 13272 6249 13338 6283
rect 13272 6215 13288 6249
rect 13322 6215 13338 6249
rect 13272 6181 13338 6215
rect 13272 6147 13288 6181
rect 13322 6147 13338 6181
rect 13272 6113 13338 6147
rect 13272 6079 13288 6113
rect 13322 6079 13338 6113
rect 13272 6045 13338 6079
rect 13272 6011 13288 6045
rect 13322 6011 13338 6045
rect 13272 5977 13338 6011
rect 13272 5943 13288 5977
rect 13322 5943 13338 5977
rect 13272 5909 13338 5943
rect 13272 5875 13288 5909
rect 13322 5875 13338 5909
rect 13272 5841 13338 5875
rect 13272 5807 13288 5841
rect 13322 5807 13338 5841
rect 13272 5773 13338 5807
rect 13272 5739 13288 5773
rect 13322 5739 13338 5773
rect 13272 5705 13338 5739
rect 13272 5671 13288 5705
rect 13322 5671 13338 5705
rect 13272 5637 13338 5671
rect 13272 5603 13288 5637
rect 13322 5603 13338 5637
rect 13272 5562 13338 5603
rect 13368 6521 13434 6562
rect 13368 6487 13384 6521
rect 13418 6487 13434 6521
rect 13368 6453 13434 6487
rect 13368 6419 13384 6453
rect 13418 6419 13434 6453
rect 13368 6385 13434 6419
rect 13368 6351 13384 6385
rect 13418 6351 13434 6385
rect 13368 6317 13434 6351
rect 13368 6283 13384 6317
rect 13418 6283 13434 6317
rect 13368 6249 13434 6283
rect 13368 6215 13384 6249
rect 13418 6215 13434 6249
rect 13368 6181 13434 6215
rect 13368 6147 13384 6181
rect 13418 6147 13434 6181
rect 13368 6113 13434 6147
rect 13368 6079 13384 6113
rect 13418 6079 13434 6113
rect 13368 6045 13434 6079
rect 13368 6011 13384 6045
rect 13418 6011 13434 6045
rect 13368 5977 13434 6011
rect 13368 5943 13384 5977
rect 13418 5943 13434 5977
rect 13368 5909 13434 5943
rect 13368 5875 13384 5909
rect 13418 5875 13434 5909
rect 13368 5841 13434 5875
rect 13368 5807 13384 5841
rect 13418 5807 13434 5841
rect 13368 5773 13434 5807
rect 13368 5739 13384 5773
rect 13418 5739 13434 5773
rect 13368 5705 13434 5739
rect 13368 5671 13384 5705
rect 13418 5671 13434 5705
rect 13368 5637 13434 5671
rect 13368 5603 13384 5637
rect 13418 5603 13434 5637
rect 13368 5562 13434 5603
rect 13464 6521 13530 6562
rect 13464 6487 13480 6521
rect 13514 6487 13530 6521
rect 13464 6453 13530 6487
rect 13464 6419 13480 6453
rect 13514 6419 13530 6453
rect 13464 6385 13530 6419
rect 13464 6351 13480 6385
rect 13514 6351 13530 6385
rect 13464 6317 13530 6351
rect 13464 6283 13480 6317
rect 13514 6283 13530 6317
rect 13464 6249 13530 6283
rect 13464 6215 13480 6249
rect 13514 6215 13530 6249
rect 13464 6181 13530 6215
rect 13464 6147 13480 6181
rect 13514 6147 13530 6181
rect 13464 6113 13530 6147
rect 13464 6079 13480 6113
rect 13514 6079 13530 6113
rect 13464 6045 13530 6079
rect 13464 6011 13480 6045
rect 13514 6011 13530 6045
rect 13464 5977 13530 6011
rect 13464 5943 13480 5977
rect 13514 5943 13530 5977
rect 13464 5909 13530 5943
rect 13464 5875 13480 5909
rect 13514 5875 13530 5909
rect 13464 5841 13530 5875
rect 13464 5807 13480 5841
rect 13514 5807 13530 5841
rect 13464 5773 13530 5807
rect 13464 5739 13480 5773
rect 13514 5739 13530 5773
rect 13464 5705 13530 5739
rect 13464 5671 13480 5705
rect 13514 5671 13530 5705
rect 13464 5637 13530 5671
rect 13464 5603 13480 5637
rect 13514 5603 13530 5637
rect 13464 5562 13530 5603
rect 13560 6521 13622 6562
rect 13560 6487 13576 6521
rect 13610 6487 13622 6521
rect 13560 6453 13622 6487
rect 13560 6419 13576 6453
rect 13610 6419 13622 6453
rect 13560 6385 13622 6419
rect 13560 6351 13576 6385
rect 13610 6351 13622 6385
rect 13560 6317 13622 6351
rect 13560 6283 13576 6317
rect 13610 6283 13622 6317
rect 13560 6249 13622 6283
rect 13560 6215 13576 6249
rect 13610 6215 13622 6249
rect 13560 6181 13622 6215
rect 13560 6147 13576 6181
rect 13610 6147 13622 6181
rect 13560 6113 13622 6147
rect 13560 6079 13576 6113
rect 13610 6079 13622 6113
rect 13560 6045 13622 6079
rect 13560 6011 13576 6045
rect 13610 6011 13622 6045
rect 13560 5977 13622 6011
rect 13560 5943 13576 5977
rect 13610 5943 13622 5977
rect 13560 5909 13622 5943
rect 13560 5875 13576 5909
rect 13610 5875 13622 5909
rect 13560 5841 13622 5875
rect 13560 5807 13576 5841
rect 13610 5807 13622 5841
rect 13560 5773 13622 5807
rect 13560 5739 13576 5773
rect 13610 5739 13622 5773
rect 13560 5705 13622 5739
rect 13560 5671 13576 5705
rect 13610 5671 13622 5705
rect 13560 5637 13622 5671
rect 13560 5603 13576 5637
rect 13610 5603 13622 5637
rect 13560 5562 13622 5603
rect 14178 6517 14240 6558
rect 14178 6483 14190 6517
rect 14224 6483 14240 6517
rect 14178 6449 14240 6483
rect 14178 6415 14190 6449
rect 14224 6415 14240 6449
rect 14178 6381 14240 6415
rect 14178 6347 14190 6381
rect 14224 6347 14240 6381
rect 14178 6313 14240 6347
rect 14178 6279 14190 6313
rect 14224 6279 14240 6313
rect 14178 6245 14240 6279
rect 14178 6211 14190 6245
rect 14224 6211 14240 6245
rect 14178 6177 14240 6211
rect 14178 6143 14190 6177
rect 14224 6143 14240 6177
rect 14178 6109 14240 6143
rect 14178 6075 14190 6109
rect 14224 6075 14240 6109
rect 14178 6041 14240 6075
rect 14178 6007 14190 6041
rect 14224 6007 14240 6041
rect 14178 5973 14240 6007
rect 14178 5939 14190 5973
rect 14224 5939 14240 5973
rect 14178 5905 14240 5939
rect 14178 5871 14190 5905
rect 14224 5871 14240 5905
rect 14178 5837 14240 5871
rect 14178 5803 14190 5837
rect 14224 5803 14240 5837
rect 14178 5769 14240 5803
rect 14178 5735 14190 5769
rect 14224 5735 14240 5769
rect 14178 5701 14240 5735
rect 14178 5667 14190 5701
rect 14224 5667 14240 5701
rect 14178 5633 14240 5667
rect 14178 5599 14190 5633
rect 14224 5599 14240 5633
rect -880 5521 -868 5555
rect -834 5521 -822 5555
rect 14178 5558 14240 5599
rect 14270 6517 14336 6558
rect 14270 6483 14286 6517
rect 14320 6483 14336 6517
rect 14270 6449 14336 6483
rect 14270 6415 14286 6449
rect 14320 6415 14336 6449
rect 14270 6381 14336 6415
rect 14270 6347 14286 6381
rect 14320 6347 14336 6381
rect 14270 6313 14336 6347
rect 14270 6279 14286 6313
rect 14320 6279 14336 6313
rect 14270 6245 14336 6279
rect 14270 6211 14286 6245
rect 14320 6211 14336 6245
rect 14270 6177 14336 6211
rect 14270 6143 14286 6177
rect 14320 6143 14336 6177
rect 14270 6109 14336 6143
rect 14270 6075 14286 6109
rect 14320 6075 14336 6109
rect 14270 6041 14336 6075
rect 14270 6007 14286 6041
rect 14320 6007 14336 6041
rect 14270 5973 14336 6007
rect 14270 5939 14286 5973
rect 14320 5939 14336 5973
rect 14270 5905 14336 5939
rect 14270 5871 14286 5905
rect 14320 5871 14336 5905
rect 14270 5837 14336 5871
rect 14270 5803 14286 5837
rect 14320 5803 14336 5837
rect 14270 5769 14336 5803
rect 14270 5735 14286 5769
rect 14320 5735 14336 5769
rect 14270 5701 14336 5735
rect 14270 5667 14286 5701
rect 14320 5667 14336 5701
rect 14270 5633 14336 5667
rect 14270 5599 14286 5633
rect 14320 5599 14336 5633
rect 14270 5558 14336 5599
rect 14366 6517 14432 6558
rect 14366 6483 14382 6517
rect 14416 6483 14432 6517
rect 14366 6449 14432 6483
rect 14366 6415 14382 6449
rect 14416 6415 14432 6449
rect 14366 6381 14432 6415
rect 14366 6347 14382 6381
rect 14416 6347 14432 6381
rect 14366 6313 14432 6347
rect 14366 6279 14382 6313
rect 14416 6279 14432 6313
rect 14366 6245 14432 6279
rect 14366 6211 14382 6245
rect 14416 6211 14432 6245
rect 14366 6177 14432 6211
rect 14366 6143 14382 6177
rect 14416 6143 14432 6177
rect 14366 6109 14432 6143
rect 14366 6075 14382 6109
rect 14416 6075 14432 6109
rect 14366 6041 14432 6075
rect 14366 6007 14382 6041
rect 14416 6007 14432 6041
rect 14366 5973 14432 6007
rect 14366 5939 14382 5973
rect 14416 5939 14432 5973
rect 14366 5905 14432 5939
rect 14366 5871 14382 5905
rect 14416 5871 14432 5905
rect 14366 5837 14432 5871
rect 14366 5803 14382 5837
rect 14416 5803 14432 5837
rect 14366 5769 14432 5803
rect 14366 5735 14382 5769
rect 14416 5735 14432 5769
rect 14366 5701 14432 5735
rect 14366 5667 14382 5701
rect 14416 5667 14432 5701
rect 14366 5633 14432 5667
rect 14366 5599 14382 5633
rect 14416 5599 14432 5633
rect 14366 5558 14432 5599
rect 14462 6517 14528 6558
rect 14462 6483 14478 6517
rect 14512 6483 14528 6517
rect 14462 6449 14528 6483
rect 14462 6415 14478 6449
rect 14512 6415 14528 6449
rect 14462 6381 14528 6415
rect 14462 6347 14478 6381
rect 14512 6347 14528 6381
rect 14462 6313 14528 6347
rect 14462 6279 14478 6313
rect 14512 6279 14528 6313
rect 14462 6245 14528 6279
rect 14462 6211 14478 6245
rect 14512 6211 14528 6245
rect 14462 6177 14528 6211
rect 14462 6143 14478 6177
rect 14512 6143 14528 6177
rect 14462 6109 14528 6143
rect 14462 6075 14478 6109
rect 14512 6075 14528 6109
rect 14462 6041 14528 6075
rect 14462 6007 14478 6041
rect 14512 6007 14528 6041
rect 14462 5973 14528 6007
rect 14462 5939 14478 5973
rect 14512 5939 14528 5973
rect 14462 5905 14528 5939
rect 14462 5871 14478 5905
rect 14512 5871 14528 5905
rect 14462 5837 14528 5871
rect 14462 5803 14478 5837
rect 14512 5803 14528 5837
rect 14462 5769 14528 5803
rect 14462 5735 14478 5769
rect 14512 5735 14528 5769
rect 14462 5701 14528 5735
rect 14462 5667 14478 5701
rect 14512 5667 14528 5701
rect 14462 5633 14528 5667
rect 14462 5599 14478 5633
rect 14512 5599 14528 5633
rect 14462 5558 14528 5599
rect 14558 6517 14624 6558
rect 14558 6483 14574 6517
rect 14608 6483 14624 6517
rect 14558 6449 14624 6483
rect 14558 6415 14574 6449
rect 14608 6415 14624 6449
rect 14558 6381 14624 6415
rect 14558 6347 14574 6381
rect 14608 6347 14624 6381
rect 14558 6313 14624 6347
rect 14558 6279 14574 6313
rect 14608 6279 14624 6313
rect 14558 6245 14624 6279
rect 14558 6211 14574 6245
rect 14608 6211 14624 6245
rect 14558 6177 14624 6211
rect 14558 6143 14574 6177
rect 14608 6143 14624 6177
rect 14558 6109 14624 6143
rect 14558 6075 14574 6109
rect 14608 6075 14624 6109
rect 14558 6041 14624 6075
rect 14558 6007 14574 6041
rect 14608 6007 14624 6041
rect 14558 5973 14624 6007
rect 14558 5939 14574 5973
rect 14608 5939 14624 5973
rect 14558 5905 14624 5939
rect 14558 5871 14574 5905
rect 14608 5871 14624 5905
rect 14558 5837 14624 5871
rect 14558 5803 14574 5837
rect 14608 5803 14624 5837
rect 14558 5769 14624 5803
rect 14558 5735 14574 5769
rect 14608 5735 14624 5769
rect 14558 5701 14624 5735
rect 14558 5667 14574 5701
rect 14608 5667 14624 5701
rect 14558 5633 14624 5667
rect 14558 5599 14574 5633
rect 14608 5599 14624 5633
rect 14558 5558 14624 5599
rect 14654 6517 14720 6558
rect 14654 6483 14670 6517
rect 14704 6483 14720 6517
rect 14654 6449 14720 6483
rect 14654 6415 14670 6449
rect 14704 6415 14720 6449
rect 14654 6381 14720 6415
rect 14654 6347 14670 6381
rect 14704 6347 14720 6381
rect 14654 6313 14720 6347
rect 14654 6279 14670 6313
rect 14704 6279 14720 6313
rect 14654 6245 14720 6279
rect 14654 6211 14670 6245
rect 14704 6211 14720 6245
rect 14654 6177 14720 6211
rect 14654 6143 14670 6177
rect 14704 6143 14720 6177
rect 14654 6109 14720 6143
rect 14654 6075 14670 6109
rect 14704 6075 14720 6109
rect 14654 6041 14720 6075
rect 14654 6007 14670 6041
rect 14704 6007 14720 6041
rect 14654 5973 14720 6007
rect 14654 5939 14670 5973
rect 14704 5939 14720 5973
rect 14654 5905 14720 5939
rect 14654 5871 14670 5905
rect 14704 5871 14720 5905
rect 14654 5837 14720 5871
rect 14654 5803 14670 5837
rect 14704 5803 14720 5837
rect 14654 5769 14720 5803
rect 14654 5735 14670 5769
rect 14704 5735 14720 5769
rect 14654 5701 14720 5735
rect 14654 5667 14670 5701
rect 14704 5667 14720 5701
rect 14654 5633 14720 5667
rect 14654 5599 14670 5633
rect 14704 5599 14720 5633
rect 14654 5558 14720 5599
rect 14750 6517 14816 6558
rect 14750 6483 14766 6517
rect 14800 6483 14816 6517
rect 14750 6449 14816 6483
rect 14750 6415 14766 6449
rect 14800 6415 14816 6449
rect 14750 6381 14816 6415
rect 14750 6347 14766 6381
rect 14800 6347 14816 6381
rect 14750 6313 14816 6347
rect 14750 6279 14766 6313
rect 14800 6279 14816 6313
rect 14750 6245 14816 6279
rect 14750 6211 14766 6245
rect 14800 6211 14816 6245
rect 14750 6177 14816 6211
rect 14750 6143 14766 6177
rect 14800 6143 14816 6177
rect 14750 6109 14816 6143
rect 14750 6075 14766 6109
rect 14800 6075 14816 6109
rect 14750 6041 14816 6075
rect 14750 6007 14766 6041
rect 14800 6007 14816 6041
rect 14750 5973 14816 6007
rect 14750 5939 14766 5973
rect 14800 5939 14816 5973
rect 14750 5905 14816 5939
rect 14750 5871 14766 5905
rect 14800 5871 14816 5905
rect 14750 5837 14816 5871
rect 14750 5803 14766 5837
rect 14800 5803 14816 5837
rect 14750 5769 14816 5803
rect 14750 5735 14766 5769
rect 14800 5735 14816 5769
rect 14750 5701 14816 5735
rect 14750 5667 14766 5701
rect 14800 5667 14816 5701
rect 14750 5633 14816 5667
rect 14750 5599 14766 5633
rect 14800 5599 14816 5633
rect 14750 5558 14816 5599
rect 14846 6517 14912 6558
rect 14846 6483 14862 6517
rect 14896 6483 14912 6517
rect 14846 6449 14912 6483
rect 14846 6415 14862 6449
rect 14896 6415 14912 6449
rect 14846 6381 14912 6415
rect 14846 6347 14862 6381
rect 14896 6347 14912 6381
rect 14846 6313 14912 6347
rect 14846 6279 14862 6313
rect 14896 6279 14912 6313
rect 14846 6245 14912 6279
rect 14846 6211 14862 6245
rect 14896 6211 14912 6245
rect 14846 6177 14912 6211
rect 14846 6143 14862 6177
rect 14896 6143 14912 6177
rect 14846 6109 14912 6143
rect 14846 6075 14862 6109
rect 14896 6075 14912 6109
rect 14846 6041 14912 6075
rect 14846 6007 14862 6041
rect 14896 6007 14912 6041
rect 14846 5973 14912 6007
rect 14846 5939 14862 5973
rect 14896 5939 14912 5973
rect 14846 5905 14912 5939
rect 14846 5871 14862 5905
rect 14896 5871 14912 5905
rect 14846 5837 14912 5871
rect 14846 5803 14862 5837
rect 14896 5803 14912 5837
rect 14846 5769 14912 5803
rect 14846 5735 14862 5769
rect 14896 5735 14912 5769
rect 14846 5701 14912 5735
rect 14846 5667 14862 5701
rect 14896 5667 14912 5701
rect 14846 5633 14912 5667
rect 14846 5599 14862 5633
rect 14896 5599 14912 5633
rect 14846 5558 14912 5599
rect 14942 6517 15004 6558
rect 14942 6483 14958 6517
rect 14992 6483 15004 6517
rect 14942 6449 15004 6483
rect 14942 6415 14958 6449
rect 14992 6415 15004 6449
rect 14942 6381 15004 6415
rect 14942 6347 14958 6381
rect 14992 6347 15004 6381
rect 14942 6313 15004 6347
rect 14942 6279 14958 6313
rect 14992 6279 15004 6313
rect 14942 6245 15004 6279
rect 14942 6211 14958 6245
rect 14992 6211 15004 6245
rect 14942 6177 15004 6211
rect 14942 6143 14958 6177
rect 14992 6143 15004 6177
rect 14942 6109 15004 6143
rect 14942 6075 14958 6109
rect 14992 6075 15004 6109
rect 14942 6041 15004 6075
rect 14942 6007 14958 6041
rect 14992 6007 15004 6041
rect 14942 5973 15004 6007
rect 14942 5939 14958 5973
rect 14992 5939 15004 5973
rect 14942 5905 15004 5939
rect 14942 5871 14958 5905
rect 14992 5871 15004 5905
rect 14942 5837 15004 5871
rect 14942 5803 14958 5837
rect 14992 5803 15004 5837
rect 14942 5769 15004 5803
rect 14942 5735 14958 5769
rect 14992 5735 15004 5769
rect 14942 5701 15004 5735
rect 14942 5667 14958 5701
rect 14992 5667 15004 5701
rect 14942 5633 15004 5667
rect 14942 5599 14958 5633
rect 14992 5599 15004 5633
rect 14942 5558 15004 5599
rect 15506 5895 15568 5926
rect 15506 5861 15518 5895
rect 15552 5861 15568 5895
rect 15506 5827 15568 5861
rect 15506 5793 15518 5827
rect 15552 5793 15568 5827
rect 15506 5759 15568 5793
rect 15506 5725 15518 5759
rect 15552 5725 15568 5759
rect 15506 5691 15568 5725
rect 15506 5657 15518 5691
rect 15552 5657 15568 5691
rect 15506 5623 15568 5657
rect 15506 5589 15518 5623
rect 15552 5589 15568 5623
rect 15506 5555 15568 5589
rect -880 5487 -822 5521
rect -880 5453 -868 5487
rect -834 5453 -822 5487
rect -880 5419 -822 5453
rect -880 5385 -868 5419
rect -834 5385 -822 5419
rect -880 5351 -822 5385
rect -880 5317 -868 5351
rect -834 5317 -822 5351
rect -880 5283 -822 5317
rect -880 5249 -868 5283
rect -834 5249 -822 5283
rect -880 5215 -822 5249
rect -880 5181 -868 5215
rect -834 5181 -822 5215
rect -880 5147 -822 5181
rect -880 5113 -868 5147
rect -834 5113 -822 5147
rect -880 5079 -822 5113
rect -880 5045 -868 5079
rect -834 5045 -822 5079
rect -880 5011 -822 5045
rect 15506 5521 15518 5555
rect 15552 5521 15568 5555
rect 15506 5487 15568 5521
rect 15506 5453 15518 5487
rect 15552 5453 15568 5487
rect 15506 5419 15568 5453
rect 15506 5385 15518 5419
rect 15552 5385 15568 5419
rect 15506 5351 15568 5385
rect 15506 5317 15518 5351
rect 15552 5317 15568 5351
rect 15506 5283 15568 5317
rect 15506 5249 15518 5283
rect 15552 5249 15568 5283
rect 15506 5215 15568 5249
rect 15506 5181 15518 5215
rect 15552 5181 15568 5215
rect 15506 5147 15568 5181
rect 15506 5113 15518 5147
rect 15552 5113 15568 5147
rect 15506 5079 15568 5113
rect 15506 5045 15518 5079
rect 15552 5045 15568 5079
rect -880 4977 -868 5011
rect -834 4977 -822 5011
rect -880 4936 -822 4977
rect 15506 5011 15568 5045
rect 1472 4903 1534 4944
rect 1472 4869 1484 4903
rect 1518 4869 1534 4903
rect 1472 4835 1534 4869
rect 1472 4801 1484 4835
rect 1518 4801 1534 4835
rect 1472 4767 1534 4801
rect 1472 4733 1484 4767
rect 1518 4733 1534 4767
rect 1472 4699 1534 4733
rect 1472 4665 1484 4699
rect 1518 4665 1534 4699
rect 1472 4631 1534 4665
rect 1472 4597 1484 4631
rect 1518 4597 1534 4631
rect 1472 4563 1534 4597
rect 1472 4529 1484 4563
rect 1518 4529 1534 4563
rect 1472 4495 1534 4529
rect 1472 4461 1484 4495
rect 1518 4461 1534 4495
rect 1472 4427 1534 4461
rect 1472 4393 1484 4427
rect 1518 4393 1534 4427
rect 1472 4359 1534 4393
rect 1472 4325 1484 4359
rect 1518 4325 1534 4359
rect 1472 4291 1534 4325
rect 1472 4257 1484 4291
rect 1518 4257 1534 4291
rect 1472 4223 1534 4257
rect 1472 4189 1484 4223
rect 1518 4189 1534 4223
rect 1472 4155 1534 4189
rect 1472 4121 1484 4155
rect 1518 4121 1534 4155
rect 1472 4087 1534 4121
rect 1472 4053 1484 4087
rect 1518 4053 1534 4087
rect 1472 4019 1534 4053
rect 1472 3985 1484 4019
rect 1518 3985 1534 4019
rect 1472 3944 1534 3985
rect 1564 4903 1630 4944
rect 1564 4869 1580 4903
rect 1614 4869 1630 4903
rect 1564 4835 1630 4869
rect 1564 4801 1580 4835
rect 1614 4801 1630 4835
rect 1564 4767 1630 4801
rect 1564 4733 1580 4767
rect 1614 4733 1630 4767
rect 1564 4699 1630 4733
rect 1564 4665 1580 4699
rect 1614 4665 1630 4699
rect 1564 4631 1630 4665
rect 1564 4597 1580 4631
rect 1614 4597 1630 4631
rect 1564 4563 1630 4597
rect 1564 4529 1580 4563
rect 1614 4529 1630 4563
rect 1564 4495 1630 4529
rect 1564 4461 1580 4495
rect 1614 4461 1630 4495
rect 1564 4427 1630 4461
rect 1564 4393 1580 4427
rect 1614 4393 1630 4427
rect 1564 4359 1630 4393
rect 1564 4325 1580 4359
rect 1614 4325 1630 4359
rect 1564 4291 1630 4325
rect 1564 4257 1580 4291
rect 1614 4257 1630 4291
rect 1564 4223 1630 4257
rect 1564 4189 1580 4223
rect 1614 4189 1630 4223
rect 1564 4155 1630 4189
rect 1564 4121 1580 4155
rect 1614 4121 1630 4155
rect 1564 4087 1630 4121
rect 1564 4053 1580 4087
rect 1614 4053 1630 4087
rect 1564 4019 1630 4053
rect 1564 3985 1580 4019
rect 1614 3985 1630 4019
rect 1564 3944 1630 3985
rect 1660 4903 1726 4944
rect 1660 4869 1676 4903
rect 1710 4869 1726 4903
rect 1660 4835 1726 4869
rect 1660 4801 1676 4835
rect 1710 4801 1726 4835
rect 1660 4767 1726 4801
rect 1660 4733 1676 4767
rect 1710 4733 1726 4767
rect 1660 4699 1726 4733
rect 1660 4665 1676 4699
rect 1710 4665 1726 4699
rect 1660 4631 1726 4665
rect 1660 4597 1676 4631
rect 1710 4597 1726 4631
rect 1660 4563 1726 4597
rect 1660 4529 1676 4563
rect 1710 4529 1726 4563
rect 1660 4495 1726 4529
rect 1660 4461 1676 4495
rect 1710 4461 1726 4495
rect 1660 4427 1726 4461
rect 1660 4393 1676 4427
rect 1710 4393 1726 4427
rect 1660 4359 1726 4393
rect 1660 4325 1676 4359
rect 1710 4325 1726 4359
rect 1660 4291 1726 4325
rect 1660 4257 1676 4291
rect 1710 4257 1726 4291
rect 1660 4223 1726 4257
rect 1660 4189 1676 4223
rect 1710 4189 1726 4223
rect 1660 4155 1726 4189
rect 1660 4121 1676 4155
rect 1710 4121 1726 4155
rect 1660 4087 1726 4121
rect 1660 4053 1676 4087
rect 1710 4053 1726 4087
rect 1660 4019 1726 4053
rect 1660 3985 1676 4019
rect 1710 3985 1726 4019
rect 1660 3944 1726 3985
rect 1756 4903 1822 4944
rect 1756 4869 1772 4903
rect 1806 4869 1822 4903
rect 1756 4835 1822 4869
rect 1756 4801 1772 4835
rect 1806 4801 1822 4835
rect 1756 4767 1822 4801
rect 1756 4733 1772 4767
rect 1806 4733 1822 4767
rect 1756 4699 1822 4733
rect 1756 4665 1772 4699
rect 1806 4665 1822 4699
rect 1756 4631 1822 4665
rect 1756 4597 1772 4631
rect 1806 4597 1822 4631
rect 1756 4563 1822 4597
rect 1756 4529 1772 4563
rect 1806 4529 1822 4563
rect 1756 4495 1822 4529
rect 1756 4461 1772 4495
rect 1806 4461 1822 4495
rect 1756 4427 1822 4461
rect 1756 4393 1772 4427
rect 1806 4393 1822 4427
rect 1756 4359 1822 4393
rect 1756 4325 1772 4359
rect 1806 4325 1822 4359
rect 1756 4291 1822 4325
rect 1756 4257 1772 4291
rect 1806 4257 1822 4291
rect 1756 4223 1822 4257
rect 1756 4189 1772 4223
rect 1806 4189 1822 4223
rect 1756 4155 1822 4189
rect 1756 4121 1772 4155
rect 1806 4121 1822 4155
rect 1756 4087 1822 4121
rect 1756 4053 1772 4087
rect 1806 4053 1822 4087
rect 1756 4019 1822 4053
rect 1756 3985 1772 4019
rect 1806 3985 1822 4019
rect 1756 3944 1822 3985
rect 1852 4903 1914 4944
rect 15506 4977 15518 5011
rect 15552 4977 15568 5011
rect 1852 4869 1868 4903
rect 1902 4869 1914 4903
rect 1852 4835 1914 4869
rect 1852 4801 1868 4835
rect 1902 4801 1914 4835
rect 1852 4767 1914 4801
rect 1852 4733 1868 4767
rect 1902 4733 1914 4767
rect 1852 4699 1914 4733
rect 1852 4665 1868 4699
rect 1902 4665 1914 4699
rect 1852 4631 1914 4665
rect 1852 4597 1868 4631
rect 1902 4597 1914 4631
rect 1852 4563 1914 4597
rect 1852 4529 1868 4563
rect 1902 4529 1914 4563
rect 1852 4495 1914 4529
rect 1852 4461 1868 4495
rect 1902 4461 1914 4495
rect 1852 4427 1914 4461
rect 1852 4393 1868 4427
rect 1902 4393 1914 4427
rect 1852 4359 1914 4393
rect 1852 4325 1868 4359
rect 1902 4325 1914 4359
rect 1852 4291 1914 4325
rect 1852 4257 1868 4291
rect 1902 4257 1914 4291
rect 1852 4223 1914 4257
rect 1852 4189 1868 4223
rect 1902 4189 1914 4223
rect 1852 4155 1914 4189
rect 1852 4121 1868 4155
rect 1902 4121 1914 4155
rect 1852 4087 1914 4121
rect 1852 4053 1868 4087
rect 1902 4053 1914 4087
rect 1852 4019 1914 4053
rect 1852 3985 1868 4019
rect 1902 3985 1914 4019
rect 1852 3944 1914 3985
rect 4428 4887 4490 4928
rect 4428 4853 4440 4887
rect 4474 4853 4490 4887
rect 4428 4819 4490 4853
rect 4428 4785 4440 4819
rect 4474 4785 4490 4819
rect 4428 4751 4490 4785
rect 4428 4717 4440 4751
rect 4474 4717 4490 4751
rect 4428 4683 4490 4717
rect 4428 4649 4440 4683
rect 4474 4649 4490 4683
rect 4428 4615 4490 4649
rect 4428 4581 4440 4615
rect 4474 4581 4490 4615
rect 4428 4547 4490 4581
rect 4428 4513 4440 4547
rect 4474 4513 4490 4547
rect 4428 4479 4490 4513
rect 4428 4445 4440 4479
rect 4474 4445 4490 4479
rect 4428 4411 4490 4445
rect 4428 4377 4440 4411
rect 4474 4377 4490 4411
rect 4428 4343 4490 4377
rect 4428 4309 4440 4343
rect 4474 4309 4490 4343
rect 4428 4275 4490 4309
rect 4428 4241 4440 4275
rect 4474 4241 4490 4275
rect 4428 4207 4490 4241
rect 4428 4173 4440 4207
rect 4474 4173 4490 4207
rect 4428 4139 4490 4173
rect 4428 4105 4440 4139
rect 4474 4105 4490 4139
rect 4428 4071 4490 4105
rect 4428 4037 4440 4071
rect 4474 4037 4490 4071
rect 4428 4003 4490 4037
rect 4428 3969 4440 4003
rect 4474 3969 4490 4003
rect 4428 3928 4490 3969
rect 4520 4887 4586 4928
rect 4520 4853 4536 4887
rect 4570 4853 4586 4887
rect 4520 4819 4586 4853
rect 4520 4785 4536 4819
rect 4570 4785 4586 4819
rect 4520 4751 4586 4785
rect 4520 4717 4536 4751
rect 4570 4717 4586 4751
rect 4520 4683 4586 4717
rect 4520 4649 4536 4683
rect 4570 4649 4586 4683
rect 4520 4615 4586 4649
rect 4520 4581 4536 4615
rect 4570 4581 4586 4615
rect 4520 4547 4586 4581
rect 4520 4513 4536 4547
rect 4570 4513 4586 4547
rect 4520 4479 4586 4513
rect 4520 4445 4536 4479
rect 4570 4445 4586 4479
rect 4520 4411 4586 4445
rect 4520 4377 4536 4411
rect 4570 4377 4586 4411
rect 4520 4343 4586 4377
rect 4520 4309 4536 4343
rect 4570 4309 4586 4343
rect 4520 4275 4586 4309
rect 4520 4241 4536 4275
rect 4570 4241 4586 4275
rect 4520 4207 4586 4241
rect 4520 4173 4536 4207
rect 4570 4173 4586 4207
rect 4520 4139 4586 4173
rect 4520 4105 4536 4139
rect 4570 4105 4586 4139
rect 4520 4071 4586 4105
rect 4520 4037 4536 4071
rect 4570 4037 4586 4071
rect 4520 4003 4586 4037
rect 4520 3969 4536 4003
rect 4570 3969 4586 4003
rect 4520 3928 4586 3969
rect 4616 4887 4682 4928
rect 4616 4853 4632 4887
rect 4666 4853 4682 4887
rect 4616 4819 4682 4853
rect 4616 4785 4632 4819
rect 4666 4785 4682 4819
rect 4616 4751 4682 4785
rect 4616 4717 4632 4751
rect 4666 4717 4682 4751
rect 4616 4683 4682 4717
rect 4616 4649 4632 4683
rect 4666 4649 4682 4683
rect 4616 4615 4682 4649
rect 4616 4581 4632 4615
rect 4666 4581 4682 4615
rect 4616 4547 4682 4581
rect 4616 4513 4632 4547
rect 4666 4513 4682 4547
rect 4616 4479 4682 4513
rect 4616 4445 4632 4479
rect 4666 4445 4682 4479
rect 4616 4411 4682 4445
rect 4616 4377 4632 4411
rect 4666 4377 4682 4411
rect 4616 4343 4682 4377
rect 4616 4309 4632 4343
rect 4666 4309 4682 4343
rect 4616 4275 4682 4309
rect 4616 4241 4632 4275
rect 4666 4241 4682 4275
rect 4616 4207 4682 4241
rect 4616 4173 4632 4207
rect 4666 4173 4682 4207
rect 4616 4139 4682 4173
rect 4616 4105 4632 4139
rect 4666 4105 4682 4139
rect 4616 4071 4682 4105
rect 4616 4037 4632 4071
rect 4666 4037 4682 4071
rect 4616 4003 4682 4037
rect 4616 3969 4632 4003
rect 4666 3969 4682 4003
rect 4616 3928 4682 3969
rect 4712 4887 4778 4928
rect 4712 4853 4728 4887
rect 4762 4853 4778 4887
rect 4712 4819 4778 4853
rect 4712 4785 4728 4819
rect 4762 4785 4778 4819
rect 4712 4751 4778 4785
rect 4712 4717 4728 4751
rect 4762 4717 4778 4751
rect 4712 4683 4778 4717
rect 4712 4649 4728 4683
rect 4762 4649 4778 4683
rect 4712 4615 4778 4649
rect 4712 4581 4728 4615
rect 4762 4581 4778 4615
rect 4712 4547 4778 4581
rect 4712 4513 4728 4547
rect 4762 4513 4778 4547
rect 4712 4479 4778 4513
rect 4712 4445 4728 4479
rect 4762 4445 4778 4479
rect 4712 4411 4778 4445
rect 4712 4377 4728 4411
rect 4762 4377 4778 4411
rect 4712 4343 4778 4377
rect 4712 4309 4728 4343
rect 4762 4309 4778 4343
rect 4712 4275 4778 4309
rect 4712 4241 4728 4275
rect 4762 4241 4778 4275
rect 4712 4207 4778 4241
rect 4712 4173 4728 4207
rect 4762 4173 4778 4207
rect 4712 4139 4778 4173
rect 4712 4105 4728 4139
rect 4762 4105 4778 4139
rect 4712 4071 4778 4105
rect 4712 4037 4728 4071
rect 4762 4037 4778 4071
rect 4712 4003 4778 4037
rect 4712 3969 4728 4003
rect 4762 3969 4778 4003
rect 4712 3928 4778 3969
rect 4808 4887 4870 4928
rect 4808 4853 4824 4887
rect 4858 4853 4870 4887
rect 4808 4819 4870 4853
rect 4808 4785 4824 4819
rect 4858 4785 4870 4819
rect 4808 4751 4870 4785
rect 4808 4717 4824 4751
rect 4858 4717 4870 4751
rect 4808 4683 4870 4717
rect 4808 4649 4824 4683
rect 4858 4649 4870 4683
rect 4808 4615 4870 4649
rect 4808 4581 4824 4615
rect 4858 4581 4870 4615
rect 4808 4547 4870 4581
rect 4808 4513 4824 4547
rect 4858 4513 4870 4547
rect 4808 4479 4870 4513
rect 4808 4445 4824 4479
rect 4858 4445 4870 4479
rect 4808 4411 4870 4445
rect 4808 4377 4824 4411
rect 4858 4377 4870 4411
rect 4808 4343 4870 4377
rect 4808 4309 4824 4343
rect 4858 4309 4870 4343
rect 4808 4275 4870 4309
rect 4808 4241 4824 4275
rect 4858 4241 4870 4275
rect 4808 4207 4870 4241
rect 4808 4173 4824 4207
rect 4858 4173 4870 4207
rect 4808 4139 4870 4173
rect 4808 4105 4824 4139
rect 4858 4105 4870 4139
rect 4808 4071 4870 4105
rect 4808 4037 4824 4071
rect 4858 4037 4870 4071
rect 4808 4003 4870 4037
rect 4808 3969 4824 4003
rect 4858 3969 4870 4003
rect 4808 3928 4870 3969
rect 7458 4887 7520 4928
rect 7458 4853 7470 4887
rect 7504 4853 7520 4887
rect 7458 4819 7520 4853
rect 7458 4785 7470 4819
rect 7504 4785 7520 4819
rect 7458 4751 7520 4785
rect 7458 4717 7470 4751
rect 7504 4717 7520 4751
rect 7458 4683 7520 4717
rect 7458 4649 7470 4683
rect 7504 4649 7520 4683
rect 7458 4615 7520 4649
rect 7458 4581 7470 4615
rect 7504 4581 7520 4615
rect 7458 4547 7520 4581
rect 7458 4513 7470 4547
rect 7504 4513 7520 4547
rect 7458 4479 7520 4513
rect 7458 4445 7470 4479
rect 7504 4445 7520 4479
rect 7458 4411 7520 4445
rect 7458 4377 7470 4411
rect 7504 4377 7520 4411
rect 7458 4343 7520 4377
rect 7458 4309 7470 4343
rect 7504 4309 7520 4343
rect 7458 4275 7520 4309
rect 7458 4241 7470 4275
rect 7504 4241 7520 4275
rect 7458 4207 7520 4241
rect 7458 4173 7470 4207
rect 7504 4173 7520 4207
rect 7458 4139 7520 4173
rect 7458 4105 7470 4139
rect 7504 4105 7520 4139
rect 7458 4071 7520 4105
rect 7458 4037 7470 4071
rect 7504 4037 7520 4071
rect 7458 4003 7520 4037
rect 7458 3969 7470 4003
rect 7504 3969 7520 4003
rect 7458 3928 7520 3969
rect 7550 4887 7616 4928
rect 7550 4853 7566 4887
rect 7600 4853 7616 4887
rect 7550 4819 7616 4853
rect 7550 4785 7566 4819
rect 7600 4785 7616 4819
rect 7550 4751 7616 4785
rect 7550 4717 7566 4751
rect 7600 4717 7616 4751
rect 7550 4683 7616 4717
rect 7550 4649 7566 4683
rect 7600 4649 7616 4683
rect 7550 4615 7616 4649
rect 7550 4581 7566 4615
rect 7600 4581 7616 4615
rect 7550 4547 7616 4581
rect 7550 4513 7566 4547
rect 7600 4513 7616 4547
rect 7550 4479 7616 4513
rect 7550 4445 7566 4479
rect 7600 4445 7616 4479
rect 7550 4411 7616 4445
rect 7550 4377 7566 4411
rect 7600 4377 7616 4411
rect 7550 4343 7616 4377
rect 7550 4309 7566 4343
rect 7600 4309 7616 4343
rect 7550 4275 7616 4309
rect 7550 4241 7566 4275
rect 7600 4241 7616 4275
rect 7550 4207 7616 4241
rect 7550 4173 7566 4207
rect 7600 4173 7616 4207
rect 7550 4139 7616 4173
rect 7550 4105 7566 4139
rect 7600 4105 7616 4139
rect 7550 4071 7616 4105
rect 7550 4037 7566 4071
rect 7600 4037 7616 4071
rect 7550 4003 7616 4037
rect 7550 3969 7566 4003
rect 7600 3969 7616 4003
rect 7550 3928 7616 3969
rect 7646 4887 7712 4928
rect 7646 4853 7662 4887
rect 7696 4853 7712 4887
rect 7646 4819 7712 4853
rect 7646 4785 7662 4819
rect 7696 4785 7712 4819
rect 7646 4751 7712 4785
rect 7646 4717 7662 4751
rect 7696 4717 7712 4751
rect 7646 4683 7712 4717
rect 7646 4649 7662 4683
rect 7696 4649 7712 4683
rect 7646 4615 7712 4649
rect 7646 4581 7662 4615
rect 7696 4581 7712 4615
rect 7646 4547 7712 4581
rect 7646 4513 7662 4547
rect 7696 4513 7712 4547
rect 7646 4479 7712 4513
rect 7646 4445 7662 4479
rect 7696 4445 7712 4479
rect 7646 4411 7712 4445
rect 7646 4377 7662 4411
rect 7696 4377 7712 4411
rect 7646 4343 7712 4377
rect 7646 4309 7662 4343
rect 7696 4309 7712 4343
rect 7646 4275 7712 4309
rect 7646 4241 7662 4275
rect 7696 4241 7712 4275
rect 7646 4207 7712 4241
rect 7646 4173 7662 4207
rect 7696 4173 7712 4207
rect 7646 4139 7712 4173
rect 7646 4105 7662 4139
rect 7696 4105 7712 4139
rect 7646 4071 7712 4105
rect 7646 4037 7662 4071
rect 7696 4037 7712 4071
rect 7646 4003 7712 4037
rect 7646 3969 7662 4003
rect 7696 3969 7712 4003
rect 7646 3928 7712 3969
rect 7742 4887 7808 4928
rect 7742 4853 7758 4887
rect 7792 4853 7808 4887
rect 7742 4819 7808 4853
rect 7742 4785 7758 4819
rect 7792 4785 7808 4819
rect 7742 4751 7808 4785
rect 7742 4717 7758 4751
rect 7792 4717 7808 4751
rect 7742 4683 7808 4717
rect 7742 4649 7758 4683
rect 7792 4649 7808 4683
rect 7742 4615 7808 4649
rect 7742 4581 7758 4615
rect 7792 4581 7808 4615
rect 7742 4547 7808 4581
rect 7742 4513 7758 4547
rect 7792 4513 7808 4547
rect 7742 4479 7808 4513
rect 7742 4445 7758 4479
rect 7792 4445 7808 4479
rect 7742 4411 7808 4445
rect 7742 4377 7758 4411
rect 7792 4377 7808 4411
rect 7742 4343 7808 4377
rect 7742 4309 7758 4343
rect 7792 4309 7808 4343
rect 7742 4275 7808 4309
rect 7742 4241 7758 4275
rect 7792 4241 7808 4275
rect 7742 4207 7808 4241
rect 7742 4173 7758 4207
rect 7792 4173 7808 4207
rect 7742 4139 7808 4173
rect 7742 4105 7758 4139
rect 7792 4105 7808 4139
rect 7742 4071 7808 4105
rect 7742 4037 7758 4071
rect 7792 4037 7808 4071
rect 7742 4003 7808 4037
rect 7742 3969 7758 4003
rect 7792 3969 7808 4003
rect 7742 3928 7808 3969
rect 7838 4887 7900 4928
rect 7838 4853 7854 4887
rect 7888 4853 7900 4887
rect 7838 4819 7900 4853
rect 7838 4785 7854 4819
rect 7888 4785 7900 4819
rect 7838 4751 7900 4785
rect 7838 4717 7854 4751
rect 7888 4717 7900 4751
rect 7838 4683 7900 4717
rect 7838 4649 7854 4683
rect 7888 4649 7900 4683
rect 7838 4615 7900 4649
rect 7838 4581 7854 4615
rect 7888 4581 7900 4615
rect 7838 4547 7900 4581
rect 7838 4513 7854 4547
rect 7888 4513 7900 4547
rect 7838 4479 7900 4513
rect 7838 4445 7854 4479
rect 7888 4445 7900 4479
rect 7838 4411 7900 4445
rect 7838 4377 7854 4411
rect 7888 4377 7900 4411
rect 7838 4343 7900 4377
rect 7838 4309 7854 4343
rect 7888 4309 7900 4343
rect 7838 4275 7900 4309
rect 7838 4241 7854 4275
rect 7888 4241 7900 4275
rect 7838 4207 7900 4241
rect 7838 4173 7854 4207
rect 7888 4173 7900 4207
rect 7838 4139 7900 4173
rect 7838 4105 7854 4139
rect 7888 4105 7900 4139
rect 7838 4071 7900 4105
rect 7838 4037 7854 4071
rect 7888 4037 7900 4071
rect 7838 4003 7900 4037
rect 7838 3969 7854 4003
rect 7888 3969 7900 4003
rect 7838 3928 7900 3969
rect 10546 4885 10608 4926
rect 10546 4851 10558 4885
rect 10592 4851 10608 4885
rect 10546 4817 10608 4851
rect 10546 4783 10558 4817
rect 10592 4783 10608 4817
rect 10546 4749 10608 4783
rect 10546 4715 10558 4749
rect 10592 4715 10608 4749
rect 10546 4681 10608 4715
rect 10546 4647 10558 4681
rect 10592 4647 10608 4681
rect 10546 4613 10608 4647
rect 10546 4579 10558 4613
rect 10592 4579 10608 4613
rect 10546 4545 10608 4579
rect 10546 4511 10558 4545
rect 10592 4511 10608 4545
rect 10546 4477 10608 4511
rect 10546 4443 10558 4477
rect 10592 4443 10608 4477
rect 10546 4409 10608 4443
rect 10546 4375 10558 4409
rect 10592 4375 10608 4409
rect 10546 4341 10608 4375
rect 10546 4307 10558 4341
rect 10592 4307 10608 4341
rect 10546 4273 10608 4307
rect 10546 4239 10558 4273
rect 10592 4239 10608 4273
rect 10546 4205 10608 4239
rect 10546 4171 10558 4205
rect 10592 4171 10608 4205
rect 10546 4137 10608 4171
rect 10546 4103 10558 4137
rect 10592 4103 10608 4137
rect 10546 4069 10608 4103
rect 10546 4035 10558 4069
rect 10592 4035 10608 4069
rect 10546 4001 10608 4035
rect 10546 3967 10558 4001
rect 10592 3967 10608 4001
rect 10546 3926 10608 3967
rect 10638 4885 10704 4926
rect 10638 4851 10654 4885
rect 10688 4851 10704 4885
rect 10638 4817 10704 4851
rect 10638 4783 10654 4817
rect 10688 4783 10704 4817
rect 10638 4749 10704 4783
rect 10638 4715 10654 4749
rect 10688 4715 10704 4749
rect 10638 4681 10704 4715
rect 10638 4647 10654 4681
rect 10688 4647 10704 4681
rect 10638 4613 10704 4647
rect 10638 4579 10654 4613
rect 10688 4579 10704 4613
rect 10638 4545 10704 4579
rect 10638 4511 10654 4545
rect 10688 4511 10704 4545
rect 10638 4477 10704 4511
rect 10638 4443 10654 4477
rect 10688 4443 10704 4477
rect 10638 4409 10704 4443
rect 10638 4375 10654 4409
rect 10688 4375 10704 4409
rect 10638 4341 10704 4375
rect 10638 4307 10654 4341
rect 10688 4307 10704 4341
rect 10638 4273 10704 4307
rect 10638 4239 10654 4273
rect 10688 4239 10704 4273
rect 10638 4205 10704 4239
rect 10638 4171 10654 4205
rect 10688 4171 10704 4205
rect 10638 4137 10704 4171
rect 10638 4103 10654 4137
rect 10688 4103 10704 4137
rect 10638 4069 10704 4103
rect 10638 4035 10654 4069
rect 10688 4035 10704 4069
rect 10638 4001 10704 4035
rect 10638 3967 10654 4001
rect 10688 3967 10704 4001
rect 10638 3926 10704 3967
rect 10734 4885 10800 4926
rect 10734 4851 10750 4885
rect 10784 4851 10800 4885
rect 10734 4817 10800 4851
rect 10734 4783 10750 4817
rect 10784 4783 10800 4817
rect 10734 4749 10800 4783
rect 10734 4715 10750 4749
rect 10784 4715 10800 4749
rect 10734 4681 10800 4715
rect 10734 4647 10750 4681
rect 10784 4647 10800 4681
rect 10734 4613 10800 4647
rect 10734 4579 10750 4613
rect 10784 4579 10800 4613
rect 10734 4545 10800 4579
rect 10734 4511 10750 4545
rect 10784 4511 10800 4545
rect 10734 4477 10800 4511
rect 10734 4443 10750 4477
rect 10784 4443 10800 4477
rect 10734 4409 10800 4443
rect 10734 4375 10750 4409
rect 10784 4375 10800 4409
rect 10734 4341 10800 4375
rect 10734 4307 10750 4341
rect 10784 4307 10800 4341
rect 10734 4273 10800 4307
rect 10734 4239 10750 4273
rect 10784 4239 10800 4273
rect 10734 4205 10800 4239
rect 10734 4171 10750 4205
rect 10784 4171 10800 4205
rect 10734 4137 10800 4171
rect 10734 4103 10750 4137
rect 10784 4103 10800 4137
rect 10734 4069 10800 4103
rect 10734 4035 10750 4069
rect 10784 4035 10800 4069
rect 10734 4001 10800 4035
rect 10734 3967 10750 4001
rect 10784 3967 10800 4001
rect 10734 3926 10800 3967
rect 10830 4885 10896 4926
rect 10830 4851 10846 4885
rect 10880 4851 10896 4885
rect 10830 4817 10896 4851
rect 10830 4783 10846 4817
rect 10880 4783 10896 4817
rect 10830 4749 10896 4783
rect 10830 4715 10846 4749
rect 10880 4715 10896 4749
rect 10830 4681 10896 4715
rect 10830 4647 10846 4681
rect 10880 4647 10896 4681
rect 10830 4613 10896 4647
rect 10830 4579 10846 4613
rect 10880 4579 10896 4613
rect 10830 4545 10896 4579
rect 10830 4511 10846 4545
rect 10880 4511 10896 4545
rect 10830 4477 10896 4511
rect 10830 4443 10846 4477
rect 10880 4443 10896 4477
rect 10830 4409 10896 4443
rect 10830 4375 10846 4409
rect 10880 4375 10896 4409
rect 10830 4341 10896 4375
rect 10830 4307 10846 4341
rect 10880 4307 10896 4341
rect 10830 4273 10896 4307
rect 10830 4239 10846 4273
rect 10880 4239 10896 4273
rect 10830 4205 10896 4239
rect 10830 4171 10846 4205
rect 10880 4171 10896 4205
rect 10830 4137 10896 4171
rect 10830 4103 10846 4137
rect 10880 4103 10896 4137
rect 10830 4069 10896 4103
rect 10830 4035 10846 4069
rect 10880 4035 10896 4069
rect 10830 4001 10896 4035
rect 10830 3967 10846 4001
rect 10880 3967 10896 4001
rect 10830 3926 10896 3967
rect 10926 4885 10988 4926
rect 15506 4943 15568 4977
rect 15506 4909 15518 4943
rect 15552 4909 15568 4943
rect 10926 4851 10942 4885
rect 10976 4851 10988 4885
rect 10926 4817 10988 4851
rect 10926 4783 10942 4817
rect 10976 4783 10988 4817
rect 10926 4749 10988 4783
rect 10926 4715 10942 4749
rect 10976 4715 10988 4749
rect 10926 4681 10988 4715
rect 10926 4647 10942 4681
rect 10976 4647 10988 4681
rect 10926 4613 10988 4647
rect 10926 4579 10942 4613
rect 10976 4579 10988 4613
rect 10926 4545 10988 4579
rect 10926 4511 10942 4545
rect 10976 4511 10988 4545
rect 10926 4477 10988 4511
rect 10926 4443 10942 4477
rect 10976 4443 10988 4477
rect 10926 4409 10988 4443
rect 10926 4375 10942 4409
rect 10976 4375 10988 4409
rect 10926 4341 10988 4375
rect 10926 4307 10942 4341
rect 10976 4307 10988 4341
rect 10926 4273 10988 4307
rect 10926 4239 10942 4273
rect 10976 4239 10988 4273
rect 10926 4205 10988 4239
rect 10926 4171 10942 4205
rect 10976 4171 10988 4205
rect 10926 4137 10988 4171
rect 10926 4103 10942 4137
rect 10976 4103 10988 4137
rect 10926 4069 10988 4103
rect 10926 4035 10942 4069
rect 10976 4035 10988 4069
rect 10926 4001 10988 4035
rect 10926 3967 10942 4001
rect 10976 3967 10988 4001
rect 10926 3926 10988 3967
rect 13702 4859 13764 4900
rect 13702 4825 13714 4859
rect 13748 4825 13764 4859
rect 13702 4791 13764 4825
rect 13702 4757 13714 4791
rect 13748 4757 13764 4791
rect 13702 4723 13764 4757
rect 13702 4689 13714 4723
rect 13748 4689 13764 4723
rect 13702 4655 13764 4689
rect 13702 4621 13714 4655
rect 13748 4621 13764 4655
rect 13702 4587 13764 4621
rect 13702 4553 13714 4587
rect 13748 4553 13764 4587
rect 13702 4519 13764 4553
rect 13702 4485 13714 4519
rect 13748 4485 13764 4519
rect 13702 4451 13764 4485
rect 13702 4417 13714 4451
rect 13748 4417 13764 4451
rect 13702 4383 13764 4417
rect 13702 4349 13714 4383
rect 13748 4349 13764 4383
rect 13702 4315 13764 4349
rect 13702 4281 13714 4315
rect 13748 4281 13764 4315
rect 13702 4247 13764 4281
rect 13702 4213 13714 4247
rect 13748 4213 13764 4247
rect 13702 4179 13764 4213
rect 13702 4145 13714 4179
rect 13748 4145 13764 4179
rect 13702 4111 13764 4145
rect 13702 4077 13714 4111
rect 13748 4077 13764 4111
rect 13702 4043 13764 4077
rect 13702 4009 13714 4043
rect 13748 4009 13764 4043
rect 13702 3975 13764 4009
rect 13702 3941 13714 3975
rect 13748 3941 13764 3975
rect 13702 3900 13764 3941
rect 13794 4859 13860 4900
rect 13794 4825 13810 4859
rect 13844 4825 13860 4859
rect 13794 4791 13860 4825
rect 13794 4757 13810 4791
rect 13844 4757 13860 4791
rect 13794 4723 13860 4757
rect 13794 4689 13810 4723
rect 13844 4689 13860 4723
rect 13794 4655 13860 4689
rect 13794 4621 13810 4655
rect 13844 4621 13860 4655
rect 13794 4587 13860 4621
rect 13794 4553 13810 4587
rect 13844 4553 13860 4587
rect 13794 4519 13860 4553
rect 13794 4485 13810 4519
rect 13844 4485 13860 4519
rect 13794 4451 13860 4485
rect 13794 4417 13810 4451
rect 13844 4417 13860 4451
rect 13794 4383 13860 4417
rect 13794 4349 13810 4383
rect 13844 4349 13860 4383
rect 13794 4315 13860 4349
rect 13794 4281 13810 4315
rect 13844 4281 13860 4315
rect 13794 4247 13860 4281
rect 13794 4213 13810 4247
rect 13844 4213 13860 4247
rect 13794 4179 13860 4213
rect 13794 4145 13810 4179
rect 13844 4145 13860 4179
rect 13794 4111 13860 4145
rect 13794 4077 13810 4111
rect 13844 4077 13860 4111
rect 13794 4043 13860 4077
rect 13794 4009 13810 4043
rect 13844 4009 13860 4043
rect 13794 3975 13860 4009
rect 13794 3941 13810 3975
rect 13844 3941 13860 3975
rect 13794 3900 13860 3941
rect 13890 4859 13956 4900
rect 13890 4825 13906 4859
rect 13940 4825 13956 4859
rect 13890 4791 13956 4825
rect 13890 4757 13906 4791
rect 13940 4757 13956 4791
rect 13890 4723 13956 4757
rect 13890 4689 13906 4723
rect 13940 4689 13956 4723
rect 13890 4655 13956 4689
rect 13890 4621 13906 4655
rect 13940 4621 13956 4655
rect 13890 4587 13956 4621
rect 13890 4553 13906 4587
rect 13940 4553 13956 4587
rect 13890 4519 13956 4553
rect 13890 4485 13906 4519
rect 13940 4485 13956 4519
rect 13890 4451 13956 4485
rect 13890 4417 13906 4451
rect 13940 4417 13956 4451
rect 13890 4383 13956 4417
rect 13890 4349 13906 4383
rect 13940 4349 13956 4383
rect 13890 4315 13956 4349
rect 13890 4281 13906 4315
rect 13940 4281 13956 4315
rect 13890 4247 13956 4281
rect 13890 4213 13906 4247
rect 13940 4213 13956 4247
rect 13890 4179 13956 4213
rect 13890 4145 13906 4179
rect 13940 4145 13956 4179
rect 13890 4111 13956 4145
rect 13890 4077 13906 4111
rect 13940 4077 13956 4111
rect 13890 4043 13956 4077
rect 13890 4009 13906 4043
rect 13940 4009 13956 4043
rect 13890 3975 13956 4009
rect 13890 3941 13906 3975
rect 13940 3941 13956 3975
rect 13890 3900 13956 3941
rect 13986 4859 14052 4900
rect 13986 4825 14002 4859
rect 14036 4825 14052 4859
rect 13986 4791 14052 4825
rect 13986 4757 14002 4791
rect 14036 4757 14052 4791
rect 13986 4723 14052 4757
rect 13986 4689 14002 4723
rect 14036 4689 14052 4723
rect 13986 4655 14052 4689
rect 13986 4621 14002 4655
rect 14036 4621 14052 4655
rect 13986 4587 14052 4621
rect 13986 4553 14002 4587
rect 14036 4553 14052 4587
rect 13986 4519 14052 4553
rect 13986 4485 14002 4519
rect 14036 4485 14052 4519
rect 13986 4451 14052 4485
rect 13986 4417 14002 4451
rect 14036 4417 14052 4451
rect 13986 4383 14052 4417
rect 13986 4349 14002 4383
rect 14036 4349 14052 4383
rect 13986 4315 14052 4349
rect 13986 4281 14002 4315
rect 14036 4281 14052 4315
rect 13986 4247 14052 4281
rect 13986 4213 14002 4247
rect 14036 4213 14052 4247
rect 13986 4179 14052 4213
rect 13986 4145 14002 4179
rect 14036 4145 14052 4179
rect 13986 4111 14052 4145
rect 13986 4077 14002 4111
rect 14036 4077 14052 4111
rect 13986 4043 14052 4077
rect 13986 4009 14002 4043
rect 14036 4009 14052 4043
rect 13986 3975 14052 4009
rect 13986 3941 14002 3975
rect 14036 3941 14052 3975
rect 13986 3900 14052 3941
rect 14082 4859 14144 4900
rect 14082 4825 14098 4859
rect 14132 4825 14144 4859
rect 14082 4791 14144 4825
rect 14082 4757 14098 4791
rect 14132 4757 14144 4791
rect 14082 4723 14144 4757
rect 14082 4689 14098 4723
rect 14132 4689 14144 4723
rect 14082 4655 14144 4689
rect 14082 4621 14098 4655
rect 14132 4621 14144 4655
rect 14082 4587 14144 4621
rect 14082 4553 14098 4587
rect 14132 4553 14144 4587
rect 14082 4519 14144 4553
rect 14082 4485 14098 4519
rect 14132 4485 14144 4519
rect 14082 4451 14144 4485
rect 14082 4417 14098 4451
rect 14132 4417 14144 4451
rect 14082 4383 14144 4417
rect 14082 4349 14098 4383
rect 14132 4349 14144 4383
rect 14082 4315 14144 4349
rect 14082 4281 14098 4315
rect 14132 4281 14144 4315
rect 14082 4247 14144 4281
rect 14082 4213 14098 4247
rect 14132 4213 14144 4247
rect 14082 4179 14144 4213
rect 14082 4145 14098 4179
rect 14132 4145 14144 4179
rect 14082 4111 14144 4145
rect 14082 4077 14098 4111
rect 14132 4077 14144 4111
rect 14082 4043 14144 4077
rect 14082 4009 14098 4043
rect 14132 4009 14144 4043
rect 14082 3975 14144 4009
rect 14082 3941 14098 3975
rect 14132 3941 14144 3975
rect 14082 3900 14144 3941
rect 15506 4875 15568 4909
rect 15506 4841 15518 4875
rect 15552 4841 15568 4875
rect 15506 4807 15568 4841
rect 15506 4773 15518 4807
rect 15552 4773 15568 4807
rect 15506 4739 15568 4773
rect 15506 4705 15518 4739
rect 15552 4705 15568 4739
rect 15506 4671 15568 4705
rect 15506 4637 15518 4671
rect 15552 4637 15568 4671
rect 15506 4603 15568 4637
rect 15506 4569 15518 4603
rect 15552 4569 15568 4603
rect 15506 4535 15568 4569
rect 15506 4501 15518 4535
rect 15552 4501 15568 4535
rect 15506 4467 15568 4501
rect 15506 4433 15518 4467
rect 15552 4433 15568 4467
rect 15506 4399 15568 4433
rect 15506 4365 15518 4399
rect 15552 4365 15568 4399
rect 15506 4331 15568 4365
rect 15506 4297 15518 4331
rect 15552 4297 15568 4331
rect 15506 4263 15568 4297
rect 15506 4229 15518 4263
rect 15552 4229 15568 4263
rect 15506 4195 15568 4229
rect 15506 4161 15518 4195
rect 15552 4161 15568 4195
rect 15506 4127 15568 4161
rect 15506 4093 15518 4127
rect 15552 4093 15568 4127
rect 15506 4059 15568 4093
rect 15506 4025 15518 4059
rect 15552 4025 15568 4059
rect 15506 3991 15568 4025
rect 15506 3957 15518 3991
rect 15552 3957 15568 3991
rect 15506 3926 15568 3957
rect 15598 5895 15664 5926
rect 15598 5861 15614 5895
rect 15648 5861 15664 5895
rect 15598 5827 15664 5861
rect 15598 5793 15614 5827
rect 15648 5793 15664 5827
rect 15598 5759 15664 5793
rect 15598 5725 15614 5759
rect 15648 5725 15664 5759
rect 15598 5691 15664 5725
rect 15598 5657 15614 5691
rect 15648 5657 15664 5691
rect 15598 5623 15664 5657
rect 15598 5589 15614 5623
rect 15648 5589 15664 5623
rect 15598 5555 15664 5589
rect 15598 5521 15614 5555
rect 15648 5521 15664 5555
rect 15598 5487 15664 5521
rect 15598 5453 15614 5487
rect 15648 5453 15664 5487
rect 15598 5419 15664 5453
rect 15598 5385 15614 5419
rect 15648 5385 15664 5419
rect 15598 5351 15664 5385
rect 15598 5317 15614 5351
rect 15648 5317 15664 5351
rect 15598 5283 15664 5317
rect 15598 5249 15614 5283
rect 15648 5249 15664 5283
rect 15598 5215 15664 5249
rect 15598 5181 15614 5215
rect 15648 5181 15664 5215
rect 15598 5147 15664 5181
rect 15598 5113 15614 5147
rect 15648 5113 15664 5147
rect 15598 5079 15664 5113
rect 15598 5045 15614 5079
rect 15648 5045 15664 5079
rect 15598 5011 15664 5045
rect 15598 4977 15614 5011
rect 15648 4977 15664 5011
rect 15598 4943 15664 4977
rect 15598 4909 15614 4943
rect 15648 4909 15664 4943
rect 15598 4875 15664 4909
rect 15598 4841 15614 4875
rect 15648 4841 15664 4875
rect 15598 4807 15664 4841
rect 15598 4773 15614 4807
rect 15648 4773 15664 4807
rect 15598 4739 15664 4773
rect 15598 4705 15614 4739
rect 15648 4705 15664 4739
rect 15598 4671 15664 4705
rect 15598 4637 15614 4671
rect 15648 4637 15664 4671
rect 15598 4603 15664 4637
rect 15598 4569 15614 4603
rect 15648 4569 15664 4603
rect 15598 4535 15664 4569
rect 15598 4501 15614 4535
rect 15648 4501 15664 4535
rect 15598 4467 15664 4501
rect 15598 4433 15614 4467
rect 15648 4433 15664 4467
rect 15598 4399 15664 4433
rect 15598 4365 15614 4399
rect 15648 4365 15664 4399
rect 15598 4331 15664 4365
rect 15598 4297 15614 4331
rect 15648 4297 15664 4331
rect 15598 4263 15664 4297
rect 15598 4229 15614 4263
rect 15648 4229 15664 4263
rect 15598 4195 15664 4229
rect 15598 4161 15614 4195
rect 15648 4161 15664 4195
rect 15598 4127 15664 4161
rect 15598 4093 15614 4127
rect 15648 4093 15664 4127
rect 15598 4059 15664 4093
rect 15598 4025 15614 4059
rect 15648 4025 15664 4059
rect 15598 3991 15664 4025
rect 15598 3957 15614 3991
rect 15648 3957 15664 3991
rect 15598 3926 15664 3957
rect 15694 5895 15756 5926
rect 15694 5861 15710 5895
rect 15744 5861 15756 5895
rect 15694 5827 15756 5861
rect 15694 5793 15710 5827
rect 15744 5793 15756 5827
rect 15694 5759 15756 5793
rect 15694 5725 15710 5759
rect 15744 5725 15756 5759
rect 15694 5691 15756 5725
rect 15694 5657 15710 5691
rect 15744 5657 15756 5691
rect 15694 5623 15756 5657
rect 15694 5589 15710 5623
rect 15744 5589 15756 5623
rect 15694 5555 15756 5589
rect 15694 5521 15710 5555
rect 15744 5521 15756 5555
rect 15694 5487 15756 5521
rect 15694 5453 15710 5487
rect 15744 5453 15756 5487
rect 15694 5419 15756 5453
rect 15694 5385 15710 5419
rect 15744 5385 15756 5419
rect 15694 5351 15756 5385
rect 15694 5317 15710 5351
rect 15744 5317 15756 5351
rect 15694 5283 15756 5317
rect 15694 5249 15710 5283
rect 15744 5249 15756 5283
rect 15694 5215 15756 5249
rect 15694 5181 15710 5215
rect 15744 5181 15756 5215
rect 15694 5147 15756 5181
rect 15694 5113 15710 5147
rect 15744 5113 15756 5147
rect 15694 5079 15756 5113
rect 15694 5045 15710 5079
rect 15744 5045 15756 5079
rect 15694 5011 15756 5045
rect 15694 4977 15710 5011
rect 15744 4977 15756 5011
rect 15694 4943 15756 4977
rect 15694 4909 15710 4943
rect 15744 4909 15756 4943
rect 15694 4875 15756 4909
rect 15694 4841 15710 4875
rect 15744 4841 15756 4875
rect 15694 4807 15756 4841
rect 15694 4773 15710 4807
rect 15744 4773 15756 4807
rect 15694 4739 15756 4773
rect 15694 4705 15710 4739
rect 15744 4705 15756 4739
rect 15694 4671 15756 4705
rect 15694 4637 15710 4671
rect 15744 4637 15756 4671
rect 15694 4603 15756 4637
rect 15694 4569 15710 4603
rect 15744 4569 15756 4603
rect 15694 4535 15756 4569
rect 15694 4501 15710 4535
rect 15744 4501 15756 4535
rect 15694 4467 15756 4501
rect 15694 4433 15710 4467
rect 15744 4433 15756 4467
rect 15694 4399 15756 4433
rect 15694 4365 15710 4399
rect 15744 4365 15756 4399
rect 15694 4331 15756 4365
rect 15694 4297 15710 4331
rect 15744 4297 15756 4331
rect 15694 4263 15756 4297
rect 15694 4229 15710 4263
rect 15744 4229 15756 4263
rect 15694 4195 15756 4229
rect 15694 4161 15710 4195
rect 15744 4161 15756 4195
rect 15694 4127 15756 4161
rect 15694 4093 15710 4127
rect 15744 4093 15756 4127
rect 15694 4059 15756 4093
rect 15694 4025 15710 4059
rect 15744 4025 15756 4059
rect 15694 3991 15756 4025
rect 15694 3957 15710 3991
rect 15744 3957 15756 3991
rect 15694 3926 15756 3957
<< ndiffc >>
rect -1686 3161 -1652 3195
rect -1686 3093 -1652 3127
rect -1686 3025 -1652 3059
rect -1686 2957 -1652 2991
rect -1686 2889 -1652 2923
rect -1686 2821 -1652 2855
rect -1686 2753 -1652 2787
rect -1686 2685 -1652 2719
rect -1686 2617 -1652 2651
rect -1686 2549 -1652 2583
rect -1686 2481 -1652 2515
rect -1686 2413 -1652 2447
rect -1686 2345 -1652 2379
rect -1686 2277 -1652 2311
rect -1590 3161 -1556 3195
rect -1590 3093 -1556 3127
rect -1590 3025 -1556 3059
rect -1590 2957 -1556 2991
rect -1590 2889 -1556 2923
rect -1590 2821 -1556 2855
rect -1590 2753 -1556 2787
rect -1590 2685 -1556 2719
rect -1590 2617 -1556 2651
rect -1590 2549 -1556 2583
rect -1590 2481 -1556 2515
rect -1590 2413 -1556 2447
rect -1590 2345 -1556 2379
rect -1590 2277 -1556 2311
rect -1494 3161 -1460 3195
rect -1494 3093 -1460 3127
rect -1494 3025 -1460 3059
rect -1494 2957 -1460 2991
rect -1494 2889 -1460 2923
rect -1494 2821 -1460 2855
rect -1494 2753 -1460 2787
rect -1494 2685 -1460 2719
rect -1494 2617 -1460 2651
rect -1494 2549 -1460 2583
rect -1494 2481 -1460 2515
rect -1494 2413 -1460 2447
rect -1494 2345 -1460 2379
rect -1494 2277 -1460 2311
rect -1398 3161 -1364 3195
rect -1398 3093 -1364 3127
rect -1398 3025 -1364 3059
rect -1398 2957 -1364 2991
rect -1398 2889 -1364 2923
rect -1398 2821 -1364 2855
rect -1398 2753 -1364 2787
rect -1398 2685 -1364 2719
rect -1398 2617 -1364 2651
rect -1398 2549 -1364 2583
rect -1398 2481 -1364 2515
rect -1398 2413 -1364 2447
rect -1398 2345 -1364 2379
rect -1398 2277 -1364 2311
rect -1302 3161 -1268 3195
rect -1302 3093 -1268 3127
rect -1302 3025 -1268 3059
rect -1302 2957 -1268 2991
rect -1302 2889 -1268 2923
rect -1302 2821 -1268 2855
rect -1302 2753 -1268 2787
rect -1302 2685 -1268 2719
rect -1302 2617 -1268 2651
rect -1302 2549 -1268 2583
rect -1302 2481 -1268 2515
rect -1302 2413 -1268 2447
rect -1302 2345 -1268 2379
rect -1302 2277 -1268 2311
rect -1206 3161 -1172 3195
rect -1206 3093 -1172 3127
rect -1206 3025 -1172 3059
rect -1206 2957 -1172 2991
rect -1206 2889 -1172 2923
rect -1206 2821 -1172 2855
rect -1206 2753 -1172 2787
rect -1206 2685 -1172 2719
rect -1206 2617 -1172 2651
rect -1206 2549 -1172 2583
rect -1206 2481 -1172 2515
rect -1206 2413 -1172 2447
rect -1206 2345 -1172 2379
rect -1206 2277 -1172 2311
rect -1110 3161 -1076 3195
rect -1110 3093 -1076 3127
rect -1110 3025 -1076 3059
rect -1110 2957 -1076 2991
rect -1110 2889 -1076 2923
rect -1110 2821 -1076 2855
rect -1110 2753 -1076 2787
rect -1110 2685 -1076 2719
rect -1110 2617 -1076 2651
rect -1110 2549 -1076 2583
rect -1110 2481 -1076 2515
rect -1110 2413 -1076 2447
rect -1110 2345 -1076 2379
rect -1110 2277 -1076 2311
rect -1014 3161 -980 3195
rect -1014 3093 -980 3127
rect -1014 3025 -980 3059
rect -1014 2957 -980 2991
rect -1014 2889 -980 2923
rect -1014 2821 -980 2855
rect -1014 2753 -980 2787
rect -1014 2685 -980 2719
rect -1014 2617 -980 2651
rect -1014 2549 -980 2583
rect -1014 2481 -980 2515
rect -1014 2413 -980 2447
rect -1014 2345 -980 2379
rect -1014 2277 -980 2311
rect -918 3161 -884 3195
rect -918 3093 -884 3127
rect -918 3025 -884 3059
rect -918 2957 -884 2991
rect -918 2889 -884 2923
rect -918 2821 -884 2855
rect -918 2753 -884 2787
rect -918 2685 -884 2719
rect -918 2617 -884 2651
rect -918 2549 -884 2583
rect -918 2481 -884 2515
rect -918 2413 -884 2447
rect -918 2345 -884 2379
rect -918 2277 -884 2311
rect 1482 2755 1516 2789
rect 1482 2687 1516 2721
rect 1482 2619 1516 2653
rect 1482 2551 1516 2585
rect 1482 2483 1516 2517
rect 1482 2415 1516 2449
rect 1482 2347 1516 2381
rect 1482 2279 1516 2313
rect 1482 2211 1516 2245
rect 1482 2143 1516 2177
rect 1482 2075 1516 2109
rect 1482 2007 1516 2041
rect 1482 1939 1516 1973
rect 1482 1871 1516 1905
rect 1578 2755 1612 2789
rect 1578 2687 1612 2721
rect 1578 2619 1612 2653
rect 1578 2551 1612 2585
rect 1578 2483 1612 2517
rect 1578 2415 1612 2449
rect 1578 2347 1612 2381
rect 1578 2279 1612 2313
rect 1578 2211 1612 2245
rect 1578 2143 1612 2177
rect 1578 2075 1612 2109
rect 1578 2007 1612 2041
rect 1578 1939 1612 1973
rect 1578 1871 1612 1905
rect 1674 2755 1708 2789
rect 1674 2687 1708 2721
rect 1674 2619 1708 2653
rect 1674 2551 1708 2585
rect 1674 2483 1708 2517
rect 1674 2415 1708 2449
rect 1674 2347 1708 2381
rect 1674 2279 1708 2313
rect 1674 2211 1708 2245
rect 1674 2143 1708 2177
rect 1674 2075 1708 2109
rect 1674 2007 1708 2041
rect 1674 1939 1708 1973
rect 1674 1871 1708 1905
rect 1770 2755 1804 2789
rect 1770 2687 1804 2721
rect 1770 2619 1804 2653
rect 1770 2551 1804 2585
rect 1770 2483 1804 2517
rect 1770 2415 1804 2449
rect 1770 2347 1804 2381
rect 1770 2279 1804 2313
rect 1770 2211 1804 2245
rect 1770 2143 1804 2177
rect 1770 2075 1804 2109
rect 1770 2007 1804 2041
rect 1770 1939 1804 1973
rect 1770 1871 1804 1905
rect 1866 2755 1900 2789
rect 1866 2687 1900 2721
rect 1866 2619 1900 2653
rect 1866 2551 1900 2585
rect 1866 2483 1900 2517
rect 1866 2415 1900 2449
rect 4438 2739 4472 2773
rect 4438 2671 4472 2705
rect 4438 2603 4472 2637
rect 4438 2535 4472 2569
rect 4438 2467 4472 2501
rect 1866 2347 1900 2381
rect 1866 2279 1900 2313
rect 4438 2399 4472 2433
rect 4438 2331 4472 2365
rect 1866 2211 1900 2245
rect 1866 2143 1900 2177
rect 1866 2075 1900 2109
rect 2500 2227 2534 2261
rect 2500 2159 2534 2193
rect 2500 2091 2534 2125
rect 2658 2227 2692 2261
rect 2658 2159 2692 2193
rect 2658 2091 2692 2125
rect 4438 2263 4472 2297
rect 4438 2195 4472 2229
rect 4438 2127 4472 2161
rect 4438 2059 4472 2093
rect 1866 2007 1900 2041
rect 1866 1939 1900 1973
rect 1866 1871 1900 1905
rect 4438 1991 4472 2025
rect 4438 1923 4472 1957
rect 4438 1855 4472 1889
rect 4534 2739 4568 2773
rect 4534 2671 4568 2705
rect 4534 2603 4568 2637
rect 4534 2535 4568 2569
rect 4534 2467 4568 2501
rect 4534 2399 4568 2433
rect 4534 2331 4568 2365
rect 4534 2263 4568 2297
rect 4534 2195 4568 2229
rect 4534 2127 4568 2161
rect 4534 2059 4568 2093
rect 4534 1991 4568 2025
rect 4534 1923 4568 1957
rect 4534 1855 4568 1889
rect 4630 2739 4664 2773
rect 4630 2671 4664 2705
rect 4630 2603 4664 2637
rect 4630 2535 4664 2569
rect 4630 2467 4664 2501
rect 4630 2399 4664 2433
rect 4630 2331 4664 2365
rect 4630 2263 4664 2297
rect 4630 2195 4664 2229
rect 4630 2127 4664 2161
rect 4630 2059 4664 2093
rect 4630 1991 4664 2025
rect 4630 1923 4664 1957
rect 4630 1855 4664 1889
rect 4726 2739 4760 2773
rect 4726 2671 4760 2705
rect 4726 2603 4760 2637
rect 4726 2535 4760 2569
rect 4726 2467 4760 2501
rect 4726 2399 4760 2433
rect 4726 2331 4760 2365
rect 4726 2263 4760 2297
rect 4726 2195 4760 2229
rect 4726 2127 4760 2161
rect 4726 2059 4760 2093
rect 4726 1991 4760 2025
rect 4726 1923 4760 1957
rect 4726 1855 4760 1889
rect 4822 2739 4856 2773
rect 4822 2671 4856 2705
rect 4822 2603 4856 2637
rect 4822 2535 4856 2569
rect 4822 2467 4856 2501
rect 7468 2739 7502 2773
rect 7468 2671 7502 2705
rect 7468 2603 7502 2637
rect 7468 2535 7502 2569
rect 7468 2467 7502 2501
rect 4822 2399 4856 2433
rect 4822 2331 4856 2365
rect 4822 2263 4856 2297
rect 7468 2399 7502 2433
rect 7468 2331 7502 2365
rect 4822 2195 4856 2229
rect 4822 2127 4856 2161
rect 4822 2059 4856 2093
rect 5500 2227 5534 2261
rect 5500 2159 5534 2193
rect 5500 2091 5534 2125
rect 5658 2227 5692 2261
rect 5658 2159 5692 2193
rect 5658 2091 5692 2125
rect 7468 2263 7502 2297
rect 7468 2195 7502 2229
rect 7468 2127 7502 2161
rect 7468 2059 7502 2093
rect 4822 1991 4856 2025
rect 4822 1923 4856 1957
rect 4822 1855 4856 1889
rect 7468 1991 7502 2025
rect 7468 1923 7502 1957
rect 7468 1855 7502 1889
rect 7564 2739 7598 2773
rect 7564 2671 7598 2705
rect 7564 2603 7598 2637
rect 7564 2535 7598 2569
rect 7564 2467 7598 2501
rect 7564 2399 7598 2433
rect 7564 2331 7598 2365
rect 7564 2263 7598 2297
rect 7564 2195 7598 2229
rect 7564 2127 7598 2161
rect 7564 2059 7598 2093
rect 7564 1991 7598 2025
rect 7564 1923 7598 1957
rect 7564 1855 7598 1889
rect 7660 2739 7694 2773
rect 7660 2671 7694 2705
rect 7660 2603 7694 2637
rect 7660 2535 7694 2569
rect 7660 2467 7694 2501
rect 7660 2399 7694 2433
rect 7660 2331 7694 2365
rect 7660 2263 7694 2297
rect 7660 2195 7694 2229
rect 7660 2127 7694 2161
rect 7660 2059 7694 2093
rect 7660 1991 7694 2025
rect 7660 1923 7694 1957
rect 7660 1855 7694 1889
rect 7756 2739 7790 2773
rect 7756 2671 7790 2705
rect 7756 2603 7790 2637
rect 7756 2535 7790 2569
rect 7756 2467 7790 2501
rect 7756 2399 7790 2433
rect 7756 2331 7790 2365
rect 7756 2263 7790 2297
rect 7756 2195 7790 2229
rect 7756 2127 7790 2161
rect 7756 2059 7790 2093
rect 7756 1991 7790 2025
rect 7756 1923 7790 1957
rect 7756 1855 7790 1889
rect 7852 2739 7886 2773
rect 7852 2671 7886 2705
rect 7852 2603 7886 2637
rect 7852 2535 7886 2569
rect 7852 2467 7886 2501
rect 10556 2737 10590 2771
rect 10556 2669 10590 2703
rect 10556 2601 10590 2635
rect 10556 2533 10590 2567
rect 10556 2465 10590 2499
rect 7852 2399 7886 2433
rect 7852 2331 7886 2365
rect 7852 2263 7886 2297
rect 10556 2397 10590 2431
rect 10556 2329 10590 2363
rect 7852 2195 7886 2229
rect 7852 2127 7886 2161
rect 7852 2059 7886 2093
rect 8500 2227 8534 2261
rect 8500 2159 8534 2193
rect 8500 2091 8534 2125
rect 8658 2227 8692 2261
rect 8658 2159 8692 2193
rect 8658 2091 8692 2125
rect 10556 2261 10590 2295
rect 10556 2193 10590 2227
rect 10556 2125 10590 2159
rect 10556 2057 10590 2091
rect 7852 1991 7886 2025
rect 7852 1923 7886 1957
rect 7852 1855 7886 1889
rect 10556 1989 10590 2023
rect 10556 1921 10590 1955
rect 10556 1853 10590 1887
rect 10652 2737 10686 2771
rect 10652 2669 10686 2703
rect 10652 2601 10686 2635
rect 10652 2533 10686 2567
rect 10652 2465 10686 2499
rect 10652 2397 10686 2431
rect 10652 2329 10686 2363
rect 10652 2261 10686 2295
rect 10652 2193 10686 2227
rect 10652 2125 10686 2159
rect 10652 2057 10686 2091
rect 10652 1989 10686 2023
rect 10652 1921 10686 1955
rect 10652 1853 10686 1887
rect 10748 2737 10782 2771
rect 10748 2669 10782 2703
rect 10748 2601 10782 2635
rect 10748 2533 10782 2567
rect 10748 2465 10782 2499
rect 10748 2397 10782 2431
rect 10748 2329 10782 2363
rect 10748 2261 10782 2295
rect 10748 2193 10782 2227
rect 10748 2125 10782 2159
rect 10748 2057 10782 2091
rect 10748 1989 10782 2023
rect 10748 1921 10782 1955
rect 10748 1853 10782 1887
rect 10844 2737 10878 2771
rect 10844 2669 10878 2703
rect 10844 2601 10878 2635
rect 10844 2533 10878 2567
rect 10844 2465 10878 2499
rect 10844 2397 10878 2431
rect 10844 2329 10878 2363
rect 10844 2261 10878 2295
rect 10844 2193 10878 2227
rect 10844 2125 10878 2159
rect 10844 2057 10878 2091
rect 10844 1989 10878 2023
rect 10844 1921 10878 1955
rect 10844 1853 10878 1887
rect 10940 2737 10974 2771
rect 10940 2669 10974 2703
rect 10940 2601 10974 2635
rect 10940 2533 10974 2567
rect 10940 2465 10974 2499
rect 13712 2711 13746 2745
rect 13712 2643 13746 2677
rect 13712 2575 13746 2609
rect 13712 2507 13746 2541
rect 10940 2397 10974 2431
rect 10940 2329 10974 2363
rect 10940 2261 10974 2295
rect 13712 2439 13746 2473
rect 13712 2371 13746 2405
rect 13712 2303 13746 2337
rect 10940 2193 10974 2227
rect 10940 2125 10974 2159
rect 10940 2057 10974 2091
rect 11500 2227 11534 2261
rect 11500 2159 11534 2193
rect 11500 2091 11534 2125
rect 11658 2227 11692 2261
rect 11658 2159 11692 2193
rect 11658 2091 11692 2125
rect 13712 2235 13746 2269
rect 13712 2167 13746 2201
rect 13712 2099 13746 2133
rect 10940 1989 10974 2023
rect 10940 1921 10974 1955
rect 10940 1853 10974 1887
rect 13712 2031 13746 2065
rect 13712 1963 13746 1997
rect 13712 1895 13746 1929
rect 13712 1827 13746 1861
rect 13808 2711 13842 2745
rect 13808 2643 13842 2677
rect 13808 2575 13842 2609
rect 13808 2507 13842 2541
rect 13808 2439 13842 2473
rect 13808 2371 13842 2405
rect 13808 2303 13842 2337
rect 13808 2235 13842 2269
rect 13808 2167 13842 2201
rect 13808 2099 13842 2133
rect 13808 2031 13842 2065
rect 13808 1963 13842 1997
rect 13808 1895 13842 1929
rect 13808 1827 13842 1861
rect 13904 2711 13938 2745
rect 13904 2643 13938 2677
rect 13904 2575 13938 2609
rect 13904 2507 13938 2541
rect 13904 2439 13938 2473
rect 13904 2371 13938 2405
rect 13904 2303 13938 2337
rect 13904 2235 13938 2269
rect 13904 2167 13938 2201
rect 13904 2099 13938 2133
rect 13904 2031 13938 2065
rect 13904 1963 13938 1997
rect 13904 1895 13938 1929
rect 13904 1827 13938 1861
rect 14000 2711 14034 2745
rect 14000 2643 14034 2677
rect 14000 2575 14034 2609
rect 14000 2507 14034 2541
rect 14000 2439 14034 2473
rect 14000 2371 14034 2405
rect 14000 2303 14034 2337
rect 14000 2235 14034 2269
rect 14000 2167 14034 2201
rect 14000 2099 14034 2133
rect 14000 2031 14034 2065
rect 14000 1963 14034 1997
rect 14000 1895 14034 1929
rect 14000 1827 14034 1861
rect 14096 2711 14130 2745
rect 14096 2643 14130 2677
rect 14096 2575 14130 2609
rect 14096 2507 14130 2541
rect 14096 2439 14130 2473
rect 14096 2371 14130 2405
rect 14096 2303 14130 2337
rect 14096 2235 14130 2269
rect 14096 2167 14130 2201
rect 14096 2099 14130 2133
rect 14500 2227 14534 2261
rect 14500 2159 14534 2193
rect 14500 2091 14534 2125
rect 14658 2227 14692 2261
rect 14658 2159 14692 2193
rect 14658 2091 14692 2125
rect 14096 2031 14130 2065
rect 14096 1963 14130 1997
rect 14096 1895 14130 1929
rect 14096 1827 14130 1861
rect 158 1193 192 1227
rect 158 1125 192 1159
rect -1686 991 -1652 1025
rect -1686 923 -1652 957
rect -1686 855 -1652 889
rect -1686 787 -1652 821
rect -1686 719 -1652 753
rect -1686 651 -1652 685
rect -1686 583 -1652 617
rect -1686 515 -1652 549
rect -1686 447 -1652 481
rect -1686 379 -1652 413
rect -1686 311 -1652 345
rect -1686 243 -1652 277
rect -1686 175 -1652 209
rect -1686 107 -1652 141
rect -1588 991 -1554 1025
rect -1588 923 -1554 957
rect -1588 855 -1554 889
rect -1588 787 -1554 821
rect -1588 719 -1554 753
rect -1588 651 -1554 685
rect -1588 583 -1554 617
rect -1588 515 -1554 549
rect -1588 447 -1554 481
rect -1588 379 -1554 413
rect -1588 311 -1554 345
rect -1588 243 -1554 277
rect -1588 175 -1554 209
rect -1588 107 -1554 141
rect -1490 991 -1456 1025
rect -1490 923 -1456 957
rect -1490 855 -1456 889
rect -1490 787 -1456 821
rect -1490 719 -1456 753
rect -1490 651 -1456 685
rect -1490 583 -1456 617
rect -1490 515 -1456 549
rect -1490 447 -1456 481
rect -1490 379 -1456 413
rect -1490 311 -1456 345
rect -1490 243 -1456 277
rect -1490 175 -1456 209
rect -1490 107 -1456 141
rect -1392 991 -1358 1025
rect -1392 923 -1358 957
rect -1392 855 -1358 889
rect -1392 787 -1358 821
rect -1392 719 -1358 753
rect -1392 651 -1358 685
rect -1392 583 -1358 617
rect -1392 515 -1358 549
rect -1392 447 -1358 481
rect -1392 379 -1358 413
rect -1392 311 -1358 345
rect -1392 243 -1358 277
rect -1392 175 -1358 209
rect -1392 107 -1358 141
rect -1294 991 -1260 1025
rect -1294 923 -1260 957
rect -1294 855 -1260 889
rect -1294 787 -1260 821
rect -1294 719 -1260 753
rect -1294 651 -1260 685
rect -1294 583 -1260 617
rect -1294 515 -1260 549
rect -1294 447 -1260 481
rect -1294 379 -1260 413
rect -1294 311 -1260 345
rect -1294 243 -1260 277
rect -1294 175 -1260 209
rect -1294 107 -1260 141
rect -1196 991 -1162 1025
rect -1196 923 -1162 957
rect -1196 855 -1162 889
rect -1196 787 -1162 821
rect -1196 719 -1162 753
rect -1196 651 -1162 685
rect -1196 583 -1162 617
rect -1196 515 -1162 549
rect -1196 447 -1162 481
rect -1196 379 -1162 413
rect -1196 311 -1162 345
rect -1196 243 -1162 277
rect -1196 175 -1162 209
rect -1196 107 -1162 141
rect -1098 991 -1064 1025
rect -1098 923 -1064 957
rect -1098 855 -1064 889
rect -1098 787 -1064 821
rect -1098 719 -1064 753
rect -1098 651 -1064 685
rect -1098 583 -1064 617
rect -1098 515 -1064 549
rect -1098 447 -1064 481
rect -1098 379 -1064 413
rect -1098 311 -1064 345
rect -1098 243 -1064 277
rect -1098 175 -1064 209
rect -1098 107 -1064 141
rect -1000 991 -966 1025
rect -1000 923 -966 957
rect -1000 855 -966 889
rect -1000 787 -966 821
rect -1000 719 -966 753
rect -1000 651 -966 685
rect -1000 583 -966 617
rect -1000 515 -966 549
rect -1000 447 -966 481
rect -1000 379 -966 413
rect -1000 311 -966 345
rect -1000 243 -966 277
rect -1000 175 -966 209
rect -1000 107 -966 141
rect -902 991 -868 1025
rect -902 923 -868 957
rect -902 855 -868 889
rect -902 787 -868 821
rect -902 719 -868 753
rect -902 651 -868 685
rect -902 583 -868 617
rect -902 515 -868 549
rect -902 447 -868 481
rect -902 379 -868 413
rect -902 311 -868 345
rect -902 243 -868 277
rect 158 1057 192 1091
rect 158 989 192 1023
rect 158 921 192 955
rect 158 853 192 887
rect 158 785 192 819
rect 158 717 192 751
rect 158 649 192 683
rect 158 581 192 615
rect 158 513 192 547
rect 158 445 192 479
rect 158 377 192 411
rect 158 309 192 343
rect 254 1193 288 1227
rect 254 1125 288 1159
rect 254 1057 288 1091
rect 254 989 288 1023
rect 254 921 288 955
rect 254 853 288 887
rect 254 785 288 819
rect 254 717 288 751
rect 254 649 288 683
rect 254 581 288 615
rect 254 513 288 547
rect 254 445 288 479
rect 254 377 288 411
rect 254 309 288 343
rect 350 1193 384 1227
rect 350 1125 384 1159
rect 350 1057 384 1091
rect 350 989 384 1023
rect 350 921 384 955
rect 350 853 384 887
rect 350 785 384 819
rect 350 717 384 751
rect 350 649 384 683
rect 350 581 384 615
rect 350 513 384 547
rect 350 445 384 479
rect 350 377 384 411
rect 350 309 384 343
rect 446 1193 480 1227
rect 446 1125 480 1159
rect 446 1057 480 1091
rect 446 989 480 1023
rect 446 921 480 955
rect 446 853 480 887
rect 446 785 480 819
rect 446 717 480 751
rect 446 649 480 683
rect 446 581 480 615
rect 446 513 480 547
rect 446 445 480 479
rect 446 377 480 411
rect 446 309 480 343
rect 542 1193 576 1227
rect 542 1125 576 1159
rect 542 1057 576 1091
rect 542 989 576 1023
rect 542 921 576 955
rect 542 853 576 887
rect 542 785 576 819
rect 542 717 576 751
rect 542 649 576 683
rect 542 581 576 615
rect 542 513 576 547
rect 542 445 576 479
rect 542 377 576 411
rect 542 309 576 343
rect 638 1193 672 1227
rect 638 1125 672 1159
rect 638 1057 672 1091
rect 638 989 672 1023
rect 638 921 672 955
rect 638 853 672 887
rect 638 785 672 819
rect 638 717 672 751
rect 638 649 672 683
rect 638 581 672 615
rect 638 513 672 547
rect 638 445 672 479
rect 638 377 672 411
rect 638 309 672 343
rect 734 1193 768 1227
rect 734 1125 768 1159
rect 734 1057 768 1091
rect 734 989 768 1023
rect 734 921 768 955
rect 734 853 768 887
rect 734 785 768 819
rect 734 717 768 751
rect 734 649 768 683
rect 734 581 768 615
rect 734 513 768 547
rect 734 445 768 479
rect 734 377 768 411
rect 734 309 768 343
rect 830 1193 864 1227
rect 830 1125 864 1159
rect 830 1057 864 1091
rect 830 989 864 1023
rect 830 921 864 955
rect 830 853 864 887
rect 830 785 864 819
rect 830 717 864 751
rect 830 649 864 683
rect 830 581 864 615
rect 830 513 864 547
rect 830 445 864 479
rect 830 377 864 411
rect 830 309 864 343
rect 926 1193 960 1227
rect 926 1125 960 1159
rect 926 1057 960 1091
rect 926 989 960 1023
rect 926 921 960 955
rect 926 853 960 887
rect 926 785 960 819
rect 926 717 960 751
rect 926 649 960 683
rect 926 581 960 615
rect 926 513 960 547
rect 926 445 960 479
rect 926 377 960 411
rect 926 309 960 343
rect 1022 1193 1056 1227
rect 1022 1125 1056 1159
rect 1022 1057 1056 1091
rect 1022 989 1056 1023
rect 1022 921 1056 955
rect 1022 853 1056 887
rect 1022 785 1056 819
rect 1022 717 1056 751
rect 1022 649 1056 683
rect 1022 581 1056 615
rect 1022 513 1056 547
rect 1022 445 1056 479
rect 1022 377 1056 411
rect 1022 309 1056 343
rect 1118 1193 1152 1227
rect 1118 1125 1152 1159
rect 1118 1057 1152 1091
rect 1118 989 1152 1023
rect 1118 921 1152 955
rect 1118 853 1152 887
rect 1118 785 1152 819
rect 1118 717 1152 751
rect 1118 649 1152 683
rect 1118 581 1152 615
rect 1118 513 1152 547
rect 1118 445 1152 479
rect 1118 377 1152 411
rect 1118 309 1152 343
rect 1214 1193 1248 1227
rect 1214 1125 1248 1159
rect 1214 1057 1248 1091
rect 1214 989 1248 1023
rect 1214 921 1248 955
rect 1214 853 1248 887
rect 1214 785 1248 819
rect 1214 717 1248 751
rect 1214 649 1248 683
rect 1214 581 1248 615
rect 1214 513 1248 547
rect 1214 445 1248 479
rect 1214 377 1248 411
rect 1214 309 1248 343
rect 1310 1193 1344 1227
rect 1310 1125 1344 1159
rect 1310 1057 1344 1091
rect 1310 989 1344 1023
rect 1310 921 1344 955
rect 1310 853 1344 887
rect 1310 785 1344 819
rect 1310 717 1344 751
rect 1310 649 1344 683
rect 1310 581 1344 615
rect 1310 513 1344 547
rect 1310 445 1344 479
rect 1310 377 1344 411
rect 1310 309 1344 343
rect 1926 1193 1960 1227
rect 1926 1125 1960 1159
rect 1926 1057 1960 1091
rect 1926 989 1960 1023
rect 1926 921 1960 955
rect 1926 853 1960 887
rect 1926 785 1960 819
rect 1926 717 1960 751
rect 1926 649 1960 683
rect 1926 581 1960 615
rect 1926 513 1960 547
rect 1926 445 1960 479
rect 1926 377 1960 411
rect 1926 309 1960 343
rect 2022 1193 2056 1227
rect 2022 1125 2056 1159
rect 2022 1057 2056 1091
rect 2022 989 2056 1023
rect 2022 921 2056 955
rect 2022 853 2056 887
rect 2022 785 2056 819
rect 2022 717 2056 751
rect 2022 649 2056 683
rect 2022 581 2056 615
rect 2022 513 2056 547
rect 2022 445 2056 479
rect 2022 377 2056 411
rect 2022 309 2056 343
rect 2118 1193 2152 1227
rect 2118 1125 2152 1159
rect 2118 1057 2152 1091
rect 2118 989 2152 1023
rect 2118 921 2152 955
rect 2118 853 2152 887
rect 2118 785 2152 819
rect 2118 717 2152 751
rect 2118 649 2152 683
rect 2118 581 2152 615
rect 2118 513 2152 547
rect 2118 445 2152 479
rect 2118 377 2152 411
rect 2118 309 2152 343
rect 2214 1193 2248 1227
rect 2214 1125 2248 1159
rect 2214 1057 2248 1091
rect 2214 989 2248 1023
rect 2214 921 2248 955
rect 2214 853 2248 887
rect 2214 785 2248 819
rect 2214 717 2248 751
rect 2214 649 2248 683
rect 2214 581 2248 615
rect 2214 513 2248 547
rect 2214 445 2248 479
rect 2214 377 2248 411
rect 2214 309 2248 343
rect 2310 1193 2344 1227
rect 2310 1125 2344 1159
rect 2310 1057 2344 1091
rect 2310 989 2344 1023
rect 2310 921 2344 955
rect 2310 853 2344 887
rect 2310 785 2344 819
rect 2310 717 2344 751
rect 2310 649 2344 683
rect 2310 581 2344 615
rect 2310 513 2344 547
rect 2310 445 2344 479
rect 2310 377 2344 411
rect 2310 309 2344 343
rect 2406 1193 2440 1227
rect 2406 1125 2440 1159
rect 2406 1057 2440 1091
rect 2406 989 2440 1023
rect 2406 921 2440 955
rect 2406 853 2440 887
rect 2406 785 2440 819
rect 2406 717 2440 751
rect 2406 649 2440 683
rect 2406 581 2440 615
rect 2406 513 2440 547
rect 2406 445 2440 479
rect 2406 377 2440 411
rect 2406 309 2440 343
rect 2502 1193 2536 1227
rect 2502 1125 2536 1159
rect 2502 1057 2536 1091
rect 2502 989 2536 1023
rect 2502 921 2536 955
rect 2502 853 2536 887
rect 2502 785 2536 819
rect 2502 717 2536 751
rect 2502 649 2536 683
rect 2502 581 2536 615
rect 2502 513 2536 547
rect 2502 445 2536 479
rect 2502 377 2536 411
rect 2502 309 2536 343
rect 2598 1193 2632 1227
rect 2598 1125 2632 1159
rect 2598 1057 2632 1091
rect 2598 989 2632 1023
rect 2598 921 2632 955
rect 2598 853 2632 887
rect 2598 785 2632 819
rect 2598 717 2632 751
rect 2598 649 2632 683
rect 2598 581 2632 615
rect 2598 513 2632 547
rect 2598 445 2632 479
rect 2598 377 2632 411
rect 2598 309 2632 343
rect 2694 1193 2728 1227
rect 2694 1125 2728 1159
rect 2694 1057 2728 1091
rect 2694 989 2728 1023
rect 2694 921 2728 955
rect 2694 853 2728 887
rect 2694 785 2728 819
rect 2694 717 2728 751
rect 2694 649 2728 683
rect 2694 581 2728 615
rect 2694 513 2728 547
rect 2694 445 2728 479
rect 2694 377 2728 411
rect 2694 309 2728 343
rect 2790 1193 2824 1227
rect 2790 1125 2824 1159
rect 2790 1057 2824 1091
rect 2790 989 2824 1023
rect 2790 921 2824 955
rect 2790 853 2824 887
rect 2790 785 2824 819
rect 2790 717 2824 751
rect 2790 649 2824 683
rect 2790 581 2824 615
rect 2790 513 2824 547
rect 2790 445 2824 479
rect 2790 377 2824 411
rect 2790 309 2824 343
rect 2886 1193 2920 1227
rect 2886 1125 2920 1159
rect 2886 1057 2920 1091
rect 2886 989 2920 1023
rect 2886 921 2920 955
rect 2886 853 2920 887
rect 2886 785 2920 819
rect 2886 717 2920 751
rect 2886 649 2920 683
rect 2886 581 2920 615
rect 2886 513 2920 547
rect 2886 445 2920 479
rect 2886 377 2920 411
rect 2886 309 2920 343
rect 2982 1193 3016 1227
rect 2982 1125 3016 1159
rect 2982 1057 3016 1091
rect 2982 989 3016 1023
rect 2982 921 3016 955
rect 2982 853 3016 887
rect 2982 785 3016 819
rect 2982 717 3016 751
rect 2982 649 3016 683
rect 2982 581 3016 615
rect 2982 513 3016 547
rect 2982 445 3016 479
rect 2982 377 3016 411
rect 2982 309 3016 343
rect 3114 1177 3148 1211
rect 3114 1109 3148 1143
rect 3114 1041 3148 1075
rect 3114 973 3148 1007
rect 3114 905 3148 939
rect 3114 837 3148 871
rect 3114 769 3148 803
rect 3114 701 3148 735
rect 3114 633 3148 667
rect 3114 565 3148 599
rect 3114 497 3148 531
rect 3114 429 3148 463
rect 3114 361 3148 395
rect 3114 293 3148 327
rect -902 175 -868 209
rect 3210 1177 3244 1211
rect 3210 1109 3244 1143
rect 3210 1041 3244 1075
rect 3210 973 3244 1007
rect 3210 905 3244 939
rect 3210 837 3244 871
rect 3210 769 3244 803
rect 3210 701 3244 735
rect 3210 633 3244 667
rect 3210 565 3244 599
rect 3210 497 3244 531
rect 3210 429 3244 463
rect 3210 361 3244 395
rect 3210 293 3244 327
rect 3306 1177 3340 1211
rect 3306 1109 3340 1143
rect 3306 1041 3340 1075
rect 3306 973 3340 1007
rect 3306 905 3340 939
rect 3306 837 3340 871
rect 3306 769 3340 803
rect 3306 701 3340 735
rect 3306 633 3340 667
rect 3306 565 3340 599
rect 3306 497 3340 531
rect 3306 429 3340 463
rect 3306 361 3340 395
rect 3306 293 3340 327
rect 3402 1177 3436 1211
rect 3402 1109 3436 1143
rect 3402 1041 3436 1075
rect 3402 973 3436 1007
rect 3402 905 3436 939
rect 3402 837 3436 871
rect 3402 769 3436 803
rect 3402 701 3436 735
rect 3402 633 3436 667
rect 3402 565 3436 599
rect 3402 497 3436 531
rect 3402 429 3436 463
rect 3402 361 3436 395
rect 3402 293 3436 327
rect 3498 1177 3532 1211
rect 3498 1109 3532 1143
rect 3498 1041 3532 1075
rect 3498 973 3532 1007
rect 3498 905 3532 939
rect 3498 837 3532 871
rect 3498 769 3532 803
rect 3498 701 3532 735
rect 3498 633 3532 667
rect 3498 565 3532 599
rect 3498 497 3532 531
rect 3498 429 3532 463
rect 3498 361 3532 395
rect 3498 293 3532 327
rect 3594 1177 3628 1211
rect 3594 1109 3628 1143
rect 3594 1041 3628 1075
rect 3594 973 3628 1007
rect 3594 905 3628 939
rect 3594 837 3628 871
rect 3594 769 3628 803
rect 3594 701 3628 735
rect 3594 633 3628 667
rect 3594 565 3628 599
rect 3594 497 3628 531
rect 3594 429 3628 463
rect 3594 361 3628 395
rect 3594 293 3628 327
rect 3690 1177 3724 1211
rect 3690 1109 3724 1143
rect 3690 1041 3724 1075
rect 3690 973 3724 1007
rect 3690 905 3724 939
rect 3690 837 3724 871
rect 3690 769 3724 803
rect 3690 701 3724 735
rect 3690 633 3724 667
rect 3690 565 3724 599
rect 3690 497 3724 531
rect 3690 429 3724 463
rect 3690 361 3724 395
rect 3690 293 3724 327
rect 3786 1177 3820 1211
rect 3786 1109 3820 1143
rect 3786 1041 3820 1075
rect 3786 973 3820 1007
rect 3786 905 3820 939
rect 3786 837 3820 871
rect 3786 769 3820 803
rect 3786 701 3820 735
rect 3786 633 3820 667
rect 3786 565 3820 599
rect 3786 497 3820 531
rect 3786 429 3820 463
rect 3786 361 3820 395
rect 3786 293 3820 327
rect 3882 1177 3916 1211
rect 3882 1109 3916 1143
rect 3882 1041 3916 1075
rect 3882 973 3916 1007
rect 3882 905 3916 939
rect 3882 837 3916 871
rect 3882 769 3916 803
rect 3882 701 3916 735
rect 3882 633 3916 667
rect 3882 565 3916 599
rect 3882 497 3916 531
rect 3882 429 3916 463
rect 3882 361 3916 395
rect 3882 293 3916 327
rect 3978 1177 4012 1211
rect 3978 1109 4012 1143
rect 3978 1041 4012 1075
rect 3978 973 4012 1007
rect 3978 905 4012 939
rect 3978 837 4012 871
rect 3978 769 4012 803
rect 3978 701 4012 735
rect 3978 633 4012 667
rect 3978 565 4012 599
rect 3978 497 4012 531
rect 3978 429 4012 463
rect 3978 361 4012 395
rect 3978 293 4012 327
rect 4074 1177 4108 1211
rect 4074 1109 4108 1143
rect 4074 1041 4108 1075
rect 4074 973 4108 1007
rect 4074 905 4108 939
rect 4074 837 4108 871
rect 4074 769 4108 803
rect 4074 701 4108 735
rect 4074 633 4108 667
rect 4074 565 4108 599
rect 4074 497 4108 531
rect 4074 429 4108 463
rect 4074 361 4108 395
rect 4074 293 4108 327
rect 4170 1177 4204 1211
rect 4170 1109 4204 1143
rect 4170 1041 4204 1075
rect 4170 973 4204 1007
rect 4170 905 4204 939
rect 4170 837 4204 871
rect 4170 769 4204 803
rect 4170 701 4204 735
rect 4170 633 4204 667
rect 4170 565 4204 599
rect 4170 497 4204 531
rect 4170 429 4204 463
rect 4170 361 4204 395
rect 4170 293 4204 327
rect 4266 1177 4300 1211
rect 4266 1109 4300 1143
rect 4266 1041 4300 1075
rect 4266 973 4300 1007
rect 4266 905 4300 939
rect 4266 837 4300 871
rect 4266 769 4300 803
rect 4266 701 4300 735
rect 4266 633 4300 667
rect 4266 565 4300 599
rect 4266 497 4300 531
rect 4266 429 4300 463
rect 4266 361 4300 395
rect 4266 293 4300 327
rect 4882 1177 4916 1211
rect 4882 1109 4916 1143
rect 4882 1041 4916 1075
rect 4882 973 4916 1007
rect 4882 905 4916 939
rect 4882 837 4916 871
rect 4882 769 4916 803
rect 4882 701 4916 735
rect 4882 633 4916 667
rect 4882 565 4916 599
rect 4882 497 4916 531
rect 4882 429 4916 463
rect 4882 361 4916 395
rect 4882 293 4916 327
rect 4978 1177 5012 1211
rect 4978 1109 5012 1143
rect 4978 1041 5012 1075
rect 4978 973 5012 1007
rect 4978 905 5012 939
rect 4978 837 5012 871
rect 4978 769 5012 803
rect 4978 701 5012 735
rect 4978 633 5012 667
rect 4978 565 5012 599
rect 4978 497 5012 531
rect 4978 429 5012 463
rect 4978 361 5012 395
rect 4978 293 5012 327
rect 5074 1177 5108 1211
rect 5074 1109 5108 1143
rect 5074 1041 5108 1075
rect 5074 973 5108 1007
rect 5074 905 5108 939
rect 5074 837 5108 871
rect 5074 769 5108 803
rect 5074 701 5108 735
rect 5074 633 5108 667
rect 5074 565 5108 599
rect 5074 497 5108 531
rect 5074 429 5108 463
rect 5074 361 5108 395
rect 5074 293 5108 327
rect 5170 1177 5204 1211
rect 5170 1109 5204 1143
rect 5170 1041 5204 1075
rect 5170 973 5204 1007
rect 5170 905 5204 939
rect 5170 837 5204 871
rect 5170 769 5204 803
rect 5170 701 5204 735
rect 5170 633 5204 667
rect 5170 565 5204 599
rect 5170 497 5204 531
rect 5170 429 5204 463
rect 5170 361 5204 395
rect 5170 293 5204 327
rect 5266 1177 5300 1211
rect 5266 1109 5300 1143
rect 5266 1041 5300 1075
rect 5266 973 5300 1007
rect 5266 905 5300 939
rect 5266 837 5300 871
rect 5266 769 5300 803
rect 5266 701 5300 735
rect 5266 633 5300 667
rect 5266 565 5300 599
rect 5266 497 5300 531
rect 5266 429 5300 463
rect 5266 361 5300 395
rect 5266 293 5300 327
rect 5362 1177 5396 1211
rect 5362 1109 5396 1143
rect 5362 1041 5396 1075
rect 5362 973 5396 1007
rect 5362 905 5396 939
rect 5362 837 5396 871
rect 5362 769 5396 803
rect 5362 701 5396 735
rect 5362 633 5396 667
rect 5362 565 5396 599
rect 5362 497 5396 531
rect 5362 429 5396 463
rect 5362 361 5396 395
rect 5362 293 5396 327
rect 5458 1177 5492 1211
rect 5458 1109 5492 1143
rect 5458 1041 5492 1075
rect 5458 973 5492 1007
rect 5458 905 5492 939
rect 5458 837 5492 871
rect 5458 769 5492 803
rect 5458 701 5492 735
rect 5458 633 5492 667
rect 5458 565 5492 599
rect 5458 497 5492 531
rect 5458 429 5492 463
rect 5458 361 5492 395
rect 5458 293 5492 327
rect 5554 1177 5588 1211
rect 5554 1109 5588 1143
rect 5554 1041 5588 1075
rect 5554 973 5588 1007
rect 5554 905 5588 939
rect 5554 837 5588 871
rect 5554 769 5588 803
rect 5554 701 5588 735
rect 5554 633 5588 667
rect 5554 565 5588 599
rect 5554 497 5588 531
rect 5554 429 5588 463
rect 5554 361 5588 395
rect 5554 293 5588 327
rect 5650 1177 5684 1211
rect 5650 1109 5684 1143
rect 5650 1041 5684 1075
rect 5650 973 5684 1007
rect 5650 905 5684 939
rect 5650 837 5684 871
rect 5650 769 5684 803
rect 5650 701 5684 735
rect 5650 633 5684 667
rect 5650 565 5684 599
rect 5650 497 5684 531
rect 5650 429 5684 463
rect 5650 361 5684 395
rect 5650 293 5684 327
rect 5746 1177 5780 1211
rect 5746 1109 5780 1143
rect 5746 1041 5780 1075
rect 5746 973 5780 1007
rect 5746 905 5780 939
rect 5746 837 5780 871
rect 5746 769 5780 803
rect 5746 701 5780 735
rect 5746 633 5780 667
rect 5746 565 5780 599
rect 5746 497 5780 531
rect 5746 429 5780 463
rect 5746 361 5780 395
rect 5746 293 5780 327
rect 5842 1177 5876 1211
rect 5842 1109 5876 1143
rect 5842 1041 5876 1075
rect 5842 973 5876 1007
rect 5842 905 5876 939
rect 5842 837 5876 871
rect 5842 769 5876 803
rect 5842 701 5876 735
rect 5842 633 5876 667
rect 5842 565 5876 599
rect 5842 497 5876 531
rect 5842 429 5876 463
rect 5842 361 5876 395
rect 5842 293 5876 327
rect 5938 1177 5972 1211
rect 5938 1109 5972 1143
rect 5938 1041 5972 1075
rect 5938 973 5972 1007
rect 5938 905 5972 939
rect 5938 837 5972 871
rect 5938 769 5972 803
rect 5938 701 5972 735
rect 5938 633 5972 667
rect 5938 565 5972 599
rect 5938 497 5972 531
rect 5938 429 5972 463
rect 5938 361 5972 395
rect 5938 293 5972 327
rect 6144 1177 6178 1211
rect 6144 1109 6178 1143
rect 6144 1041 6178 1075
rect 6144 973 6178 1007
rect 6144 905 6178 939
rect 6144 837 6178 871
rect 6144 769 6178 803
rect 6144 701 6178 735
rect 6144 633 6178 667
rect 6144 565 6178 599
rect 6144 497 6178 531
rect 6144 429 6178 463
rect 6144 361 6178 395
rect 6144 293 6178 327
rect 6240 1177 6274 1211
rect 6240 1109 6274 1143
rect 6240 1041 6274 1075
rect 6240 973 6274 1007
rect 6240 905 6274 939
rect 6240 837 6274 871
rect 6240 769 6274 803
rect 6240 701 6274 735
rect 6240 633 6274 667
rect 6240 565 6274 599
rect 6240 497 6274 531
rect 6240 429 6274 463
rect 6240 361 6274 395
rect 6240 293 6274 327
rect 6336 1177 6370 1211
rect 6336 1109 6370 1143
rect 6336 1041 6370 1075
rect 6336 973 6370 1007
rect 6336 905 6370 939
rect 6336 837 6370 871
rect 6336 769 6370 803
rect 6336 701 6370 735
rect 6336 633 6370 667
rect 6336 565 6370 599
rect 6336 497 6370 531
rect 6336 429 6370 463
rect 6336 361 6370 395
rect 6336 293 6370 327
rect 6432 1177 6466 1211
rect 6432 1109 6466 1143
rect 6432 1041 6466 1075
rect 6432 973 6466 1007
rect 6432 905 6466 939
rect 6432 837 6466 871
rect 6432 769 6466 803
rect 6432 701 6466 735
rect 6432 633 6466 667
rect 6432 565 6466 599
rect 6432 497 6466 531
rect 6432 429 6466 463
rect 6432 361 6466 395
rect 6432 293 6466 327
rect 6528 1177 6562 1211
rect 6528 1109 6562 1143
rect 6528 1041 6562 1075
rect 6528 973 6562 1007
rect 6528 905 6562 939
rect 6528 837 6562 871
rect 6528 769 6562 803
rect 6528 701 6562 735
rect 6528 633 6562 667
rect 6528 565 6562 599
rect 6528 497 6562 531
rect 6528 429 6562 463
rect 6528 361 6562 395
rect 6528 293 6562 327
rect 6624 1177 6658 1211
rect 6624 1109 6658 1143
rect 6624 1041 6658 1075
rect 6624 973 6658 1007
rect 6624 905 6658 939
rect 6624 837 6658 871
rect 6624 769 6658 803
rect 6624 701 6658 735
rect 6624 633 6658 667
rect 6624 565 6658 599
rect 6624 497 6658 531
rect 6624 429 6658 463
rect 6624 361 6658 395
rect 6624 293 6658 327
rect 6720 1177 6754 1211
rect 6720 1109 6754 1143
rect 6720 1041 6754 1075
rect 6720 973 6754 1007
rect 6720 905 6754 939
rect 6720 837 6754 871
rect 6720 769 6754 803
rect 6720 701 6754 735
rect 6720 633 6754 667
rect 6720 565 6754 599
rect 6720 497 6754 531
rect 6720 429 6754 463
rect 6720 361 6754 395
rect 6720 293 6754 327
rect 6816 1177 6850 1211
rect 6816 1109 6850 1143
rect 6816 1041 6850 1075
rect 6816 973 6850 1007
rect 6816 905 6850 939
rect 6816 837 6850 871
rect 6816 769 6850 803
rect 6816 701 6850 735
rect 6816 633 6850 667
rect 6816 565 6850 599
rect 6816 497 6850 531
rect 6816 429 6850 463
rect 6816 361 6850 395
rect 6816 293 6850 327
rect 6912 1177 6946 1211
rect 6912 1109 6946 1143
rect 6912 1041 6946 1075
rect 6912 973 6946 1007
rect 6912 905 6946 939
rect 6912 837 6946 871
rect 6912 769 6946 803
rect 6912 701 6946 735
rect 6912 633 6946 667
rect 6912 565 6946 599
rect 6912 497 6946 531
rect 6912 429 6946 463
rect 6912 361 6946 395
rect 6912 293 6946 327
rect 7008 1177 7042 1211
rect 7008 1109 7042 1143
rect 7008 1041 7042 1075
rect 7008 973 7042 1007
rect 7008 905 7042 939
rect 7008 837 7042 871
rect 7008 769 7042 803
rect 7008 701 7042 735
rect 7008 633 7042 667
rect 7008 565 7042 599
rect 7008 497 7042 531
rect 7008 429 7042 463
rect 7008 361 7042 395
rect 7008 293 7042 327
rect 7104 1177 7138 1211
rect 7104 1109 7138 1143
rect 7104 1041 7138 1075
rect 7104 973 7138 1007
rect 7104 905 7138 939
rect 7104 837 7138 871
rect 7104 769 7138 803
rect 7104 701 7138 735
rect 7104 633 7138 667
rect 7104 565 7138 599
rect 7104 497 7138 531
rect 7104 429 7138 463
rect 7104 361 7138 395
rect 7104 293 7138 327
rect 7200 1177 7234 1211
rect 7200 1109 7234 1143
rect 7200 1041 7234 1075
rect 7200 973 7234 1007
rect 7200 905 7234 939
rect 7200 837 7234 871
rect 7200 769 7234 803
rect 7200 701 7234 735
rect 7200 633 7234 667
rect 7200 565 7234 599
rect 7200 497 7234 531
rect 7200 429 7234 463
rect 7200 361 7234 395
rect 7200 293 7234 327
rect 7296 1177 7330 1211
rect 7296 1109 7330 1143
rect 7296 1041 7330 1075
rect 7296 973 7330 1007
rect 7296 905 7330 939
rect 7296 837 7330 871
rect 7296 769 7330 803
rect 7296 701 7330 735
rect 7296 633 7330 667
rect 7296 565 7330 599
rect 7296 497 7330 531
rect 7296 429 7330 463
rect 7296 361 7330 395
rect 7296 293 7330 327
rect 7912 1177 7946 1211
rect 7912 1109 7946 1143
rect 7912 1041 7946 1075
rect 7912 973 7946 1007
rect 7912 905 7946 939
rect 7912 837 7946 871
rect 7912 769 7946 803
rect 7912 701 7946 735
rect 7912 633 7946 667
rect 7912 565 7946 599
rect 7912 497 7946 531
rect 7912 429 7946 463
rect 7912 361 7946 395
rect 7912 293 7946 327
rect 8008 1177 8042 1211
rect 8008 1109 8042 1143
rect 8008 1041 8042 1075
rect 8008 973 8042 1007
rect 8008 905 8042 939
rect 8008 837 8042 871
rect 8008 769 8042 803
rect 8008 701 8042 735
rect 8008 633 8042 667
rect 8008 565 8042 599
rect 8008 497 8042 531
rect 8008 429 8042 463
rect 8008 361 8042 395
rect 8008 293 8042 327
rect 8104 1177 8138 1211
rect 8104 1109 8138 1143
rect 8104 1041 8138 1075
rect 8104 973 8138 1007
rect 8104 905 8138 939
rect 8104 837 8138 871
rect 8104 769 8138 803
rect 8104 701 8138 735
rect 8104 633 8138 667
rect 8104 565 8138 599
rect 8104 497 8138 531
rect 8104 429 8138 463
rect 8104 361 8138 395
rect 8104 293 8138 327
rect 8200 1177 8234 1211
rect 8200 1109 8234 1143
rect 8200 1041 8234 1075
rect 8200 973 8234 1007
rect 8200 905 8234 939
rect 8200 837 8234 871
rect 8200 769 8234 803
rect 8200 701 8234 735
rect 8200 633 8234 667
rect 8200 565 8234 599
rect 8200 497 8234 531
rect 8200 429 8234 463
rect 8200 361 8234 395
rect 8200 293 8234 327
rect 8296 1177 8330 1211
rect 8296 1109 8330 1143
rect 8296 1041 8330 1075
rect 8296 973 8330 1007
rect 8296 905 8330 939
rect 8296 837 8330 871
rect 8296 769 8330 803
rect 8296 701 8330 735
rect 8296 633 8330 667
rect 8296 565 8330 599
rect 8296 497 8330 531
rect 8296 429 8330 463
rect 8296 361 8330 395
rect 8296 293 8330 327
rect 8392 1177 8426 1211
rect 8392 1109 8426 1143
rect 8392 1041 8426 1075
rect 8392 973 8426 1007
rect 8392 905 8426 939
rect 8392 837 8426 871
rect 8392 769 8426 803
rect 8392 701 8426 735
rect 8392 633 8426 667
rect 8392 565 8426 599
rect 8392 497 8426 531
rect 8392 429 8426 463
rect 8392 361 8426 395
rect 8392 293 8426 327
rect 8488 1177 8522 1211
rect 8488 1109 8522 1143
rect 8488 1041 8522 1075
rect 8488 973 8522 1007
rect 8488 905 8522 939
rect 8488 837 8522 871
rect 8488 769 8522 803
rect 8488 701 8522 735
rect 8488 633 8522 667
rect 8488 565 8522 599
rect 8488 497 8522 531
rect 8488 429 8522 463
rect 8488 361 8522 395
rect 8488 293 8522 327
rect 8584 1177 8618 1211
rect 8584 1109 8618 1143
rect 8584 1041 8618 1075
rect 8584 973 8618 1007
rect 8584 905 8618 939
rect 8584 837 8618 871
rect 8584 769 8618 803
rect 8584 701 8618 735
rect 8584 633 8618 667
rect 8584 565 8618 599
rect 8584 497 8618 531
rect 8584 429 8618 463
rect 8584 361 8618 395
rect 8584 293 8618 327
rect 8680 1177 8714 1211
rect 8680 1109 8714 1143
rect 8680 1041 8714 1075
rect 8680 973 8714 1007
rect 8680 905 8714 939
rect 8680 837 8714 871
rect 8680 769 8714 803
rect 8680 701 8714 735
rect 8680 633 8714 667
rect 8680 565 8714 599
rect 8680 497 8714 531
rect 8680 429 8714 463
rect 8680 361 8714 395
rect 8680 293 8714 327
rect 8776 1177 8810 1211
rect 8776 1109 8810 1143
rect 8776 1041 8810 1075
rect 8776 973 8810 1007
rect 8776 905 8810 939
rect 8776 837 8810 871
rect 8776 769 8810 803
rect 8776 701 8810 735
rect 8776 633 8810 667
rect 8776 565 8810 599
rect 8776 497 8810 531
rect 8776 429 8810 463
rect 8776 361 8810 395
rect 8776 293 8810 327
rect 8872 1177 8906 1211
rect 8872 1109 8906 1143
rect 8872 1041 8906 1075
rect 8872 973 8906 1007
rect 8872 905 8906 939
rect 8872 837 8906 871
rect 8872 769 8906 803
rect 8872 701 8906 735
rect 8872 633 8906 667
rect 8872 565 8906 599
rect 8872 497 8906 531
rect 8872 429 8906 463
rect 8872 361 8906 395
rect 8872 293 8906 327
rect 8968 1177 9002 1211
rect 8968 1109 9002 1143
rect 8968 1041 9002 1075
rect 8968 973 9002 1007
rect 8968 905 9002 939
rect 8968 837 9002 871
rect 8968 769 9002 803
rect 8968 701 9002 735
rect 8968 633 9002 667
rect 8968 565 9002 599
rect 8968 497 9002 531
rect 8968 429 9002 463
rect 8968 361 9002 395
rect 8968 293 9002 327
rect 9232 1175 9266 1209
rect 9232 1107 9266 1141
rect 9232 1039 9266 1073
rect 9232 971 9266 1005
rect 9232 903 9266 937
rect 9232 835 9266 869
rect 9232 767 9266 801
rect 9232 699 9266 733
rect 9232 631 9266 665
rect 9232 563 9266 597
rect 9232 495 9266 529
rect 9232 427 9266 461
rect 9232 359 9266 393
rect 9232 291 9266 325
rect -902 107 -868 141
rect 9328 1175 9362 1209
rect 9328 1107 9362 1141
rect 9328 1039 9362 1073
rect 9328 971 9362 1005
rect 9328 903 9362 937
rect 9328 835 9362 869
rect 9328 767 9362 801
rect 9328 699 9362 733
rect 9328 631 9362 665
rect 9328 563 9362 597
rect 9328 495 9362 529
rect 9328 427 9362 461
rect 9328 359 9362 393
rect 9328 291 9362 325
rect 9424 1175 9458 1209
rect 9424 1107 9458 1141
rect 9424 1039 9458 1073
rect 9424 971 9458 1005
rect 9424 903 9458 937
rect 9424 835 9458 869
rect 9424 767 9458 801
rect 9424 699 9458 733
rect 9424 631 9458 665
rect 9424 563 9458 597
rect 9424 495 9458 529
rect 9424 427 9458 461
rect 9424 359 9458 393
rect 9424 291 9458 325
rect 9520 1175 9554 1209
rect 9520 1107 9554 1141
rect 9520 1039 9554 1073
rect 9520 971 9554 1005
rect 9520 903 9554 937
rect 9520 835 9554 869
rect 9520 767 9554 801
rect 9520 699 9554 733
rect 9520 631 9554 665
rect 9520 563 9554 597
rect 9520 495 9554 529
rect 9520 427 9554 461
rect 9520 359 9554 393
rect 9520 291 9554 325
rect 9616 1175 9650 1209
rect 9616 1107 9650 1141
rect 9616 1039 9650 1073
rect 9616 971 9650 1005
rect 9616 903 9650 937
rect 9616 835 9650 869
rect 9616 767 9650 801
rect 9616 699 9650 733
rect 9616 631 9650 665
rect 9616 563 9650 597
rect 9616 495 9650 529
rect 9616 427 9650 461
rect 9616 359 9650 393
rect 9616 291 9650 325
rect 9712 1175 9746 1209
rect 9712 1107 9746 1141
rect 9712 1039 9746 1073
rect 9712 971 9746 1005
rect 9712 903 9746 937
rect 9712 835 9746 869
rect 9712 767 9746 801
rect 9712 699 9746 733
rect 9712 631 9746 665
rect 9712 563 9746 597
rect 9712 495 9746 529
rect 9712 427 9746 461
rect 9712 359 9746 393
rect 9712 291 9746 325
rect 9808 1175 9842 1209
rect 9808 1107 9842 1141
rect 9808 1039 9842 1073
rect 9808 971 9842 1005
rect 9808 903 9842 937
rect 9808 835 9842 869
rect 9808 767 9842 801
rect 9808 699 9842 733
rect 9808 631 9842 665
rect 9808 563 9842 597
rect 9808 495 9842 529
rect 9808 427 9842 461
rect 9808 359 9842 393
rect 9808 291 9842 325
rect 9904 1175 9938 1209
rect 9904 1107 9938 1141
rect 9904 1039 9938 1073
rect 9904 971 9938 1005
rect 9904 903 9938 937
rect 9904 835 9938 869
rect 9904 767 9938 801
rect 9904 699 9938 733
rect 9904 631 9938 665
rect 9904 563 9938 597
rect 9904 495 9938 529
rect 9904 427 9938 461
rect 9904 359 9938 393
rect 9904 291 9938 325
rect 10000 1175 10034 1209
rect 10000 1107 10034 1141
rect 10000 1039 10034 1073
rect 10000 971 10034 1005
rect 10000 903 10034 937
rect 10000 835 10034 869
rect 10000 767 10034 801
rect 10000 699 10034 733
rect 10000 631 10034 665
rect 10000 563 10034 597
rect 10000 495 10034 529
rect 10000 427 10034 461
rect 10000 359 10034 393
rect 10000 291 10034 325
rect 10096 1175 10130 1209
rect 10096 1107 10130 1141
rect 10096 1039 10130 1073
rect 10096 971 10130 1005
rect 10096 903 10130 937
rect 10096 835 10130 869
rect 10096 767 10130 801
rect 10096 699 10130 733
rect 10096 631 10130 665
rect 10096 563 10130 597
rect 10096 495 10130 529
rect 10096 427 10130 461
rect 10096 359 10130 393
rect 10096 291 10130 325
rect 10192 1175 10226 1209
rect 10192 1107 10226 1141
rect 10192 1039 10226 1073
rect 10192 971 10226 1005
rect 10192 903 10226 937
rect 10192 835 10226 869
rect 10192 767 10226 801
rect 10192 699 10226 733
rect 10192 631 10226 665
rect 10192 563 10226 597
rect 10192 495 10226 529
rect 10192 427 10226 461
rect 10192 359 10226 393
rect 10192 291 10226 325
rect 10288 1175 10322 1209
rect 10288 1107 10322 1141
rect 10288 1039 10322 1073
rect 10288 971 10322 1005
rect 10288 903 10322 937
rect 10288 835 10322 869
rect 10288 767 10322 801
rect 10288 699 10322 733
rect 10288 631 10322 665
rect 10288 563 10322 597
rect 10288 495 10322 529
rect 10288 427 10322 461
rect 10288 359 10322 393
rect 10288 291 10322 325
rect 10384 1175 10418 1209
rect 10384 1107 10418 1141
rect 10384 1039 10418 1073
rect 10384 971 10418 1005
rect 10384 903 10418 937
rect 10384 835 10418 869
rect 10384 767 10418 801
rect 10384 699 10418 733
rect 10384 631 10418 665
rect 10384 563 10418 597
rect 10384 495 10418 529
rect 10384 427 10418 461
rect 10384 359 10418 393
rect 10384 291 10418 325
rect 11000 1175 11034 1209
rect 11000 1107 11034 1141
rect 11000 1039 11034 1073
rect 11000 971 11034 1005
rect 11000 903 11034 937
rect 11000 835 11034 869
rect 11000 767 11034 801
rect 11000 699 11034 733
rect 11000 631 11034 665
rect 11000 563 11034 597
rect 11000 495 11034 529
rect 11000 427 11034 461
rect 11000 359 11034 393
rect 11000 291 11034 325
rect 11096 1175 11130 1209
rect 11096 1107 11130 1141
rect 11096 1039 11130 1073
rect 11096 971 11130 1005
rect 11096 903 11130 937
rect 11096 835 11130 869
rect 11096 767 11130 801
rect 11096 699 11130 733
rect 11096 631 11130 665
rect 11096 563 11130 597
rect 11096 495 11130 529
rect 11096 427 11130 461
rect 11096 359 11130 393
rect 11096 291 11130 325
rect 11192 1175 11226 1209
rect 11192 1107 11226 1141
rect 11192 1039 11226 1073
rect 11192 971 11226 1005
rect 11192 903 11226 937
rect 11192 835 11226 869
rect 11192 767 11226 801
rect 11192 699 11226 733
rect 11192 631 11226 665
rect 11192 563 11226 597
rect 11192 495 11226 529
rect 11192 427 11226 461
rect 11192 359 11226 393
rect 11192 291 11226 325
rect 11288 1175 11322 1209
rect 11288 1107 11322 1141
rect 11288 1039 11322 1073
rect 11288 971 11322 1005
rect 11288 903 11322 937
rect 11288 835 11322 869
rect 11288 767 11322 801
rect 11288 699 11322 733
rect 11288 631 11322 665
rect 11288 563 11322 597
rect 11288 495 11322 529
rect 11288 427 11322 461
rect 11288 359 11322 393
rect 11288 291 11322 325
rect 11384 1175 11418 1209
rect 11384 1107 11418 1141
rect 11384 1039 11418 1073
rect 11384 971 11418 1005
rect 11384 903 11418 937
rect 11384 835 11418 869
rect 11384 767 11418 801
rect 11384 699 11418 733
rect 11384 631 11418 665
rect 11384 563 11418 597
rect 11384 495 11418 529
rect 11384 427 11418 461
rect 11384 359 11418 393
rect 11384 291 11418 325
rect 11480 1175 11514 1209
rect 11480 1107 11514 1141
rect 11480 1039 11514 1073
rect 11480 971 11514 1005
rect 11480 903 11514 937
rect 11480 835 11514 869
rect 11480 767 11514 801
rect 11480 699 11514 733
rect 11480 631 11514 665
rect 11480 563 11514 597
rect 11480 495 11514 529
rect 11480 427 11514 461
rect 11480 359 11514 393
rect 11480 291 11514 325
rect 11576 1175 11610 1209
rect 11576 1107 11610 1141
rect 11576 1039 11610 1073
rect 11576 971 11610 1005
rect 11576 903 11610 937
rect 11576 835 11610 869
rect 11576 767 11610 801
rect 11576 699 11610 733
rect 11576 631 11610 665
rect 11576 563 11610 597
rect 11576 495 11610 529
rect 11576 427 11610 461
rect 11576 359 11610 393
rect 11576 291 11610 325
rect 11672 1175 11706 1209
rect 11672 1107 11706 1141
rect 11672 1039 11706 1073
rect 11672 971 11706 1005
rect 11672 903 11706 937
rect 11672 835 11706 869
rect 11672 767 11706 801
rect 11672 699 11706 733
rect 11672 631 11706 665
rect 11672 563 11706 597
rect 11672 495 11706 529
rect 11672 427 11706 461
rect 11672 359 11706 393
rect 11672 291 11706 325
rect 11768 1175 11802 1209
rect 11768 1107 11802 1141
rect 11768 1039 11802 1073
rect 11768 971 11802 1005
rect 11768 903 11802 937
rect 11768 835 11802 869
rect 11768 767 11802 801
rect 11768 699 11802 733
rect 11768 631 11802 665
rect 11768 563 11802 597
rect 11768 495 11802 529
rect 11768 427 11802 461
rect 11768 359 11802 393
rect 11768 291 11802 325
rect 11864 1175 11898 1209
rect 11864 1107 11898 1141
rect 11864 1039 11898 1073
rect 11864 971 11898 1005
rect 11864 903 11898 937
rect 11864 835 11898 869
rect 11864 767 11898 801
rect 11864 699 11898 733
rect 11864 631 11898 665
rect 11864 563 11898 597
rect 11864 495 11898 529
rect 11864 427 11898 461
rect 11864 359 11898 393
rect 11864 291 11898 325
rect 11960 1175 11994 1209
rect 11960 1107 11994 1141
rect 11960 1039 11994 1073
rect 11960 971 11994 1005
rect 11960 903 11994 937
rect 11960 835 11994 869
rect 11960 767 11994 801
rect 11960 699 11994 733
rect 11960 631 11994 665
rect 11960 563 11994 597
rect 11960 495 11994 529
rect 11960 427 11994 461
rect 11960 359 11994 393
rect 11960 291 11994 325
rect 15422 1227 15456 1261
rect 12056 1175 12090 1209
rect 12056 1107 12090 1141
rect 12056 1039 12090 1073
rect 12056 971 12090 1005
rect 12056 903 12090 937
rect 12056 835 12090 869
rect 12056 767 12090 801
rect 12056 699 12090 733
rect 12056 631 12090 665
rect 12056 563 12090 597
rect 12056 495 12090 529
rect 12056 427 12090 461
rect 12056 359 12090 393
rect 12056 291 12090 325
rect 12388 1149 12422 1183
rect 12388 1081 12422 1115
rect 12388 1013 12422 1047
rect 12388 945 12422 979
rect 12388 877 12422 911
rect 12388 809 12422 843
rect 12388 741 12422 775
rect 12388 673 12422 707
rect 12388 605 12422 639
rect 12388 537 12422 571
rect 12388 469 12422 503
rect 12388 401 12422 435
rect 12388 333 12422 367
rect 12388 265 12422 299
rect 12484 1149 12518 1183
rect 12484 1081 12518 1115
rect 12484 1013 12518 1047
rect 12484 945 12518 979
rect 12484 877 12518 911
rect 12484 809 12518 843
rect 12484 741 12518 775
rect 12484 673 12518 707
rect 12484 605 12518 639
rect 12484 537 12518 571
rect 12484 469 12518 503
rect 12484 401 12518 435
rect 12484 333 12518 367
rect 12484 265 12518 299
rect 12580 1149 12614 1183
rect 12580 1081 12614 1115
rect 12580 1013 12614 1047
rect 12580 945 12614 979
rect 12580 877 12614 911
rect 12580 809 12614 843
rect 12580 741 12614 775
rect 12580 673 12614 707
rect 12580 605 12614 639
rect 12580 537 12614 571
rect 12580 469 12614 503
rect 12580 401 12614 435
rect 12580 333 12614 367
rect 12580 265 12614 299
rect 12676 1149 12710 1183
rect 12676 1081 12710 1115
rect 12676 1013 12710 1047
rect 12676 945 12710 979
rect 12676 877 12710 911
rect 12676 809 12710 843
rect 12676 741 12710 775
rect 12676 673 12710 707
rect 12676 605 12710 639
rect 12676 537 12710 571
rect 12676 469 12710 503
rect 12676 401 12710 435
rect 12676 333 12710 367
rect 12676 265 12710 299
rect 12772 1149 12806 1183
rect 12772 1081 12806 1115
rect 12772 1013 12806 1047
rect 12772 945 12806 979
rect 12772 877 12806 911
rect 12772 809 12806 843
rect 12772 741 12806 775
rect 12772 673 12806 707
rect 12772 605 12806 639
rect 12772 537 12806 571
rect 12772 469 12806 503
rect 12772 401 12806 435
rect 12772 333 12806 367
rect 12772 265 12806 299
rect 12868 1149 12902 1183
rect 12868 1081 12902 1115
rect 12868 1013 12902 1047
rect 12868 945 12902 979
rect 12868 877 12902 911
rect 12868 809 12902 843
rect 12868 741 12902 775
rect 12868 673 12902 707
rect 12868 605 12902 639
rect 12868 537 12902 571
rect 12868 469 12902 503
rect 12868 401 12902 435
rect 12868 333 12902 367
rect 12868 265 12902 299
rect 12964 1149 12998 1183
rect 12964 1081 12998 1115
rect 12964 1013 12998 1047
rect 12964 945 12998 979
rect 12964 877 12998 911
rect 12964 809 12998 843
rect 12964 741 12998 775
rect 12964 673 12998 707
rect 12964 605 12998 639
rect 12964 537 12998 571
rect 12964 469 12998 503
rect 12964 401 12998 435
rect 12964 333 12998 367
rect 12964 265 12998 299
rect 13060 1149 13094 1183
rect 13060 1081 13094 1115
rect 13060 1013 13094 1047
rect 13060 945 13094 979
rect 13060 877 13094 911
rect 13060 809 13094 843
rect 13060 741 13094 775
rect 13060 673 13094 707
rect 13060 605 13094 639
rect 13060 537 13094 571
rect 13060 469 13094 503
rect 13060 401 13094 435
rect 13060 333 13094 367
rect 13060 265 13094 299
rect 13156 1149 13190 1183
rect 13156 1081 13190 1115
rect 13156 1013 13190 1047
rect 13156 945 13190 979
rect 13156 877 13190 911
rect 13156 809 13190 843
rect 13156 741 13190 775
rect 13156 673 13190 707
rect 13156 605 13190 639
rect 13156 537 13190 571
rect 13156 469 13190 503
rect 13156 401 13190 435
rect 13156 333 13190 367
rect 13156 265 13190 299
rect 13252 1149 13286 1183
rect 13252 1081 13286 1115
rect 13252 1013 13286 1047
rect 13252 945 13286 979
rect 13252 877 13286 911
rect 13252 809 13286 843
rect 13252 741 13286 775
rect 13252 673 13286 707
rect 13252 605 13286 639
rect 13252 537 13286 571
rect 13252 469 13286 503
rect 13252 401 13286 435
rect 13252 333 13286 367
rect 13252 265 13286 299
rect 13348 1149 13382 1183
rect 13348 1081 13382 1115
rect 13348 1013 13382 1047
rect 13348 945 13382 979
rect 13348 877 13382 911
rect 13348 809 13382 843
rect 13348 741 13382 775
rect 13348 673 13382 707
rect 13348 605 13382 639
rect 13348 537 13382 571
rect 13348 469 13382 503
rect 13348 401 13382 435
rect 13348 333 13382 367
rect 13348 265 13382 299
rect 13444 1149 13478 1183
rect 13444 1081 13478 1115
rect 13444 1013 13478 1047
rect 13444 945 13478 979
rect 13444 877 13478 911
rect 13444 809 13478 843
rect 13444 741 13478 775
rect 13444 673 13478 707
rect 13444 605 13478 639
rect 13444 537 13478 571
rect 13444 469 13478 503
rect 13444 401 13478 435
rect 13444 333 13478 367
rect 13444 265 13478 299
rect 13540 1149 13574 1183
rect 13540 1081 13574 1115
rect 13540 1013 13574 1047
rect 13540 945 13574 979
rect 13540 877 13574 911
rect 13540 809 13574 843
rect 13540 741 13574 775
rect 13540 673 13574 707
rect 13540 605 13574 639
rect 13540 537 13574 571
rect 13540 469 13574 503
rect 13540 401 13574 435
rect 13540 333 13574 367
rect 13540 265 13574 299
rect 14156 1149 14190 1183
rect 14156 1081 14190 1115
rect 14156 1013 14190 1047
rect 14156 945 14190 979
rect 14156 877 14190 911
rect 14156 809 14190 843
rect 14156 741 14190 775
rect 14156 673 14190 707
rect 14156 605 14190 639
rect 14156 537 14190 571
rect 14156 469 14190 503
rect 14156 401 14190 435
rect 14156 333 14190 367
rect 14156 265 14190 299
rect 14252 1149 14286 1183
rect 14252 1081 14286 1115
rect 14252 1013 14286 1047
rect 14252 945 14286 979
rect 14252 877 14286 911
rect 14252 809 14286 843
rect 14252 741 14286 775
rect 14252 673 14286 707
rect 14252 605 14286 639
rect 14252 537 14286 571
rect 14252 469 14286 503
rect 14252 401 14286 435
rect 14252 333 14286 367
rect 14252 265 14286 299
rect 14348 1149 14382 1183
rect 14348 1081 14382 1115
rect 14348 1013 14382 1047
rect 14348 945 14382 979
rect 14348 877 14382 911
rect 14348 809 14382 843
rect 14348 741 14382 775
rect 14348 673 14382 707
rect 14348 605 14382 639
rect 14348 537 14382 571
rect 14348 469 14382 503
rect 14348 401 14382 435
rect 14348 333 14382 367
rect 14348 265 14382 299
rect 14444 1149 14478 1183
rect 14444 1081 14478 1115
rect 14444 1013 14478 1047
rect 14444 945 14478 979
rect 14444 877 14478 911
rect 14444 809 14478 843
rect 14444 741 14478 775
rect 14444 673 14478 707
rect 14444 605 14478 639
rect 14444 537 14478 571
rect 14444 469 14478 503
rect 14444 401 14478 435
rect 14444 333 14478 367
rect 14444 265 14478 299
rect 14540 1149 14574 1183
rect 14540 1081 14574 1115
rect 14540 1013 14574 1047
rect 14540 945 14574 979
rect 14540 877 14574 911
rect 14540 809 14574 843
rect 14540 741 14574 775
rect 14540 673 14574 707
rect 14540 605 14574 639
rect 14540 537 14574 571
rect 14540 469 14574 503
rect 14540 401 14574 435
rect 14540 333 14574 367
rect 14540 265 14574 299
rect 14636 1149 14670 1183
rect 14636 1081 14670 1115
rect 14636 1013 14670 1047
rect 14636 945 14670 979
rect 14636 877 14670 911
rect 14636 809 14670 843
rect 14636 741 14670 775
rect 14636 673 14670 707
rect 14636 605 14670 639
rect 14636 537 14670 571
rect 14636 469 14670 503
rect 14636 401 14670 435
rect 14636 333 14670 367
rect 14636 265 14670 299
rect 14732 1149 14766 1183
rect 14732 1081 14766 1115
rect 14732 1013 14766 1047
rect 14732 945 14766 979
rect 14732 877 14766 911
rect 14732 809 14766 843
rect 14732 741 14766 775
rect 14732 673 14766 707
rect 14732 605 14766 639
rect 14732 537 14766 571
rect 14732 469 14766 503
rect 14732 401 14766 435
rect 14732 333 14766 367
rect 14732 265 14766 299
rect 14828 1149 14862 1183
rect 14828 1081 14862 1115
rect 14828 1013 14862 1047
rect 14828 945 14862 979
rect 14828 877 14862 911
rect 14828 809 14862 843
rect 14828 741 14862 775
rect 14828 673 14862 707
rect 14828 605 14862 639
rect 14828 537 14862 571
rect 14828 469 14862 503
rect 14828 401 14862 435
rect 14828 333 14862 367
rect 14828 265 14862 299
rect 14924 1149 14958 1183
rect 14924 1081 14958 1115
rect 14924 1013 14958 1047
rect 14924 945 14958 979
rect 14924 877 14958 911
rect 14924 809 14958 843
rect 14924 741 14958 775
rect 14924 673 14958 707
rect 14924 605 14958 639
rect 14924 537 14958 571
rect 14924 469 14958 503
rect 14924 401 14958 435
rect 14924 333 14958 367
rect 14924 265 14958 299
rect 15020 1149 15054 1183
rect 15020 1081 15054 1115
rect 15020 1013 15054 1047
rect 15020 945 15054 979
rect 15020 877 15054 911
rect 15020 809 15054 843
rect 15020 741 15054 775
rect 15020 673 15054 707
rect 15020 605 15054 639
rect 15020 537 15054 571
rect 15020 469 15054 503
rect 15020 401 15054 435
rect 15020 333 15054 367
rect 15020 265 15054 299
rect 15116 1149 15150 1183
rect 15116 1081 15150 1115
rect 15116 1013 15150 1047
rect 15116 945 15150 979
rect 15116 877 15150 911
rect 15116 809 15150 843
rect 15116 741 15150 775
rect 15116 673 15150 707
rect 15116 605 15150 639
rect 15116 537 15150 571
rect 15116 469 15150 503
rect 15116 401 15150 435
rect 15116 333 15150 367
rect 15116 265 15150 299
rect 15212 1149 15246 1183
rect 15212 1081 15246 1115
rect 15212 1013 15246 1047
rect 15212 945 15246 979
rect 15212 877 15246 911
rect 15212 809 15246 843
rect 15212 741 15246 775
rect 15212 673 15246 707
rect 15212 605 15246 639
rect 15212 537 15246 571
rect 15212 469 15246 503
rect 15212 401 15246 435
rect 15212 333 15246 367
rect 15212 265 15246 299
rect 15422 1159 15456 1193
rect 15422 1091 15456 1125
rect 15422 1023 15456 1057
rect 15422 955 15456 989
rect 15422 887 15456 921
rect 15422 819 15456 853
rect 15422 751 15456 785
rect 15422 683 15456 717
rect 15422 615 15456 649
rect 15422 547 15456 581
rect 15422 479 15456 513
rect 15422 411 15456 445
rect 15422 343 15456 377
rect 15422 275 15456 309
rect 15422 207 15456 241
rect 15422 139 15456 173
rect 15510 1227 15544 1261
rect 15510 1159 15544 1193
rect 15510 1091 15544 1125
rect 15510 1023 15544 1057
rect 15510 955 15544 989
rect 15510 887 15544 921
rect 15510 819 15544 853
rect 15510 751 15544 785
rect 15510 683 15544 717
rect 15510 615 15544 649
rect 15510 547 15544 581
rect 15510 479 15544 513
rect 15510 411 15544 445
rect 15510 343 15544 377
rect 15510 275 15544 309
rect 15510 207 15544 241
rect 15510 139 15544 173
<< pdiffc >>
rect 194 6531 228 6565
rect 194 6463 228 6497
rect 194 6395 228 6429
rect 194 6327 228 6361
rect 194 6259 228 6293
rect 194 6191 228 6225
rect 194 6123 228 6157
rect 194 6055 228 6089
rect 194 5987 228 6021
rect -1652 5861 -1618 5895
rect -1652 5793 -1618 5827
rect -1652 5725 -1618 5759
rect -1652 5657 -1618 5691
rect -1652 5589 -1618 5623
rect -1652 5521 -1618 5555
rect -1652 5453 -1618 5487
rect -1652 5385 -1618 5419
rect -1652 5317 -1618 5351
rect -1652 5249 -1618 5283
rect -1652 5181 -1618 5215
rect -1652 5113 -1618 5147
rect -1652 5045 -1618 5079
rect -1652 4977 -1618 5011
rect -1554 5861 -1520 5895
rect -1554 5793 -1520 5827
rect -1554 5725 -1520 5759
rect -1554 5657 -1520 5691
rect -1554 5589 -1520 5623
rect -1554 5521 -1520 5555
rect -1554 5453 -1520 5487
rect -1554 5385 -1520 5419
rect -1554 5317 -1520 5351
rect -1554 5249 -1520 5283
rect -1554 5181 -1520 5215
rect -1554 5113 -1520 5147
rect -1554 5045 -1520 5079
rect -1554 4977 -1520 5011
rect -1456 5861 -1422 5895
rect -1456 5793 -1422 5827
rect -1456 5725 -1422 5759
rect -1456 5657 -1422 5691
rect -1456 5589 -1422 5623
rect -1456 5521 -1422 5555
rect -1456 5453 -1422 5487
rect -1456 5385 -1422 5419
rect -1456 5317 -1422 5351
rect -1456 5249 -1422 5283
rect -1456 5181 -1422 5215
rect -1456 5113 -1422 5147
rect -1456 5045 -1422 5079
rect -1456 4977 -1422 5011
rect -1358 5861 -1324 5895
rect -1358 5793 -1324 5827
rect -1358 5725 -1324 5759
rect -1358 5657 -1324 5691
rect -1358 5589 -1324 5623
rect -1358 5521 -1324 5555
rect -1358 5453 -1324 5487
rect -1358 5385 -1324 5419
rect -1358 5317 -1324 5351
rect -1358 5249 -1324 5283
rect -1358 5181 -1324 5215
rect -1358 5113 -1324 5147
rect -1358 5045 -1324 5079
rect -1358 4977 -1324 5011
rect -1260 5861 -1226 5895
rect -1260 5793 -1226 5827
rect -1260 5725 -1226 5759
rect -1260 5657 -1226 5691
rect -1260 5589 -1226 5623
rect -1260 5521 -1226 5555
rect -1260 5453 -1226 5487
rect -1260 5385 -1226 5419
rect -1260 5317 -1226 5351
rect -1260 5249 -1226 5283
rect -1260 5181 -1226 5215
rect -1260 5113 -1226 5147
rect -1260 5045 -1226 5079
rect -1260 4977 -1226 5011
rect -1162 5861 -1128 5895
rect -1162 5793 -1128 5827
rect -1162 5725 -1128 5759
rect -1162 5657 -1128 5691
rect -1162 5589 -1128 5623
rect -1162 5521 -1128 5555
rect -1162 5453 -1128 5487
rect -1162 5385 -1128 5419
rect -1162 5317 -1128 5351
rect -1162 5249 -1128 5283
rect -1162 5181 -1128 5215
rect -1162 5113 -1128 5147
rect -1162 5045 -1128 5079
rect -1162 4977 -1128 5011
rect -1064 5861 -1030 5895
rect -1064 5793 -1030 5827
rect -1064 5725 -1030 5759
rect -1064 5657 -1030 5691
rect -1064 5589 -1030 5623
rect -1064 5521 -1030 5555
rect -1064 5453 -1030 5487
rect -1064 5385 -1030 5419
rect -1064 5317 -1030 5351
rect -1064 5249 -1030 5283
rect -1064 5181 -1030 5215
rect -1064 5113 -1030 5147
rect -1064 5045 -1030 5079
rect -1064 4977 -1030 5011
rect -966 5861 -932 5895
rect -966 5793 -932 5827
rect -966 5725 -932 5759
rect -966 5657 -932 5691
rect -966 5589 -932 5623
rect -966 5521 -932 5555
rect -966 5453 -932 5487
rect -966 5385 -932 5419
rect -966 5317 -932 5351
rect -966 5249 -932 5283
rect -966 5181 -932 5215
rect -966 5113 -932 5147
rect -966 5045 -932 5079
rect -966 4977 -932 5011
rect -868 5861 -834 5895
rect -868 5793 -834 5827
rect -868 5725 -834 5759
rect -868 5657 -834 5691
rect -868 5589 -834 5623
rect 194 5919 228 5953
rect 194 5851 228 5885
rect 194 5783 228 5817
rect 194 5715 228 5749
rect 194 5647 228 5681
rect 290 6531 324 6565
rect 290 6463 324 6497
rect 290 6395 324 6429
rect 290 6327 324 6361
rect 290 6259 324 6293
rect 290 6191 324 6225
rect 290 6123 324 6157
rect 290 6055 324 6089
rect 290 5987 324 6021
rect 290 5919 324 5953
rect 290 5851 324 5885
rect 290 5783 324 5817
rect 290 5715 324 5749
rect 290 5647 324 5681
rect 386 6531 420 6565
rect 386 6463 420 6497
rect 386 6395 420 6429
rect 386 6327 420 6361
rect 386 6259 420 6293
rect 386 6191 420 6225
rect 386 6123 420 6157
rect 386 6055 420 6089
rect 386 5987 420 6021
rect 386 5919 420 5953
rect 386 5851 420 5885
rect 386 5783 420 5817
rect 386 5715 420 5749
rect 386 5647 420 5681
rect 482 6531 516 6565
rect 482 6463 516 6497
rect 482 6395 516 6429
rect 482 6327 516 6361
rect 482 6259 516 6293
rect 482 6191 516 6225
rect 482 6123 516 6157
rect 482 6055 516 6089
rect 482 5987 516 6021
rect 482 5919 516 5953
rect 482 5851 516 5885
rect 482 5783 516 5817
rect 482 5715 516 5749
rect 482 5647 516 5681
rect 578 6531 612 6565
rect 578 6463 612 6497
rect 578 6395 612 6429
rect 578 6327 612 6361
rect 578 6259 612 6293
rect 578 6191 612 6225
rect 578 6123 612 6157
rect 578 6055 612 6089
rect 578 5987 612 6021
rect 578 5919 612 5953
rect 578 5851 612 5885
rect 578 5783 612 5817
rect 578 5715 612 5749
rect 578 5647 612 5681
rect 674 6531 708 6565
rect 674 6463 708 6497
rect 674 6395 708 6429
rect 674 6327 708 6361
rect 674 6259 708 6293
rect 674 6191 708 6225
rect 674 6123 708 6157
rect 674 6055 708 6089
rect 674 5987 708 6021
rect 674 5919 708 5953
rect 674 5851 708 5885
rect 674 5783 708 5817
rect 674 5715 708 5749
rect 674 5647 708 5681
rect 770 6531 804 6565
rect 770 6463 804 6497
rect 770 6395 804 6429
rect 770 6327 804 6361
rect 770 6259 804 6293
rect 770 6191 804 6225
rect 770 6123 804 6157
rect 770 6055 804 6089
rect 770 5987 804 6021
rect 770 5919 804 5953
rect 770 5851 804 5885
rect 770 5783 804 5817
rect 770 5715 804 5749
rect 770 5647 804 5681
rect 866 6531 900 6565
rect 866 6463 900 6497
rect 866 6395 900 6429
rect 866 6327 900 6361
rect 866 6259 900 6293
rect 866 6191 900 6225
rect 866 6123 900 6157
rect 866 6055 900 6089
rect 866 5987 900 6021
rect 866 5919 900 5953
rect 866 5851 900 5885
rect 866 5783 900 5817
rect 866 5715 900 5749
rect 866 5647 900 5681
rect 962 6531 996 6565
rect 962 6463 996 6497
rect 962 6395 996 6429
rect 962 6327 996 6361
rect 962 6259 996 6293
rect 962 6191 996 6225
rect 962 6123 996 6157
rect 962 6055 996 6089
rect 962 5987 996 6021
rect 962 5919 996 5953
rect 962 5851 996 5885
rect 962 5783 996 5817
rect 962 5715 996 5749
rect 962 5647 996 5681
rect 1058 6531 1092 6565
rect 1058 6463 1092 6497
rect 1058 6395 1092 6429
rect 1058 6327 1092 6361
rect 1058 6259 1092 6293
rect 1058 6191 1092 6225
rect 1058 6123 1092 6157
rect 1058 6055 1092 6089
rect 1058 5987 1092 6021
rect 1058 5919 1092 5953
rect 1058 5851 1092 5885
rect 1058 5783 1092 5817
rect 1058 5715 1092 5749
rect 1058 5647 1092 5681
rect 1154 6531 1188 6565
rect 1154 6463 1188 6497
rect 1154 6395 1188 6429
rect 1154 6327 1188 6361
rect 1154 6259 1188 6293
rect 1154 6191 1188 6225
rect 1154 6123 1188 6157
rect 1154 6055 1188 6089
rect 1154 5987 1188 6021
rect 1154 5919 1188 5953
rect 1154 5851 1188 5885
rect 1154 5783 1188 5817
rect 1154 5715 1188 5749
rect 1154 5647 1188 5681
rect 1250 6531 1284 6565
rect 1250 6463 1284 6497
rect 1250 6395 1284 6429
rect 1250 6327 1284 6361
rect 1250 6259 1284 6293
rect 1250 6191 1284 6225
rect 1250 6123 1284 6157
rect 1250 6055 1284 6089
rect 1250 5987 1284 6021
rect 1250 5919 1284 5953
rect 1250 5851 1284 5885
rect 1250 5783 1284 5817
rect 1250 5715 1284 5749
rect 1250 5647 1284 5681
rect 1346 6531 1380 6565
rect 1346 6463 1380 6497
rect 1346 6395 1380 6429
rect 1346 6327 1380 6361
rect 1346 6259 1380 6293
rect 1346 6191 1380 6225
rect 1346 6123 1380 6157
rect 1346 6055 1380 6089
rect 1346 5987 1380 6021
rect 1346 5919 1380 5953
rect 1346 5851 1380 5885
rect 1346 5783 1380 5817
rect 1346 5715 1380 5749
rect 1346 5647 1380 5681
rect 1960 6527 1994 6561
rect 1960 6459 1994 6493
rect 1960 6391 1994 6425
rect 1960 6323 1994 6357
rect 1960 6255 1994 6289
rect 1960 6187 1994 6221
rect 1960 6119 1994 6153
rect 1960 6051 1994 6085
rect 1960 5983 1994 6017
rect 1960 5915 1994 5949
rect 1960 5847 1994 5881
rect 1960 5779 1994 5813
rect 1960 5711 1994 5745
rect 1960 5643 1994 5677
rect 2056 6527 2090 6561
rect 2056 6459 2090 6493
rect 2056 6391 2090 6425
rect 2056 6323 2090 6357
rect 2056 6255 2090 6289
rect 2056 6187 2090 6221
rect 2056 6119 2090 6153
rect 2056 6051 2090 6085
rect 2056 5983 2090 6017
rect 2056 5915 2090 5949
rect 2056 5847 2090 5881
rect 2056 5779 2090 5813
rect 2056 5711 2090 5745
rect 2056 5643 2090 5677
rect 2152 6527 2186 6561
rect 2152 6459 2186 6493
rect 2152 6391 2186 6425
rect 2152 6323 2186 6357
rect 2152 6255 2186 6289
rect 2152 6187 2186 6221
rect 2152 6119 2186 6153
rect 2152 6051 2186 6085
rect 2152 5983 2186 6017
rect 2152 5915 2186 5949
rect 2152 5847 2186 5881
rect 2152 5779 2186 5813
rect 2152 5711 2186 5745
rect 2152 5643 2186 5677
rect 2248 6527 2282 6561
rect 2248 6459 2282 6493
rect 2248 6391 2282 6425
rect 2248 6323 2282 6357
rect 2248 6255 2282 6289
rect 2248 6187 2282 6221
rect 2248 6119 2282 6153
rect 2248 6051 2282 6085
rect 2248 5983 2282 6017
rect 2248 5915 2282 5949
rect 2248 5847 2282 5881
rect 2248 5779 2282 5813
rect 2248 5711 2282 5745
rect 2248 5643 2282 5677
rect 2344 6527 2378 6561
rect 2344 6459 2378 6493
rect 2344 6391 2378 6425
rect 2344 6323 2378 6357
rect 2344 6255 2378 6289
rect 2344 6187 2378 6221
rect 2344 6119 2378 6153
rect 2344 6051 2378 6085
rect 2344 5983 2378 6017
rect 2344 5915 2378 5949
rect 2344 5847 2378 5881
rect 2344 5779 2378 5813
rect 2344 5711 2378 5745
rect 2344 5643 2378 5677
rect 2440 6527 2474 6561
rect 2440 6459 2474 6493
rect 2440 6391 2474 6425
rect 2440 6323 2474 6357
rect 2440 6255 2474 6289
rect 2440 6187 2474 6221
rect 2440 6119 2474 6153
rect 2440 6051 2474 6085
rect 2440 5983 2474 6017
rect 2440 5915 2474 5949
rect 2440 5847 2474 5881
rect 2440 5779 2474 5813
rect 2440 5711 2474 5745
rect 2440 5643 2474 5677
rect 2536 6527 2570 6561
rect 2536 6459 2570 6493
rect 2536 6391 2570 6425
rect 2536 6323 2570 6357
rect 2536 6255 2570 6289
rect 2536 6187 2570 6221
rect 2536 6119 2570 6153
rect 2536 6051 2570 6085
rect 2536 5983 2570 6017
rect 2536 5915 2570 5949
rect 2536 5847 2570 5881
rect 2536 5779 2570 5813
rect 2536 5711 2570 5745
rect 2536 5643 2570 5677
rect 2632 6527 2666 6561
rect 2632 6459 2666 6493
rect 2632 6391 2666 6425
rect 2632 6323 2666 6357
rect 2632 6255 2666 6289
rect 2632 6187 2666 6221
rect 2632 6119 2666 6153
rect 2632 6051 2666 6085
rect 2632 5983 2666 6017
rect 2632 5915 2666 5949
rect 2632 5847 2666 5881
rect 2632 5779 2666 5813
rect 2632 5711 2666 5745
rect 2632 5643 2666 5677
rect 2728 6527 2762 6561
rect 2728 6459 2762 6493
rect 2728 6391 2762 6425
rect 2728 6323 2762 6357
rect 2728 6255 2762 6289
rect 2728 6187 2762 6221
rect 2728 6119 2762 6153
rect 2728 6051 2762 6085
rect 2728 5983 2762 6017
rect 2728 5915 2762 5949
rect 2728 5847 2762 5881
rect 2728 5779 2762 5813
rect 2728 5711 2762 5745
rect 2728 5643 2762 5677
rect 3150 6515 3184 6549
rect 3150 6447 3184 6481
rect 3150 6379 3184 6413
rect 3150 6311 3184 6345
rect 3150 6243 3184 6277
rect 3150 6175 3184 6209
rect 3150 6107 3184 6141
rect 3150 6039 3184 6073
rect 3150 5971 3184 6005
rect 3150 5903 3184 5937
rect 3150 5835 3184 5869
rect 3150 5767 3184 5801
rect 3150 5699 3184 5733
rect 3150 5631 3184 5665
rect 3246 6515 3280 6549
rect 3246 6447 3280 6481
rect 3246 6379 3280 6413
rect 3246 6311 3280 6345
rect 3246 6243 3280 6277
rect 3246 6175 3280 6209
rect 3246 6107 3280 6141
rect 3246 6039 3280 6073
rect 3246 5971 3280 6005
rect 3246 5903 3280 5937
rect 3246 5835 3280 5869
rect 3246 5767 3280 5801
rect 3246 5699 3280 5733
rect 3246 5631 3280 5665
rect 3342 6515 3376 6549
rect 3342 6447 3376 6481
rect 3342 6379 3376 6413
rect 3342 6311 3376 6345
rect 3342 6243 3376 6277
rect 3342 6175 3376 6209
rect 3342 6107 3376 6141
rect 3342 6039 3376 6073
rect 3342 5971 3376 6005
rect 3342 5903 3376 5937
rect 3342 5835 3376 5869
rect 3342 5767 3376 5801
rect 3342 5699 3376 5733
rect 3342 5631 3376 5665
rect 3438 6515 3472 6549
rect 3438 6447 3472 6481
rect 3438 6379 3472 6413
rect 3438 6311 3472 6345
rect 3438 6243 3472 6277
rect 3438 6175 3472 6209
rect 3438 6107 3472 6141
rect 3438 6039 3472 6073
rect 3438 5971 3472 6005
rect 3438 5903 3472 5937
rect 3438 5835 3472 5869
rect 3438 5767 3472 5801
rect 3438 5699 3472 5733
rect 3438 5631 3472 5665
rect 3534 6515 3568 6549
rect 3534 6447 3568 6481
rect 3534 6379 3568 6413
rect 3534 6311 3568 6345
rect 3534 6243 3568 6277
rect 3534 6175 3568 6209
rect 3534 6107 3568 6141
rect 3534 6039 3568 6073
rect 3534 5971 3568 6005
rect 3534 5903 3568 5937
rect 3534 5835 3568 5869
rect 3534 5767 3568 5801
rect 3534 5699 3568 5733
rect 3534 5631 3568 5665
rect 3630 6515 3664 6549
rect 3630 6447 3664 6481
rect 3630 6379 3664 6413
rect 3630 6311 3664 6345
rect 3630 6243 3664 6277
rect 3630 6175 3664 6209
rect 3630 6107 3664 6141
rect 3630 6039 3664 6073
rect 3630 5971 3664 6005
rect 3630 5903 3664 5937
rect 3630 5835 3664 5869
rect 3630 5767 3664 5801
rect 3630 5699 3664 5733
rect 3630 5631 3664 5665
rect 3726 6515 3760 6549
rect 3726 6447 3760 6481
rect 3726 6379 3760 6413
rect 3726 6311 3760 6345
rect 3726 6243 3760 6277
rect 3726 6175 3760 6209
rect 3726 6107 3760 6141
rect 3726 6039 3760 6073
rect 3726 5971 3760 6005
rect 3726 5903 3760 5937
rect 3726 5835 3760 5869
rect 3726 5767 3760 5801
rect 3726 5699 3760 5733
rect 3726 5631 3760 5665
rect 3822 6515 3856 6549
rect 3822 6447 3856 6481
rect 3822 6379 3856 6413
rect 3822 6311 3856 6345
rect 3822 6243 3856 6277
rect 3822 6175 3856 6209
rect 3822 6107 3856 6141
rect 3822 6039 3856 6073
rect 3822 5971 3856 6005
rect 3822 5903 3856 5937
rect 3822 5835 3856 5869
rect 3822 5767 3856 5801
rect 3822 5699 3856 5733
rect 3822 5631 3856 5665
rect 3918 6515 3952 6549
rect 3918 6447 3952 6481
rect 3918 6379 3952 6413
rect 3918 6311 3952 6345
rect 3918 6243 3952 6277
rect 3918 6175 3952 6209
rect 3918 6107 3952 6141
rect 3918 6039 3952 6073
rect 3918 5971 3952 6005
rect 3918 5903 3952 5937
rect 3918 5835 3952 5869
rect 3918 5767 3952 5801
rect 3918 5699 3952 5733
rect 3918 5631 3952 5665
rect 4014 6515 4048 6549
rect 4014 6447 4048 6481
rect 4014 6379 4048 6413
rect 4014 6311 4048 6345
rect 4014 6243 4048 6277
rect 4014 6175 4048 6209
rect 4014 6107 4048 6141
rect 4014 6039 4048 6073
rect 4014 5971 4048 6005
rect 4014 5903 4048 5937
rect 4014 5835 4048 5869
rect 4014 5767 4048 5801
rect 4014 5699 4048 5733
rect 4014 5631 4048 5665
rect 4110 6515 4144 6549
rect 4110 6447 4144 6481
rect 4110 6379 4144 6413
rect 4110 6311 4144 6345
rect 4110 6243 4144 6277
rect 4110 6175 4144 6209
rect 4110 6107 4144 6141
rect 4110 6039 4144 6073
rect 4110 5971 4144 6005
rect 4110 5903 4144 5937
rect 4110 5835 4144 5869
rect 4110 5767 4144 5801
rect 4110 5699 4144 5733
rect 4110 5631 4144 5665
rect 4206 6515 4240 6549
rect 4206 6447 4240 6481
rect 4206 6379 4240 6413
rect 4206 6311 4240 6345
rect 4206 6243 4240 6277
rect 4206 6175 4240 6209
rect 4206 6107 4240 6141
rect 4206 6039 4240 6073
rect 4206 5971 4240 6005
rect 4206 5903 4240 5937
rect 4206 5835 4240 5869
rect 4206 5767 4240 5801
rect 4206 5699 4240 5733
rect 4206 5631 4240 5665
rect 4302 6515 4336 6549
rect 4302 6447 4336 6481
rect 4302 6379 4336 6413
rect 4302 6311 4336 6345
rect 4302 6243 4336 6277
rect 4302 6175 4336 6209
rect 4302 6107 4336 6141
rect 4302 6039 4336 6073
rect 4302 5971 4336 6005
rect 4302 5903 4336 5937
rect 4302 5835 4336 5869
rect 4302 5767 4336 5801
rect 4302 5699 4336 5733
rect 4302 5631 4336 5665
rect 4916 6511 4950 6545
rect 4916 6443 4950 6477
rect 4916 6375 4950 6409
rect 4916 6307 4950 6341
rect 4916 6239 4950 6273
rect 4916 6171 4950 6205
rect 4916 6103 4950 6137
rect 4916 6035 4950 6069
rect 4916 5967 4950 6001
rect 4916 5899 4950 5933
rect 4916 5831 4950 5865
rect 4916 5763 4950 5797
rect 4916 5695 4950 5729
rect 4916 5627 4950 5661
rect 5012 6511 5046 6545
rect 5012 6443 5046 6477
rect 5012 6375 5046 6409
rect 5012 6307 5046 6341
rect 5012 6239 5046 6273
rect 5012 6171 5046 6205
rect 5012 6103 5046 6137
rect 5012 6035 5046 6069
rect 5012 5967 5046 6001
rect 5012 5899 5046 5933
rect 5012 5831 5046 5865
rect 5012 5763 5046 5797
rect 5012 5695 5046 5729
rect 5012 5627 5046 5661
rect 5108 6511 5142 6545
rect 5108 6443 5142 6477
rect 5108 6375 5142 6409
rect 5108 6307 5142 6341
rect 5108 6239 5142 6273
rect 5108 6171 5142 6205
rect 5108 6103 5142 6137
rect 5108 6035 5142 6069
rect 5108 5967 5142 6001
rect 5108 5899 5142 5933
rect 5108 5831 5142 5865
rect 5108 5763 5142 5797
rect 5108 5695 5142 5729
rect 5108 5627 5142 5661
rect 5204 6511 5238 6545
rect 5204 6443 5238 6477
rect 5204 6375 5238 6409
rect 5204 6307 5238 6341
rect 5204 6239 5238 6273
rect 5204 6171 5238 6205
rect 5204 6103 5238 6137
rect 5204 6035 5238 6069
rect 5204 5967 5238 6001
rect 5204 5899 5238 5933
rect 5204 5831 5238 5865
rect 5204 5763 5238 5797
rect 5204 5695 5238 5729
rect 5204 5627 5238 5661
rect 5300 6511 5334 6545
rect 5300 6443 5334 6477
rect 5300 6375 5334 6409
rect 5300 6307 5334 6341
rect 5300 6239 5334 6273
rect 5300 6171 5334 6205
rect 5300 6103 5334 6137
rect 5300 6035 5334 6069
rect 5300 5967 5334 6001
rect 5300 5899 5334 5933
rect 5300 5831 5334 5865
rect 5300 5763 5334 5797
rect 5300 5695 5334 5729
rect 5300 5627 5334 5661
rect 5396 6511 5430 6545
rect 5396 6443 5430 6477
rect 5396 6375 5430 6409
rect 5396 6307 5430 6341
rect 5396 6239 5430 6273
rect 5396 6171 5430 6205
rect 5396 6103 5430 6137
rect 5396 6035 5430 6069
rect 5396 5967 5430 6001
rect 5396 5899 5430 5933
rect 5396 5831 5430 5865
rect 5396 5763 5430 5797
rect 5396 5695 5430 5729
rect 5396 5627 5430 5661
rect 5492 6511 5526 6545
rect 5492 6443 5526 6477
rect 5492 6375 5526 6409
rect 5492 6307 5526 6341
rect 5492 6239 5526 6273
rect 5492 6171 5526 6205
rect 5492 6103 5526 6137
rect 5492 6035 5526 6069
rect 5492 5967 5526 6001
rect 5492 5899 5526 5933
rect 5492 5831 5526 5865
rect 5492 5763 5526 5797
rect 5492 5695 5526 5729
rect 5492 5627 5526 5661
rect 5588 6511 5622 6545
rect 5588 6443 5622 6477
rect 5588 6375 5622 6409
rect 5588 6307 5622 6341
rect 5588 6239 5622 6273
rect 5588 6171 5622 6205
rect 5588 6103 5622 6137
rect 5588 6035 5622 6069
rect 5588 5967 5622 6001
rect 5588 5899 5622 5933
rect 5588 5831 5622 5865
rect 5588 5763 5622 5797
rect 5588 5695 5622 5729
rect 5588 5627 5622 5661
rect 5684 6511 5718 6545
rect 5684 6443 5718 6477
rect 5684 6375 5718 6409
rect 5684 6307 5718 6341
rect 5684 6239 5718 6273
rect 5684 6171 5718 6205
rect 5684 6103 5718 6137
rect 5684 6035 5718 6069
rect 5684 5967 5718 6001
rect 5684 5899 5718 5933
rect 5684 5831 5718 5865
rect 5684 5763 5718 5797
rect 5684 5695 5718 5729
rect 5684 5627 5718 5661
rect 6180 6515 6214 6549
rect 6180 6447 6214 6481
rect 6180 6379 6214 6413
rect 6180 6311 6214 6345
rect 6180 6243 6214 6277
rect 6180 6175 6214 6209
rect 6180 6107 6214 6141
rect 6180 6039 6214 6073
rect 6180 5971 6214 6005
rect 6180 5903 6214 5937
rect 6180 5835 6214 5869
rect 6180 5767 6214 5801
rect 6180 5699 6214 5733
rect 6180 5631 6214 5665
rect 6276 6515 6310 6549
rect 6276 6447 6310 6481
rect 6276 6379 6310 6413
rect 6276 6311 6310 6345
rect 6276 6243 6310 6277
rect 6276 6175 6310 6209
rect 6276 6107 6310 6141
rect 6276 6039 6310 6073
rect 6276 5971 6310 6005
rect 6276 5903 6310 5937
rect 6276 5835 6310 5869
rect 6276 5767 6310 5801
rect 6276 5699 6310 5733
rect 6276 5631 6310 5665
rect 6372 6515 6406 6549
rect 6372 6447 6406 6481
rect 6372 6379 6406 6413
rect 6372 6311 6406 6345
rect 6372 6243 6406 6277
rect 6372 6175 6406 6209
rect 6372 6107 6406 6141
rect 6372 6039 6406 6073
rect 6372 5971 6406 6005
rect 6372 5903 6406 5937
rect 6372 5835 6406 5869
rect 6372 5767 6406 5801
rect 6372 5699 6406 5733
rect 6372 5631 6406 5665
rect 6468 6515 6502 6549
rect 6468 6447 6502 6481
rect 6468 6379 6502 6413
rect 6468 6311 6502 6345
rect 6468 6243 6502 6277
rect 6468 6175 6502 6209
rect 6468 6107 6502 6141
rect 6468 6039 6502 6073
rect 6468 5971 6502 6005
rect 6468 5903 6502 5937
rect 6468 5835 6502 5869
rect 6468 5767 6502 5801
rect 6468 5699 6502 5733
rect 6468 5631 6502 5665
rect 6564 6515 6598 6549
rect 6564 6447 6598 6481
rect 6564 6379 6598 6413
rect 6564 6311 6598 6345
rect 6564 6243 6598 6277
rect 6564 6175 6598 6209
rect 6564 6107 6598 6141
rect 6564 6039 6598 6073
rect 6564 5971 6598 6005
rect 6564 5903 6598 5937
rect 6564 5835 6598 5869
rect 6564 5767 6598 5801
rect 6564 5699 6598 5733
rect 6564 5631 6598 5665
rect 6660 6515 6694 6549
rect 6660 6447 6694 6481
rect 6660 6379 6694 6413
rect 6660 6311 6694 6345
rect 6660 6243 6694 6277
rect 6660 6175 6694 6209
rect 6660 6107 6694 6141
rect 6660 6039 6694 6073
rect 6660 5971 6694 6005
rect 6660 5903 6694 5937
rect 6660 5835 6694 5869
rect 6660 5767 6694 5801
rect 6660 5699 6694 5733
rect 6660 5631 6694 5665
rect 6756 6515 6790 6549
rect 6756 6447 6790 6481
rect 6756 6379 6790 6413
rect 6756 6311 6790 6345
rect 6756 6243 6790 6277
rect 6756 6175 6790 6209
rect 6756 6107 6790 6141
rect 6756 6039 6790 6073
rect 6756 5971 6790 6005
rect 6756 5903 6790 5937
rect 6756 5835 6790 5869
rect 6756 5767 6790 5801
rect 6756 5699 6790 5733
rect 6756 5631 6790 5665
rect 6852 6515 6886 6549
rect 6852 6447 6886 6481
rect 6852 6379 6886 6413
rect 6852 6311 6886 6345
rect 6852 6243 6886 6277
rect 6852 6175 6886 6209
rect 6852 6107 6886 6141
rect 6852 6039 6886 6073
rect 6852 5971 6886 6005
rect 6852 5903 6886 5937
rect 6852 5835 6886 5869
rect 6852 5767 6886 5801
rect 6852 5699 6886 5733
rect 6852 5631 6886 5665
rect 6948 6515 6982 6549
rect 6948 6447 6982 6481
rect 6948 6379 6982 6413
rect 6948 6311 6982 6345
rect 6948 6243 6982 6277
rect 6948 6175 6982 6209
rect 6948 6107 6982 6141
rect 6948 6039 6982 6073
rect 6948 5971 6982 6005
rect 6948 5903 6982 5937
rect 6948 5835 6982 5869
rect 6948 5767 6982 5801
rect 6948 5699 6982 5733
rect 6948 5631 6982 5665
rect 7044 6515 7078 6549
rect 7044 6447 7078 6481
rect 7044 6379 7078 6413
rect 7044 6311 7078 6345
rect 7044 6243 7078 6277
rect 7044 6175 7078 6209
rect 7044 6107 7078 6141
rect 7044 6039 7078 6073
rect 7044 5971 7078 6005
rect 7044 5903 7078 5937
rect 7044 5835 7078 5869
rect 7044 5767 7078 5801
rect 7044 5699 7078 5733
rect 7044 5631 7078 5665
rect 7140 6515 7174 6549
rect 7140 6447 7174 6481
rect 7140 6379 7174 6413
rect 7140 6311 7174 6345
rect 7140 6243 7174 6277
rect 7140 6175 7174 6209
rect 7140 6107 7174 6141
rect 7140 6039 7174 6073
rect 7140 5971 7174 6005
rect 7140 5903 7174 5937
rect 7140 5835 7174 5869
rect 7140 5767 7174 5801
rect 7140 5699 7174 5733
rect 7140 5631 7174 5665
rect 7236 6515 7270 6549
rect 7236 6447 7270 6481
rect 7236 6379 7270 6413
rect 7236 6311 7270 6345
rect 7236 6243 7270 6277
rect 7236 6175 7270 6209
rect 7236 6107 7270 6141
rect 7236 6039 7270 6073
rect 7236 5971 7270 6005
rect 7236 5903 7270 5937
rect 7236 5835 7270 5869
rect 7236 5767 7270 5801
rect 7236 5699 7270 5733
rect 7236 5631 7270 5665
rect 7332 6515 7366 6549
rect 7332 6447 7366 6481
rect 7332 6379 7366 6413
rect 7332 6311 7366 6345
rect 7332 6243 7366 6277
rect 7332 6175 7366 6209
rect 7332 6107 7366 6141
rect 7332 6039 7366 6073
rect 7332 5971 7366 6005
rect 7332 5903 7366 5937
rect 7332 5835 7366 5869
rect 7332 5767 7366 5801
rect 7332 5699 7366 5733
rect 7332 5631 7366 5665
rect 7946 6511 7980 6545
rect 7946 6443 7980 6477
rect 7946 6375 7980 6409
rect 7946 6307 7980 6341
rect 7946 6239 7980 6273
rect 7946 6171 7980 6205
rect 7946 6103 7980 6137
rect 7946 6035 7980 6069
rect 7946 5967 7980 6001
rect 7946 5899 7980 5933
rect 7946 5831 7980 5865
rect 7946 5763 7980 5797
rect 7946 5695 7980 5729
rect 7946 5627 7980 5661
rect 8042 6511 8076 6545
rect 8042 6443 8076 6477
rect 8042 6375 8076 6409
rect 8042 6307 8076 6341
rect 8042 6239 8076 6273
rect 8042 6171 8076 6205
rect 8042 6103 8076 6137
rect 8042 6035 8076 6069
rect 8042 5967 8076 6001
rect 8042 5899 8076 5933
rect 8042 5831 8076 5865
rect 8042 5763 8076 5797
rect 8042 5695 8076 5729
rect 8042 5627 8076 5661
rect 8138 6511 8172 6545
rect 8138 6443 8172 6477
rect 8138 6375 8172 6409
rect 8138 6307 8172 6341
rect 8138 6239 8172 6273
rect 8138 6171 8172 6205
rect 8138 6103 8172 6137
rect 8138 6035 8172 6069
rect 8138 5967 8172 6001
rect 8138 5899 8172 5933
rect 8138 5831 8172 5865
rect 8138 5763 8172 5797
rect 8138 5695 8172 5729
rect 8138 5627 8172 5661
rect 8234 6511 8268 6545
rect 8234 6443 8268 6477
rect 8234 6375 8268 6409
rect 8234 6307 8268 6341
rect 8234 6239 8268 6273
rect 8234 6171 8268 6205
rect 8234 6103 8268 6137
rect 8234 6035 8268 6069
rect 8234 5967 8268 6001
rect 8234 5899 8268 5933
rect 8234 5831 8268 5865
rect 8234 5763 8268 5797
rect 8234 5695 8268 5729
rect 8234 5627 8268 5661
rect 8330 6511 8364 6545
rect 8330 6443 8364 6477
rect 8330 6375 8364 6409
rect 8330 6307 8364 6341
rect 8330 6239 8364 6273
rect 8330 6171 8364 6205
rect 8330 6103 8364 6137
rect 8330 6035 8364 6069
rect 8330 5967 8364 6001
rect 8330 5899 8364 5933
rect 8330 5831 8364 5865
rect 8330 5763 8364 5797
rect 8330 5695 8364 5729
rect 8330 5627 8364 5661
rect 8426 6511 8460 6545
rect 8426 6443 8460 6477
rect 8426 6375 8460 6409
rect 8426 6307 8460 6341
rect 8426 6239 8460 6273
rect 8426 6171 8460 6205
rect 8426 6103 8460 6137
rect 8426 6035 8460 6069
rect 8426 5967 8460 6001
rect 8426 5899 8460 5933
rect 8426 5831 8460 5865
rect 8426 5763 8460 5797
rect 8426 5695 8460 5729
rect 8426 5627 8460 5661
rect 8522 6511 8556 6545
rect 8522 6443 8556 6477
rect 8522 6375 8556 6409
rect 8522 6307 8556 6341
rect 8522 6239 8556 6273
rect 8522 6171 8556 6205
rect 8522 6103 8556 6137
rect 8522 6035 8556 6069
rect 8522 5967 8556 6001
rect 8522 5899 8556 5933
rect 8522 5831 8556 5865
rect 8522 5763 8556 5797
rect 8522 5695 8556 5729
rect 8522 5627 8556 5661
rect 8618 6511 8652 6545
rect 8618 6443 8652 6477
rect 8618 6375 8652 6409
rect 8618 6307 8652 6341
rect 8618 6239 8652 6273
rect 8618 6171 8652 6205
rect 8618 6103 8652 6137
rect 8618 6035 8652 6069
rect 8618 5967 8652 6001
rect 8618 5899 8652 5933
rect 8618 5831 8652 5865
rect 8618 5763 8652 5797
rect 8618 5695 8652 5729
rect 8618 5627 8652 5661
rect 8714 6511 8748 6545
rect 8714 6443 8748 6477
rect 8714 6375 8748 6409
rect 8714 6307 8748 6341
rect 8714 6239 8748 6273
rect 8714 6171 8748 6205
rect 8714 6103 8748 6137
rect 8714 6035 8748 6069
rect 8714 5967 8748 6001
rect 8714 5899 8748 5933
rect 8714 5831 8748 5865
rect 8714 5763 8748 5797
rect 8714 5695 8748 5729
rect 8714 5627 8748 5661
rect 9268 6513 9302 6547
rect 9268 6445 9302 6479
rect 9268 6377 9302 6411
rect 9268 6309 9302 6343
rect 9268 6241 9302 6275
rect 9268 6173 9302 6207
rect 9268 6105 9302 6139
rect 9268 6037 9302 6071
rect 9268 5969 9302 6003
rect 9268 5901 9302 5935
rect 9268 5833 9302 5867
rect 9268 5765 9302 5799
rect 9268 5697 9302 5731
rect 9268 5629 9302 5663
rect 9364 6513 9398 6547
rect 9364 6445 9398 6479
rect 9364 6377 9398 6411
rect 9364 6309 9398 6343
rect 9364 6241 9398 6275
rect 9364 6173 9398 6207
rect 9364 6105 9398 6139
rect 9364 6037 9398 6071
rect 9364 5969 9398 6003
rect 9364 5901 9398 5935
rect 9364 5833 9398 5867
rect 9364 5765 9398 5799
rect 9364 5697 9398 5731
rect 9364 5629 9398 5663
rect 9460 6513 9494 6547
rect 9460 6445 9494 6479
rect 9460 6377 9494 6411
rect 9460 6309 9494 6343
rect 9460 6241 9494 6275
rect 9460 6173 9494 6207
rect 9460 6105 9494 6139
rect 9460 6037 9494 6071
rect 9460 5969 9494 6003
rect 9460 5901 9494 5935
rect 9460 5833 9494 5867
rect 9460 5765 9494 5799
rect 9460 5697 9494 5731
rect 9460 5629 9494 5663
rect 9556 6513 9590 6547
rect 9556 6445 9590 6479
rect 9556 6377 9590 6411
rect 9556 6309 9590 6343
rect 9556 6241 9590 6275
rect 9556 6173 9590 6207
rect 9556 6105 9590 6139
rect 9556 6037 9590 6071
rect 9556 5969 9590 6003
rect 9556 5901 9590 5935
rect 9556 5833 9590 5867
rect 9556 5765 9590 5799
rect 9556 5697 9590 5731
rect 9556 5629 9590 5663
rect 9652 6513 9686 6547
rect 9652 6445 9686 6479
rect 9652 6377 9686 6411
rect 9652 6309 9686 6343
rect 9652 6241 9686 6275
rect 9652 6173 9686 6207
rect 9652 6105 9686 6139
rect 9652 6037 9686 6071
rect 9652 5969 9686 6003
rect 9652 5901 9686 5935
rect 9652 5833 9686 5867
rect 9652 5765 9686 5799
rect 9652 5697 9686 5731
rect 9652 5629 9686 5663
rect 9748 6513 9782 6547
rect 9748 6445 9782 6479
rect 9748 6377 9782 6411
rect 9748 6309 9782 6343
rect 9748 6241 9782 6275
rect 9748 6173 9782 6207
rect 9748 6105 9782 6139
rect 9748 6037 9782 6071
rect 9748 5969 9782 6003
rect 9748 5901 9782 5935
rect 9748 5833 9782 5867
rect 9748 5765 9782 5799
rect 9748 5697 9782 5731
rect 9748 5629 9782 5663
rect 9844 6513 9878 6547
rect 9844 6445 9878 6479
rect 9844 6377 9878 6411
rect 9844 6309 9878 6343
rect 9844 6241 9878 6275
rect 9844 6173 9878 6207
rect 9844 6105 9878 6139
rect 9844 6037 9878 6071
rect 9844 5969 9878 6003
rect 9844 5901 9878 5935
rect 9844 5833 9878 5867
rect 9844 5765 9878 5799
rect 9844 5697 9878 5731
rect 9844 5629 9878 5663
rect 9940 6513 9974 6547
rect 9940 6445 9974 6479
rect 9940 6377 9974 6411
rect 9940 6309 9974 6343
rect 9940 6241 9974 6275
rect 9940 6173 9974 6207
rect 9940 6105 9974 6139
rect 9940 6037 9974 6071
rect 9940 5969 9974 6003
rect 9940 5901 9974 5935
rect 9940 5833 9974 5867
rect 9940 5765 9974 5799
rect 9940 5697 9974 5731
rect 9940 5629 9974 5663
rect 10036 6513 10070 6547
rect 10036 6445 10070 6479
rect 10036 6377 10070 6411
rect 10036 6309 10070 6343
rect 10036 6241 10070 6275
rect 10036 6173 10070 6207
rect 10036 6105 10070 6139
rect 10036 6037 10070 6071
rect 10036 5969 10070 6003
rect 10036 5901 10070 5935
rect 10036 5833 10070 5867
rect 10036 5765 10070 5799
rect 10036 5697 10070 5731
rect 10036 5629 10070 5663
rect 10132 6513 10166 6547
rect 10132 6445 10166 6479
rect 10132 6377 10166 6411
rect 10132 6309 10166 6343
rect 10132 6241 10166 6275
rect 10132 6173 10166 6207
rect 10132 6105 10166 6139
rect 10132 6037 10166 6071
rect 10132 5969 10166 6003
rect 10132 5901 10166 5935
rect 10132 5833 10166 5867
rect 10132 5765 10166 5799
rect 10132 5697 10166 5731
rect 10132 5629 10166 5663
rect 10228 6513 10262 6547
rect 10228 6445 10262 6479
rect 10228 6377 10262 6411
rect 10228 6309 10262 6343
rect 10228 6241 10262 6275
rect 10228 6173 10262 6207
rect 10228 6105 10262 6139
rect 10228 6037 10262 6071
rect 10228 5969 10262 6003
rect 10228 5901 10262 5935
rect 10228 5833 10262 5867
rect 10228 5765 10262 5799
rect 10228 5697 10262 5731
rect 10228 5629 10262 5663
rect 10324 6513 10358 6547
rect 10324 6445 10358 6479
rect 10324 6377 10358 6411
rect 10324 6309 10358 6343
rect 10324 6241 10358 6275
rect 10324 6173 10358 6207
rect 10324 6105 10358 6139
rect 10324 6037 10358 6071
rect 10324 5969 10358 6003
rect 10324 5901 10358 5935
rect 10324 5833 10358 5867
rect 10324 5765 10358 5799
rect 10324 5697 10358 5731
rect 10324 5629 10358 5663
rect 10420 6513 10454 6547
rect 10420 6445 10454 6479
rect 10420 6377 10454 6411
rect 10420 6309 10454 6343
rect 10420 6241 10454 6275
rect 10420 6173 10454 6207
rect 10420 6105 10454 6139
rect 10420 6037 10454 6071
rect 10420 5969 10454 6003
rect 10420 5901 10454 5935
rect 10420 5833 10454 5867
rect 10420 5765 10454 5799
rect 10420 5697 10454 5731
rect 10420 5629 10454 5663
rect 11034 6509 11068 6543
rect 11034 6441 11068 6475
rect 11034 6373 11068 6407
rect 11034 6305 11068 6339
rect 11034 6237 11068 6271
rect 11034 6169 11068 6203
rect 11034 6101 11068 6135
rect 11034 6033 11068 6067
rect 11034 5965 11068 5999
rect 11034 5897 11068 5931
rect 11034 5829 11068 5863
rect 11034 5761 11068 5795
rect 11034 5693 11068 5727
rect 11034 5625 11068 5659
rect 11130 6509 11164 6543
rect 11130 6441 11164 6475
rect 11130 6373 11164 6407
rect 11130 6305 11164 6339
rect 11130 6237 11164 6271
rect 11130 6169 11164 6203
rect 11130 6101 11164 6135
rect 11130 6033 11164 6067
rect 11130 5965 11164 5999
rect 11130 5897 11164 5931
rect 11130 5829 11164 5863
rect 11130 5761 11164 5795
rect 11130 5693 11164 5727
rect 11130 5625 11164 5659
rect 11226 6509 11260 6543
rect 11226 6441 11260 6475
rect 11226 6373 11260 6407
rect 11226 6305 11260 6339
rect 11226 6237 11260 6271
rect 11226 6169 11260 6203
rect 11226 6101 11260 6135
rect 11226 6033 11260 6067
rect 11226 5965 11260 5999
rect 11226 5897 11260 5931
rect 11226 5829 11260 5863
rect 11226 5761 11260 5795
rect 11226 5693 11260 5727
rect 11226 5625 11260 5659
rect 11322 6509 11356 6543
rect 11322 6441 11356 6475
rect 11322 6373 11356 6407
rect 11322 6305 11356 6339
rect 11322 6237 11356 6271
rect 11322 6169 11356 6203
rect 11322 6101 11356 6135
rect 11322 6033 11356 6067
rect 11322 5965 11356 5999
rect 11322 5897 11356 5931
rect 11322 5829 11356 5863
rect 11322 5761 11356 5795
rect 11322 5693 11356 5727
rect 11322 5625 11356 5659
rect 11418 6509 11452 6543
rect 11418 6441 11452 6475
rect 11418 6373 11452 6407
rect 11418 6305 11452 6339
rect 11418 6237 11452 6271
rect 11418 6169 11452 6203
rect 11418 6101 11452 6135
rect 11418 6033 11452 6067
rect 11418 5965 11452 5999
rect 11418 5897 11452 5931
rect 11418 5829 11452 5863
rect 11418 5761 11452 5795
rect 11418 5693 11452 5727
rect 11418 5625 11452 5659
rect 11514 6509 11548 6543
rect 11514 6441 11548 6475
rect 11514 6373 11548 6407
rect 11514 6305 11548 6339
rect 11514 6237 11548 6271
rect 11514 6169 11548 6203
rect 11514 6101 11548 6135
rect 11514 6033 11548 6067
rect 11514 5965 11548 5999
rect 11514 5897 11548 5931
rect 11514 5829 11548 5863
rect 11514 5761 11548 5795
rect 11514 5693 11548 5727
rect 11514 5625 11548 5659
rect 11610 6509 11644 6543
rect 11610 6441 11644 6475
rect 11610 6373 11644 6407
rect 11610 6305 11644 6339
rect 11610 6237 11644 6271
rect 11610 6169 11644 6203
rect 11610 6101 11644 6135
rect 11610 6033 11644 6067
rect 11610 5965 11644 5999
rect 11610 5897 11644 5931
rect 11610 5829 11644 5863
rect 11610 5761 11644 5795
rect 11610 5693 11644 5727
rect 11610 5625 11644 5659
rect 11706 6509 11740 6543
rect 11706 6441 11740 6475
rect 11706 6373 11740 6407
rect 11706 6305 11740 6339
rect 11706 6237 11740 6271
rect 11706 6169 11740 6203
rect 11706 6101 11740 6135
rect 11706 6033 11740 6067
rect 11706 5965 11740 5999
rect 11706 5897 11740 5931
rect 11706 5829 11740 5863
rect 11706 5761 11740 5795
rect 11706 5693 11740 5727
rect 11706 5625 11740 5659
rect 11802 6509 11836 6543
rect 11802 6441 11836 6475
rect 11802 6373 11836 6407
rect 11802 6305 11836 6339
rect 11802 6237 11836 6271
rect 11802 6169 11836 6203
rect 11802 6101 11836 6135
rect 11802 6033 11836 6067
rect 11802 5965 11836 5999
rect 11802 5897 11836 5931
rect 11802 5829 11836 5863
rect 11802 5761 11836 5795
rect 11802 5693 11836 5727
rect 11802 5625 11836 5659
rect 12424 6487 12458 6521
rect 12424 6419 12458 6453
rect 12424 6351 12458 6385
rect 12424 6283 12458 6317
rect 12424 6215 12458 6249
rect 12424 6147 12458 6181
rect 12424 6079 12458 6113
rect 12424 6011 12458 6045
rect 12424 5943 12458 5977
rect 12424 5875 12458 5909
rect 12424 5807 12458 5841
rect 12424 5739 12458 5773
rect 12424 5671 12458 5705
rect 12424 5603 12458 5637
rect 12520 6487 12554 6521
rect 12520 6419 12554 6453
rect 12520 6351 12554 6385
rect 12520 6283 12554 6317
rect 12520 6215 12554 6249
rect 12520 6147 12554 6181
rect 12520 6079 12554 6113
rect 12520 6011 12554 6045
rect 12520 5943 12554 5977
rect 12520 5875 12554 5909
rect 12520 5807 12554 5841
rect 12520 5739 12554 5773
rect 12520 5671 12554 5705
rect 12520 5603 12554 5637
rect 12616 6487 12650 6521
rect 12616 6419 12650 6453
rect 12616 6351 12650 6385
rect 12616 6283 12650 6317
rect 12616 6215 12650 6249
rect 12616 6147 12650 6181
rect 12616 6079 12650 6113
rect 12616 6011 12650 6045
rect 12616 5943 12650 5977
rect 12616 5875 12650 5909
rect 12616 5807 12650 5841
rect 12616 5739 12650 5773
rect 12616 5671 12650 5705
rect 12616 5603 12650 5637
rect 12712 6487 12746 6521
rect 12712 6419 12746 6453
rect 12712 6351 12746 6385
rect 12712 6283 12746 6317
rect 12712 6215 12746 6249
rect 12712 6147 12746 6181
rect 12712 6079 12746 6113
rect 12712 6011 12746 6045
rect 12712 5943 12746 5977
rect 12712 5875 12746 5909
rect 12712 5807 12746 5841
rect 12712 5739 12746 5773
rect 12712 5671 12746 5705
rect 12712 5603 12746 5637
rect 12808 6487 12842 6521
rect 12808 6419 12842 6453
rect 12808 6351 12842 6385
rect 12808 6283 12842 6317
rect 12808 6215 12842 6249
rect 12808 6147 12842 6181
rect 12808 6079 12842 6113
rect 12808 6011 12842 6045
rect 12808 5943 12842 5977
rect 12808 5875 12842 5909
rect 12808 5807 12842 5841
rect 12808 5739 12842 5773
rect 12808 5671 12842 5705
rect 12808 5603 12842 5637
rect 12904 6487 12938 6521
rect 12904 6419 12938 6453
rect 12904 6351 12938 6385
rect 12904 6283 12938 6317
rect 12904 6215 12938 6249
rect 12904 6147 12938 6181
rect 12904 6079 12938 6113
rect 12904 6011 12938 6045
rect 12904 5943 12938 5977
rect 12904 5875 12938 5909
rect 12904 5807 12938 5841
rect 12904 5739 12938 5773
rect 12904 5671 12938 5705
rect 12904 5603 12938 5637
rect 13000 6487 13034 6521
rect 13000 6419 13034 6453
rect 13000 6351 13034 6385
rect 13000 6283 13034 6317
rect 13000 6215 13034 6249
rect 13000 6147 13034 6181
rect 13000 6079 13034 6113
rect 13000 6011 13034 6045
rect 13000 5943 13034 5977
rect 13000 5875 13034 5909
rect 13000 5807 13034 5841
rect 13000 5739 13034 5773
rect 13000 5671 13034 5705
rect 13000 5603 13034 5637
rect 13096 6487 13130 6521
rect 13096 6419 13130 6453
rect 13096 6351 13130 6385
rect 13096 6283 13130 6317
rect 13096 6215 13130 6249
rect 13096 6147 13130 6181
rect 13096 6079 13130 6113
rect 13096 6011 13130 6045
rect 13096 5943 13130 5977
rect 13096 5875 13130 5909
rect 13096 5807 13130 5841
rect 13096 5739 13130 5773
rect 13096 5671 13130 5705
rect 13096 5603 13130 5637
rect 13192 6487 13226 6521
rect 13192 6419 13226 6453
rect 13192 6351 13226 6385
rect 13192 6283 13226 6317
rect 13192 6215 13226 6249
rect 13192 6147 13226 6181
rect 13192 6079 13226 6113
rect 13192 6011 13226 6045
rect 13192 5943 13226 5977
rect 13192 5875 13226 5909
rect 13192 5807 13226 5841
rect 13192 5739 13226 5773
rect 13192 5671 13226 5705
rect 13192 5603 13226 5637
rect 13288 6487 13322 6521
rect 13288 6419 13322 6453
rect 13288 6351 13322 6385
rect 13288 6283 13322 6317
rect 13288 6215 13322 6249
rect 13288 6147 13322 6181
rect 13288 6079 13322 6113
rect 13288 6011 13322 6045
rect 13288 5943 13322 5977
rect 13288 5875 13322 5909
rect 13288 5807 13322 5841
rect 13288 5739 13322 5773
rect 13288 5671 13322 5705
rect 13288 5603 13322 5637
rect 13384 6487 13418 6521
rect 13384 6419 13418 6453
rect 13384 6351 13418 6385
rect 13384 6283 13418 6317
rect 13384 6215 13418 6249
rect 13384 6147 13418 6181
rect 13384 6079 13418 6113
rect 13384 6011 13418 6045
rect 13384 5943 13418 5977
rect 13384 5875 13418 5909
rect 13384 5807 13418 5841
rect 13384 5739 13418 5773
rect 13384 5671 13418 5705
rect 13384 5603 13418 5637
rect 13480 6487 13514 6521
rect 13480 6419 13514 6453
rect 13480 6351 13514 6385
rect 13480 6283 13514 6317
rect 13480 6215 13514 6249
rect 13480 6147 13514 6181
rect 13480 6079 13514 6113
rect 13480 6011 13514 6045
rect 13480 5943 13514 5977
rect 13480 5875 13514 5909
rect 13480 5807 13514 5841
rect 13480 5739 13514 5773
rect 13480 5671 13514 5705
rect 13480 5603 13514 5637
rect 13576 6487 13610 6521
rect 13576 6419 13610 6453
rect 13576 6351 13610 6385
rect 13576 6283 13610 6317
rect 13576 6215 13610 6249
rect 13576 6147 13610 6181
rect 13576 6079 13610 6113
rect 13576 6011 13610 6045
rect 13576 5943 13610 5977
rect 13576 5875 13610 5909
rect 13576 5807 13610 5841
rect 13576 5739 13610 5773
rect 13576 5671 13610 5705
rect 13576 5603 13610 5637
rect 14190 6483 14224 6517
rect 14190 6415 14224 6449
rect 14190 6347 14224 6381
rect 14190 6279 14224 6313
rect 14190 6211 14224 6245
rect 14190 6143 14224 6177
rect 14190 6075 14224 6109
rect 14190 6007 14224 6041
rect 14190 5939 14224 5973
rect 14190 5871 14224 5905
rect 14190 5803 14224 5837
rect 14190 5735 14224 5769
rect 14190 5667 14224 5701
rect 14190 5599 14224 5633
rect -868 5521 -834 5555
rect 14286 6483 14320 6517
rect 14286 6415 14320 6449
rect 14286 6347 14320 6381
rect 14286 6279 14320 6313
rect 14286 6211 14320 6245
rect 14286 6143 14320 6177
rect 14286 6075 14320 6109
rect 14286 6007 14320 6041
rect 14286 5939 14320 5973
rect 14286 5871 14320 5905
rect 14286 5803 14320 5837
rect 14286 5735 14320 5769
rect 14286 5667 14320 5701
rect 14286 5599 14320 5633
rect 14382 6483 14416 6517
rect 14382 6415 14416 6449
rect 14382 6347 14416 6381
rect 14382 6279 14416 6313
rect 14382 6211 14416 6245
rect 14382 6143 14416 6177
rect 14382 6075 14416 6109
rect 14382 6007 14416 6041
rect 14382 5939 14416 5973
rect 14382 5871 14416 5905
rect 14382 5803 14416 5837
rect 14382 5735 14416 5769
rect 14382 5667 14416 5701
rect 14382 5599 14416 5633
rect 14478 6483 14512 6517
rect 14478 6415 14512 6449
rect 14478 6347 14512 6381
rect 14478 6279 14512 6313
rect 14478 6211 14512 6245
rect 14478 6143 14512 6177
rect 14478 6075 14512 6109
rect 14478 6007 14512 6041
rect 14478 5939 14512 5973
rect 14478 5871 14512 5905
rect 14478 5803 14512 5837
rect 14478 5735 14512 5769
rect 14478 5667 14512 5701
rect 14478 5599 14512 5633
rect 14574 6483 14608 6517
rect 14574 6415 14608 6449
rect 14574 6347 14608 6381
rect 14574 6279 14608 6313
rect 14574 6211 14608 6245
rect 14574 6143 14608 6177
rect 14574 6075 14608 6109
rect 14574 6007 14608 6041
rect 14574 5939 14608 5973
rect 14574 5871 14608 5905
rect 14574 5803 14608 5837
rect 14574 5735 14608 5769
rect 14574 5667 14608 5701
rect 14574 5599 14608 5633
rect 14670 6483 14704 6517
rect 14670 6415 14704 6449
rect 14670 6347 14704 6381
rect 14670 6279 14704 6313
rect 14670 6211 14704 6245
rect 14670 6143 14704 6177
rect 14670 6075 14704 6109
rect 14670 6007 14704 6041
rect 14670 5939 14704 5973
rect 14670 5871 14704 5905
rect 14670 5803 14704 5837
rect 14670 5735 14704 5769
rect 14670 5667 14704 5701
rect 14670 5599 14704 5633
rect 14766 6483 14800 6517
rect 14766 6415 14800 6449
rect 14766 6347 14800 6381
rect 14766 6279 14800 6313
rect 14766 6211 14800 6245
rect 14766 6143 14800 6177
rect 14766 6075 14800 6109
rect 14766 6007 14800 6041
rect 14766 5939 14800 5973
rect 14766 5871 14800 5905
rect 14766 5803 14800 5837
rect 14766 5735 14800 5769
rect 14766 5667 14800 5701
rect 14766 5599 14800 5633
rect 14862 6483 14896 6517
rect 14862 6415 14896 6449
rect 14862 6347 14896 6381
rect 14862 6279 14896 6313
rect 14862 6211 14896 6245
rect 14862 6143 14896 6177
rect 14862 6075 14896 6109
rect 14862 6007 14896 6041
rect 14862 5939 14896 5973
rect 14862 5871 14896 5905
rect 14862 5803 14896 5837
rect 14862 5735 14896 5769
rect 14862 5667 14896 5701
rect 14862 5599 14896 5633
rect 14958 6483 14992 6517
rect 14958 6415 14992 6449
rect 14958 6347 14992 6381
rect 14958 6279 14992 6313
rect 14958 6211 14992 6245
rect 14958 6143 14992 6177
rect 14958 6075 14992 6109
rect 14958 6007 14992 6041
rect 14958 5939 14992 5973
rect 14958 5871 14992 5905
rect 14958 5803 14992 5837
rect 14958 5735 14992 5769
rect 14958 5667 14992 5701
rect 14958 5599 14992 5633
rect 15518 5861 15552 5895
rect 15518 5793 15552 5827
rect 15518 5725 15552 5759
rect 15518 5657 15552 5691
rect 15518 5589 15552 5623
rect -868 5453 -834 5487
rect -868 5385 -834 5419
rect -868 5317 -834 5351
rect -868 5249 -834 5283
rect -868 5181 -834 5215
rect -868 5113 -834 5147
rect -868 5045 -834 5079
rect 15518 5521 15552 5555
rect 15518 5453 15552 5487
rect 15518 5385 15552 5419
rect 15518 5317 15552 5351
rect 15518 5249 15552 5283
rect 15518 5181 15552 5215
rect 15518 5113 15552 5147
rect 15518 5045 15552 5079
rect -868 4977 -834 5011
rect 1484 4869 1518 4903
rect 1484 4801 1518 4835
rect 1484 4733 1518 4767
rect 1484 4665 1518 4699
rect 1484 4597 1518 4631
rect 1484 4529 1518 4563
rect 1484 4461 1518 4495
rect 1484 4393 1518 4427
rect 1484 4325 1518 4359
rect 1484 4257 1518 4291
rect 1484 4189 1518 4223
rect 1484 4121 1518 4155
rect 1484 4053 1518 4087
rect 1484 3985 1518 4019
rect 1580 4869 1614 4903
rect 1580 4801 1614 4835
rect 1580 4733 1614 4767
rect 1580 4665 1614 4699
rect 1580 4597 1614 4631
rect 1580 4529 1614 4563
rect 1580 4461 1614 4495
rect 1580 4393 1614 4427
rect 1580 4325 1614 4359
rect 1580 4257 1614 4291
rect 1580 4189 1614 4223
rect 1580 4121 1614 4155
rect 1580 4053 1614 4087
rect 1580 3985 1614 4019
rect 1676 4869 1710 4903
rect 1676 4801 1710 4835
rect 1676 4733 1710 4767
rect 1676 4665 1710 4699
rect 1676 4597 1710 4631
rect 1676 4529 1710 4563
rect 1676 4461 1710 4495
rect 1676 4393 1710 4427
rect 1676 4325 1710 4359
rect 1676 4257 1710 4291
rect 1676 4189 1710 4223
rect 1676 4121 1710 4155
rect 1676 4053 1710 4087
rect 1676 3985 1710 4019
rect 1772 4869 1806 4903
rect 1772 4801 1806 4835
rect 1772 4733 1806 4767
rect 1772 4665 1806 4699
rect 1772 4597 1806 4631
rect 1772 4529 1806 4563
rect 1772 4461 1806 4495
rect 1772 4393 1806 4427
rect 1772 4325 1806 4359
rect 1772 4257 1806 4291
rect 1772 4189 1806 4223
rect 1772 4121 1806 4155
rect 1772 4053 1806 4087
rect 1772 3985 1806 4019
rect 15518 4977 15552 5011
rect 1868 4869 1902 4903
rect 1868 4801 1902 4835
rect 1868 4733 1902 4767
rect 1868 4665 1902 4699
rect 1868 4597 1902 4631
rect 1868 4529 1902 4563
rect 1868 4461 1902 4495
rect 1868 4393 1902 4427
rect 1868 4325 1902 4359
rect 1868 4257 1902 4291
rect 1868 4189 1902 4223
rect 1868 4121 1902 4155
rect 1868 4053 1902 4087
rect 1868 3985 1902 4019
rect 4440 4853 4474 4887
rect 4440 4785 4474 4819
rect 4440 4717 4474 4751
rect 4440 4649 4474 4683
rect 4440 4581 4474 4615
rect 4440 4513 4474 4547
rect 4440 4445 4474 4479
rect 4440 4377 4474 4411
rect 4440 4309 4474 4343
rect 4440 4241 4474 4275
rect 4440 4173 4474 4207
rect 4440 4105 4474 4139
rect 4440 4037 4474 4071
rect 4440 3969 4474 4003
rect 4536 4853 4570 4887
rect 4536 4785 4570 4819
rect 4536 4717 4570 4751
rect 4536 4649 4570 4683
rect 4536 4581 4570 4615
rect 4536 4513 4570 4547
rect 4536 4445 4570 4479
rect 4536 4377 4570 4411
rect 4536 4309 4570 4343
rect 4536 4241 4570 4275
rect 4536 4173 4570 4207
rect 4536 4105 4570 4139
rect 4536 4037 4570 4071
rect 4536 3969 4570 4003
rect 4632 4853 4666 4887
rect 4632 4785 4666 4819
rect 4632 4717 4666 4751
rect 4632 4649 4666 4683
rect 4632 4581 4666 4615
rect 4632 4513 4666 4547
rect 4632 4445 4666 4479
rect 4632 4377 4666 4411
rect 4632 4309 4666 4343
rect 4632 4241 4666 4275
rect 4632 4173 4666 4207
rect 4632 4105 4666 4139
rect 4632 4037 4666 4071
rect 4632 3969 4666 4003
rect 4728 4853 4762 4887
rect 4728 4785 4762 4819
rect 4728 4717 4762 4751
rect 4728 4649 4762 4683
rect 4728 4581 4762 4615
rect 4728 4513 4762 4547
rect 4728 4445 4762 4479
rect 4728 4377 4762 4411
rect 4728 4309 4762 4343
rect 4728 4241 4762 4275
rect 4728 4173 4762 4207
rect 4728 4105 4762 4139
rect 4728 4037 4762 4071
rect 4728 3969 4762 4003
rect 4824 4853 4858 4887
rect 4824 4785 4858 4819
rect 4824 4717 4858 4751
rect 4824 4649 4858 4683
rect 4824 4581 4858 4615
rect 4824 4513 4858 4547
rect 4824 4445 4858 4479
rect 4824 4377 4858 4411
rect 4824 4309 4858 4343
rect 4824 4241 4858 4275
rect 4824 4173 4858 4207
rect 4824 4105 4858 4139
rect 4824 4037 4858 4071
rect 4824 3969 4858 4003
rect 7470 4853 7504 4887
rect 7470 4785 7504 4819
rect 7470 4717 7504 4751
rect 7470 4649 7504 4683
rect 7470 4581 7504 4615
rect 7470 4513 7504 4547
rect 7470 4445 7504 4479
rect 7470 4377 7504 4411
rect 7470 4309 7504 4343
rect 7470 4241 7504 4275
rect 7470 4173 7504 4207
rect 7470 4105 7504 4139
rect 7470 4037 7504 4071
rect 7470 3969 7504 4003
rect 7566 4853 7600 4887
rect 7566 4785 7600 4819
rect 7566 4717 7600 4751
rect 7566 4649 7600 4683
rect 7566 4581 7600 4615
rect 7566 4513 7600 4547
rect 7566 4445 7600 4479
rect 7566 4377 7600 4411
rect 7566 4309 7600 4343
rect 7566 4241 7600 4275
rect 7566 4173 7600 4207
rect 7566 4105 7600 4139
rect 7566 4037 7600 4071
rect 7566 3969 7600 4003
rect 7662 4853 7696 4887
rect 7662 4785 7696 4819
rect 7662 4717 7696 4751
rect 7662 4649 7696 4683
rect 7662 4581 7696 4615
rect 7662 4513 7696 4547
rect 7662 4445 7696 4479
rect 7662 4377 7696 4411
rect 7662 4309 7696 4343
rect 7662 4241 7696 4275
rect 7662 4173 7696 4207
rect 7662 4105 7696 4139
rect 7662 4037 7696 4071
rect 7662 3969 7696 4003
rect 7758 4853 7792 4887
rect 7758 4785 7792 4819
rect 7758 4717 7792 4751
rect 7758 4649 7792 4683
rect 7758 4581 7792 4615
rect 7758 4513 7792 4547
rect 7758 4445 7792 4479
rect 7758 4377 7792 4411
rect 7758 4309 7792 4343
rect 7758 4241 7792 4275
rect 7758 4173 7792 4207
rect 7758 4105 7792 4139
rect 7758 4037 7792 4071
rect 7758 3969 7792 4003
rect 7854 4853 7888 4887
rect 7854 4785 7888 4819
rect 7854 4717 7888 4751
rect 7854 4649 7888 4683
rect 7854 4581 7888 4615
rect 7854 4513 7888 4547
rect 7854 4445 7888 4479
rect 7854 4377 7888 4411
rect 7854 4309 7888 4343
rect 7854 4241 7888 4275
rect 7854 4173 7888 4207
rect 7854 4105 7888 4139
rect 7854 4037 7888 4071
rect 7854 3969 7888 4003
rect 10558 4851 10592 4885
rect 10558 4783 10592 4817
rect 10558 4715 10592 4749
rect 10558 4647 10592 4681
rect 10558 4579 10592 4613
rect 10558 4511 10592 4545
rect 10558 4443 10592 4477
rect 10558 4375 10592 4409
rect 10558 4307 10592 4341
rect 10558 4239 10592 4273
rect 10558 4171 10592 4205
rect 10558 4103 10592 4137
rect 10558 4035 10592 4069
rect 10558 3967 10592 4001
rect 10654 4851 10688 4885
rect 10654 4783 10688 4817
rect 10654 4715 10688 4749
rect 10654 4647 10688 4681
rect 10654 4579 10688 4613
rect 10654 4511 10688 4545
rect 10654 4443 10688 4477
rect 10654 4375 10688 4409
rect 10654 4307 10688 4341
rect 10654 4239 10688 4273
rect 10654 4171 10688 4205
rect 10654 4103 10688 4137
rect 10654 4035 10688 4069
rect 10654 3967 10688 4001
rect 10750 4851 10784 4885
rect 10750 4783 10784 4817
rect 10750 4715 10784 4749
rect 10750 4647 10784 4681
rect 10750 4579 10784 4613
rect 10750 4511 10784 4545
rect 10750 4443 10784 4477
rect 10750 4375 10784 4409
rect 10750 4307 10784 4341
rect 10750 4239 10784 4273
rect 10750 4171 10784 4205
rect 10750 4103 10784 4137
rect 10750 4035 10784 4069
rect 10750 3967 10784 4001
rect 10846 4851 10880 4885
rect 10846 4783 10880 4817
rect 10846 4715 10880 4749
rect 10846 4647 10880 4681
rect 10846 4579 10880 4613
rect 10846 4511 10880 4545
rect 10846 4443 10880 4477
rect 10846 4375 10880 4409
rect 10846 4307 10880 4341
rect 10846 4239 10880 4273
rect 10846 4171 10880 4205
rect 10846 4103 10880 4137
rect 10846 4035 10880 4069
rect 10846 3967 10880 4001
rect 15518 4909 15552 4943
rect 10942 4851 10976 4885
rect 10942 4783 10976 4817
rect 10942 4715 10976 4749
rect 10942 4647 10976 4681
rect 10942 4579 10976 4613
rect 10942 4511 10976 4545
rect 10942 4443 10976 4477
rect 10942 4375 10976 4409
rect 10942 4307 10976 4341
rect 10942 4239 10976 4273
rect 10942 4171 10976 4205
rect 10942 4103 10976 4137
rect 10942 4035 10976 4069
rect 10942 3967 10976 4001
rect 13714 4825 13748 4859
rect 13714 4757 13748 4791
rect 13714 4689 13748 4723
rect 13714 4621 13748 4655
rect 13714 4553 13748 4587
rect 13714 4485 13748 4519
rect 13714 4417 13748 4451
rect 13714 4349 13748 4383
rect 13714 4281 13748 4315
rect 13714 4213 13748 4247
rect 13714 4145 13748 4179
rect 13714 4077 13748 4111
rect 13714 4009 13748 4043
rect 13714 3941 13748 3975
rect 13810 4825 13844 4859
rect 13810 4757 13844 4791
rect 13810 4689 13844 4723
rect 13810 4621 13844 4655
rect 13810 4553 13844 4587
rect 13810 4485 13844 4519
rect 13810 4417 13844 4451
rect 13810 4349 13844 4383
rect 13810 4281 13844 4315
rect 13810 4213 13844 4247
rect 13810 4145 13844 4179
rect 13810 4077 13844 4111
rect 13810 4009 13844 4043
rect 13810 3941 13844 3975
rect 13906 4825 13940 4859
rect 13906 4757 13940 4791
rect 13906 4689 13940 4723
rect 13906 4621 13940 4655
rect 13906 4553 13940 4587
rect 13906 4485 13940 4519
rect 13906 4417 13940 4451
rect 13906 4349 13940 4383
rect 13906 4281 13940 4315
rect 13906 4213 13940 4247
rect 13906 4145 13940 4179
rect 13906 4077 13940 4111
rect 13906 4009 13940 4043
rect 13906 3941 13940 3975
rect 14002 4825 14036 4859
rect 14002 4757 14036 4791
rect 14002 4689 14036 4723
rect 14002 4621 14036 4655
rect 14002 4553 14036 4587
rect 14002 4485 14036 4519
rect 14002 4417 14036 4451
rect 14002 4349 14036 4383
rect 14002 4281 14036 4315
rect 14002 4213 14036 4247
rect 14002 4145 14036 4179
rect 14002 4077 14036 4111
rect 14002 4009 14036 4043
rect 14002 3941 14036 3975
rect 14098 4825 14132 4859
rect 14098 4757 14132 4791
rect 14098 4689 14132 4723
rect 14098 4621 14132 4655
rect 14098 4553 14132 4587
rect 14098 4485 14132 4519
rect 14098 4417 14132 4451
rect 14098 4349 14132 4383
rect 14098 4281 14132 4315
rect 14098 4213 14132 4247
rect 14098 4145 14132 4179
rect 14098 4077 14132 4111
rect 14098 4009 14132 4043
rect 14098 3941 14132 3975
rect 15518 4841 15552 4875
rect 15518 4773 15552 4807
rect 15518 4705 15552 4739
rect 15518 4637 15552 4671
rect 15518 4569 15552 4603
rect 15518 4501 15552 4535
rect 15518 4433 15552 4467
rect 15518 4365 15552 4399
rect 15518 4297 15552 4331
rect 15518 4229 15552 4263
rect 15518 4161 15552 4195
rect 15518 4093 15552 4127
rect 15518 4025 15552 4059
rect 15518 3957 15552 3991
rect 15614 5861 15648 5895
rect 15614 5793 15648 5827
rect 15614 5725 15648 5759
rect 15614 5657 15648 5691
rect 15614 5589 15648 5623
rect 15614 5521 15648 5555
rect 15614 5453 15648 5487
rect 15614 5385 15648 5419
rect 15614 5317 15648 5351
rect 15614 5249 15648 5283
rect 15614 5181 15648 5215
rect 15614 5113 15648 5147
rect 15614 5045 15648 5079
rect 15614 4977 15648 5011
rect 15614 4909 15648 4943
rect 15614 4841 15648 4875
rect 15614 4773 15648 4807
rect 15614 4705 15648 4739
rect 15614 4637 15648 4671
rect 15614 4569 15648 4603
rect 15614 4501 15648 4535
rect 15614 4433 15648 4467
rect 15614 4365 15648 4399
rect 15614 4297 15648 4331
rect 15614 4229 15648 4263
rect 15614 4161 15648 4195
rect 15614 4093 15648 4127
rect 15614 4025 15648 4059
rect 15614 3957 15648 3991
rect 15710 5861 15744 5895
rect 15710 5793 15744 5827
rect 15710 5725 15744 5759
rect 15710 5657 15744 5691
rect 15710 5589 15744 5623
rect 15710 5521 15744 5555
rect 15710 5453 15744 5487
rect 15710 5385 15744 5419
rect 15710 5317 15744 5351
rect 15710 5249 15744 5283
rect 15710 5181 15744 5215
rect 15710 5113 15744 5147
rect 15710 5045 15744 5079
rect 15710 4977 15744 5011
rect 15710 4909 15744 4943
rect 15710 4841 15744 4875
rect 15710 4773 15744 4807
rect 15710 4705 15744 4739
rect 15710 4637 15744 4671
rect 15710 4569 15744 4603
rect 15710 4501 15744 4535
rect 15710 4433 15744 4467
rect 15710 4365 15744 4399
rect 15710 4297 15744 4331
rect 15710 4229 15744 4263
rect 15710 4161 15744 4195
rect 15710 4093 15744 4127
rect 15710 4025 15744 4059
rect 15710 3957 15744 3991
<< psubdiff >>
rect -2308 833 -1944 884
rect -2308 255 -2279 833
rect -1973 255 -1944 833
rect -2308 204 -1944 255
<< nsubdiff >>
rect -2310 7123 -1942 7156
rect -2310 6477 -2279 7123
rect -1973 6477 -1942 7123
rect -2310 6444 -1942 6477
<< psubdiffcont >>
rect -2279 255 -1973 833
<< nsubdiffcont >>
rect -2279 6477 -1973 7123
<< poly >>
rect 272 6807 338 6823
rect 272 6773 288 6807
rect 322 6773 338 6807
rect 272 6757 338 6773
rect 2712 6803 2778 6819
rect 2712 6769 2728 6803
rect 2762 6769 2778 6803
rect 290 6702 320 6757
rect 2712 6753 2778 6769
rect 3228 6791 3294 6807
rect 3228 6757 3244 6791
rect 3278 6757 3294 6791
rect 2730 6706 2760 6753
rect 3228 6741 3294 6757
rect 5668 6787 5734 6803
rect 5668 6753 5684 6787
rect 5718 6753 5734 6787
rect 290 6674 370 6702
rect 2682 6696 2760 6706
rect 244 6644 1330 6674
rect 244 6606 274 6644
rect 340 6606 370 6644
rect 436 6606 466 6644
rect 532 6606 562 6644
rect 628 6606 658 6644
rect 724 6606 754 6644
rect 820 6606 850 6644
rect 916 6606 946 6644
rect 1012 6606 1042 6644
rect 1108 6606 1138 6644
rect 1204 6606 1234 6644
rect 1300 6606 1330 6644
rect 2010 6666 2760 6696
rect 3246 6686 3276 6741
rect 5668 6737 5734 6753
rect 6258 6791 6324 6807
rect 6258 6757 6274 6791
rect 6308 6757 6324 6791
rect 6258 6741 6324 6757
rect 8698 6787 8764 6803
rect 8698 6753 8714 6787
rect 8748 6753 8764 6787
rect 5686 6690 5716 6737
rect -1606 5936 -1566 5962
rect -1508 5936 -1468 5962
rect -1410 5936 -1370 5962
rect -1312 5936 -1272 5962
rect -1214 5936 -1174 5962
rect -1116 5936 -1076 5962
rect -1018 5936 -978 5962
rect -920 5936 -880 5962
rect 2010 6602 2040 6666
rect 2106 6602 2136 6666
rect 2202 6602 2232 6666
rect 2298 6602 2328 6666
rect 2394 6602 2424 6666
rect 2490 6602 2520 6666
rect 2586 6602 2616 6666
rect 2682 6602 2712 6666
rect 3246 6658 3326 6686
rect 5638 6680 5716 6690
rect 3200 6628 4286 6658
rect 244 5580 274 5606
rect 340 5580 370 5606
rect 436 5580 466 5606
rect 532 5580 562 5606
rect 628 5580 658 5606
rect 724 5580 754 5606
rect 820 5580 850 5606
rect 916 5580 946 5606
rect 1012 5580 1042 5606
rect 1108 5580 1138 5606
rect 1204 5580 1234 5606
rect 1300 5580 1330 5606
rect 3200 6590 3230 6628
rect 3296 6590 3326 6628
rect 3392 6590 3422 6628
rect 3488 6590 3518 6628
rect 3584 6590 3614 6628
rect 3680 6590 3710 6628
rect 3776 6590 3806 6628
rect 3872 6590 3902 6628
rect 3968 6590 3998 6628
rect 4064 6590 4094 6628
rect 4160 6590 4190 6628
rect 4256 6590 4286 6628
rect 4966 6650 5716 6680
rect 6276 6686 6306 6741
rect 8698 6737 8764 6753
rect 9346 6789 9412 6805
rect 9346 6755 9362 6789
rect 9396 6755 9412 6789
rect 9346 6739 9412 6755
rect 11786 6785 11852 6801
rect 11786 6751 11802 6785
rect 11836 6751 11852 6785
rect 8716 6690 8746 6737
rect 6276 6658 6356 6686
rect 8668 6680 8746 6690
rect 2010 5576 2040 5602
rect 2106 5576 2136 5602
rect 2202 5576 2232 5602
rect 2298 5576 2328 5602
rect 2394 5576 2424 5602
rect 2490 5576 2520 5602
rect 2586 5576 2616 5602
rect 2682 5576 2712 5602
rect 4966 6586 4996 6650
rect 5062 6586 5092 6650
rect 5158 6586 5188 6650
rect 5254 6586 5284 6650
rect 5350 6586 5380 6650
rect 5446 6586 5476 6650
rect 5542 6586 5572 6650
rect 5638 6586 5668 6650
rect 6230 6628 7316 6658
rect 6230 6590 6260 6628
rect 6326 6590 6356 6628
rect 6422 6590 6452 6628
rect 6518 6590 6548 6628
rect 6614 6590 6644 6628
rect 6710 6590 6740 6628
rect 6806 6590 6836 6628
rect 6902 6590 6932 6628
rect 6998 6590 7028 6628
rect 7094 6590 7124 6628
rect 7190 6590 7220 6628
rect 7286 6590 7316 6628
rect 7996 6650 8746 6680
rect 9364 6684 9394 6739
rect 11786 6735 11852 6751
rect 12502 6763 12568 6779
rect 11804 6688 11834 6735
rect 12502 6729 12518 6763
rect 12552 6729 12568 6763
rect 12502 6713 12568 6729
rect 14942 6759 15008 6775
rect 14942 6725 14958 6759
rect 14992 6725 15008 6759
rect 9364 6656 9444 6684
rect 11756 6678 11834 6688
rect 3200 5564 3230 5590
rect 3296 5564 3326 5590
rect 3392 5564 3422 5590
rect 3488 5564 3518 5590
rect 3584 5564 3614 5590
rect 3680 5564 3710 5590
rect 3776 5564 3806 5590
rect 3872 5564 3902 5590
rect 3968 5564 3998 5590
rect 4064 5564 4094 5590
rect 4160 5564 4190 5590
rect 4256 5564 4286 5590
rect 7996 6586 8026 6650
rect 8092 6586 8122 6650
rect 8188 6586 8218 6650
rect 8284 6586 8314 6650
rect 8380 6586 8410 6650
rect 8476 6586 8506 6650
rect 8572 6586 8602 6650
rect 8668 6586 8698 6650
rect 9318 6626 10404 6656
rect 9318 6588 9348 6626
rect 9414 6588 9444 6626
rect 9510 6588 9540 6626
rect 9606 6588 9636 6626
rect 9702 6588 9732 6626
rect 9798 6588 9828 6626
rect 9894 6588 9924 6626
rect 9990 6588 10020 6626
rect 10086 6588 10116 6626
rect 10182 6588 10212 6626
rect 10278 6588 10308 6626
rect 10374 6588 10404 6626
rect 11084 6648 11834 6678
rect 12520 6658 12550 6713
rect 14942 6709 15008 6725
rect 14960 6662 14990 6709
rect 4966 5560 4996 5586
rect 5062 5560 5092 5586
rect 5158 5560 5188 5586
rect 5254 5560 5284 5586
rect 5350 5560 5380 5586
rect 5446 5560 5476 5586
rect 5542 5560 5572 5586
rect 5638 5560 5668 5586
rect 6230 5564 6260 5590
rect 6326 5564 6356 5590
rect 6422 5564 6452 5590
rect 6518 5564 6548 5590
rect 6614 5564 6644 5590
rect 6710 5564 6740 5590
rect 6806 5564 6836 5590
rect 6902 5564 6932 5590
rect 6998 5564 7028 5590
rect 7094 5564 7124 5590
rect 7190 5564 7220 5590
rect 7286 5564 7316 5590
rect 11084 6584 11114 6648
rect 11180 6584 11210 6648
rect 11276 6584 11306 6648
rect 11372 6584 11402 6648
rect 11468 6584 11498 6648
rect 11564 6584 11594 6648
rect 11660 6584 11690 6648
rect 11756 6584 11786 6648
rect 12520 6630 12600 6658
rect 14912 6652 14990 6662
rect 12474 6600 13560 6630
rect 7996 5560 8026 5586
rect 8092 5560 8122 5586
rect 8188 5560 8218 5586
rect 8284 5560 8314 5586
rect 8380 5560 8410 5586
rect 8476 5560 8506 5586
rect 8572 5560 8602 5586
rect 8668 5560 8698 5586
rect 9318 5562 9348 5588
rect 9414 5562 9444 5588
rect 9510 5562 9540 5588
rect 9606 5562 9636 5588
rect 9702 5562 9732 5588
rect 9798 5562 9828 5588
rect 9894 5562 9924 5588
rect 9990 5562 10020 5588
rect 10086 5562 10116 5588
rect 10182 5562 10212 5588
rect 10278 5562 10308 5588
rect 10374 5562 10404 5588
rect 12474 6562 12504 6600
rect 12570 6562 12600 6600
rect 12666 6562 12696 6600
rect 12762 6562 12792 6600
rect 12858 6562 12888 6600
rect 12954 6562 12984 6600
rect 13050 6562 13080 6600
rect 13146 6562 13176 6600
rect 13242 6562 13272 6600
rect 13338 6562 13368 6600
rect 13434 6562 13464 6600
rect 13530 6562 13560 6600
rect 14240 6622 14990 6652
rect 11084 5558 11114 5584
rect 11180 5558 11210 5584
rect 11276 5558 11306 5584
rect 11372 5558 11402 5584
rect 11468 5558 11498 5584
rect 11564 5558 11594 5584
rect 11660 5558 11690 5584
rect 11756 5558 11786 5584
rect 14240 6558 14270 6622
rect 14336 6558 14366 6622
rect 14432 6558 14462 6622
rect 14528 6558 14558 6622
rect 14624 6558 14654 6622
rect 14720 6558 14750 6622
rect 14816 6558 14846 6622
rect 14912 6558 14942 6622
rect 12474 5536 12504 5562
rect 12570 5536 12600 5562
rect 12666 5536 12696 5562
rect 12762 5536 12792 5562
rect 12858 5536 12888 5562
rect 12954 5536 12984 5562
rect 13050 5536 13080 5562
rect 13146 5536 13176 5562
rect 13242 5536 13272 5562
rect 13338 5536 13368 5562
rect 13434 5536 13464 5562
rect 13530 5536 13560 5562
rect 15568 5926 15598 5952
rect 15664 5926 15694 5952
rect 14240 5532 14270 5558
rect 14336 5532 14366 5558
rect 14432 5532 14462 5558
rect 14528 5532 14558 5558
rect 14624 5532 14654 5558
rect 14720 5532 14750 5558
rect 14816 5532 14846 5558
rect 14912 5532 14942 5558
rect 1534 4990 1852 5020
rect 1534 4944 1564 4990
rect 1630 4944 1660 4990
rect 1726 4944 1756 4990
rect 1822 4944 1852 4990
rect 4490 4974 4808 5004
rect -1606 4866 -1566 4936
rect -1508 4866 -1468 4936
rect -1410 4868 -1370 4936
rect -1412 4866 -1370 4868
rect -1312 4866 -1272 4936
rect -1214 4866 -1174 4936
rect -1116 4866 -1076 4936
rect -1018 4866 -978 4936
rect -920 4866 -880 4936
rect -1606 4828 -880 4866
rect -1070 4785 -1030 4828
rect -1083 4769 -1017 4785
rect -1083 4735 -1067 4769
rect -1033 4735 -1017 4769
rect -1083 4719 -1017 4735
rect 4490 4928 4520 4974
rect 4586 4928 4616 4974
rect 4682 4928 4712 4974
rect 4778 4928 4808 4974
rect 7520 4974 7838 5004
rect 7520 4928 7550 4974
rect 7616 4928 7646 4974
rect 7712 4928 7742 4974
rect 7808 4928 7838 4974
rect 10608 4972 10926 5002
rect 1534 3874 1564 3944
rect 1630 3918 1660 3944
rect 1726 3874 1756 3944
rect 1822 3918 1852 3944
rect 10608 4926 10638 4972
rect 10704 4926 10734 4972
rect 10800 4926 10830 4972
rect 10896 4926 10926 4972
rect 13764 4946 14082 4976
rect 1534 3844 1612 3874
rect 1726 3844 1804 3874
rect 1582 3793 1612 3844
rect 1774 3793 1804 3844
rect 4490 3858 4520 3928
rect 4586 3902 4616 3928
rect 4682 3858 4712 3928
rect 4778 3902 4808 3928
rect 7520 3858 7550 3928
rect 7616 3902 7646 3928
rect 7712 3858 7742 3928
rect 7808 3902 7838 3928
rect 13764 4900 13794 4946
rect 13860 4900 13890 4946
rect 13956 4900 13986 4946
rect 14052 4900 14082 4946
rect 4490 3828 4568 3858
rect 4682 3828 4760 3858
rect 7520 3828 7598 3858
rect 7712 3828 7790 3858
rect 1564 3777 1630 3793
rect 1564 3743 1580 3777
rect 1614 3743 1630 3777
rect 1564 3727 1630 3743
rect 1756 3777 1822 3793
rect 4538 3777 4568 3828
rect 4730 3777 4760 3828
rect 7568 3777 7598 3828
rect 7760 3777 7790 3828
rect 10608 3856 10638 3926
rect 10704 3900 10734 3926
rect 10800 3856 10830 3926
rect 10896 3900 10926 3926
rect 10608 3826 10686 3856
rect 10800 3826 10878 3856
rect 1756 3743 1772 3777
rect 1806 3743 1822 3777
rect 1756 3727 1822 3743
rect 4520 3761 4586 3777
rect 4520 3727 4536 3761
rect 4570 3727 4586 3761
rect 4520 3711 4586 3727
rect 4712 3761 4778 3777
rect 4712 3727 4728 3761
rect 4762 3727 4778 3761
rect 4712 3711 4778 3727
rect 7550 3761 7616 3777
rect 7550 3727 7566 3761
rect 7600 3727 7616 3761
rect 7550 3711 7616 3727
rect 7742 3761 7808 3777
rect 10656 3775 10686 3826
rect 10848 3775 10878 3826
rect 13764 3830 13794 3900
rect 13860 3874 13890 3900
rect 13956 3830 13986 3900
rect 14052 3874 14082 3900
rect 15568 3876 15598 3926
rect 15664 3876 15694 3926
rect 15568 3846 15694 3876
rect 13764 3800 13842 3830
rect 13956 3800 14034 3830
rect 7742 3727 7758 3761
rect 7792 3727 7808 3761
rect 7742 3711 7808 3727
rect 10638 3759 10704 3775
rect 10638 3725 10654 3759
rect 10688 3725 10704 3759
rect 10638 3709 10704 3725
rect 10830 3759 10896 3775
rect 10830 3725 10846 3759
rect 10880 3725 10896 3759
rect 13812 3749 13842 3800
rect 14004 3749 14034 3800
rect 15568 3795 15598 3846
rect 15550 3779 15616 3795
rect 10830 3709 10896 3725
rect 13794 3733 13860 3749
rect 13794 3699 13810 3733
rect 13844 3699 13860 3733
rect 13794 3683 13860 3699
rect 13986 3733 14052 3749
rect 13986 3699 14002 3733
rect 14036 3699 14052 3733
rect 15550 3745 15566 3779
rect 15600 3745 15616 3779
rect 15550 3729 15616 3745
rect 13986 3683 14052 3699
rect -1606 3428 -1540 3444
rect -1606 3394 -1590 3428
rect -1556 3394 -1540 3428
rect -1606 3378 -1540 3394
rect -1590 3336 -1560 3378
rect -1636 3300 -934 3336
rect -1636 3236 -1606 3300
rect -1540 3236 -1510 3300
rect -1444 3236 -1414 3300
rect -1348 3236 -1318 3300
rect -1252 3236 -1222 3300
rect -1156 3236 -1126 3300
rect -1060 3236 -1030 3300
rect -964 3236 -934 3300
rect 1562 3002 1628 3018
rect 1562 2968 1578 3002
rect 1612 2968 1628 3002
rect 1562 2952 1628 2968
rect 1598 2922 1628 2952
rect 4518 2986 4584 3002
rect 4518 2952 4534 2986
rect 4568 2952 4584 2986
rect 4518 2936 4584 2952
rect 7548 2986 7614 3002
rect 7548 2952 7564 2986
rect 7598 2952 7614 2986
rect 7548 2936 7614 2952
rect 1598 2892 1658 2922
rect 4554 2906 4584 2936
rect 7584 2906 7614 2936
rect 10636 2984 10702 3000
rect 10636 2950 10652 2984
rect 10686 2950 10702 2984
rect 10636 2934 10702 2950
rect 1532 2862 1850 2892
rect 4554 2876 4614 2906
rect 7584 2876 7644 2906
rect 10672 2904 10702 2934
rect 13792 2958 13858 2974
rect 13792 2924 13808 2958
rect 13842 2924 13858 2958
rect 13792 2908 13858 2924
rect 1532 2830 1562 2862
rect 1628 2830 1658 2862
rect 1724 2854 1850 2862
rect 1724 2830 1754 2854
rect 1820 2830 1850 2854
rect 4488 2846 4806 2876
rect -1636 2210 -1606 2236
rect -1540 2210 -1510 2236
rect -1444 2210 -1414 2236
rect -1348 2210 -1318 2236
rect -1252 2210 -1222 2236
rect -1156 2210 -1126 2236
rect -1060 2210 -1030 2236
rect -964 2210 -934 2236
rect 4488 2814 4518 2846
rect 4584 2814 4614 2846
rect 4680 2838 4806 2846
rect 4680 2814 4710 2838
rect 4776 2814 4806 2838
rect 7518 2846 7836 2876
rect 10672 2874 10732 2904
rect 13828 2878 13858 2908
rect 7518 2814 7548 2846
rect 7614 2814 7644 2846
rect 7710 2838 7836 2846
rect 7710 2814 7740 2838
rect 7806 2814 7836 2838
rect 10606 2844 10924 2874
rect 13828 2848 13888 2878
rect 2546 2428 2646 2444
rect 2546 2394 2579 2428
rect 2613 2394 2646 2428
rect 2546 2276 2646 2394
rect 2546 2050 2646 2076
rect 1532 1804 1562 1830
rect 1628 1804 1658 1830
rect 1724 1804 1754 1830
rect 1820 1804 1850 1830
rect 5546 2428 5646 2444
rect 5546 2394 5579 2428
rect 5613 2394 5646 2428
rect 5546 2276 5646 2394
rect 5546 2050 5646 2076
rect 10606 2812 10636 2844
rect 10702 2812 10732 2844
rect 10798 2836 10924 2844
rect 10798 2812 10828 2836
rect 10894 2812 10924 2836
rect 13762 2818 14080 2848
rect 8546 2428 8646 2444
rect 8546 2394 8579 2428
rect 8613 2394 8646 2428
rect 8546 2276 8646 2394
rect 8546 2050 8646 2076
rect 4488 1788 4518 1814
rect 4584 1788 4614 1814
rect 4680 1788 4710 1814
rect 4776 1788 4806 1814
rect 7518 1788 7548 1814
rect 7614 1788 7644 1814
rect 7710 1788 7740 1814
rect 7806 1788 7836 1814
rect 13762 2786 13792 2818
rect 13858 2786 13888 2818
rect 13954 2810 14080 2818
rect 13954 2786 13984 2810
rect 14050 2786 14080 2810
rect 11546 2428 11646 2444
rect 11546 2394 11579 2428
rect 11613 2394 11646 2428
rect 11546 2276 11646 2394
rect 11546 2050 11646 2076
rect 10606 1786 10636 1812
rect 10702 1786 10732 1812
rect 10798 1786 10828 1812
rect 10894 1786 10924 1812
rect 14546 2428 14646 2444
rect 14546 2394 14579 2428
rect 14613 2394 14646 2428
rect 14546 2276 14646 2394
rect 14546 2050 14646 2076
rect 13762 1760 13792 1786
rect 13858 1760 13888 1786
rect 13954 1760 13984 1786
rect 14050 1760 14080 1786
rect 15450 1492 15516 1508
rect 15450 1458 15466 1492
rect 15500 1458 15516 1492
rect 15450 1442 15516 1458
rect -1111 1298 -1045 1314
rect -1111 1264 -1095 1298
rect -1061 1264 -1045 1298
rect -1111 1248 -1045 1264
rect -915 1298 -849 1314
rect -915 1264 -899 1298
rect -865 1264 -849 1298
rect 208 1306 1294 1336
rect 208 1268 238 1306
rect 304 1268 334 1306
rect 400 1268 430 1306
rect 496 1268 526 1306
rect 592 1268 622 1306
rect 688 1268 718 1306
rect 784 1268 814 1306
rect 880 1268 910 1306
rect 976 1268 1006 1306
rect 1072 1268 1102 1306
rect 1168 1268 1198 1306
rect 1264 1268 1294 1306
rect 1976 1310 2966 1340
rect 1976 1268 2006 1310
rect 2072 1268 2102 1310
rect 2168 1268 2198 1310
rect 2264 1268 2294 1310
rect 2360 1268 2390 1310
rect 2456 1268 2486 1310
rect 2552 1268 2582 1310
rect 2648 1268 2678 1310
rect 2744 1268 2774 1310
rect 2840 1268 2870 1310
rect 2936 1268 2966 1310
rect 3164 1290 4250 1320
rect -915 1248 -849 1264
rect -1100 1180 -1060 1248
rect -904 1180 -864 1248
rect -1640 1140 -858 1180
rect -1640 1066 -1600 1140
rect -1542 1066 -1502 1140
rect -1444 1066 -1404 1140
rect -1346 1066 -1306 1140
rect -1248 1066 -1208 1140
rect -1150 1066 -1110 1140
rect -1052 1066 -1012 1140
rect -954 1066 -914 1140
rect 3164 1252 3194 1290
rect 3260 1252 3290 1290
rect 3356 1252 3386 1290
rect 3452 1252 3482 1290
rect 3548 1252 3578 1290
rect 3644 1252 3674 1290
rect 3740 1252 3770 1290
rect 3836 1252 3866 1290
rect 3932 1252 3962 1290
rect 4028 1252 4058 1290
rect 4124 1252 4154 1290
rect 4220 1252 4250 1290
rect 4932 1294 5922 1324
rect 4932 1252 4962 1294
rect 5028 1252 5058 1294
rect 5124 1252 5154 1294
rect 5220 1252 5250 1294
rect 5316 1252 5346 1294
rect 5412 1252 5442 1294
rect 5508 1252 5538 1294
rect 5604 1252 5634 1294
rect 5700 1252 5730 1294
rect 5796 1252 5826 1294
rect 5892 1252 5922 1294
rect 6194 1290 7280 1320
rect 6194 1252 6224 1290
rect 6290 1252 6320 1290
rect 6386 1252 6416 1290
rect 6482 1252 6512 1290
rect 6578 1252 6608 1290
rect 6674 1252 6704 1290
rect 6770 1252 6800 1290
rect 6866 1252 6896 1290
rect 6962 1252 6992 1290
rect 7058 1252 7088 1290
rect 7154 1252 7184 1290
rect 7250 1252 7280 1290
rect 7962 1294 8952 1324
rect 7962 1252 7992 1294
rect 8058 1252 8088 1294
rect 8154 1252 8184 1294
rect 8250 1252 8280 1294
rect 8346 1252 8376 1294
rect 8442 1252 8472 1294
rect 8538 1252 8568 1294
rect 8634 1252 8664 1294
rect 8730 1252 8760 1294
rect 8826 1252 8856 1294
rect 8922 1252 8952 1294
rect 9282 1288 10368 1318
rect 208 214 238 268
rect 304 242 334 268
rect 400 242 430 268
rect 496 242 526 268
rect 592 242 622 268
rect 688 242 718 268
rect 784 242 814 268
rect 880 242 910 268
rect 976 242 1006 268
rect 1072 242 1102 268
rect 1168 242 1198 268
rect 1264 242 1294 268
rect 1976 242 2006 268
rect 2072 242 2102 268
rect 2168 242 2198 268
rect 2264 242 2294 268
rect 2360 242 2390 268
rect 2456 242 2486 268
rect 2552 242 2582 268
rect 2648 242 2678 268
rect 176 184 238 214
rect 2744 208 2774 268
rect 2840 242 2870 268
rect 2936 242 2966 268
rect 9282 1250 9312 1288
rect 9378 1250 9408 1288
rect 9474 1250 9504 1288
rect 9570 1250 9600 1288
rect 9666 1250 9696 1288
rect 9762 1250 9792 1288
rect 9858 1250 9888 1288
rect 9954 1250 9984 1288
rect 10050 1250 10080 1288
rect 10146 1250 10176 1288
rect 10242 1250 10272 1288
rect 10338 1250 10368 1288
rect 11050 1292 12040 1322
rect 15468 1300 15498 1442
rect 11050 1250 11080 1292
rect 11146 1250 11176 1292
rect 11242 1250 11272 1292
rect 11338 1250 11368 1292
rect 11434 1250 11464 1292
rect 11530 1250 11560 1292
rect 11626 1250 11656 1292
rect 11722 1250 11752 1292
rect 11818 1250 11848 1292
rect 11914 1250 11944 1292
rect 12010 1250 12040 1292
rect 12438 1262 13524 1292
rect 176 146 206 184
rect 2744 178 2802 208
rect 3164 198 3194 252
rect 3260 226 3290 252
rect 3356 226 3386 252
rect 3452 226 3482 252
rect 3548 226 3578 252
rect 3644 226 3674 252
rect 3740 226 3770 252
rect 3836 226 3866 252
rect 3932 226 3962 252
rect 4028 226 4058 252
rect 4124 226 4154 252
rect 4220 226 4250 252
rect 4932 226 4962 252
rect 5028 226 5058 252
rect 5124 226 5154 252
rect 5220 226 5250 252
rect 5316 226 5346 252
rect 5412 226 5442 252
rect 5508 226 5538 252
rect 5604 226 5634 252
rect 140 130 206 146
rect 140 96 156 130
rect 190 96 206 130
rect 140 80 206 96
rect 2772 146 2802 178
rect 3132 168 3194 198
rect 5700 192 5730 252
rect 5796 226 5826 252
rect 5892 226 5922 252
rect 6194 198 6224 252
rect 6290 226 6320 252
rect 6386 226 6416 252
rect 6482 226 6512 252
rect 6578 226 6608 252
rect 6674 226 6704 252
rect 6770 226 6800 252
rect 6866 226 6896 252
rect 6962 226 6992 252
rect 7058 226 7088 252
rect 7154 226 7184 252
rect 7250 226 7280 252
rect 7962 226 7992 252
rect 8058 226 8088 252
rect 8154 226 8184 252
rect 8250 226 8280 252
rect 8346 226 8376 252
rect 8442 226 8472 252
rect 8538 226 8568 252
rect 8634 226 8664 252
rect 2772 130 2838 146
rect 3132 130 3162 168
rect 5700 162 5758 192
rect 2772 96 2788 130
rect 2822 96 2838 130
rect 2772 80 2838 96
rect 3096 114 3162 130
rect 3096 80 3112 114
rect 3146 80 3162 114
rect -1640 40 -1600 66
rect -1542 40 -1502 66
rect -1444 40 -1404 66
rect -1346 40 -1306 66
rect -1248 40 -1208 66
rect -1150 40 -1110 66
rect -1052 40 -1012 66
rect -954 40 -914 66
rect 3096 64 3162 80
rect 5728 130 5758 162
rect 6162 168 6224 198
rect 8730 192 8760 252
rect 8826 226 8856 252
rect 8922 226 8952 252
rect 12438 1224 12468 1262
rect 12534 1224 12564 1262
rect 12630 1224 12660 1262
rect 12726 1224 12756 1262
rect 12822 1224 12852 1262
rect 12918 1224 12948 1262
rect 13014 1224 13044 1262
rect 13110 1224 13140 1262
rect 13206 1224 13236 1262
rect 13302 1224 13332 1262
rect 13398 1224 13428 1262
rect 13494 1224 13524 1262
rect 14206 1266 15196 1296
rect 14206 1224 14236 1266
rect 14302 1224 14332 1266
rect 14398 1224 14428 1266
rect 14494 1224 14524 1266
rect 14590 1224 14620 1266
rect 14686 1224 14716 1266
rect 14782 1224 14812 1266
rect 14878 1224 14908 1266
rect 14974 1224 15004 1266
rect 15070 1224 15100 1266
rect 15166 1224 15196 1266
rect 9282 196 9312 250
rect 9378 224 9408 250
rect 9474 224 9504 250
rect 9570 224 9600 250
rect 9666 224 9696 250
rect 9762 224 9792 250
rect 9858 224 9888 250
rect 9954 224 9984 250
rect 10050 224 10080 250
rect 10146 224 10176 250
rect 10242 224 10272 250
rect 10338 224 10368 250
rect 11050 224 11080 250
rect 11146 224 11176 250
rect 11242 224 11272 250
rect 11338 224 11368 250
rect 11434 224 11464 250
rect 11530 224 11560 250
rect 11626 224 11656 250
rect 11722 224 11752 250
rect 6162 130 6192 168
rect 8730 162 8788 192
rect 5728 114 5794 130
rect 5728 80 5744 114
rect 5778 80 5794 114
rect 5728 64 5794 80
rect 6126 114 6192 130
rect 6126 80 6142 114
rect 6176 80 6192 114
rect 6126 64 6192 80
rect 8758 130 8788 162
rect 9250 166 9312 196
rect 11818 190 11848 250
rect 11914 224 11944 250
rect 12010 224 12040 250
rect 8758 114 8824 130
rect 9250 128 9280 166
rect 11818 160 11876 190
rect 12438 170 12468 224
rect 12534 198 12564 224
rect 12630 198 12660 224
rect 12726 198 12756 224
rect 12822 198 12852 224
rect 12918 198 12948 224
rect 13014 198 13044 224
rect 13110 198 13140 224
rect 13206 198 13236 224
rect 13302 198 13332 224
rect 13398 198 13428 224
rect 13494 198 13524 224
rect 14206 198 14236 224
rect 14302 198 14332 224
rect 14398 198 14428 224
rect 14494 198 14524 224
rect 14590 198 14620 224
rect 14686 198 14716 224
rect 14782 198 14812 224
rect 14878 198 14908 224
rect 8758 80 8774 114
rect 8808 80 8824 114
rect 8758 64 8824 80
rect 9214 112 9280 128
rect 9214 78 9230 112
rect 9264 78 9280 112
rect 9214 62 9280 78
rect 11846 128 11876 160
rect 12406 140 12468 170
rect 14974 164 15004 224
rect 15070 198 15100 224
rect 15166 198 15196 224
rect 11846 112 11912 128
rect 11846 78 11862 112
rect 11896 78 11912 112
rect 12406 102 12436 140
rect 14974 134 15032 164
rect 11846 62 11912 78
rect 12370 86 12436 102
rect 12370 52 12386 86
rect 12420 52 12436 86
rect 12370 36 12436 52
rect 15002 102 15032 134
rect 15002 86 15068 102
rect 15002 52 15018 86
rect 15052 52 15068 86
rect 15468 74 15498 100
rect 15002 36 15068 52
<< polycont >>
rect 288 6773 322 6807
rect 2728 6769 2762 6803
rect 3244 6757 3278 6791
rect 5684 6753 5718 6787
rect 6274 6757 6308 6791
rect 8714 6753 8748 6787
rect 9362 6755 9396 6789
rect 11802 6751 11836 6785
rect 12518 6729 12552 6763
rect 14958 6725 14992 6759
rect -1067 4735 -1033 4769
rect 1580 3743 1614 3777
rect 1772 3743 1806 3777
rect 4536 3727 4570 3761
rect 4728 3727 4762 3761
rect 7566 3727 7600 3761
rect 7758 3727 7792 3761
rect 10654 3725 10688 3759
rect 10846 3725 10880 3759
rect 13810 3699 13844 3733
rect 14002 3699 14036 3733
rect 15566 3745 15600 3779
rect -1590 3394 -1556 3428
rect 1578 2968 1612 3002
rect 4534 2952 4568 2986
rect 7564 2952 7598 2986
rect 10652 2950 10686 2984
rect 13808 2924 13842 2958
rect 2579 2394 2613 2428
rect 5579 2394 5613 2428
rect 8579 2394 8613 2428
rect 11579 2394 11613 2428
rect 14579 2394 14613 2428
rect 15466 1458 15500 1492
rect -1095 1264 -1061 1298
rect -899 1264 -865 1298
rect 156 96 190 130
rect 2788 96 2822 130
rect 3112 80 3146 114
rect 5744 80 5778 114
rect 6142 80 6176 114
rect 8774 80 8808 114
rect 9230 78 9264 112
rect 11862 78 11896 112
rect 12386 52 12420 86
rect 15018 52 15052 86
<< locali >>
rect -2310 7123 -1942 7148
rect -2310 6477 -2279 7123
rect -1973 6728 -1942 7123
rect 272 6773 288 6807
rect 322 6773 338 6807
rect 764 6728 798 6858
rect 2712 6769 2728 6803
rect 2762 6769 2778 6803
rect 3228 6757 3244 6791
rect 3278 6757 3294 6791
rect -1973 6644 1392 6728
rect 2440 6702 2474 6754
rect 1960 6668 2768 6702
rect 3720 6684 3754 6842
rect 5668 6753 5684 6787
rect 5718 6753 5734 6787
rect 6258 6757 6274 6791
rect 6308 6757 6324 6791
rect 5396 6686 5430 6738
rect -1973 6477 -1942 6644
rect -2310 6452 -1942 6477
rect -1188 6042 -1102 6644
rect 194 6591 228 6644
rect 194 6519 228 6531
rect 194 6447 228 6463
rect 194 6375 228 6395
rect 194 6303 228 6327
rect 194 6231 228 6259
rect 194 6159 228 6191
rect 194 6089 228 6123
rect -1652 6006 -834 6042
rect -1652 5921 -1618 6006
rect -1652 5849 -1618 5861
rect -1652 5777 -1618 5793
rect -1652 5705 -1618 5725
rect -1652 5633 -1618 5657
rect -1652 5561 -1618 5589
rect -1652 5489 -1618 5521
rect -1652 5419 -1618 5453
rect -1652 5351 -1618 5383
rect -1652 5283 -1618 5311
rect -1652 5215 -1618 5239
rect -1652 5147 -1618 5167
rect -1652 5079 -1618 5095
rect -1652 5011 -1618 5023
rect -1652 4932 -1618 4951
rect -1554 5921 -1520 5938
rect -1554 5849 -1520 5861
rect -1554 5777 -1520 5793
rect -1554 5705 -1520 5725
rect -1554 5633 -1520 5657
rect -1554 5561 -1520 5589
rect -1554 5489 -1520 5521
rect -1554 5419 -1520 5453
rect -1554 5351 -1520 5383
rect -1554 5283 -1520 5311
rect -1554 5215 -1520 5239
rect -1554 5147 -1520 5167
rect -1554 5079 -1520 5095
rect -1554 5011 -1520 5023
rect -1554 4876 -1520 4951
rect -1456 5921 -1422 6006
rect -1456 5849 -1422 5861
rect -1456 5777 -1422 5793
rect -1456 5705 -1422 5725
rect -1456 5633 -1422 5657
rect -1456 5561 -1422 5589
rect -1456 5489 -1422 5521
rect -1456 5419 -1422 5453
rect -1456 5351 -1422 5383
rect -1456 5283 -1422 5311
rect -1456 5215 -1422 5239
rect -1456 5147 -1422 5167
rect -1456 5079 -1422 5095
rect -1456 5011 -1422 5023
rect -1456 4932 -1422 4951
rect -1358 5921 -1324 5938
rect -1358 5849 -1324 5861
rect -1358 5777 -1324 5793
rect -1358 5705 -1324 5725
rect -1358 5633 -1324 5657
rect -1358 5561 -1324 5589
rect -1358 5489 -1324 5521
rect -1358 5419 -1324 5453
rect -1358 5351 -1324 5383
rect -1358 5283 -1324 5311
rect -1358 5215 -1324 5239
rect -1358 5147 -1324 5167
rect -1358 5079 -1324 5095
rect -1358 5011 -1324 5023
rect -1358 4876 -1324 4951
rect -1260 5921 -1226 6006
rect -1260 5849 -1226 5861
rect -1260 5777 -1226 5793
rect -1260 5705 -1226 5725
rect -1260 5633 -1226 5657
rect -1260 5561 -1226 5589
rect -1260 5489 -1226 5521
rect -1260 5419 -1226 5453
rect -1260 5351 -1226 5383
rect -1260 5283 -1226 5311
rect -1260 5215 -1226 5239
rect -1260 5147 -1226 5167
rect -1260 5079 -1226 5095
rect -1260 5011 -1226 5023
rect -1260 4932 -1226 4951
rect -1162 5921 -1128 5938
rect -1162 5849 -1128 5861
rect -1162 5777 -1128 5793
rect -1162 5705 -1128 5725
rect -1162 5633 -1128 5657
rect -1162 5561 -1128 5589
rect -1162 5489 -1128 5521
rect -1162 5419 -1128 5453
rect -1162 5351 -1128 5383
rect -1162 5283 -1128 5311
rect -1162 5215 -1128 5239
rect -1162 5147 -1128 5167
rect -1162 5079 -1128 5095
rect -1162 5011 -1128 5023
rect -1162 4876 -1128 4951
rect -1064 5921 -1030 6006
rect -1064 5849 -1030 5861
rect -1064 5777 -1030 5793
rect -1064 5705 -1030 5725
rect -1064 5633 -1030 5657
rect -1064 5561 -1030 5589
rect -1064 5489 -1030 5521
rect -1064 5419 -1030 5453
rect -1064 5351 -1030 5383
rect -1064 5283 -1030 5311
rect -1064 5215 -1030 5239
rect -1064 5147 -1030 5167
rect -1064 5079 -1030 5095
rect -1064 5011 -1030 5023
rect -1064 4932 -1030 4951
rect -966 5921 -932 5938
rect -966 5849 -932 5861
rect -966 5777 -932 5793
rect -966 5705 -932 5725
rect -966 5633 -932 5657
rect -966 5561 -932 5589
rect -966 5489 -932 5521
rect -966 5419 -932 5453
rect -966 5351 -932 5383
rect -966 5283 -932 5311
rect -966 5215 -932 5239
rect -966 5147 -932 5167
rect -966 5079 -932 5095
rect -966 5011 -932 5023
rect -966 4876 -932 4951
rect -868 5921 -834 6006
rect -868 5849 -834 5861
rect -868 5777 -834 5793
rect -868 5705 -834 5725
rect -868 5633 -834 5657
rect 194 6021 228 6053
rect 194 5953 228 5981
rect 194 5885 228 5909
rect 194 5817 228 5837
rect 194 5749 228 5765
rect 194 5681 228 5693
rect 194 5602 228 5621
rect 290 6591 324 6608
rect 290 6519 324 6531
rect 290 6447 324 6463
rect 290 6375 324 6395
rect 290 6303 324 6327
rect 290 6231 324 6259
rect 290 6159 324 6191
rect 290 6089 324 6123
rect 290 6021 324 6053
rect 290 5953 324 5981
rect 290 5885 324 5909
rect 290 5817 324 5837
rect 290 5749 324 5765
rect 290 5681 324 5693
rect -868 5561 -834 5589
rect -868 5489 -834 5521
rect 290 5550 324 5621
rect 386 6591 420 6644
rect 386 6519 420 6531
rect 386 6447 420 6463
rect 386 6375 420 6395
rect 386 6303 420 6327
rect 386 6231 420 6259
rect 386 6159 420 6191
rect 386 6089 420 6123
rect 386 6021 420 6053
rect 386 5953 420 5981
rect 386 5885 420 5909
rect 386 5817 420 5837
rect 386 5749 420 5765
rect 386 5681 420 5693
rect 386 5604 420 5621
rect 482 6591 516 6608
rect 482 6519 516 6531
rect 482 6447 516 6463
rect 482 6375 516 6395
rect 482 6303 516 6327
rect 482 6231 516 6259
rect 482 6159 516 6191
rect 482 6089 516 6123
rect 482 6021 516 6053
rect 482 5953 516 5981
rect 482 5885 516 5909
rect 482 5817 516 5837
rect 482 5749 516 5765
rect 482 5681 516 5693
rect 482 5550 516 5621
rect 578 6591 612 6644
rect 578 6519 612 6531
rect 578 6447 612 6463
rect 578 6375 612 6395
rect 578 6303 612 6327
rect 578 6231 612 6259
rect 578 6159 612 6191
rect 578 6089 612 6123
rect 578 6021 612 6053
rect 578 5953 612 5981
rect 578 5885 612 5909
rect 578 5817 612 5837
rect 578 5749 612 5765
rect 578 5681 612 5693
rect 578 5604 612 5621
rect 674 6591 708 6608
rect 674 6519 708 6531
rect 674 6447 708 6463
rect 674 6375 708 6395
rect 674 6303 708 6327
rect 674 6231 708 6259
rect 674 6159 708 6191
rect 674 6089 708 6123
rect 674 6021 708 6053
rect 674 5953 708 5981
rect 674 5885 708 5909
rect 674 5817 708 5837
rect 674 5749 708 5765
rect 674 5681 708 5693
rect 674 5550 708 5621
rect 770 6591 804 6644
rect 770 6519 804 6531
rect 770 6447 804 6463
rect 770 6375 804 6395
rect 770 6303 804 6327
rect 770 6231 804 6259
rect 770 6159 804 6191
rect 770 6089 804 6123
rect 770 6021 804 6053
rect 770 5953 804 5981
rect 770 5885 804 5909
rect 770 5817 804 5837
rect 770 5749 804 5765
rect 770 5681 804 5693
rect 770 5604 804 5621
rect 866 6591 900 6608
rect 866 6519 900 6531
rect 866 6447 900 6463
rect 866 6375 900 6395
rect 866 6303 900 6327
rect 866 6231 900 6259
rect 866 6159 900 6191
rect 866 6089 900 6123
rect 866 6021 900 6053
rect 866 5953 900 5981
rect 866 5885 900 5909
rect 866 5817 900 5837
rect 866 5749 900 5765
rect 866 5681 900 5693
rect 866 5550 900 5621
rect 962 6591 996 6644
rect 962 6519 996 6531
rect 962 6447 996 6463
rect 962 6375 996 6395
rect 962 6303 996 6327
rect 962 6231 996 6259
rect 962 6159 996 6191
rect 962 6089 996 6123
rect 962 6021 996 6053
rect 962 5953 996 5981
rect 962 5885 996 5909
rect 962 5817 996 5837
rect 962 5749 996 5765
rect 962 5681 996 5693
rect 962 5604 996 5621
rect 1058 6591 1092 6608
rect 1058 6519 1092 6531
rect 1058 6447 1092 6463
rect 1058 6375 1092 6395
rect 1058 6303 1092 6327
rect 1058 6231 1092 6259
rect 1058 6159 1092 6191
rect 1058 6089 1092 6123
rect 1058 6021 1092 6053
rect 1058 5953 1092 5981
rect 1058 5885 1092 5909
rect 1058 5817 1092 5837
rect 1058 5749 1092 5765
rect 1058 5681 1092 5693
rect 1058 5550 1092 5621
rect 1154 6591 1188 6644
rect 1154 6519 1188 6531
rect 1154 6447 1188 6463
rect 1154 6375 1188 6395
rect 1154 6303 1188 6327
rect 1154 6231 1188 6259
rect 1154 6159 1188 6191
rect 1154 6089 1188 6123
rect 1154 6021 1188 6053
rect 1154 5953 1188 5981
rect 1154 5885 1188 5909
rect 1154 5817 1188 5837
rect 1154 5749 1188 5765
rect 1154 5681 1188 5693
rect 1154 5604 1188 5621
rect 1250 6591 1284 6608
rect 1250 6519 1284 6531
rect 1250 6447 1284 6463
rect 1250 6375 1284 6395
rect 1250 6303 1284 6327
rect 1250 6231 1284 6259
rect 1250 6159 1284 6191
rect 1250 6089 1284 6123
rect 1250 6021 1284 6053
rect 1250 5953 1284 5981
rect 1250 5885 1284 5909
rect 1250 5817 1284 5837
rect 1250 5749 1284 5765
rect 1250 5681 1284 5693
rect 1250 5550 1284 5621
rect 1346 6591 1380 6644
rect 1346 6519 1380 6531
rect 1346 6447 1380 6463
rect 1346 6375 1380 6395
rect 1346 6303 1380 6327
rect 1346 6231 1380 6259
rect 1346 6159 1380 6191
rect 1346 6089 1380 6123
rect 1346 6021 1380 6053
rect 1346 5953 1380 5981
rect 1346 5885 1380 5909
rect 1346 5817 1380 5837
rect 1346 5749 1380 5765
rect 1346 5681 1380 5693
rect 1346 5604 1380 5621
rect 1960 6587 1994 6668
rect 1960 6515 1994 6527
rect 1960 6443 1994 6459
rect 1960 6371 1994 6391
rect 1960 6299 1994 6323
rect 1960 6227 1994 6255
rect 1960 6155 1994 6187
rect 1960 6085 1994 6119
rect 1960 6017 1994 6049
rect 1960 5949 1994 5977
rect 1960 5881 1994 5905
rect 1960 5813 1994 5833
rect 1960 5745 1994 5761
rect 1960 5677 1994 5689
rect 1960 5598 1994 5617
rect 2056 6587 2090 6604
rect 2056 6515 2090 6527
rect 2056 6443 2090 6459
rect 2056 6371 2090 6391
rect 2056 6299 2090 6323
rect 2056 6227 2090 6255
rect 2056 6155 2090 6187
rect 2056 6085 2090 6119
rect 2056 6017 2090 6049
rect 2056 5949 2090 5977
rect 2056 5881 2090 5905
rect 2056 5813 2090 5833
rect 2056 5745 2090 5761
rect 2056 5677 2090 5689
rect 290 5516 1284 5550
rect 2056 5548 2090 5617
rect 2152 6587 2186 6668
rect 2152 6515 2186 6527
rect 2152 6443 2186 6459
rect 2152 6371 2186 6391
rect 2152 6299 2186 6323
rect 2152 6227 2186 6255
rect 2152 6155 2186 6187
rect 2152 6085 2186 6119
rect 2152 6017 2186 6049
rect 2152 5949 2186 5977
rect 2152 5881 2186 5905
rect 2152 5813 2186 5833
rect 2152 5745 2186 5761
rect 2152 5677 2186 5689
rect 2152 5598 2186 5617
rect 2248 6587 2282 6604
rect 2248 6515 2282 6527
rect 2248 6443 2282 6459
rect 2248 6371 2282 6391
rect 2248 6299 2282 6323
rect 2248 6227 2282 6255
rect 2248 6155 2282 6187
rect 2248 6085 2282 6119
rect 2248 6017 2282 6049
rect 2248 5949 2282 5977
rect 2248 5881 2282 5905
rect 2248 5813 2282 5833
rect 2248 5745 2282 5761
rect 2248 5677 2282 5689
rect 2248 5548 2282 5617
rect 2344 6587 2378 6668
rect 2344 6515 2378 6527
rect 2344 6443 2378 6459
rect 2344 6371 2378 6391
rect 2344 6299 2378 6323
rect 2344 6227 2378 6255
rect 2344 6155 2378 6187
rect 2344 6085 2378 6119
rect 2344 6017 2378 6049
rect 2344 5949 2378 5977
rect 2344 5881 2378 5905
rect 2344 5813 2378 5833
rect 2344 5745 2378 5761
rect 2344 5677 2378 5689
rect 2344 5598 2378 5617
rect 2440 6587 2474 6604
rect 2440 6515 2474 6527
rect 2440 6443 2474 6459
rect 2440 6371 2474 6391
rect 2440 6299 2474 6323
rect 2440 6227 2474 6255
rect 2440 6155 2474 6187
rect 2440 6085 2474 6119
rect 2440 6017 2474 6049
rect 2440 5949 2474 5977
rect 2440 5881 2474 5905
rect 2440 5813 2474 5833
rect 2440 5745 2474 5761
rect 2440 5677 2474 5689
rect 2440 5548 2474 5617
rect 2536 6587 2570 6668
rect 2536 6515 2570 6527
rect 2536 6443 2570 6459
rect 2536 6371 2570 6391
rect 2536 6299 2570 6323
rect 2536 6227 2570 6255
rect 2536 6155 2570 6187
rect 2536 6085 2570 6119
rect 2536 6017 2570 6049
rect 2536 5949 2570 5977
rect 2536 5881 2570 5905
rect 2536 5813 2570 5833
rect 2536 5745 2570 5761
rect 2536 5677 2570 5689
rect 2536 5598 2570 5617
rect 2632 6587 2666 6604
rect 2632 6515 2666 6527
rect 2632 6443 2666 6459
rect 2632 6371 2666 6391
rect 2632 6299 2666 6323
rect 2632 6227 2666 6255
rect 2632 6155 2666 6187
rect 2632 6085 2666 6119
rect 2632 6017 2666 6049
rect 2632 5949 2666 5977
rect 2632 5881 2666 5905
rect 2632 5813 2666 5833
rect 2632 5745 2666 5761
rect 2632 5677 2666 5689
rect 2632 5548 2666 5617
rect 2728 6587 2762 6668
rect 2728 6515 2762 6527
rect 2728 6443 2762 6459
rect 2728 6371 2762 6391
rect 2728 6299 2762 6323
rect 2728 6227 2762 6255
rect 2728 6155 2762 6187
rect 2728 6085 2762 6119
rect 2728 6017 2762 6049
rect 2728 5949 2762 5977
rect 2728 5881 2762 5905
rect 2728 5813 2762 5833
rect 2728 5745 2762 5761
rect 2728 5677 2762 5689
rect 2728 5600 2762 5617
rect 3150 6650 4344 6684
rect 4916 6652 5724 6686
rect 6750 6684 6784 6842
rect 8698 6753 8714 6787
rect 8748 6753 8764 6787
rect 9346 6755 9362 6789
rect 9396 6755 9412 6789
rect 8426 6686 8460 6738
rect 3150 6575 3184 6650
rect 3150 6503 3184 6515
rect 3150 6431 3184 6447
rect 3150 6359 3184 6379
rect 3150 6287 3184 6311
rect 3150 6215 3184 6243
rect 3150 6143 3184 6175
rect 3150 6073 3184 6107
rect 3150 6005 3184 6037
rect 3150 5937 3184 5965
rect 3150 5869 3184 5893
rect 3150 5801 3184 5821
rect 3150 5733 3184 5749
rect 3150 5665 3184 5677
rect 3150 5586 3184 5605
rect 3246 6575 3280 6592
rect 3246 6503 3280 6515
rect 3246 6431 3280 6447
rect 3246 6359 3280 6379
rect 3246 6287 3280 6311
rect 3246 6215 3280 6243
rect 3246 6143 3280 6175
rect 3246 6073 3280 6107
rect 3246 6005 3280 6037
rect 3246 5937 3280 5965
rect 3246 5869 3280 5893
rect 3246 5801 3280 5821
rect 3246 5733 3280 5749
rect 3246 5665 3280 5677
rect -868 5419 -834 5453
rect -868 5351 -834 5383
rect 880 5406 914 5516
rect 2056 5514 2666 5548
rect 3246 5534 3280 5605
rect 3342 6575 3376 6650
rect 3342 6503 3376 6515
rect 3342 6431 3376 6447
rect 3342 6359 3376 6379
rect 3342 6287 3376 6311
rect 3342 6215 3376 6243
rect 3342 6143 3376 6175
rect 3342 6073 3376 6107
rect 3342 6005 3376 6037
rect 3342 5937 3376 5965
rect 3342 5869 3376 5893
rect 3342 5801 3376 5821
rect 3342 5733 3376 5749
rect 3342 5665 3376 5677
rect 3342 5588 3376 5605
rect 3438 6575 3472 6592
rect 3438 6503 3472 6515
rect 3438 6431 3472 6447
rect 3438 6359 3472 6379
rect 3438 6287 3472 6311
rect 3438 6215 3472 6243
rect 3438 6143 3472 6175
rect 3438 6073 3472 6107
rect 3438 6005 3472 6037
rect 3438 5937 3472 5965
rect 3438 5869 3472 5893
rect 3438 5801 3472 5821
rect 3438 5733 3472 5749
rect 3438 5665 3472 5677
rect 3438 5534 3472 5605
rect 3534 6575 3568 6650
rect 3534 6503 3568 6515
rect 3534 6431 3568 6447
rect 3534 6359 3568 6379
rect 3534 6287 3568 6311
rect 3534 6215 3568 6243
rect 3534 6143 3568 6175
rect 3534 6073 3568 6107
rect 3534 6005 3568 6037
rect 3534 5937 3568 5965
rect 3534 5869 3568 5893
rect 3534 5801 3568 5821
rect 3534 5733 3568 5749
rect 3534 5665 3568 5677
rect 3534 5588 3568 5605
rect 3630 6575 3664 6592
rect 3630 6503 3664 6515
rect 3630 6431 3664 6447
rect 3630 6359 3664 6379
rect 3630 6287 3664 6311
rect 3630 6215 3664 6243
rect 3630 6143 3664 6175
rect 3630 6073 3664 6107
rect 3630 6005 3664 6037
rect 3630 5937 3664 5965
rect 3630 5869 3664 5893
rect 3630 5801 3664 5821
rect 3630 5733 3664 5749
rect 3630 5665 3664 5677
rect 3630 5534 3664 5605
rect 3726 6575 3760 6650
rect 3726 6503 3760 6515
rect 3726 6431 3760 6447
rect 3726 6359 3760 6379
rect 3726 6287 3760 6311
rect 3726 6215 3760 6243
rect 3726 6143 3760 6175
rect 3726 6073 3760 6107
rect 3726 6005 3760 6037
rect 3726 5937 3760 5965
rect 3726 5869 3760 5893
rect 3726 5801 3760 5821
rect 3726 5733 3760 5749
rect 3726 5665 3760 5677
rect 3726 5588 3760 5605
rect 3822 6575 3856 6592
rect 3822 6503 3856 6515
rect 3822 6431 3856 6447
rect 3822 6359 3856 6379
rect 3822 6287 3856 6311
rect 3822 6215 3856 6243
rect 3822 6143 3856 6175
rect 3822 6073 3856 6107
rect 3822 6005 3856 6037
rect 3822 5937 3856 5965
rect 3822 5869 3856 5893
rect 3822 5801 3856 5821
rect 3822 5733 3856 5749
rect 3822 5665 3856 5677
rect 3822 5534 3856 5605
rect 3918 6575 3952 6650
rect 3918 6503 3952 6515
rect 3918 6431 3952 6447
rect 3918 6359 3952 6379
rect 3918 6287 3952 6311
rect 3918 6215 3952 6243
rect 3918 6143 3952 6175
rect 3918 6073 3952 6107
rect 3918 6005 3952 6037
rect 3918 5937 3952 5965
rect 3918 5869 3952 5893
rect 3918 5801 3952 5821
rect 3918 5733 3952 5749
rect 3918 5665 3952 5677
rect 3918 5588 3952 5605
rect 4014 6575 4048 6592
rect 4014 6503 4048 6515
rect 4014 6431 4048 6447
rect 4014 6359 4048 6379
rect 4014 6287 4048 6311
rect 4014 6215 4048 6243
rect 4014 6143 4048 6175
rect 4014 6073 4048 6107
rect 4014 6005 4048 6037
rect 4014 5937 4048 5965
rect 4014 5869 4048 5893
rect 4014 5801 4048 5821
rect 4014 5733 4048 5749
rect 4014 5665 4048 5677
rect 4014 5534 4048 5605
rect 4110 6575 4144 6650
rect 4110 6503 4144 6515
rect 4110 6431 4144 6447
rect 4110 6359 4144 6379
rect 4110 6287 4144 6311
rect 4110 6215 4144 6243
rect 4110 6143 4144 6175
rect 4110 6073 4144 6107
rect 4110 6005 4144 6037
rect 4110 5937 4144 5965
rect 4110 5869 4144 5893
rect 4110 5801 4144 5821
rect 4110 5733 4144 5749
rect 4110 5665 4144 5677
rect 4110 5588 4144 5605
rect 4206 6575 4240 6592
rect 4206 6503 4240 6515
rect 4206 6431 4240 6447
rect 4206 6359 4240 6379
rect 4206 6287 4240 6311
rect 4206 6215 4240 6243
rect 4206 6143 4240 6175
rect 4206 6073 4240 6107
rect 4206 6005 4240 6037
rect 4206 5937 4240 5965
rect 4206 5869 4240 5893
rect 4206 5801 4240 5821
rect 4206 5733 4240 5749
rect 4206 5665 4240 5677
rect 4206 5534 4240 5605
rect 4302 6575 4336 6650
rect 4302 6503 4336 6515
rect 4302 6431 4336 6447
rect 4302 6359 4336 6379
rect 4302 6287 4336 6311
rect 4302 6215 4336 6243
rect 4302 6143 4336 6175
rect 4302 6073 4336 6107
rect 4302 6005 4336 6037
rect 4302 5937 4336 5965
rect 4302 5869 4336 5893
rect 4302 5801 4336 5821
rect 4302 5733 4336 5749
rect 4302 5665 4336 5677
rect 4302 5588 4336 5605
rect 4916 6571 4950 6652
rect 4916 6499 4950 6511
rect 4916 6427 4950 6443
rect 4916 6355 4950 6375
rect 4916 6283 4950 6307
rect 4916 6211 4950 6239
rect 4916 6139 4950 6171
rect 4916 6069 4950 6103
rect 4916 6001 4950 6033
rect 4916 5933 4950 5961
rect 4916 5865 4950 5889
rect 4916 5797 4950 5817
rect 4916 5729 4950 5745
rect 4916 5661 4950 5673
rect 4916 5582 4950 5601
rect 5012 6571 5046 6588
rect 5012 6499 5046 6511
rect 5012 6427 5046 6443
rect 5012 6355 5046 6375
rect 5012 6283 5046 6307
rect 5012 6211 5046 6239
rect 5012 6139 5046 6171
rect 5012 6069 5046 6103
rect 5012 6001 5046 6033
rect 5012 5933 5046 5961
rect 5012 5865 5046 5889
rect 5012 5797 5046 5817
rect 5012 5729 5046 5745
rect 5012 5661 5046 5673
rect 2344 5410 2378 5514
rect 3246 5500 4240 5534
rect 5012 5532 5046 5601
rect 5108 6571 5142 6652
rect 5108 6499 5142 6511
rect 5108 6427 5142 6443
rect 5108 6355 5142 6375
rect 5108 6283 5142 6307
rect 5108 6211 5142 6239
rect 5108 6139 5142 6171
rect 5108 6069 5142 6103
rect 5108 6001 5142 6033
rect 5108 5933 5142 5961
rect 5108 5865 5142 5889
rect 5108 5797 5142 5817
rect 5108 5729 5142 5745
rect 5108 5661 5142 5673
rect 5108 5582 5142 5601
rect 5204 6571 5238 6588
rect 5204 6499 5238 6511
rect 5204 6427 5238 6443
rect 5204 6355 5238 6375
rect 5204 6283 5238 6307
rect 5204 6211 5238 6239
rect 5204 6139 5238 6171
rect 5204 6069 5238 6103
rect 5204 6001 5238 6033
rect 5204 5933 5238 5961
rect 5204 5865 5238 5889
rect 5204 5797 5238 5817
rect 5204 5729 5238 5745
rect 5204 5661 5238 5673
rect 5204 5532 5238 5601
rect 5300 6571 5334 6652
rect 5300 6499 5334 6511
rect 5300 6427 5334 6443
rect 5300 6355 5334 6375
rect 5300 6283 5334 6307
rect 5300 6211 5334 6239
rect 5300 6139 5334 6171
rect 5300 6069 5334 6103
rect 5300 6001 5334 6033
rect 5300 5933 5334 5961
rect 5300 5865 5334 5889
rect 5300 5797 5334 5817
rect 5300 5729 5334 5745
rect 5300 5661 5334 5673
rect 5300 5582 5334 5601
rect 5396 6571 5430 6588
rect 5396 6499 5430 6511
rect 5396 6427 5430 6443
rect 5396 6355 5430 6375
rect 5396 6283 5430 6307
rect 5396 6211 5430 6239
rect 5396 6139 5430 6171
rect 5396 6069 5430 6103
rect 5396 6001 5430 6033
rect 5396 5933 5430 5961
rect 5396 5865 5430 5889
rect 5396 5797 5430 5817
rect 5396 5729 5430 5745
rect 5396 5661 5430 5673
rect 5396 5532 5430 5601
rect 5492 6571 5526 6652
rect 5492 6499 5526 6511
rect 5492 6427 5526 6443
rect 5492 6355 5526 6375
rect 5492 6283 5526 6307
rect 5492 6211 5526 6239
rect 5492 6139 5526 6171
rect 5492 6069 5526 6103
rect 5492 6001 5526 6033
rect 5492 5933 5526 5961
rect 5492 5865 5526 5889
rect 5492 5797 5526 5817
rect 5492 5729 5526 5745
rect 5492 5661 5526 5673
rect 5492 5582 5526 5601
rect 5588 6571 5622 6588
rect 5588 6499 5622 6511
rect 5588 6427 5622 6443
rect 5588 6355 5622 6375
rect 5588 6283 5622 6307
rect 5588 6211 5622 6239
rect 5588 6139 5622 6171
rect 5588 6069 5622 6103
rect 5588 6001 5622 6033
rect 5588 5933 5622 5961
rect 5588 5865 5622 5889
rect 5588 5797 5622 5817
rect 5588 5729 5622 5745
rect 5588 5661 5622 5673
rect 5588 5532 5622 5601
rect 5684 6571 5718 6652
rect 5684 6499 5718 6511
rect 5684 6427 5718 6443
rect 5684 6355 5718 6375
rect 5684 6283 5718 6307
rect 5684 6211 5718 6239
rect 5684 6139 5718 6171
rect 5684 6069 5718 6103
rect 5684 6001 5718 6033
rect 5684 5933 5718 5961
rect 5684 5865 5718 5889
rect 5684 5797 5718 5817
rect 5684 5729 5718 5745
rect 5684 5661 5718 5673
rect 5684 5584 5718 5601
rect 6180 6650 7374 6684
rect 7946 6652 8754 6686
rect 9838 6682 9872 6840
rect 11786 6751 11802 6785
rect 11836 6751 11852 6785
rect 11514 6684 11548 6736
rect 12502 6729 12518 6763
rect 12552 6729 12568 6763
rect 6180 6575 6214 6650
rect 6180 6503 6214 6515
rect 6180 6431 6214 6447
rect 6180 6359 6214 6379
rect 6180 6287 6214 6311
rect 6180 6215 6214 6243
rect 6180 6143 6214 6175
rect 6180 6073 6214 6107
rect 6180 6005 6214 6037
rect 6180 5937 6214 5965
rect 6180 5869 6214 5893
rect 6180 5801 6214 5821
rect 6180 5733 6214 5749
rect 6180 5665 6214 5677
rect 6180 5586 6214 5605
rect 6276 6575 6310 6592
rect 6276 6503 6310 6515
rect 6276 6431 6310 6447
rect 6276 6359 6310 6379
rect 6276 6287 6310 6311
rect 6276 6215 6310 6243
rect 6276 6143 6310 6175
rect 6276 6073 6310 6107
rect 6276 6005 6310 6037
rect 6276 5937 6310 5965
rect 6276 5869 6310 5893
rect 6276 5801 6310 5821
rect 6276 5733 6310 5749
rect 6276 5665 6310 5677
rect 3836 5390 3870 5500
rect 5012 5498 5622 5532
rect 6276 5534 6310 5605
rect 6372 6575 6406 6650
rect 6372 6503 6406 6515
rect 6372 6431 6406 6447
rect 6372 6359 6406 6379
rect 6372 6287 6406 6311
rect 6372 6215 6406 6243
rect 6372 6143 6406 6175
rect 6372 6073 6406 6107
rect 6372 6005 6406 6037
rect 6372 5937 6406 5965
rect 6372 5869 6406 5893
rect 6372 5801 6406 5821
rect 6372 5733 6406 5749
rect 6372 5665 6406 5677
rect 6372 5588 6406 5605
rect 6468 6575 6502 6592
rect 6468 6503 6502 6515
rect 6468 6431 6502 6447
rect 6468 6359 6502 6379
rect 6468 6287 6502 6311
rect 6468 6215 6502 6243
rect 6468 6143 6502 6175
rect 6468 6073 6502 6107
rect 6468 6005 6502 6037
rect 6468 5937 6502 5965
rect 6468 5869 6502 5893
rect 6468 5801 6502 5821
rect 6468 5733 6502 5749
rect 6468 5665 6502 5677
rect 6468 5534 6502 5605
rect 6564 6575 6598 6650
rect 6564 6503 6598 6515
rect 6564 6431 6598 6447
rect 6564 6359 6598 6379
rect 6564 6287 6598 6311
rect 6564 6215 6598 6243
rect 6564 6143 6598 6175
rect 6564 6073 6598 6107
rect 6564 6005 6598 6037
rect 6564 5937 6598 5965
rect 6564 5869 6598 5893
rect 6564 5801 6598 5821
rect 6564 5733 6598 5749
rect 6564 5665 6598 5677
rect 6564 5588 6598 5605
rect 6660 6575 6694 6592
rect 6660 6503 6694 6515
rect 6660 6431 6694 6447
rect 6660 6359 6694 6379
rect 6660 6287 6694 6311
rect 6660 6215 6694 6243
rect 6660 6143 6694 6175
rect 6660 6073 6694 6107
rect 6660 6005 6694 6037
rect 6660 5937 6694 5965
rect 6660 5869 6694 5893
rect 6660 5801 6694 5821
rect 6660 5733 6694 5749
rect 6660 5665 6694 5677
rect 6660 5534 6694 5605
rect 6756 6575 6790 6650
rect 6756 6503 6790 6515
rect 6756 6431 6790 6447
rect 6756 6359 6790 6379
rect 6756 6287 6790 6311
rect 6756 6215 6790 6243
rect 6756 6143 6790 6175
rect 6756 6073 6790 6107
rect 6756 6005 6790 6037
rect 6756 5937 6790 5965
rect 6756 5869 6790 5893
rect 6756 5801 6790 5821
rect 6756 5733 6790 5749
rect 6756 5665 6790 5677
rect 6756 5588 6790 5605
rect 6852 6575 6886 6592
rect 6852 6503 6886 6515
rect 6852 6431 6886 6447
rect 6852 6359 6886 6379
rect 6852 6287 6886 6311
rect 6852 6215 6886 6243
rect 6852 6143 6886 6175
rect 6852 6073 6886 6107
rect 6852 6005 6886 6037
rect 6852 5937 6886 5965
rect 6852 5869 6886 5893
rect 6852 5801 6886 5821
rect 6852 5733 6886 5749
rect 6852 5665 6886 5677
rect 6852 5534 6886 5605
rect 6948 6575 6982 6650
rect 6948 6503 6982 6515
rect 6948 6431 6982 6447
rect 6948 6359 6982 6379
rect 6948 6287 6982 6311
rect 6948 6215 6982 6243
rect 6948 6143 6982 6175
rect 6948 6073 6982 6107
rect 6948 6005 6982 6037
rect 6948 5937 6982 5965
rect 6948 5869 6982 5893
rect 6948 5801 6982 5821
rect 6948 5733 6982 5749
rect 6948 5665 6982 5677
rect 6948 5588 6982 5605
rect 7044 6575 7078 6592
rect 7044 6503 7078 6515
rect 7044 6431 7078 6447
rect 7044 6359 7078 6379
rect 7044 6287 7078 6311
rect 7044 6215 7078 6243
rect 7044 6143 7078 6175
rect 7044 6073 7078 6107
rect 7044 6005 7078 6037
rect 7044 5937 7078 5965
rect 7044 5869 7078 5893
rect 7044 5801 7078 5821
rect 7044 5733 7078 5749
rect 7044 5665 7078 5677
rect 7044 5534 7078 5605
rect 7140 6575 7174 6650
rect 7140 6503 7174 6515
rect 7140 6431 7174 6447
rect 7140 6359 7174 6379
rect 7140 6287 7174 6311
rect 7140 6215 7174 6243
rect 7140 6143 7174 6175
rect 7140 6073 7174 6107
rect 7140 6005 7174 6037
rect 7140 5937 7174 5965
rect 7140 5869 7174 5893
rect 7140 5801 7174 5821
rect 7140 5733 7174 5749
rect 7140 5665 7174 5677
rect 7140 5588 7174 5605
rect 7236 6575 7270 6592
rect 7236 6503 7270 6515
rect 7236 6431 7270 6447
rect 7236 6359 7270 6379
rect 7236 6287 7270 6311
rect 7236 6215 7270 6243
rect 7236 6143 7270 6175
rect 7236 6073 7270 6107
rect 7236 6005 7270 6037
rect 7236 5937 7270 5965
rect 7236 5869 7270 5893
rect 7236 5801 7270 5821
rect 7236 5733 7270 5749
rect 7236 5665 7270 5677
rect 7236 5534 7270 5605
rect 7332 6575 7366 6650
rect 7332 6503 7366 6515
rect 7332 6431 7366 6447
rect 7332 6359 7366 6379
rect 7332 6287 7366 6311
rect 7332 6215 7366 6243
rect 7332 6143 7366 6175
rect 7332 6073 7366 6107
rect 7332 6005 7366 6037
rect 7332 5937 7366 5965
rect 7332 5869 7366 5893
rect 7332 5801 7366 5821
rect 7332 5733 7366 5749
rect 7332 5665 7366 5677
rect 7332 5588 7366 5605
rect 7946 6571 7980 6652
rect 7946 6499 7980 6511
rect 7946 6427 7980 6443
rect 7946 6355 7980 6375
rect 7946 6283 7980 6307
rect 7946 6211 7980 6239
rect 7946 6139 7980 6171
rect 7946 6069 7980 6103
rect 7946 6001 7980 6033
rect 7946 5933 7980 5961
rect 7946 5865 7980 5889
rect 7946 5797 7980 5817
rect 7946 5729 7980 5745
rect 7946 5661 7980 5673
rect 7946 5582 7980 5601
rect 8042 6571 8076 6588
rect 8042 6499 8076 6511
rect 8042 6427 8076 6443
rect 8042 6355 8076 6375
rect 8042 6283 8076 6307
rect 8042 6211 8076 6239
rect 8042 6139 8076 6171
rect 8042 6069 8076 6103
rect 8042 6001 8076 6033
rect 8042 5933 8076 5961
rect 8042 5865 8076 5889
rect 8042 5797 8076 5817
rect 8042 5729 8076 5745
rect 8042 5661 8076 5673
rect 6276 5500 7270 5534
rect 8042 5532 8076 5601
rect 8138 6571 8172 6652
rect 8138 6499 8172 6511
rect 8138 6427 8172 6443
rect 8138 6355 8172 6375
rect 8138 6283 8172 6307
rect 8138 6211 8172 6239
rect 8138 6139 8172 6171
rect 8138 6069 8172 6103
rect 8138 6001 8172 6033
rect 8138 5933 8172 5961
rect 8138 5865 8172 5889
rect 8138 5797 8172 5817
rect 8138 5729 8172 5745
rect 8138 5661 8172 5673
rect 8138 5582 8172 5601
rect 8234 6571 8268 6588
rect 8234 6499 8268 6511
rect 8234 6427 8268 6443
rect 8234 6355 8268 6375
rect 8234 6283 8268 6307
rect 8234 6211 8268 6239
rect 8234 6139 8268 6171
rect 8234 6069 8268 6103
rect 8234 6001 8268 6033
rect 8234 5933 8268 5961
rect 8234 5865 8268 5889
rect 8234 5797 8268 5817
rect 8234 5729 8268 5745
rect 8234 5661 8268 5673
rect 8234 5532 8268 5601
rect 8330 6571 8364 6652
rect 8330 6499 8364 6511
rect 8330 6427 8364 6443
rect 8330 6355 8364 6375
rect 8330 6283 8364 6307
rect 8330 6211 8364 6239
rect 8330 6139 8364 6171
rect 8330 6069 8364 6103
rect 8330 6001 8364 6033
rect 8330 5933 8364 5961
rect 8330 5865 8364 5889
rect 8330 5797 8364 5817
rect 8330 5729 8364 5745
rect 8330 5661 8364 5673
rect 8330 5582 8364 5601
rect 8426 6571 8460 6588
rect 8426 6499 8460 6511
rect 8426 6427 8460 6443
rect 8426 6355 8460 6375
rect 8426 6283 8460 6307
rect 8426 6211 8460 6239
rect 8426 6139 8460 6171
rect 8426 6069 8460 6103
rect 8426 6001 8460 6033
rect 8426 5933 8460 5961
rect 8426 5865 8460 5889
rect 8426 5797 8460 5817
rect 8426 5729 8460 5745
rect 8426 5661 8460 5673
rect 8426 5532 8460 5601
rect 8522 6571 8556 6652
rect 8522 6499 8556 6511
rect 8522 6427 8556 6443
rect 8522 6355 8556 6375
rect 8522 6283 8556 6307
rect 8522 6211 8556 6239
rect 8522 6139 8556 6171
rect 8522 6069 8556 6103
rect 8522 6001 8556 6033
rect 8522 5933 8556 5961
rect 8522 5865 8556 5889
rect 8522 5797 8556 5817
rect 8522 5729 8556 5745
rect 8522 5661 8556 5673
rect 8522 5582 8556 5601
rect 8618 6571 8652 6588
rect 8618 6499 8652 6511
rect 8618 6427 8652 6443
rect 8618 6355 8652 6375
rect 8618 6283 8652 6307
rect 8618 6211 8652 6239
rect 8618 6139 8652 6171
rect 8618 6069 8652 6103
rect 8618 6001 8652 6033
rect 8618 5933 8652 5961
rect 8618 5865 8652 5889
rect 8618 5797 8652 5817
rect 8618 5729 8652 5745
rect 8618 5661 8652 5673
rect 8618 5532 8652 5601
rect 8714 6571 8748 6652
rect 8714 6499 8748 6511
rect 8714 6427 8748 6443
rect 8714 6355 8748 6375
rect 8714 6283 8748 6307
rect 8714 6211 8748 6239
rect 8714 6139 8748 6171
rect 8714 6069 8748 6103
rect 8714 6001 8748 6033
rect 8714 5933 8748 5961
rect 8714 5865 8748 5889
rect 8714 5797 8748 5817
rect 8714 5729 8748 5745
rect 8714 5661 8748 5673
rect 8714 5584 8748 5601
rect 9268 6648 10462 6682
rect 11034 6650 11842 6684
rect 12994 6656 13028 6814
rect 14942 6725 14958 6759
rect 14992 6725 15008 6759
rect 14670 6658 14704 6710
rect 9268 6573 9302 6648
rect 9268 6501 9302 6513
rect 9268 6429 9302 6445
rect 9268 6357 9302 6377
rect 9268 6285 9302 6309
rect 9268 6213 9302 6241
rect 9268 6141 9302 6173
rect 9268 6071 9302 6105
rect 9268 6003 9302 6035
rect 9268 5935 9302 5963
rect 9268 5867 9302 5891
rect 9268 5799 9302 5819
rect 9268 5731 9302 5747
rect 9268 5663 9302 5675
rect 9268 5584 9302 5603
rect 9364 6573 9398 6590
rect 9364 6501 9398 6513
rect 9364 6429 9398 6445
rect 9364 6357 9398 6377
rect 9364 6285 9398 6309
rect 9364 6213 9398 6241
rect 9364 6141 9398 6173
rect 9364 6071 9398 6105
rect 9364 6003 9398 6035
rect 9364 5935 9398 5963
rect 9364 5867 9398 5891
rect 9364 5799 9398 5819
rect 9364 5731 9398 5747
rect 9364 5663 9398 5675
rect 5300 5394 5334 5498
rect 6866 5390 6900 5500
rect 8042 5498 8652 5532
rect 9364 5532 9398 5603
rect 9460 6573 9494 6648
rect 9460 6501 9494 6513
rect 9460 6429 9494 6445
rect 9460 6357 9494 6377
rect 9460 6285 9494 6309
rect 9460 6213 9494 6241
rect 9460 6141 9494 6173
rect 9460 6071 9494 6105
rect 9460 6003 9494 6035
rect 9460 5935 9494 5963
rect 9460 5867 9494 5891
rect 9460 5799 9494 5819
rect 9460 5731 9494 5747
rect 9460 5663 9494 5675
rect 9460 5586 9494 5603
rect 9556 6573 9590 6590
rect 9556 6501 9590 6513
rect 9556 6429 9590 6445
rect 9556 6357 9590 6377
rect 9556 6285 9590 6309
rect 9556 6213 9590 6241
rect 9556 6141 9590 6173
rect 9556 6071 9590 6105
rect 9556 6003 9590 6035
rect 9556 5935 9590 5963
rect 9556 5867 9590 5891
rect 9556 5799 9590 5819
rect 9556 5731 9590 5747
rect 9556 5663 9590 5675
rect 9556 5532 9590 5603
rect 9652 6573 9686 6648
rect 9652 6501 9686 6513
rect 9652 6429 9686 6445
rect 9652 6357 9686 6377
rect 9652 6285 9686 6309
rect 9652 6213 9686 6241
rect 9652 6141 9686 6173
rect 9652 6071 9686 6105
rect 9652 6003 9686 6035
rect 9652 5935 9686 5963
rect 9652 5867 9686 5891
rect 9652 5799 9686 5819
rect 9652 5731 9686 5747
rect 9652 5663 9686 5675
rect 9652 5586 9686 5603
rect 9748 6573 9782 6590
rect 9748 6501 9782 6513
rect 9748 6429 9782 6445
rect 9748 6357 9782 6377
rect 9748 6285 9782 6309
rect 9748 6213 9782 6241
rect 9748 6141 9782 6173
rect 9748 6071 9782 6105
rect 9748 6003 9782 6035
rect 9748 5935 9782 5963
rect 9748 5867 9782 5891
rect 9748 5799 9782 5819
rect 9748 5731 9782 5747
rect 9748 5663 9782 5675
rect 9748 5532 9782 5603
rect 9844 6573 9878 6648
rect 9844 6501 9878 6513
rect 9844 6429 9878 6445
rect 9844 6357 9878 6377
rect 9844 6285 9878 6309
rect 9844 6213 9878 6241
rect 9844 6141 9878 6173
rect 9844 6071 9878 6105
rect 9844 6003 9878 6035
rect 9844 5935 9878 5963
rect 9844 5867 9878 5891
rect 9844 5799 9878 5819
rect 9844 5731 9878 5747
rect 9844 5663 9878 5675
rect 9844 5586 9878 5603
rect 9940 6573 9974 6590
rect 9940 6501 9974 6513
rect 9940 6429 9974 6445
rect 9940 6357 9974 6377
rect 9940 6285 9974 6309
rect 9940 6213 9974 6241
rect 9940 6141 9974 6173
rect 9940 6071 9974 6105
rect 9940 6003 9974 6035
rect 9940 5935 9974 5963
rect 9940 5867 9974 5891
rect 9940 5799 9974 5819
rect 9940 5731 9974 5747
rect 9940 5663 9974 5675
rect 9940 5532 9974 5603
rect 10036 6573 10070 6648
rect 10036 6501 10070 6513
rect 10036 6429 10070 6445
rect 10036 6357 10070 6377
rect 10036 6285 10070 6309
rect 10036 6213 10070 6241
rect 10036 6141 10070 6173
rect 10036 6071 10070 6105
rect 10036 6003 10070 6035
rect 10036 5935 10070 5963
rect 10036 5867 10070 5891
rect 10036 5799 10070 5819
rect 10036 5731 10070 5747
rect 10036 5663 10070 5675
rect 10036 5586 10070 5603
rect 10132 6573 10166 6590
rect 10132 6501 10166 6513
rect 10132 6429 10166 6445
rect 10132 6357 10166 6377
rect 10132 6285 10166 6309
rect 10132 6213 10166 6241
rect 10132 6141 10166 6173
rect 10132 6071 10166 6105
rect 10132 6003 10166 6035
rect 10132 5935 10166 5963
rect 10132 5867 10166 5891
rect 10132 5799 10166 5819
rect 10132 5731 10166 5747
rect 10132 5663 10166 5675
rect 10132 5532 10166 5603
rect 10228 6573 10262 6648
rect 10228 6501 10262 6513
rect 10228 6429 10262 6445
rect 10228 6357 10262 6377
rect 10228 6285 10262 6309
rect 10228 6213 10262 6241
rect 10228 6141 10262 6173
rect 10228 6071 10262 6105
rect 10228 6003 10262 6035
rect 10228 5935 10262 5963
rect 10228 5867 10262 5891
rect 10228 5799 10262 5819
rect 10228 5731 10262 5747
rect 10228 5663 10262 5675
rect 10228 5586 10262 5603
rect 10324 6573 10358 6590
rect 10324 6501 10358 6513
rect 10324 6429 10358 6445
rect 10324 6357 10358 6377
rect 10324 6285 10358 6309
rect 10324 6213 10358 6241
rect 10324 6141 10358 6173
rect 10324 6071 10358 6105
rect 10324 6003 10358 6035
rect 10324 5935 10358 5963
rect 10324 5867 10358 5891
rect 10324 5799 10358 5819
rect 10324 5731 10358 5747
rect 10324 5663 10358 5675
rect 10324 5532 10358 5603
rect 10420 6573 10454 6648
rect 10420 6501 10454 6513
rect 10420 6429 10454 6445
rect 10420 6357 10454 6377
rect 10420 6285 10454 6309
rect 10420 6213 10454 6241
rect 10420 6141 10454 6173
rect 10420 6071 10454 6105
rect 10420 6003 10454 6035
rect 10420 5935 10454 5963
rect 10420 5867 10454 5891
rect 10420 5799 10454 5819
rect 10420 5731 10454 5747
rect 10420 5663 10454 5675
rect 10420 5586 10454 5603
rect 11034 6569 11068 6650
rect 11034 6497 11068 6509
rect 11034 6425 11068 6441
rect 11034 6353 11068 6373
rect 11034 6281 11068 6305
rect 11034 6209 11068 6237
rect 11034 6137 11068 6169
rect 11034 6067 11068 6101
rect 11034 5999 11068 6031
rect 11034 5931 11068 5959
rect 11034 5863 11068 5887
rect 11034 5795 11068 5815
rect 11034 5727 11068 5743
rect 11034 5659 11068 5671
rect 11034 5580 11068 5599
rect 11130 6569 11164 6586
rect 11130 6497 11164 6509
rect 11130 6425 11164 6441
rect 11130 6353 11164 6373
rect 11130 6281 11164 6305
rect 11130 6209 11164 6237
rect 11130 6137 11164 6169
rect 11130 6067 11164 6101
rect 11130 5999 11164 6031
rect 11130 5931 11164 5959
rect 11130 5863 11164 5887
rect 11130 5795 11164 5815
rect 11130 5727 11164 5743
rect 11130 5659 11164 5671
rect 9364 5498 10358 5532
rect 11130 5530 11164 5599
rect 11226 6569 11260 6650
rect 11226 6497 11260 6509
rect 11226 6425 11260 6441
rect 11226 6353 11260 6373
rect 11226 6281 11260 6305
rect 11226 6209 11260 6237
rect 11226 6137 11260 6169
rect 11226 6067 11260 6101
rect 11226 5999 11260 6031
rect 11226 5931 11260 5959
rect 11226 5863 11260 5887
rect 11226 5795 11260 5815
rect 11226 5727 11260 5743
rect 11226 5659 11260 5671
rect 11226 5580 11260 5599
rect 11322 6569 11356 6586
rect 11322 6497 11356 6509
rect 11322 6425 11356 6441
rect 11322 6353 11356 6373
rect 11322 6281 11356 6305
rect 11322 6209 11356 6237
rect 11322 6137 11356 6169
rect 11322 6067 11356 6101
rect 11322 5999 11356 6031
rect 11322 5931 11356 5959
rect 11322 5863 11356 5887
rect 11322 5795 11356 5815
rect 11322 5727 11356 5743
rect 11322 5659 11356 5671
rect 11322 5530 11356 5599
rect 11418 6569 11452 6650
rect 11418 6497 11452 6509
rect 11418 6425 11452 6441
rect 11418 6353 11452 6373
rect 11418 6281 11452 6305
rect 11418 6209 11452 6237
rect 11418 6137 11452 6169
rect 11418 6067 11452 6101
rect 11418 5999 11452 6031
rect 11418 5931 11452 5959
rect 11418 5863 11452 5887
rect 11418 5795 11452 5815
rect 11418 5727 11452 5743
rect 11418 5659 11452 5671
rect 11418 5580 11452 5599
rect 11514 6569 11548 6586
rect 11514 6497 11548 6509
rect 11514 6425 11548 6441
rect 11514 6353 11548 6373
rect 11514 6281 11548 6305
rect 11514 6209 11548 6237
rect 11514 6137 11548 6169
rect 11514 6067 11548 6101
rect 11514 5999 11548 6031
rect 11514 5931 11548 5959
rect 11514 5863 11548 5887
rect 11514 5795 11548 5815
rect 11514 5727 11548 5743
rect 11514 5659 11548 5671
rect 11514 5530 11548 5599
rect 11610 6569 11644 6650
rect 11610 6497 11644 6509
rect 11610 6425 11644 6441
rect 11610 6353 11644 6373
rect 11610 6281 11644 6305
rect 11610 6209 11644 6237
rect 11610 6137 11644 6169
rect 11610 6067 11644 6101
rect 11610 5999 11644 6031
rect 11610 5931 11644 5959
rect 11610 5863 11644 5887
rect 11610 5795 11644 5815
rect 11610 5727 11644 5743
rect 11610 5659 11644 5671
rect 11610 5580 11644 5599
rect 11706 6569 11740 6586
rect 11706 6497 11740 6509
rect 11706 6425 11740 6441
rect 11706 6353 11740 6373
rect 11706 6281 11740 6305
rect 11706 6209 11740 6237
rect 11706 6137 11740 6169
rect 11706 6067 11740 6101
rect 11706 5999 11740 6031
rect 11706 5931 11740 5959
rect 11706 5863 11740 5887
rect 11706 5795 11740 5815
rect 11706 5727 11740 5743
rect 11706 5659 11740 5671
rect 11706 5530 11740 5599
rect 11802 6569 11836 6650
rect 11802 6497 11836 6509
rect 11802 6425 11836 6441
rect 11802 6353 11836 6373
rect 11802 6281 11836 6305
rect 11802 6209 11836 6237
rect 11802 6137 11836 6169
rect 11802 6067 11836 6101
rect 11802 5999 11836 6031
rect 11802 5931 11836 5959
rect 11802 5863 11836 5887
rect 11802 5795 11836 5815
rect 11802 5727 11836 5743
rect 11802 5659 11836 5671
rect 11802 5582 11836 5599
rect 12424 6622 13618 6656
rect 14190 6624 14998 6658
rect 12424 6547 12458 6622
rect 12424 6475 12458 6487
rect 12424 6403 12458 6419
rect 12424 6331 12458 6351
rect 12424 6259 12458 6283
rect 12424 6187 12458 6215
rect 12424 6115 12458 6147
rect 12424 6045 12458 6079
rect 12424 5977 12458 6009
rect 12424 5909 12458 5937
rect 12424 5841 12458 5865
rect 12424 5773 12458 5793
rect 12424 5705 12458 5721
rect 12424 5637 12458 5649
rect 12424 5558 12458 5577
rect 12520 6547 12554 6564
rect 12520 6475 12554 6487
rect 12520 6403 12554 6419
rect 12520 6331 12554 6351
rect 12520 6259 12554 6283
rect 12520 6187 12554 6215
rect 12520 6115 12554 6147
rect 12520 6045 12554 6079
rect 12520 5977 12554 6009
rect 12520 5909 12554 5937
rect 12520 5841 12554 5865
rect 12520 5773 12554 5793
rect 12520 5705 12554 5721
rect 12520 5637 12554 5649
rect 8330 5394 8364 5498
rect 9954 5388 9988 5498
rect 11130 5496 11740 5530
rect 12520 5506 12554 5577
rect 12616 6547 12650 6622
rect 12616 6475 12650 6487
rect 12616 6403 12650 6419
rect 12616 6331 12650 6351
rect 12616 6259 12650 6283
rect 12616 6187 12650 6215
rect 12616 6115 12650 6147
rect 12616 6045 12650 6079
rect 12616 5977 12650 6009
rect 12616 5909 12650 5937
rect 12616 5841 12650 5865
rect 12616 5773 12650 5793
rect 12616 5705 12650 5721
rect 12616 5637 12650 5649
rect 12616 5560 12650 5577
rect 12712 6547 12746 6564
rect 12712 6475 12746 6487
rect 12712 6403 12746 6419
rect 12712 6331 12746 6351
rect 12712 6259 12746 6283
rect 12712 6187 12746 6215
rect 12712 6115 12746 6147
rect 12712 6045 12746 6079
rect 12712 5977 12746 6009
rect 12712 5909 12746 5937
rect 12712 5841 12746 5865
rect 12712 5773 12746 5793
rect 12712 5705 12746 5721
rect 12712 5637 12746 5649
rect 12712 5506 12746 5577
rect 12808 6547 12842 6622
rect 12808 6475 12842 6487
rect 12808 6403 12842 6419
rect 12808 6331 12842 6351
rect 12808 6259 12842 6283
rect 12808 6187 12842 6215
rect 12808 6115 12842 6147
rect 12808 6045 12842 6079
rect 12808 5977 12842 6009
rect 12808 5909 12842 5937
rect 12808 5841 12842 5865
rect 12808 5773 12842 5793
rect 12808 5705 12842 5721
rect 12808 5637 12842 5649
rect 12808 5560 12842 5577
rect 12904 6547 12938 6564
rect 12904 6475 12938 6487
rect 12904 6403 12938 6419
rect 12904 6331 12938 6351
rect 12904 6259 12938 6283
rect 12904 6187 12938 6215
rect 12904 6115 12938 6147
rect 12904 6045 12938 6079
rect 12904 5977 12938 6009
rect 12904 5909 12938 5937
rect 12904 5841 12938 5865
rect 12904 5773 12938 5793
rect 12904 5705 12938 5721
rect 12904 5637 12938 5649
rect 12904 5506 12938 5577
rect 13000 6547 13034 6622
rect 13000 6475 13034 6487
rect 13000 6403 13034 6419
rect 13000 6331 13034 6351
rect 13000 6259 13034 6283
rect 13000 6187 13034 6215
rect 13000 6115 13034 6147
rect 13000 6045 13034 6079
rect 13000 5977 13034 6009
rect 13000 5909 13034 5937
rect 13000 5841 13034 5865
rect 13000 5773 13034 5793
rect 13000 5705 13034 5721
rect 13000 5637 13034 5649
rect 13000 5560 13034 5577
rect 13096 6547 13130 6564
rect 13096 6475 13130 6487
rect 13096 6403 13130 6419
rect 13096 6331 13130 6351
rect 13096 6259 13130 6283
rect 13096 6187 13130 6215
rect 13096 6115 13130 6147
rect 13096 6045 13130 6079
rect 13096 5977 13130 6009
rect 13096 5909 13130 5937
rect 13096 5841 13130 5865
rect 13096 5773 13130 5793
rect 13096 5705 13130 5721
rect 13096 5637 13130 5649
rect 13096 5506 13130 5577
rect 13192 6547 13226 6622
rect 13192 6475 13226 6487
rect 13192 6403 13226 6419
rect 13192 6331 13226 6351
rect 13192 6259 13226 6283
rect 13192 6187 13226 6215
rect 13192 6115 13226 6147
rect 13192 6045 13226 6079
rect 13192 5977 13226 6009
rect 13192 5909 13226 5937
rect 13192 5841 13226 5865
rect 13192 5773 13226 5793
rect 13192 5705 13226 5721
rect 13192 5637 13226 5649
rect 13192 5560 13226 5577
rect 13288 6547 13322 6564
rect 13288 6475 13322 6487
rect 13288 6403 13322 6419
rect 13288 6331 13322 6351
rect 13288 6259 13322 6283
rect 13288 6187 13322 6215
rect 13288 6115 13322 6147
rect 13288 6045 13322 6079
rect 13288 5977 13322 6009
rect 13288 5909 13322 5937
rect 13288 5841 13322 5865
rect 13288 5773 13322 5793
rect 13288 5705 13322 5721
rect 13288 5637 13322 5649
rect 13288 5506 13322 5577
rect 13384 6547 13418 6622
rect 13384 6475 13418 6487
rect 13384 6403 13418 6419
rect 13384 6331 13418 6351
rect 13384 6259 13418 6283
rect 13384 6187 13418 6215
rect 13384 6115 13418 6147
rect 13384 6045 13418 6079
rect 13384 5977 13418 6009
rect 13384 5909 13418 5937
rect 13384 5841 13418 5865
rect 13384 5773 13418 5793
rect 13384 5705 13418 5721
rect 13384 5637 13418 5649
rect 13384 5560 13418 5577
rect 13480 6547 13514 6564
rect 13480 6475 13514 6487
rect 13480 6403 13514 6419
rect 13480 6331 13514 6351
rect 13480 6259 13514 6283
rect 13480 6187 13514 6215
rect 13480 6115 13514 6147
rect 13480 6045 13514 6079
rect 13480 5977 13514 6009
rect 13480 5909 13514 5937
rect 13480 5841 13514 5865
rect 13480 5773 13514 5793
rect 13480 5705 13514 5721
rect 13480 5637 13514 5649
rect 13480 5506 13514 5577
rect 13576 6547 13610 6622
rect 13576 6475 13610 6487
rect 13576 6403 13610 6419
rect 13576 6331 13610 6351
rect 13576 6259 13610 6283
rect 13576 6187 13610 6215
rect 13576 6115 13610 6147
rect 13576 6045 13610 6079
rect 13576 5977 13610 6009
rect 13576 5909 13610 5937
rect 13576 5841 13610 5865
rect 13576 5773 13610 5793
rect 13576 5705 13610 5721
rect 13576 5637 13610 5649
rect 13576 5560 13610 5577
rect 14190 6543 14224 6624
rect 14190 6471 14224 6483
rect 14190 6399 14224 6415
rect 14190 6327 14224 6347
rect 14190 6255 14224 6279
rect 14190 6183 14224 6211
rect 14190 6111 14224 6143
rect 14190 6041 14224 6075
rect 14190 5973 14224 6005
rect 14190 5905 14224 5933
rect 14190 5837 14224 5861
rect 14190 5769 14224 5789
rect 14190 5701 14224 5717
rect 14190 5633 14224 5645
rect 14190 5554 14224 5573
rect 14286 6543 14320 6560
rect 14286 6471 14320 6483
rect 14286 6399 14320 6415
rect 14286 6327 14320 6347
rect 14286 6255 14320 6279
rect 14286 6183 14320 6211
rect 14286 6111 14320 6143
rect 14286 6041 14320 6075
rect 14286 5973 14320 6005
rect 14286 5905 14320 5933
rect 14286 5837 14320 5861
rect 14286 5769 14320 5789
rect 14286 5701 14320 5717
rect 14286 5633 14320 5645
rect 11418 5392 11452 5496
rect 12520 5472 13514 5506
rect 14286 5504 14320 5573
rect 14382 6543 14416 6624
rect 14382 6471 14416 6483
rect 14382 6399 14416 6415
rect 14382 6327 14416 6347
rect 14382 6255 14416 6279
rect 14382 6183 14416 6211
rect 14382 6111 14416 6143
rect 14382 6041 14416 6075
rect 14382 5973 14416 6005
rect 14382 5905 14416 5933
rect 14382 5837 14416 5861
rect 14382 5769 14416 5789
rect 14382 5701 14416 5717
rect 14382 5633 14416 5645
rect 14382 5554 14416 5573
rect 14478 6543 14512 6560
rect 14478 6471 14512 6483
rect 14478 6399 14512 6415
rect 14478 6327 14512 6347
rect 14478 6255 14512 6279
rect 14478 6183 14512 6211
rect 14478 6111 14512 6143
rect 14478 6041 14512 6075
rect 14478 5973 14512 6005
rect 14478 5905 14512 5933
rect 14478 5837 14512 5861
rect 14478 5769 14512 5789
rect 14478 5701 14512 5717
rect 14478 5633 14512 5645
rect 14478 5504 14512 5573
rect 14574 6543 14608 6624
rect 14574 6471 14608 6483
rect 14574 6399 14608 6415
rect 14574 6327 14608 6347
rect 14574 6255 14608 6279
rect 14574 6183 14608 6211
rect 14574 6111 14608 6143
rect 14574 6041 14608 6075
rect 14574 5973 14608 6005
rect 14574 5905 14608 5933
rect 14574 5837 14608 5861
rect 14574 5769 14608 5789
rect 14574 5701 14608 5717
rect 14574 5633 14608 5645
rect 14574 5554 14608 5573
rect 14670 6543 14704 6560
rect 14670 6471 14704 6483
rect 14670 6399 14704 6415
rect 14670 6327 14704 6347
rect 14670 6255 14704 6279
rect 14670 6183 14704 6211
rect 14670 6111 14704 6143
rect 14670 6041 14704 6075
rect 14670 5973 14704 6005
rect 14670 5905 14704 5933
rect 14670 5837 14704 5861
rect 14670 5769 14704 5789
rect 14670 5701 14704 5717
rect 14670 5633 14704 5645
rect 14670 5504 14704 5573
rect 14766 6543 14800 6624
rect 14766 6471 14800 6483
rect 14766 6399 14800 6415
rect 14766 6327 14800 6347
rect 14766 6255 14800 6279
rect 14766 6183 14800 6211
rect 14766 6111 14800 6143
rect 14766 6041 14800 6075
rect 14766 5973 14800 6005
rect 14766 5905 14800 5933
rect 14766 5837 14800 5861
rect 14766 5769 14800 5789
rect 14766 5701 14800 5717
rect 14766 5633 14800 5645
rect 14766 5554 14800 5573
rect 14862 6543 14896 6560
rect 14862 6471 14896 6483
rect 14862 6399 14896 6415
rect 14862 6327 14896 6347
rect 14862 6255 14896 6279
rect 14862 6183 14896 6211
rect 14862 6111 14896 6143
rect 14862 6041 14896 6075
rect 14862 5973 14896 6005
rect 14862 5905 14896 5933
rect 14862 5837 14896 5861
rect 14862 5769 14896 5789
rect 14862 5701 14896 5717
rect 14862 5633 14896 5645
rect 14862 5504 14896 5573
rect 14958 6543 14992 6624
rect 14958 6471 14992 6483
rect 14958 6399 14992 6415
rect 14958 6327 14992 6347
rect 14958 6255 14992 6279
rect 14958 6183 14992 6211
rect 14958 6111 14992 6143
rect 14958 6041 14992 6075
rect 15614 6032 15648 6148
rect 14958 5973 14992 6005
rect 14958 5905 14992 5933
rect 14958 5837 14992 5861
rect 14958 5769 14992 5789
rect 14958 5701 14992 5717
rect 14958 5633 14992 5645
rect 14958 5556 14992 5573
rect 15518 5996 15744 6032
rect 15518 5895 15552 5996
rect 15518 5827 15552 5845
rect 15518 5759 15552 5773
rect 15518 5691 15552 5701
rect 15518 5623 15552 5629
rect 13110 5362 13144 5472
rect 14286 5470 14896 5504
rect 15518 5555 15552 5557
rect 15518 5519 15552 5521
rect 14574 5366 14608 5470
rect 15518 5447 15552 5453
rect 15518 5375 15552 5385
rect -868 5283 -834 5311
rect -868 5215 -834 5239
rect -868 5147 -834 5167
rect 15518 5303 15552 5317
rect 15518 5231 15552 5249
rect 15518 5159 15552 5181
rect -868 5079 -834 5095
rect 1580 5028 1614 5090
rect -868 5011 -834 5023
rect 1482 4994 1908 5028
rect 4536 5012 4570 5074
rect 7566 5012 7600 5074
rect 15518 5087 15552 5113
rect -868 4934 -834 4951
rect -1554 4842 -932 4876
rect 1484 4929 1518 4994
rect 1484 4857 1518 4869
rect -1162 4840 -1124 4842
rect -1158 4768 -1124 4840
rect 1484 4785 1518 4801
rect -1083 4768 -1067 4769
rect -1158 4735 -1067 4768
rect -1033 4735 -1017 4769
rect -1158 4734 -1068 4735
rect 1484 4713 1518 4733
rect 1484 4641 1518 4665
rect 1484 4569 1518 4597
rect 1484 4497 1518 4529
rect 1484 4427 1518 4461
rect 1484 4359 1518 4391
rect 1484 4291 1518 4319
rect 1484 4223 1518 4247
rect 1484 4155 1518 4175
rect 1484 4087 1518 4103
rect 1484 4019 1518 4031
rect 1484 3940 1518 3959
rect 1580 4929 1614 4946
rect 1580 4857 1614 4869
rect 1580 4785 1614 4801
rect 1580 4713 1614 4733
rect 1580 4641 1614 4665
rect 1580 4569 1614 4597
rect 1580 4497 1614 4529
rect 1580 4427 1614 4461
rect 1580 4359 1614 4391
rect 1580 4291 1614 4319
rect 1580 4223 1614 4247
rect 1580 4155 1614 4175
rect 1580 4087 1614 4103
rect 1580 4019 1614 4031
rect 1580 3884 1614 3959
rect 1676 4929 1710 4994
rect 1676 4857 1710 4869
rect 1676 4785 1710 4801
rect 1676 4713 1710 4733
rect 1676 4641 1710 4665
rect 1676 4569 1710 4597
rect 1676 4497 1710 4529
rect 1676 4427 1710 4461
rect 1676 4359 1710 4391
rect 1676 4291 1710 4319
rect 1676 4223 1710 4247
rect 1676 4155 1710 4175
rect 1676 4087 1710 4103
rect 1676 4019 1710 4031
rect 1676 3940 1710 3959
rect 1772 4929 1806 4946
rect 1772 4857 1806 4869
rect 1772 4785 1806 4801
rect 1772 4713 1806 4733
rect 1772 4641 1806 4665
rect 1772 4569 1806 4597
rect 1772 4497 1806 4529
rect 1772 4427 1806 4461
rect 1772 4359 1806 4391
rect 1772 4291 1806 4319
rect 1772 4223 1806 4247
rect 1772 4155 1806 4175
rect 1772 4087 1806 4103
rect 1772 4019 1806 4031
rect 1676 3884 1710 3886
rect 1772 3884 1806 3959
rect 1868 4929 1902 4994
rect 4438 4978 4864 5012
rect 7468 4978 7894 5012
rect 10654 5010 10688 5072
rect 1868 4857 1902 4869
rect 1868 4785 1902 4801
rect 1868 4713 1902 4733
rect 1868 4641 1902 4665
rect 1868 4569 1902 4597
rect 1868 4497 1902 4529
rect 1868 4427 1902 4461
rect 1868 4359 1902 4391
rect 1868 4291 1902 4319
rect 1868 4223 1902 4247
rect 1868 4155 1902 4175
rect 1868 4087 1902 4103
rect 1868 4019 1902 4031
rect 1868 3940 1902 3959
rect 4440 4913 4474 4978
rect 4440 4841 4474 4853
rect 4440 4769 4474 4785
rect 4440 4697 4474 4717
rect 4440 4625 4474 4649
rect 4440 4553 4474 4581
rect 4440 4481 4474 4513
rect 4440 4411 4474 4445
rect 4440 4343 4474 4375
rect 4440 4275 4474 4303
rect 4440 4207 4474 4231
rect 4440 4139 4474 4159
rect 4440 4071 4474 4087
rect 4440 4003 4474 4015
rect 4440 3924 4474 3943
rect 4536 4913 4570 4930
rect 4536 4841 4570 4853
rect 4536 4769 4570 4785
rect 4536 4697 4570 4717
rect 4536 4625 4570 4649
rect 4536 4553 4570 4581
rect 4536 4481 4570 4513
rect 4536 4411 4570 4445
rect 4536 4343 4570 4375
rect 4536 4275 4570 4303
rect 4536 4207 4570 4231
rect 4536 4139 4570 4159
rect 4536 4071 4570 4087
rect 4536 4003 4570 4015
rect 1580 3850 1806 3884
rect 4536 3868 4570 3943
rect 4632 4913 4666 4978
rect 4632 4841 4666 4853
rect 4632 4769 4666 4785
rect 4632 4697 4666 4717
rect 4632 4625 4666 4649
rect 4632 4553 4666 4581
rect 4632 4481 4666 4513
rect 4632 4411 4666 4445
rect 4632 4343 4666 4375
rect 4632 4275 4666 4303
rect 4632 4207 4666 4231
rect 4632 4139 4666 4159
rect 4632 4071 4666 4087
rect 4632 4003 4666 4015
rect 4632 3924 4666 3943
rect 4728 4913 4762 4930
rect 4728 4841 4762 4853
rect 4728 4769 4762 4785
rect 4728 4697 4762 4717
rect 4728 4625 4762 4649
rect 4728 4553 4762 4581
rect 4728 4481 4762 4513
rect 4728 4411 4762 4445
rect 4728 4343 4762 4375
rect 4728 4275 4762 4303
rect 4728 4207 4762 4231
rect 4728 4139 4762 4159
rect 4728 4071 4762 4087
rect 4728 4003 4762 4015
rect 4632 3868 4666 3870
rect 4728 3868 4762 3943
rect 4824 4913 4858 4978
rect 4824 4841 4858 4853
rect 4824 4769 4858 4785
rect 4824 4697 4858 4717
rect 4824 4625 4858 4649
rect 4824 4553 4858 4581
rect 4824 4481 4858 4513
rect 4824 4411 4858 4445
rect 4824 4343 4858 4375
rect 4824 4275 4858 4303
rect 4824 4207 4858 4231
rect 4824 4139 4858 4159
rect 4824 4071 4858 4087
rect 4824 4003 4858 4015
rect 4824 3924 4858 3943
rect 7470 4913 7504 4978
rect 7470 4841 7504 4853
rect 7470 4769 7504 4785
rect 7470 4697 7504 4717
rect 7470 4625 7504 4649
rect 7470 4553 7504 4581
rect 7470 4481 7504 4513
rect 7470 4411 7504 4445
rect 7470 4343 7504 4375
rect 7470 4275 7504 4303
rect 7470 4207 7504 4231
rect 7470 4139 7504 4159
rect 7470 4071 7504 4087
rect 7470 4003 7504 4015
rect 7470 3924 7504 3943
rect 7566 4913 7600 4930
rect 7566 4841 7600 4853
rect 7566 4769 7600 4785
rect 7566 4697 7600 4717
rect 7566 4625 7600 4649
rect 7566 4553 7600 4581
rect 7566 4481 7600 4513
rect 7566 4411 7600 4445
rect 7566 4343 7600 4375
rect 7566 4275 7600 4303
rect 7566 4207 7600 4231
rect 7566 4139 7600 4159
rect 7566 4071 7600 4087
rect 7566 4003 7600 4015
rect 1564 3743 1580 3777
rect 1614 3743 1630 3777
rect 1676 3754 1710 3850
rect 4536 3834 4762 3868
rect 7566 3868 7600 3943
rect 7662 4913 7696 4978
rect 7662 4841 7696 4853
rect 7662 4769 7696 4785
rect 7662 4697 7696 4717
rect 7662 4625 7696 4649
rect 7662 4553 7696 4581
rect 7662 4481 7696 4513
rect 7662 4411 7696 4445
rect 7662 4343 7696 4375
rect 7662 4275 7696 4303
rect 7662 4207 7696 4231
rect 7662 4139 7696 4159
rect 7662 4071 7696 4087
rect 7662 4003 7696 4015
rect 7662 3924 7696 3943
rect 7758 4913 7792 4930
rect 7758 4841 7792 4853
rect 7758 4769 7792 4785
rect 7758 4697 7792 4717
rect 7758 4625 7792 4649
rect 7758 4553 7792 4581
rect 7758 4481 7792 4513
rect 7758 4411 7792 4445
rect 7758 4343 7792 4375
rect 7758 4275 7792 4303
rect 7758 4207 7792 4231
rect 7758 4139 7792 4159
rect 7758 4071 7792 4087
rect 7758 4003 7792 4015
rect 7662 3868 7696 3870
rect 7758 3868 7792 3943
rect 7854 4913 7888 4978
rect 10556 4976 10982 5010
rect 13810 4984 13844 5046
rect 15518 5015 15552 5045
rect 7854 4841 7888 4853
rect 7854 4769 7888 4785
rect 7854 4697 7888 4717
rect 7854 4625 7888 4649
rect 7854 4553 7888 4581
rect 7854 4481 7888 4513
rect 7854 4411 7888 4445
rect 7854 4343 7888 4375
rect 7854 4275 7888 4303
rect 7854 4207 7888 4231
rect 7854 4139 7888 4159
rect 7854 4071 7888 4087
rect 7854 4003 7888 4015
rect 7854 3924 7888 3943
rect 10558 4911 10592 4976
rect 10558 4839 10592 4851
rect 10558 4767 10592 4783
rect 10558 4695 10592 4715
rect 10558 4623 10592 4647
rect 10558 4551 10592 4579
rect 10558 4479 10592 4511
rect 10558 4409 10592 4443
rect 10558 4341 10592 4373
rect 10558 4273 10592 4301
rect 10558 4205 10592 4229
rect 10558 4137 10592 4157
rect 10558 4069 10592 4085
rect 10558 4001 10592 4013
rect 10558 3922 10592 3941
rect 10654 4911 10688 4928
rect 10654 4839 10688 4851
rect 10654 4767 10688 4783
rect 10654 4695 10688 4715
rect 10654 4623 10688 4647
rect 10654 4551 10688 4579
rect 10654 4479 10688 4511
rect 10654 4409 10688 4443
rect 10654 4341 10688 4373
rect 10654 4273 10688 4301
rect 10654 4205 10688 4229
rect 10654 4137 10688 4157
rect 10654 4069 10688 4085
rect 10654 4001 10688 4013
rect 7566 3834 7792 3868
rect 10654 3866 10688 3941
rect 10750 4911 10784 4976
rect 10750 4839 10784 4851
rect 10750 4767 10784 4783
rect 10750 4695 10784 4715
rect 10750 4623 10784 4647
rect 10750 4551 10784 4579
rect 10750 4479 10784 4511
rect 10750 4409 10784 4443
rect 10750 4341 10784 4373
rect 10750 4273 10784 4301
rect 10750 4205 10784 4229
rect 10750 4137 10784 4157
rect 10750 4069 10784 4085
rect 10750 4001 10784 4013
rect 10750 3922 10784 3941
rect 10846 4911 10880 4928
rect 10846 4839 10880 4851
rect 10846 4767 10880 4783
rect 10846 4695 10880 4715
rect 10846 4623 10880 4647
rect 10846 4551 10880 4579
rect 10846 4479 10880 4511
rect 10846 4409 10880 4443
rect 10846 4341 10880 4373
rect 10846 4273 10880 4301
rect 10846 4205 10880 4229
rect 10846 4137 10880 4157
rect 10846 4069 10880 4085
rect 10846 4001 10880 4013
rect 10750 3866 10784 3868
rect 10846 3866 10880 3941
rect 10942 4911 10976 4976
rect 13712 4950 14138 4984
rect 10942 4839 10976 4851
rect 10942 4767 10976 4783
rect 10942 4695 10976 4715
rect 10942 4623 10976 4647
rect 10942 4551 10976 4579
rect 10942 4479 10976 4511
rect 10942 4409 10976 4443
rect 10942 4341 10976 4373
rect 10942 4273 10976 4301
rect 10942 4205 10976 4229
rect 10942 4137 10976 4157
rect 10942 4069 10976 4085
rect 10942 4001 10976 4013
rect 10942 3922 10976 3941
rect 13714 4885 13748 4950
rect 13714 4813 13748 4825
rect 13714 4741 13748 4757
rect 13714 4669 13748 4689
rect 13714 4597 13748 4621
rect 13714 4525 13748 4553
rect 13714 4453 13748 4485
rect 13714 4383 13748 4417
rect 13714 4315 13748 4347
rect 13714 4247 13748 4275
rect 13714 4179 13748 4203
rect 13714 4111 13748 4131
rect 13714 4043 13748 4059
rect 13714 3975 13748 3987
rect 13714 3896 13748 3915
rect 13810 4885 13844 4902
rect 13810 4813 13844 4825
rect 13810 4741 13844 4757
rect 13810 4669 13844 4689
rect 13810 4597 13844 4621
rect 13810 4525 13844 4553
rect 13810 4453 13844 4485
rect 13810 4383 13844 4417
rect 13810 4315 13844 4347
rect 13810 4247 13844 4275
rect 13810 4179 13844 4203
rect 13810 4111 13844 4131
rect 13810 4043 13844 4059
rect 13810 3975 13844 3987
rect 1756 3743 1772 3777
rect 1806 3743 1822 3777
rect 4520 3727 4536 3761
rect 4570 3727 4586 3761
rect 4632 3738 4666 3834
rect 4712 3727 4728 3761
rect 4762 3727 4778 3761
rect 7550 3727 7566 3761
rect 7600 3727 7616 3761
rect 7662 3738 7696 3834
rect 10654 3832 10880 3866
rect 13810 3840 13844 3915
rect 13906 4885 13940 4950
rect 13906 4813 13940 4825
rect 13906 4741 13940 4757
rect 13906 4669 13940 4689
rect 13906 4597 13940 4621
rect 13906 4525 13940 4553
rect 13906 4453 13940 4485
rect 13906 4383 13940 4417
rect 13906 4315 13940 4347
rect 13906 4247 13940 4275
rect 13906 4179 13940 4203
rect 13906 4111 13940 4131
rect 13906 4043 13940 4059
rect 13906 3975 13940 3987
rect 13906 3896 13940 3915
rect 14002 4885 14036 4902
rect 14002 4813 14036 4825
rect 14002 4741 14036 4757
rect 14002 4669 14036 4689
rect 14002 4597 14036 4621
rect 14002 4525 14036 4553
rect 14002 4453 14036 4485
rect 14002 4383 14036 4417
rect 14002 4315 14036 4347
rect 14002 4247 14036 4275
rect 14002 4179 14036 4203
rect 14002 4111 14036 4131
rect 14002 4043 14036 4059
rect 14002 3975 14036 3987
rect 13906 3840 13940 3842
rect 14002 3840 14036 3915
rect 14098 4885 14132 4950
rect 14098 4813 14132 4825
rect 14098 4741 14132 4757
rect 14098 4669 14132 4689
rect 14098 4597 14132 4621
rect 14098 4525 14132 4553
rect 14098 4453 14132 4485
rect 14098 4383 14132 4417
rect 14098 4315 14132 4347
rect 14098 4247 14132 4275
rect 14098 4179 14132 4203
rect 14098 4111 14132 4131
rect 14098 4043 14132 4059
rect 14098 3975 14132 3987
rect 15518 4943 15552 4977
rect 15518 4875 15552 4909
rect 15518 4807 15552 4837
rect 15518 4739 15552 4765
rect 15518 4671 15552 4693
rect 15518 4603 15552 4621
rect 15518 4535 15552 4549
rect 15518 4467 15552 4477
rect 15518 4399 15552 4405
rect 15518 4331 15552 4333
rect 15518 4295 15552 4297
rect 15518 4223 15552 4229
rect 15518 4151 15552 4161
rect 15518 4079 15552 4093
rect 15518 4007 15552 4025
rect 15518 3918 15552 3957
rect 15614 5895 15648 5930
rect 15614 5827 15648 5845
rect 15614 5759 15648 5773
rect 15614 5691 15648 5701
rect 15614 5623 15648 5629
rect 15614 5555 15648 5557
rect 15614 5519 15648 5521
rect 15614 5447 15648 5453
rect 15614 5375 15648 5385
rect 15614 5303 15648 5317
rect 15614 5231 15648 5249
rect 15614 5159 15648 5181
rect 15614 5087 15648 5113
rect 15614 5015 15648 5045
rect 15614 4943 15648 4977
rect 15614 4875 15648 4909
rect 15614 4807 15648 4837
rect 15614 4739 15648 4765
rect 15614 4671 15648 4693
rect 15614 4603 15648 4621
rect 15614 4535 15648 4549
rect 15614 4467 15648 4477
rect 15614 4399 15648 4405
rect 15614 4331 15648 4333
rect 15614 4295 15648 4297
rect 15614 4223 15648 4229
rect 15614 4151 15648 4161
rect 15614 4079 15648 4093
rect 15614 4007 15648 4025
rect 14098 3896 14132 3915
rect 15614 3884 15648 3957
rect 15710 5895 15744 5996
rect 15710 5827 15744 5845
rect 15710 5759 15744 5773
rect 15710 5691 15744 5701
rect 15710 5623 15744 5629
rect 15710 5555 15744 5557
rect 15710 5519 15744 5521
rect 15710 5447 15744 5453
rect 15710 5375 15744 5385
rect 15710 5303 15744 5317
rect 15710 5231 15744 5249
rect 15710 5159 15744 5181
rect 15710 5087 15744 5113
rect 15710 5015 15744 5045
rect 15710 4943 15744 4977
rect 15710 4875 15744 4909
rect 15710 4807 15744 4837
rect 15710 4739 15744 4765
rect 15710 4671 15744 4693
rect 15710 4603 15744 4621
rect 15710 4535 15744 4549
rect 15710 4467 15744 4477
rect 15710 4399 15744 4405
rect 15710 4331 15744 4333
rect 15710 4295 15744 4297
rect 15710 4223 15744 4229
rect 15710 4151 15744 4161
rect 15710 4079 15744 4093
rect 15710 4007 15744 4025
rect 15710 3922 15744 3957
rect 15614 3850 15744 3884
rect 7742 3727 7758 3761
rect 7792 3727 7808 3761
rect 10638 3725 10654 3759
rect 10688 3725 10704 3759
rect 10750 3736 10784 3832
rect 13810 3806 14036 3840
rect 10830 3725 10846 3759
rect 10880 3725 10896 3759
rect 13794 3699 13810 3733
rect 13844 3699 13860 3733
rect 13906 3710 13940 3806
rect 15550 3779 15616 3780
rect 15550 3745 15566 3779
rect 15600 3745 15616 3779
rect 15550 3744 15616 3745
rect 15710 3760 15744 3850
rect 13986 3699 14002 3733
rect 14036 3699 14052 3733
rect -1606 3394 -1590 3428
rect -1556 3394 -1540 3428
rect -1590 3290 -1110 3324
rect -1076 3290 -980 3324
rect -1686 3221 -1652 3240
rect -1686 3149 -1652 3161
rect -1686 3077 -1652 3093
rect -1686 3005 -1652 3025
rect -1686 2933 -1652 2957
rect -1686 2861 -1652 2889
rect -1686 2789 -1652 2821
rect -1686 2719 -1652 2753
rect -1686 2651 -1652 2683
rect -1686 2583 -1652 2611
rect -1686 2515 -1652 2539
rect -1686 2447 -1652 2467
rect -1686 2379 -1652 2395
rect -1686 2311 -1652 2323
rect -1686 2172 -1652 2251
rect -1590 3221 -1556 3290
rect -1590 3149 -1556 3161
rect -1590 3077 -1556 3093
rect -1590 3005 -1556 3025
rect -1590 2933 -1556 2957
rect -1590 2861 -1556 2889
rect -1590 2789 -1556 2821
rect -1590 2719 -1556 2753
rect -1590 2651 -1556 2683
rect -1590 2583 -1556 2611
rect -1590 2515 -1556 2539
rect -1590 2447 -1556 2467
rect -1590 2379 -1556 2395
rect -1590 2311 -1556 2323
rect -1590 2232 -1556 2251
rect -1494 3221 -1460 3240
rect -1494 3149 -1460 3161
rect -1494 3077 -1460 3093
rect -1494 3005 -1460 3025
rect -1494 2933 -1460 2957
rect -1494 2861 -1460 2889
rect -1494 2789 -1460 2821
rect -1494 2719 -1460 2753
rect -1494 2651 -1460 2683
rect -1494 2583 -1460 2611
rect -1494 2515 -1460 2539
rect -1494 2447 -1460 2467
rect -1494 2379 -1460 2395
rect -1494 2311 -1460 2323
rect -1494 2172 -1460 2251
rect -1398 3221 -1364 3290
rect -1398 3149 -1364 3161
rect -1398 3077 -1364 3093
rect -1398 3005 -1364 3025
rect -1398 2933 -1364 2957
rect -1398 2861 -1364 2889
rect -1398 2789 -1364 2821
rect -1398 2719 -1364 2753
rect -1398 2651 -1364 2683
rect -1398 2583 -1364 2611
rect -1398 2515 -1364 2539
rect -1398 2447 -1364 2467
rect -1398 2379 -1364 2395
rect -1398 2311 -1364 2323
rect -1398 2232 -1364 2251
rect -1302 3221 -1268 3240
rect -1302 3149 -1268 3161
rect -1302 3077 -1268 3093
rect -1302 3005 -1268 3025
rect -1302 2933 -1268 2957
rect -1302 2861 -1268 2889
rect -1302 2789 -1268 2821
rect -1302 2719 -1268 2753
rect -1302 2651 -1268 2683
rect -1302 2583 -1268 2611
rect -1302 2515 -1268 2539
rect -1302 2447 -1268 2467
rect -1302 2379 -1268 2395
rect -1302 2311 -1268 2323
rect -1302 2172 -1268 2251
rect -1206 3221 -1172 3290
rect -1206 3149 -1172 3161
rect -1206 3077 -1172 3093
rect -1206 3005 -1172 3025
rect -1206 2933 -1172 2957
rect -1206 2861 -1172 2889
rect -1206 2789 -1172 2821
rect -1206 2719 -1172 2753
rect -1206 2651 -1172 2683
rect -1206 2583 -1172 2611
rect -1206 2515 -1172 2539
rect -1206 2447 -1172 2467
rect -1206 2379 -1172 2395
rect -1206 2311 -1172 2323
rect -1206 2232 -1172 2251
rect -1110 3221 -1076 3240
rect -1110 3149 -1076 3161
rect -1110 3077 -1076 3093
rect -1110 3005 -1076 3025
rect -1110 2933 -1076 2957
rect -1110 2861 -1076 2889
rect -1110 2789 -1076 2821
rect -1110 2719 -1076 2753
rect -1110 2651 -1076 2683
rect -1110 2583 -1076 2611
rect -1110 2515 -1076 2539
rect -1110 2447 -1076 2467
rect -1110 2379 -1076 2395
rect -1110 2311 -1076 2323
rect -1110 2172 -1076 2251
rect -1014 3221 -980 3290
rect -1014 3149 -980 3161
rect -1014 3077 -980 3093
rect -1014 3005 -980 3025
rect -1014 2933 -980 2957
rect -1014 2861 -980 2889
rect -1014 2789 -980 2821
rect -1014 2719 -980 2753
rect -1014 2651 -980 2683
rect -1014 2583 -980 2611
rect -1014 2515 -980 2539
rect -1014 2447 -980 2467
rect -1014 2379 -980 2395
rect -1014 2311 -980 2323
rect -1014 2232 -980 2251
rect -918 3221 -884 3240
rect -918 3149 -884 3161
rect -918 3077 -884 3093
rect -918 3005 -884 3025
rect 1562 2968 1578 3002
rect 1612 2968 1628 3002
rect -918 2933 -884 2957
rect 1674 2906 1708 2960
rect 4518 2952 4534 2986
rect 4568 2952 4584 2986
rect 7548 2952 7564 2986
rect 7598 2952 7614 2986
rect -918 2861 -884 2889
rect 1578 2872 1804 2906
rect 4630 2890 4664 2944
rect 10636 2950 10652 2984
rect 10686 2950 10702 2984
rect 7660 2890 7694 2944
rect -918 2789 -884 2821
rect -918 2719 -884 2753
rect -918 2651 -884 2683
rect -918 2583 -884 2611
rect -918 2515 -884 2539
rect -918 2447 -884 2467
rect -918 2379 -884 2395
rect -918 2311 -884 2323
rect -918 2172 -884 2251
rect -1686 2138 -1097 2172
rect -1063 2138 -884 2172
rect 1482 2815 1516 2832
rect 1482 2743 1516 2755
rect 1482 2671 1516 2687
rect 1482 2599 1516 2619
rect 1482 2527 1516 2551
rect 1482 2455 1516 2483
rect 1482 2383 1516 2415
rect 1482 2313 1516 2347
rect 1482 2245 1516 2277
rect 1482 2177 1516 2205
rect 1482 2109 1516 2133
rect 1482 2041 1516 2061
rect 1482 1973 1516 1989
rect 1482 1905 1516 1917
rect 1482 1780 1516 1845
rect 1578 2815 1612 2872
rect 1674 2868 1708 2872
rect 1578 2743 1612 2755
rect 1578 2671 1612 2687
rect 1578 2599 1612 2619
rect 1578 2527 1612 2551
rect 1578 2455 1612 2483
rect 1578 2383 1612 2415
rect 1578 2313 1612 2347
rect 1578 2245 1612 2277
rect 1578 2177 1612 2205
rect 1578 2109 1612 2133
rect 1578 2041 1612 2061
rect 1578 1973 1612 1989
rect 1578 1905 1612 1917
rect 1578 1826 1612 1845
rect 1674 2815 1708 2832
rect 1674 2743 1708 2755
rect 1674 2671 1708 2687
rect 1674 2599 1708 2619
rect 1674 2527 1708 2551
rect 1674 2455 1708 2483
rect 1674 2383 1708 2415
rect 1674 2313 1708 2347
rect 1674 2245 1708 2277
rect 1674 2177 1708 2205
rect 1674 2109 1708 2133
rect 1674 2041 1708 2061
rect 1674 1973 1708 1989
rect 1674 1905 1708 1917
rect 1674 1780 1708 1845
rect 1770 2815 1804 2872
rect 4534 2856 4760 2890
rect 1770 2743 1804 2755
rect 1770 2671 1804 2687
rect 1770 2599 1804 2619
rect 1770 2527 1804 2551
rect 1770 2455 1804 2483
rect 1770 2383 1804 2415
rect 1770 2313 1804 2347
rect 1770 2245 1804 2277
rect 1770 2177 1804 2205
rect 1770 2109 1804 2133
rect 1770 2041 1804 2061
rect 1770 1973 1804 1989
rect 1770 1905 1804 1917
rect 1770 1828 1804 1845
rect 1866 2815 1900 2832
rect 1866 2743 1900 2755
rect 1866 2671 1900 2687
rect 1866 2599 1900 2619
rect 1866 2527 1900 2551
rect 1866 2455 1900 2483
rect 4438 2799 4472 2816
rect 4438 2727 4472 2739
rect 4438 2655 4472 2671
rect 4438 2583 4472 2603
rect 4438 2511 4472 2535
rect 4438 2439 4472 2467
rect 1866 2383 1900 2415
rect 2546 2394 2579 2428
rect 2613 2394 2646 2428
rect 4438 2367 4472 2399
rect 1866 2313 1900 2347
rect 2426 2316 2692 2350
rect 1866 2245 1900 2277
rect 1866 2177 1900 2205
rect 1866 2109 1900 2133
rect 1866 2041 1900 2061
rect 1866 1973 1900 1989
rect 1866 1905 1900 1917
rect 2500 2261 2534 2280
rect 2500 2193 2534 2195
rect 2500 2157 2534 2159
rect 2500 1912 2534 2091
rect 2658 2261 2692 2316
rect 2658 2193 2692 2195
rect 2658 2157 2692 2159
rect 2658 2072 2692 2091
rect 4438 2297 4472 2331
rect 4438 2229 4472 2261
rect 4438 2161 4472 2189
rect 4438 2093 4472 2117
rect 1866 1780 1900 1845
rect 1482 1746 1900 1780
rect 2102 1878 2534 1912
rect 4438 2025 4472 2045
rect 4438 1957 4472 1973
rect 4438 1889 4472 1901
rect 1578 1696 1612 1746
rect 2102 1522 2136 1878
rect 4438 1764 4472 1829
rect 4534 2799 4568 2856
rect 4630 2852 4664 2856
rect 4534 2727 4568 2739
rect 4534 2655 4568 2671
rect 4534 2583 4568 2603
rect 4534 2511 4568 2535
rect 4534 2439 4568 2467
rect 4534 2367 4568 2399
rect 4534 2297 4568 2331
rect 4534 2229 4568 2261
rect 4534 2161 4568 2189
rect 4534 2093 4568 2117
rect 4534 2025 4568 2045
rect 4534 1957 4568 1973
rect 4534 1889 4568 1901
rect 4534 1810 4568 1829
rect 4630 2799 4664 2816
rect 4630 2727 4664 2739
rect 4630 2655 4664 2671
rect 4630 2583 4664 2603
rect 4630 2511 4664 2535
rect 4630 2439 4664 2467
rect 4630 2367 4664 2399
rect 4630 2297 4664 2331
rect 4630 2229 4664 2261
rect 4630 2161 4664 2189
rect 4630 2093 4664 2117
rect 4630 2025 4664 2045
rect 4630 1957 4664 1973
rect 4630 1889 4664 1901
rect 4630 1764 4664 1829
rect 4726 2799 4760 2856
rect 7564 2856 7790 2890
rect 10748 2888 10782 2942
rect 13792 2924 13808 2958
rect 13842 2924 13858 2958
rect 4726 2727 4760 2739
rect 4726 2655 4760 2671
rect 4726 2583 4760 2603
rect 4726 2511 4760 2535
rect 4726 2439 4760 2467
rect 4726 2367 4760 2399
rect 4726 2297 4760 2331
rect 4726 2229 4760 2261
rect 4726 2161 4760 2189
rect 4726 2093 4760 2117
rect 4726 2025 4760 2045
rect 4726 1957 4760 1973
rect 4726 1889 4760 1901
rect 4726 1812 4760 1829
rect 4822 2799 4856 2816
rect 4822 2727 4856 2739
rect 4822 2655 4856 2671
rect 4822 2583 4856 2603
rect 4822 2511 4856 2535
rect 4822 2439 4856 2467
rect 7468 2799 7502 2816
rect 7468 2727 7502 2739
rect 7468 2655 7502 2671
rect 7468 2583 7502 2603
rect 7468 2511 7502 2535
rect 7468 2439 7502 2467
rect 4822 2367 4856 2399
rect 5546 2394 5579 2428
rect 5613 2394 5646 2428
rect 7468 2367 7502 2399
rect 4822 2297 4856 2331
rect 5426 2316 5692 2350
rect 4822 2229 4856 2261
rect 4822 2161 4856 2189
rect 4822 2093 4856 2117
rect 4822 2025 4856 2045
rect 4822 1957 4856 1973
rect 4822 1889 4856 1901
rect 4822 1764 4856 1829
rect 5500 2261 5534 2280
rect 5500 2193 5534 2195
rect 5500 2157 5534 2159
rect 5500 1788 5534 2091
rect 5658 2261 5692 2316
rect 5658 2193 5692 2195
rect 5658 2157 5692 2159
rect 5658 2070 5692 2091
rect 7468 2297 7502 2331
rect 7468 2229 7502 2261
rect 7468 2161 7502 2189
rect 7468 2093 7502 2117
rect 4438 1730 4856 1764
rect 4974 1754 5534 1788
rect 7468 2025 7502 2045
rect 7468 1957 7502 1973
rect 7468 1889 7502 1901
rect 7468 1764 7502 1829
rect 7564 2799 7598 2856
rect 7660 2852 7694 2856
rect 7564 2727 7598 2739
rect 7564 2655 7598 2671
rect 7564 2583 7598 2603
rect 7564 2511 7598 2535
rect 7564 2439 7598 2467
rect 7564 2367 7598 2399
rect 7564 2297 7598 2331
rect 7564 2229 7598 2261
rect 7564 2161 7598 2189
rect 7564 2093 7598 2117
rect 7564 2025 7598 2045
rect 7564 1957 7598 1973
rect 7564 1889 7598 1901
rect 7564 1810 7598 1829
rect 7660 2799 7694 2816
rect 7660 2727 7694 2739
rect 7660 2655 7694 2671
rect 7660 2583 7694 2603
rect 7660 2511 7694 2535
rect 7660 2439 7694 2467
rect 7660 2367 7694 2399
rect 7660 2297 7694 2331
rect 7660 2229 7694 2261
rect 7660 2161 7694 2189
rect 7660 2093 7694 2117
rect 7660 2025 7694 2045
rect 7660 1957 7694 1973
rect 7660 1889 7694 1901
rect 7660 1764 7694 1829
rect 7756 2799 7790 2856
rect 10652 2854 10878 2888
rect 13904 2862 13938 2916
rect 7756 2727 7790 2739
rect 7756 2655 7790 2671
rect 7756 2583 7790 2603
rect 7756 2511 7790 2535
rect 7756 2439 7790 2467
rect 7756 2367 7790 2399
rect 7756 2297 7790 2331
rect 7756 2229 7790 2261
rect 7756 2161 7790 2189
rect 7756 2093 7790 2117
rect 7756 2025 7790 2045
rect 7756 1957 7790 1973
rect 7756 1889 7790 1901
rect 7756 1812 7790 1829
rect 7852 2799 7886 2816
rect 7852 2727 7886 2739
rect 7852 2655 7886 2671
rect 7852 2583 7886 2603
rect 7852 2511 7886 2535
rect 7852 2439 7886 2467
rect 10556 2797 10590 2814
rect 10556 2725 10590 2737
rect 10556 2653 10590 2669
rect 10556 2581 10590 2601
rect 10556 2509 10590 2533
rect 10556 2437 10590 2465
rect 7852 2367 7886 2399
rect 8546 2394 8579 2428
rect 8613 2394 8646 2428
rect 10556 2365 10590 2397
rect 7852 2297 7886 2331
rect 8426 2316 8692 2350
rect 7852 2229 7886 2261
rect 7852 2161 7886 2189
rect 7852 2093 7886 2117
rect 7852 2025 7886 2045
rect 7852 1957 7886 1973
rect 7852 1889 7886 1901
rect 7852 1764 7886 1829
rect 8500 2261 8534 2280
rect 8500 2193 8534 2195
rect 8500 2157 8534 2159
rect 8500 1802 8534 2091
rect 8658 2261 8692 2316
rect 8658 2193 8692 2195
rect 8658 2157 8692 2159
rect 8658 2070 8692 2091
rect 10556 2295 10590 2329
rect 10556 2227 10590 2259
rect 10556 2159 10590 2187
rect 10556 2091 10590 2115
rect 4534 1680 4568 1730
rect 1664 1488 2136 1522
rect 4974 1490 5008 1754
rect 7468 1730 7886 1764
rect 8002 1768 8534 1802
rect 10556 2023 10590 2043
rect 10556 1955 10590 1971
rect 10556 1887 10590 1899
rect 7564 1680 7598 1730
rect 8002 1496 8036 1768
rect 10556 1762 10590 1827
rect 10652 2797 10686 2854
rect 10748 2850 10782 2854
rect 10652 2725 10686 2737
rect 10652 2653 10686 2669
rect 10652 2581 10686 2601
rect 10652 2509 10686 2533
rect 10652 2437 10686 2465
rect 10652 2365 10686 2397
rect 10652 2295 10686 2329
rect 10652 2227 10686 2259
rect 10652 2159 10686 2187
rect 10652 2091 10686 2115
rect 10652 2023 10686 2043
rect 10652 1955 10686 1971
rect 10652 1887 10686 1899
rect 10652 1808 10686 1827
rect 10748 2797 10782 2814
rect 10748 2725 10782 2737
rect 10748 2653 10782 2669
rect 10748 2581 10782 2601
rect 10748 2509 10782 2533
rect 10748 2437 10782 2465
rect 10748 2365 10782 2397
rect 10748 2295 10782 2329
rect 10748 2227 10782 2259
rect 10748 2159 10782 2187
rect 10748 2091 10782 2115
rect 10748 2023 10782 2043
rect 10748 1955 10782 1971
rect 10748 1887 10782 1899
rect 10748 1762 10782 1827
rect 10844 2797 10878 2854
rect 13808 2828 14034 2862
rect 10844 2725 10878 2737
rect 10844 2653 10878 2669
rect 10844 2581 10878 2601
rect 10844 2509 10878 2533
rect 10844 2437 10878 2465
rect 10844 2365 10878 2397
rect 10844 2295 10878 2329
rect 10844 2227 10878 2259
rect 10844 2159 10878 2187
rect 10844 2091 10878 2115
rect 10844 2023 10878 2043
rect 10844 1955 10878 1971
rect 10844 1887 10878 1899
rect 10844 1810 10878 1827
rect 10940 2797 10974 2814
rect 10940 2725 10974 2737
rect 10940 2653 10974 2669
rect 10940 2581 10974 2601
rect 10940 2509 10974 2533
rect 10940 2437 10974 2465
rect 13712 2771 13746 2788
rect 13712 2699 13746 2711
rect 13712 2627 13746 2643
rect 13712 2555 13746 2575
rect 13712 2483 13746 2507
rect 10940 2365 10974 2397
rect 11546 2394 11579 2428
rect 11613 2394 11646 2428
rect 13712 2411 13746 2439
rect 10940 2295 10974 2329
rect 11426 2316 11692 2350
rect 10940 2227 10974 2259
rect 10940 2159 10974 2187
rect 10940 2091 10974 2115
rect 10940 2023 10974 2043
rect 10940 1955 10974 1971
rect 10940 1887 10974 1899
rect 10940 1762 10974 1827
rect 10556 1728 10974 1762
rect 11500 2261 11534 2280
rect 11500 2193 11534 2195
rect 11500 2157 11534 2159
rect 10652 1678 10686 1728
rect 11500 1690 11534 2091
rect 11658 2261 11692 2316
rect 11658 2193 11692 2195
rect 11658 2157 11692 2159
rect 11658 2068 11692 2091
rect 13712 2339 13746 2371
rect 13712 2269 13746 2303
rect 13712 2201 13746 2233
rect 13712 2133 13746 2161
rect 13712 2065 13746 2089
rect 13712 1997 13746 2017
rect 13712 1929 13746 1945
rect 13712 1861 13746 1873
rect 13712 1736 13746 1801
rect 13808 2771 13842 2828
rect 13904 2824 13938 2828
rect 13808 2699 13842 2711
rect 13808 2627 13842 2643
rect 13808 2555 13842 2575
rect 13808 2483 13842 2507
rect 13808 2411 13842 2439
rect 13808 2339 13842 2371
rect 13808 2269 13842 2303
rect 13808 2201 13842 2233
rect 13808 2133 13842 2161
rect 13808 2065 13842 2089
rect 13808 1997 13842 2017
rect 13808 1929 13842 1945
rect 13808 1861 13842 1873
rect 13808 1782 13842 1801
rect 13904 2771 13938 2788
rect 13904 2699 13938 2711
rect 13904 2627 13938 2643
rect 13904 2555 13938 2575
rect 13904 2483 13938 2507
rect 13904 2411 13938 2439
rect 13904 2339 13938 2371
rect 13904 2269 13938 2303
rect 13904 2201 13938 2233
rect 13904 2133 13938 2161
rect 13904 2065 13938 2089
rect 13904 1997 13938 2017
rect 13904 1929 13938 1945
rect 13904 1861 13938 1873
rect 13904 1736 13938 1801
rect 14000 2771 14034 2828
rect 14000 2699 14034 2711
rect 14000 2627 14034 2643
rect 14000 2555 14034 2575
rect 14000 2483 14034 2507
rect 14000 2411 14034 2439
rect 14000 2339 14034 2371
rect 14000 2269 14034 2303
rect 14000 2201 14034 2233
rect 14000 2133 14034 2161
rect 14000 2065 14034 2089
rect 14000 1997 14034 2017
rect 14000 1929 14034 1945
rect 14000 1861 14034 1873
rect 14000 1784 14034 1801
rect 14096 2771 14130 2788
rect 14096 2699 14130 2711
rect 14096 2627 14130 2643
rect 14096 2555 14130 2575
rect 14096 2483 14130 2507
rect 14096 2411 14130 2439
rect 14546 2394 14579 2428
rect 14613 2394 14646 2428
rect 14096 2339 14130 2371
rect 14426 2316 14692 2350
rect 14096 2269 14130 2303
rect 14096 2201 14130 2233
rect 14096 2133 14130 2161
rect 14096 2065 14130 2089
rect 14096 1997 14130 2017
rect 14096 1929 14130 1945
rect 14096 1861 14130 1873
rect 14096 1736 14130 1801
rect 13712 1702 14130 1736
rect 14500 2261 14534 2280
rect 14500 2193 14534 2195
rect 14500 2157 14534 2159
rect 10966 1656 11534 1690
rect 10966 1498 11000 1656
rect 13808 1652 13842 1702
rect 14500 1638 14534 2091
rect 14658 2261 14692 2316
rect 14658 2193 14692 2195
rect 14658 2157 14692 2159
rect 14658 2070 14692 2091
rect 734 1346 768 1424
rect 252 1312 1248 1346
rect -1200 1264 -1095 1298
rect -1061 1264 -1045 1298
rect -915 1264 -899 1298
rect -865 1264 -849 1298
rect -1200 1178 -1166 1264
rect 158 1253 192 1272
rect 158 1181 192 1193
rect -1588 1144 -966 1178
rect -1686 1051 -1652 1072
rect -1686 979 -1652 991
rect -1686 907 -1652 923
rect -2308 833 -1944 876
rect -2308 255 -2279 833
rect -1973 255 -1944 833
rect -2308 236 -1944 255
rect -1686 835 -1652 855
rect -1686 763 -1652 787
rect -1686 691 -1652 719
rect -1686 619 -1652 651
rect -1686 549 -1652 583
rect -1686 481 -1652 513
rect -1686 413 -1652 441
rect -1686 345 -1652 369
rect -1686 277 -1652 297
rect -2308 212 -1942 236
rect -2026 -18 -1942 212
rect -1686 209 -1652 225
rect -1686 141 -1652 153
rect -1686 -18 -1652 81
rect -1588 1051 -1554 1144
rect -1588 979 -1554 991
rect -1588 907 -1554 923
rect -1588 835 -1554 855
rect -1588 763 -1554 787
rect -1588 691 -1554 719
rect -1588 619 -1554 651
rect -1588 549 -1554 583
rect -1588 481 -1554 513
rect -1588 413 -1554 441
rect -1588 345 -1554 369
rect -1588 277 -1554 297
rect -1588 209 -1554 225
rect -1588 141 -1554 153
rect -1588 60 -1554 81
rect -1490 1051 -1456 1068
rect -1490 979 -1456 991
rect -1490 907 -1456 923
rect -1490 835 -1456 855
rect -1490 763 -1456 787
rect -1490 691 -1456 719
rect -1490 619 -1456 651
rect -1490 549 -1456 583
rect -1490 481 -1456 513
rect -1490 413 -1456 441
rect -1490 345 -1456 369
rect -1490 277 -1456 297
rect -1490 209 -1456 225
rect -1490 141 -1456 153
rect -1490 -18 -1456 81
rect -1392 1051 -1358 1144
rect -1392 979 -1358 991
rect -1392 907 -1358 923
rect -1392 835 -1358 855
rect -1392 763 -1358 787
rect -1392 691 -1358 719
rect -1392 619 -1358 651
rect -1392 549 -1358 583
rect -1392 481 -1358 513
rect -1392 413 -1358 441
rect -1392 345 -1358 369
rect -1392 277 -1358 297
rect -1392 209 -1358 225
rect -1392 141 -1358 153
rect -1392 60 -1358 81
rect -1294 1051 -1260 1068
rect -1294 979 -1260 991
rect -1294 907 -1260 923
rect -1294 835 -1260 855
rect -1294 763 -1260 787
rect -1294 691 -1260 719
rect -1294 619 -1260 651
rect -1294 549 -1260 583
rect -1294 481 -1260 513
rect -1294 413 -1260 441
rect -1294 345 -1260 369
rect -1294 277 -1260 297
rect -1294 209 -1260 225
rect -1294 141 -1260 153
rect -1294 -18 -1260 81
rect -1196 1051 -1162 1144
rect -1196 979 -1162 991
rect -1196 907 -1162 923
rect -1196 835 -1162 855
rect -1196 763 -1162 787
rect -1196 691 -1162 719
rect -1196 619 -1162 651
rect -1196 549 -1162 583
rect -1196 481 -1162 513
rect -1196 413 -1162 441
rect -1196 345 -1162 369
rect -1196 277 -1162 297
rect -1196 209 -1162 225
rect -1196 141 -1162 153
rect -1196 60 -1162 81
rect -1098 1051 -1064 1068
rect -1098 979 -1064 991
rect -1098 907 -1064 923
rect -1098 835 -1064 855
rect -1098 763 -1064 787
rect -1098 691 -1064 719
rect -1098 619 -1064 651
rect -1098 549 -1064 583
rect -1098 481 -1064 513
rect -1098 413 -1064 441
rect -1098 345 -1064 369
rect -1098 277 -1064 297
rect -1098 209 -1064 225
rect -1098 141 -1064 153
rect -1098 -18 -1064 81
rect -1000 1051 -966 1144
rect 158 1109 192 1125
rect -1000 979 -966 991
rect -1000 907 -966 923
rect -1000 835 -966 855
rect -1000 763 -966 787
rect -1000 691 -966 719
rect -1000 619 -966 651
rect -1000 549 -966 583
rect -1000 481 -966 513
rect -1000 413 -966 441
rect -1000 345 -966 369
rect -1000 277 -966 297
rect -1000 209 -966 225
rect -1000 141 -966 153
rect -1000 60 -966 81
rect -902 1051 -868 1070
rect -902 979 -868 991
rect -902 907 -868 923
rect -902 835 -868 855
rect -902 763 -868 787
rect -902 691 -868 719
rect -902 619 -868 651
rect -902 549 -868 583
rect -902 481 -868 513
rect -902 413 -868 441
rect -902 345 -868 369
rect -902 277 -868 297
rect -902 209 -868 225
rect 158 1037 192 1057
rect 158 965 192 989
rect 158 893 192 921
rect 158 821 192 853
rect 158 751 192 785
rect 158 683 192 715
rect 158 615 192 643
rect 158 547 192 571
rect 158 479 192 499
rect 158 411 192 427
rect 158 343 192 355
rect 158 214 192 283
rect 254 1253 288 1312
rect 254 1181 288 1193
rect 254 1109 288 1125
rect 254 1037 288 1057
rect 254 965 288 989
rect 254 893 288 921
rect 254 821 288 853
rect 254 751 288 785
rect 254 683 288 715
rect 254 615 288 643
rect 254 547 288 571
rect 254 479 288 499
rect 254 411 288 427
rect 254 343 288 355
rect 254 264 288 283
rect 350 1253 384 1270
rect 350 1181 384 1193
rect 350 1109 384 1125
rect 350 1037 384 1057
rect 350 965 384 989
rect 350 893 384 921
rect 350 821 384 853
rect 350 751 384 785
rect 350 683 384 715
rect 350 615 384 643
rect 350 547 384 571
rect 350 479 384 499
rect 350 411 384 427
rect 350 343 384 355
rect 350 214 384 283
rect 446 1253 480 1312
rect 446 1181 480 1193
rect 446 1109 480 1125
rect 446 1037 480 1057
rect 446 965 480 989
rect 446 893 480 921
rect 446 821 480 853
rect 446 751 480 785
rect 446 683 480 715
rect 446 615 480 643
rect 446 547 480 571
rect 446 479 480 499
rect 446 411 480 427
rect 446 343 480 355
rect 446 264 480 283
rect 542 1253 576 1270
rect 542 1181 576 1193
rect 542 1109 576 1125
rect 542 1037 576 1057
rect 542 965 576 989
rect 542 893 576 921
rect 542 821 576 853
rect 542 751 576 785
rect 542 683 576 715
rect 542 615 576 643
rect 542 547 576 571
rect 542 479 576 499
rect 542 411 576 427
rect 542 343 576 355
rect 542 214 576 283
rect 638 1253 672 1312
rect 638 1181 672 1193
rect 638 1109 672 1125
rect 638 1037 672 1057
rect 638 965 672 989
rect 638 893 672 921
rect 638 821 672 853
rect 638 751 672 785
rect 638 683 672 715
rect 638 615 672 643
rect 638 547 672 571
rect 638 479 672 499
rect 638 411 672 427
rect 638 343 672 355
rect 638 264 672 283
rect 734 1253 768 1270
rect 734 1181 768 1193
rect 734 1109 768 1125
rect 734 1037 768 1057
rect 734 965 768 989
rect 734 893 768 921
rect 734 821 768 853
rect 734 751 768 785
rect 734 683 768 715
rect 734 615 768 643
rect 734 547 768 571
rect 734 479 768 499
rect 734 411 768 427
rect 734 343 768 355
rect 734 214 768 283
rect 830 1253 864 1312
rect 830 1181 864 1193
rect 830 1109 864 1125
rect 830 1037 864 1057
rect 830 965 864 989
rect 830 893 864 921
rect 830 821 864 853
rect 830 751 864 785
rect 830 683 864 715
rect 830 615 864 643
rect 830 547 864 571
rect 830 479 864 499
rect 830 411 864 427
rect 830 343 864 355
rect 830 264 864 283
rect 926 1253 960 1270
rect 926 1181 960 1193
rect 926 1109 960 1125
rect 926 1037 960 1057
rect 926 965 960 989
rect 926 893 960 921
rect 926 821 960 853
rect 926 751 960 785
rect 926 683 960 715
rect 926 615 960 643
rect 926 547 960 571
rect 926 479 960 499
rect 926 411 960 427
rect 926 343 960 355
rect 926 214 960 283
rect 1022 1253 1056 1312
rect 1022 1181 1056 1193
rect 1022 1109 1056 1125
rect 1022 1037 1056 1057
rect 1022 965 1056 989
rect 1022 893 1056 921
rect 1022 821 1056 853
rect 1022 751 1056 785
rect 1022 683 1056 715
rect 1022 615 1056 643
rect 1022 547 1056 571
rect 1022 479 1056 499
rect 1022 411 1056 427
rect 1022 343 1056 355
rect 1022 264 1056 283
rect 1118 1253 1152 1270
rect 1118 1181 1152 1193
rect 1118 1109 1152 1125
rect 1118 1037 1152 1057
rect 1118 965 1152 989
rect 1118 893 1152 921
rect 1118 821 1152 853
rect 1118 751 1152 785
rect 1118 683 1152 715
rect 1118 615 1152 643
rect 1118 547 1152 571
rect 1118 479 1152 499
rect 1118 411 1152 427
rect 1118 343 1152 355
rect 1118 214 1152 283
rect 1214 1253 1248 1312
rect 1214 1181 1248 1193
rect 1214 1109 1248 1125
rect 1214 1037 1248 1057
rect 1214 965 1248 989
rect 1214 893 1248 921
rect 1214 821 1248 853
rect 1214 751 1248 785
rect 1214 683 1248 715
rect 1214 615 1248 643
rect 1214 547 1248 571
rect 1214 479 1248 499
rect 1214 411 1248 427
rect 1214 343 1248 355
rect 1214 266 1248 283
rect 1310 1253 1344 1270
rect 1310 1181 1344 1193
rect 1310 1109 1344 1125
rect 1310 1037 1344 1057
rect 1310 965 1344 989
rect 1310 893 1344 921
rect 1310 821 1344 853
rect 1310 751 1344 785
rect 1310 683 1344 715
rect 1310 615 1344 643
rect 1310 547 1344 571
rect 1310 479 1344 499
rect 1310 411 1344 427
rect 1310 343 1344 355
rect 1310 214 1344 283
rect 158 180 1344 214
rect -902 141 -868 153
rect 140 96 156 130
rect 190 96 206 130
rect -902 -18 -868 81
rect 626 -18 722 180
rect 830 120 864 180
rect 1664 24 1698 1488
rect 4664 1456 5008 1490
rect 7664 1462 8036 1496
rect 10664 1464 11000 1498
rect 14152 1604 14534 1638
rect 2400 1368 2434 1418
rect 2022 1334 3016 1368
rect 1926 1253 1960 1272
rect 1926 1181 1960 1193
rect 1926 1109 1960 1125
rect 1926 1037 1960 1057
rect 1926 965 1960 989
rect 1926 893 1960 921
rect 1926 821 1960 853
rect 1926 751 1960 785
rect 1926 683 1960 715
rect 1926 615 1960 643
rect 1926 547 1960 571
rect 1926 479 1960 499
rect 1926 411 1960 427
rect 1926 343 1960 355
rect 1926 216 1960 283
rect 2022 1253 2056 1334
rect 2022 1181 2056 1193
rect 2022 1109 2056 1125
rect 2022 1037 2056 1057
rect 2022 965 2056 989
rect 2022 893 2056 921
rect 2022 821 2056 853
rect 2022 751 2056 785
rect 2022 683 2056 715
rect 2022 615 2056 643
rect 2022 547 2056 571
rect 2022 479 2056 499
rect 2022 411 2056 427
rect 2022 343 2056 355
rect 2022 264 2056 283
rect 2118 1253 2152 1272
rect 2118 1181 2152 1193
rect 2118 1109 2152 1125
rect 2118 1037 2152 1057
rect 2118 965 2152 989
rect 2118 893 2152 921
rect 2118 821 2152 853
rect 2118 751 2152 785
rect 2118 683 2152 715
rect 2118 615 2152 643
rect 2118 547 2152 571
rect 2118 479 2152 499
rect 2118 411 2152 427
rect 2118 343 2152 355
rect 2118 216 2152 283
rect 2214 1253 2248 1334
rect 2214 1181 2248 1193
rect 2214 1109 2248 1125
rect 2214 1037 2248 1057
rect 2214 965 2248 989
rect 2214 893 2248 921
rect 2214 821 2248 853
rect 2214 751 2248 785
rect 2214 683 2248 715
rect 2214 615 2248 643
rect 2214 547 2248 571
rect 2214 479 2248 499
rect 2214 411 2248 427
rect 2214 343 2248 355
rect 2214 264 2248 283
rect 2310 1253 2344 1272
rect 2310 1181 2344 1193
rect 2310 1109 2344 1125
rect 2310 1037 2344 1057
rect 2310 965 2344 989
rect 2310 893 2344 921
rect 2310 821 2344 853
rect 2310 751 2344 785
rect 2310 683 2344 715
rect 2310 615 2344 643
rect 2310 547 2344 571
rect 2310 479 2344 499
rect 2310 411 2344 427
rect 2310 343 2344 355
rect 2310 216 2344 283
rect 2406 1253 2440 1334
rect 2406 1181 2440 1193
rect 2406 1109 2440 1125
rect 2406 1037 2440 1057
rect 2406 965 2440 989
rect 2406 893 2440 921
rect 2406 821 2440 853
rect 2406 751 2440 785
rect 2406 683 2440 715
rect 2406 615 2440 643
rect 2406 547 2440 571
rect 2406 479 2440 499
rect 2406 411 2440 427
rect 2406 343 2440 355
rect 2406 264 2440 283
rect 2502 1253 2536 1272
rect 2502 1181 2536 1193
rect 2502 1109 2536 1125
rect 2502 1037 2536 1057
rect 2502 965 2536 989
rect 2502 893 2536 921
rect 2502 821 2536 853
rect 2502 751 2536 785
rect 2502 683 2536 715
rect 2502 615 2536 643
rect 2502 547 2536 571
rect 2502 479 2536 499
rect 2502 411 2536 427
rect 2502 343 2536 355
rect 2502 216 2536 283
rect 2598 1253 2632 1334
rect 2598 1181 2632 1193
rect 2598 1109 2632 1125
rect 2598 1037 2632 1057
rect 2598 965 2632 989
rect 2598 893 2632 921
rect 2598 821 2632 853
rect 2598 751 2632 785
rect 2598 683 2632 715
rect 2598 615 2632 643
rect 2598 547 2632 571
rect 2598 479 2632 499
rect 2598 411 2632 427
rect 2598 343 2632 355
rect 2598 266 2632 283
rect 2694 1253 2728 1272
rect 2694 1181 2728 1193
rect 2694 1109 2728 1125
rect 2694 1037 2728 1057
rect 2694 965 2728 989
rect 2694 893 2728 921
rect 2694 821 2728 853
rect 2694 751 2728 785
rect 2694 683 2728 715
rect 2694 615 2728 643
rect 2694 547 2728 571
rect 2694 479 2728 499
rect 2694 411 2728 427
rect 2694 343 2728 355
rect 2694 216 2728 283
rect 2790 1253 2824 1334
rect 2790 1181 2824 1193
rect 2790 1109 2824 1125
rect 2790 1037 2824 1057
rect 2790 965 2824 989
rect 2790 893 2824 921
rect 2790 821 2824 853
rect 2790 751 2824 785
rect 2790 683 2824 715
rect 2790 615 2824 643
rect 2790 547 2824 571
rect 2790 479 2824 499
rect 2790 411 2824 427
rect 2790 343 2824 355
rect 2790 266 2824 283
rect 2886 1253 2920 1272
rect 2886 1181 2920 1193
rect 2886 1109 2920 1125
rect 2886 1037 2920 1057
rect 2886 965 2920 989
rect 2886 893 2920 921
rect 2886 821 2920 853
rect 2886 751 2920 785
rect 2886 683 2920 715
rect 2886 615 2920 643
rect 2886 547 2920 571
rect 2886 479 2920 499
rect 2886 411 2920 427
rect 2886 343 2920 355
rect 2886 216 2920 283
rect 2982 1253 3016 1334
rect 3690 1330 3724 1408
rect 3208 1296 4204 1330
rect 2982 1181 3016 1193
rect 2982 1109 3016 1125
rect 2982 1037 3016 1057
rect 2982 965 3016 989
rect 2982 893 3016 921
rect 2982 821 3016 853
rect 2982 751 3016 785
rect 2982 683 3016 715
rect 2982 615 3016 643
rect 2982 547 3016 571
rect 2982 479 3016 499
rect 2982 411 3016 427
rect 2982 343 3016 355
rect 2982 266 3016 283
rect 3114 1237 3148 1256
rect 3114 1165 3148 1177
rect 3114 1093 3148 1109
rect 3114 1021 3148 1041
rect 3114 949 3148 973
rect 3114 877 3148 905
rect 3114 805 3148 837
rect 3114 735 3148 769
rect 3114 667 3148 699
rect 3114 599 3148 627
rect 3114 531 3148 555
rect 3114 463 3148 483
rect 3114 395 3148 411
rect 3114 327 3148 339
rect 1926 182 2920 216
rect 3114 198 3148 267
rect 3210 1237 3244 1296
rect 3210 1165 3244 1177
rect 3210 1093 3244 1109
rect 3210 1021 3244 1041
rect 3210 949 3244 973
rect 3210 877 3244 905
rect 3210 805 3244 837
rect 3210 735 3244 769
rect 3210 667 3244 699
rect 3210 599 3244 627
rect 3210 531 3244 555
rect 3210 463 3244 483
rect 3210 395 3244 411
rect 3210 327 3244 339
rect 3210 248 3244 267
rect 3306 1237 3340 1254
rect 3306 1165 3340 1177
rect 3306 1093 3340 1109
rect 3306 1021 3340 1041
rect 3306 949 3340 973
rect 3306 877 3340 905
rect 3306 805 3340 837
rect 3306 735 3340 769
rect 3306 667 3340 699
rect 3306 599 3340 627
rect 3306 531 3340 555
rect 3306 463 3340 483
rect 3306 395 3340 411
rect 3306 327 3340 339
rect 3306 198 3340 267
rect 3402 1237 3436 1296
rect 3402 1165 3436 1177
rect 3402 1093 3436 1109
rect 3402 1021 3436 1041
rect 3402 949 3436 973
rect 3402 877 3436 905
rect 3402 805 3436 837
rect 3402 735 3436 769
rect 3402 667 3436 699
rect 3402 599 3436 627
rect 3402 531 3436 555
rect 3402 463 3436 483
rect 3402 395 3436 411
rect 3402 327 3436 339
rect 3402 248 3436 267
rect 3498 1237 3532 1254
rect 3498 1165 3532 1177
rect 3498 1093 3532 1109
rect 3498 1021 3532 1041
rect 3498 949 3532 973
rect 3498 877 3532 905
rect 3498 805 3532 837
rect 3498 735 3532 769
rect 3498 667 3532 699
rect 3498 599 3532 627
rect 3498 531 3532 555
rect 3498 463 3532 483
rect 3498 395 3532 411
rect 3498 327 3532 339
rect 3498 198 3532 267
rect 3594 1237 3628 1296
rect 3594 1165 3628 1177
rect 3594 1093 3628 1109
rect 3594 1021 3628 1041
rect 3594 949 3628 973
rect 3594 877 3628 905
rect 3594 805 3628 837
rect 3594 735 3628 769
rect 3594 667 3628 699
rect 3594 599 3628 627
rect 3594 531 3628 555
rect 3594 463 3628 483
rect 3594 395 3628 411
rect 3594 327 3628 339
rect 3594 248 3628 267
rect 3690 1237 3724 1254
rect 3690 1165 3724 1177
rect 3690 1093 3724 1109
rect 3690 1021 3724 1041
rect 3690 949 3724 973
rect 3690 877 3724 905
rect 3690 805 3724 837
rect 3690 735 3724 769
rect 3690 667 3724 699
rect 3690 599 3724 627
rect 3690 531 3724 555
rect 3690 463 3724 483
rect 3690 395 3724 411
rect 3690 327 3724 339
rect 3690 198 3724 267
rect 3786 1237 3820 1296
rect 3786 1165 3820 1177
rect 3786 1093 3820 1109
rect 3786 1021 3820 1041
rect 3786 949 3820 973
rect 3786 877 3820 905
rect 3786 805 3820 837
rect 3786 735 3820 769
rect 3786 667 3820 699
rect 3786 599 3820 627
rect 3786 531 3820 555
rect 3786 463 3820 483
rect 3786 395 3820 411
rect 3786 327 3820 339
rect 3786 248 3820 267
rect 3882 1237 3916 1254
rect 3882 1165 3916 1177
rect 3882 1093 3916 1109
rect 3882 1021 3916 1041
rect 3882 949 3916 973
rect 3882 877 3916 905
rect 3882 805 3916 837
rect 3882 735 3916 769
rect 3882 667 3916 699
rect 3882 599 3916 627
rect 3882 531 3916 555
rect 3882 463 3916 483
rect 3882 395 3916 411
rect 3882 327 3916 339
rect 3882 198 3916 267
rect 3978 1237 4012 1296
rect 3978 1165 4012 1177
rect 3978 1093 4012 1109
rect 3978 1021 4012 1041
rect 3978 949 4012 973
rect 3978 877 4012 905
rect 3978 805 4012 837
rect 3978 735 4012 769
rect 3978 667 4012 699
rect 3978 599 4012 627
rect 3978 531 4012 555
rect 3978 463 4012 483
rect 3978 395 4012 411
rect 3978 327 4012 339
rect 3978 248 4012 267
rect 4074 1237 4108 1254
rect 4074 1165 4108 1177
rect 4074 1093 4108 1109
rect 4074 1021 4108 1041
rect 4074 949 4108 973
rect 4074 877 4108 905
rect 4074 805 4108 837
rect 4074 735 4108 769
rect 4074 667 4108 699
rect 4074 599 4108 627
rect 4074 531 4108 555
rect 4074 463 4108 483
rect 4074 395 4108 411
rect 4074 327 4108 339
rect 4074 198 4108 267
rect 4170 1237 4204 1296
rect 4170 1165 4204 1177
rect 4170 1093 4204 1109
rect 4170 1021 4204 1041
rect 4170 949 4204 973
rect 4170 877 4204 905
rect 4170 805 4204 837
rect 4170 735 4204 769
rect 4170 667 4204 699
rect 4170 599 4204 627
rect 4170 531 4204 555
rect 4170 463 4204 483
rect 4170 395 4204 411
rect 4170 327 4204 339
rect 4170 250 4204 267
rect 4266 1237 4300 1254
rect 4266 1165 4300 1177
rect 4266 1093 4300 1109
rect 4266 1021 4300 1041
rect 4266 949 4300 973
rect 4266 877 4300 905
rect 4266 805 4300 837
rect 4266 735 4300 769
rect 4266 667 4300 699
rect 4266 599 4300 627
rect 4266 531 4300 555
rect 4266 463 4300 483
rect 4266 395 4300 411
rect 4266 327 4300 339
rect 4266 198 4300 267
rect 2494 146 2528 182
rect 3114 164 4300 198
rect 2772 96 2788 130
rect 2822 96 2838 130
rect 3096 80 3112 114
rect 3146 80 3162 114
rect 3786 104 3820 164
rect 4664 16 4698 1456
rect 5356 1352 5390 1402
rect 4978 1318 5972 1352
rect 6720 1330 6754 1408
rect 4882 1237 4916 1256
rect 4882 1165 4916 1177
rect 4882 1093 4916 1109
rect 4882 1021 4916 1041
rect 4882 949 4916 973
rect 4882 877 4916 905
rect 4882 805 4916 837
rect 4882 735 4916 769
rect 4882 667 4916 699
rect 4882 599 4916 627
rect 4882 531 4916 555
rect 4882 463 4916 483
rect 4882 395 4916 411
rect 4882 327 4916 339
rect 4882 200 4916 267
rect 4978 1237 5012 1318
rect 4978 1165 5012 1177
rect 4978 1093 5012 1109
rect 4978 1021 5012 1041
rect 4978 949 5012 973
rect 4978 877 5012 905
rect 4978 805 5012 837
rect 4978 735 5012 769
rect 4978 667 5012 699
rect 4978 599 5012 627
rect 4978 531 5012 555
rect 4978 463 5012 483
rect 4978 395 5012 411
rect 4978 327 5012 339
rect 4978 248 5012 267
rect 5074 1237 5108 1256
rect 5074 1165 5108 1177
rect 5074 1093 5108 1109
rect 5074 1021 5108 1041
rect 5074 949 5108 973
rect 5074 877 5108 905
rect 5074 805 5108 837
rect 5074 735 5108 769
rect 5074 667 5108 699
rect 5074 599 5108 627
rect 5074 531 5108 555
rect 5074 463 5108 483
rect 5074 395 5108 411
rect 5074 327 5108 339
rect 5074 200 5108 267
rect 5170 1237 5204 1318
rect 5170 1165 5204 1177
rect 5170 1093 5204 1109
rect 5170 1021 5204 1041
rect 5170 949 5204 973
rect 5170 877 5204 905
rect 5170 805 5204 837
rect 5170 735 5204 769
rect 5170 667 5204 699
rect 5170 599 5204 627
rect 5170 531 5204 555
rect 5170 463 5204 483
rect 5170 395 5204 411
rect 5170 327 5204 339
rect 5170 248 5204 267
rect 5266 1237 5300 1256
rect 5266 1165 5300 1177
rect 5266 1093 5300 1109
rect 5266 1021 5300 1041
rect 5266 949 5300 973
rect 5266 877 5300 905
rect 5266 805 5300 837
rect 5266 735 5300 769
rect 5266 667 5300 699
rect 5266 599 5300 627
rect 5266 531 5300 555
rect 5266 463 5300 483
rect 5266 395 5300 411
rect 5266 327 5300 339
rect 5266 200 5300 267
rect 5362 1237 5396 1318
rect 5362 1165 5396 1177
rect 5362 1093 5396 1109
rect 5362 1021 5396 1041
rect 5362 949 5396 973
rect 5362 877 5396 905
rect 5362 805 5396 837
rect 5362 735 5396 769
rect 5362 667 5396 699
rect 5362 599 5396 627
rect 5362 531 5396 555
rect 5362 463 5396 483
rect 5362 395 5396 411
rect 5362 327 5396 339
rect 5362 248 5396 267
rect 5458 1237 5492 1256
rect 5458 1165 5492 1177
rect 5458 1093 5492 1109
rect 5458 1021 5492 1041
rect 5458 949 5492 973
rect 5458 877 5492 905
rect 5458 805 5492 837
rect 5458 735 5492 769
rect 5458 667 5492 699
rect 5458 599 5492 627
rect 5458 531 5492 555
rect 5458 463 5492 483
rect 5458 395 5492 411
rect 5458 327 5492 339
rect 5458 200 5492 267
rect 5554 1237 5588 1318
rect 5554 1165 5588 1177
rect 5554 1093 5588 1109
rect 5554 1021 5588 1041
rect 5554 949 5588 973
rect 5554 877 5588 905
rect 5554 805 5588 837
rect 5554 735 5588 769
rect 5554 667 5588 699
rect 5554 599 5588 627
rect 5554 531 5588 555
rect 5554 463 5588 483
rect 5554 395 5588 411
rect 5554 327 5588 339
rect 5554 250 5588 267
rect 5650 1237 5684 1256
rect 5650 1165 5684 1177
rect 5650 1093 5684 1109
rect 5650 1021 5684 1041
rect 5650 949 5684 973
rect 5650 877 5684 905
rect 5650 805 5684 837
rect 5650 735 5684 769
rect 5650 667 5684 699
rect 5650 599 5684 627
rect 5650 531 5684 555
rect 5650 463 5684 483
rect 5650 395 5684 411
rect 5650 327 5684 339
rect 5650 200 5684 267
rect 5746 1237 5780 1318
rect 5746 1165 5780 1177
rect 5746 1093 5780 1109
rect 5746 1021 5780 1041
rect 5746 949 5780 973
rect 5746 877 5780 905
rect 5746 805 5780 837
rect 5746 735 5780 769
rect 5746 667 5780 699
rect 5746 599 5780 627
rect 5746 531 5780 555
rect 5746 463 5780 483
rect 5746 395 5780 411
rect 5746 327 5780 339
rect 5746 250 5780 267
rect 5842 1237 5876 1256
rect 5842 1165 5876 1177
rect 5842 1093 5876 1109
rect 5842 1021 5876 1041
rect 5842 949 5876 973
rect 5842 877 5876 905
rect 5842 805 5876 837
rect 5842 735 5876 769
rect 5842 667 5876 699
rect 5842 599 5876 627
rect 5842 531 5876 555
rect 5842 463 5876 483
rect 5842 395 5876 411
rect 5842 327 5876 339
rect 5842 200 5876 267
rect 5938 1237 5972 1318
rect 6238 1296 7234 1330
rect 5938 1165 5972 1177
rect 5938 1093 5972 1109
rect 5938 1021 5972 1041
rect 5938 949 5972 973
rect 5938 877 5972 905
rect 5938 805 5972 837
rect 5938 735 5972 769
rect 5938 667 5972 699
rect 5938 599 5972 627
rect 5938 531 5972 555
rect 5938 463 5972 483
rect 5938 395 5972 411
rect 5938 327 5972 339
rect 5938 250 5972 267
rect 6144 1237 6178 1256
rect 6144 1165 6178 1177
rect 6144 1093 6178 1109
rect 6144 1021 6178 1041
rect 6144 949 6178 973
rect 6144 877 6178 905
rect 6144 805 6178 837
rect 6144 735 6178 769
rect 6144 667 6178 699
rect 6144 599 6178 627
rect 6144 531 6178 555
rect 6144 463 6178 483
rect 6144 395 6178 411
rect 6144 327 6178 339
rect 4882 166 5876 200
rect 6144 198 6178 267
rect 6240 1237 6274 1296
rect 6240 1165 6274 1177
rect 6240 1093 6274 1109
rect 6240 1021 6274 1041
rect 6240 949 6274 973
rect 6240 877 6274 905
rect 6240 805 6274 837
rect 6240 735 6274 769
rect 6240 667 6274 699
rect 6240 599 6274 627
rect 6240 531 6274 555
rect 6240 463 6274 483
rect 6240 395 6274 411
rect 6240 327 6274 339
rect 6240 248 6274 267
rect 6336 1237 6370 1254
rect 6336 1165 6370 1177
rect 6336 1093 6370 1109
rect 6336 1021 6370 1041
rect 6336 949 6370 973
rect 6336 877 6370 905
rect 6336 805 6370 837
rect 6336 735 6370 769
rect 6336 667 6370 699
rect 6336 599 6370 627
rect 6336 531 6370 555
rect 6336 463 6370 483
rect 6336 395 6370 411
rect 6336 327 6370 339
rect 6336 198 6370 267
rect 6432 1237 6466 1296
rect 6432 1165 6466 1177
rect 6432 1093 6466 1109
rect 6432 1021 6466 1041
rect 6432 949 6466 973
rect 6432 877 6466 905
rect 6432 805 6466 837
rect 6432 735 6466 769
rect 6432 667 6466 699
rect 6432 599 6466 627
rect 6432 531 6466 555
rect 6432 463 6466 483
rect 6432 395 6466 411
rect 6432 327 6466 339
rect 6432 248 6466 267
rect 6528 1237 6562 1254
rect 6528 1165 6562 1177
rect 6528 1093 6562 1109
rect 6528 1021 6562 1041
rect 6528 949 6562 973
rect 6528 877 6562 905
rect 6528 805 6562 837
rect 6528 735 6562 769
rect 6528 667 6562 699
rect 6528 599 6562 627
rect 6528 531 6562 555
rect 6528 463 6562 483
rect 6528 395 6562 411
rect 6528 327 6562 339
rect 6528 198 6562 267
rect 6624 1237 6658 1296
rect 6624 1165 6658 1177
rect 6624 1093 6658 1109
rect 6624 1021 6658 1041
rect 6624 949 6658 973
rect 6624 877 6658 905
rect 6624 805 6658 837
rect 6624 735 6658 769
rect 6624 667 6658 699
rect 6624 599 6658 627
rect 6624 531 6658 555
rect 6624 463 6658 483
rect 6624 395 6658 411
rect 6624 327 6658 339
rect 6624 248 6658 267
rect 6720 1237 6754 1254
rect 6720 1165 6754 1177
rect 6720 1093 6754 1109
rect 6720 1021 6754 1041
rect 6720 949 6754 973
rect 6720 877 6754 905
rect 6720 805 6754 837
rect 6720 735 6754 769
rect 6720 667 6754 699
rect 6720 599 6754 627
rect 6720 531 6754 555
rect 6720 463 6754 483
rect 6720 395 6754 411
rect 6720 327 6754 339
rect 6720 198 6754 267
rect 6816 1237 6850 1296
rect 6816 1165 6850 1177
rect 6816 1093 6850 1109
rect 6816 1021 6850 1041
rect 6816 949 6850 973
rect 6816 877 6850 905
rect 6816 805 6850 837
rect 6816 735 6850 769
rect 6816 667 6850 699
rect 6816 599 6850 627
rect 6816 531 6850 555
rect 6816 463 6850 483
rect 6816 395 6850 411
rect 6816 327 6850 339
rect 6816 248 6850 267
rect 6912 1237 6946 1254
rect 6912 1165 6946 1177
rect 6912 1093 6946 1109
rect 6912 1021 6946 1041
rect 6912 949 6946 973
rect 6912 877 6946 905
rect 6912 805 6946 837
rect 6912 735 6946 769
rect 6912 667 6946 699
rect 6912 599 6946 627
rect 6912 531 6946 555
rect 6912 463 6946 483
rect 6912 395 6946 411
rect 6912 327 6946 339
rect 6912 198 6946 267
rect 7008 1237 7042 1296
rect 7008 1165 7042 1177
rect 7008 1093 7042 1109
rect 7008 1021 7042 1041
rect 7008 949 7042 973
rect 7008 877 7042 905
rect 7008 805 7042 837
rect 7008 735 7042 769
rect 7008 667 7042 699
rect 7008 599 7042 627
rect 7008 531 7042 555
rect 7008 463 7042 483
rect 7008 395 7042 411
rect 7008 327 7042 339
rect 7008 248 7042 267
rect 7104 1237 7138 1254
rect 7104 1165 7138 1177
rect 7104 1093 7138 1109
rect 7104 1021 7138 1041
rect 7104 949 7138 973
rect 7104 877 7138 905
rect 7104 805 7138 837
rect 7104 735 7138 769
rect 7104 667 7138 699
rect 7104 599 7138 627
rect 7104 531 7138 555
rect 7104 463 7138 483
rect 7104 395 7138 411
rect 7104 327 7138 339
rect 7104 198 7138 267
rect 7200 1237 7234 1296
rect 7200 1165 7234 1177
rect 7200 1093 7234 1109
rect 7200 1021 7234 1041
rect 7200 949 7234 973
rect 7200 877 7234 905
rect 7200 805 7234 837
rect 7200 735 7234 769
rect 7200 667 7234 699
rect 7200 599 7234 627
rect 7200 531 7234 555
rect 7200 463 7234 483
rect 7200 395 7234 411
rect 7200 327 7234 339
rect 7200 250 7234 267
rect 7296 1237 7330 1254
rect 7296 1165 7330 1177
rect 7296 1093 7330 1109
rect 7296 1021 7330 1041
rect 7296 949 7330 973
rect 7296 877 7330 905
rect 7296 805 7330 837
rect 7296 735 7330 769
rect 7296 667 7330 699
rect 7296 599 7330 627
rect 7296 531 7330 555
rect 7296 463 7330 483
rect 7296 395 7330 411
rect 7296 327 7330 339
rect 7296 198 7330 267
rect 5450 130 5484 166
rect 6144 164 7330 198
rect 5728 80 5744 114
rect 5778 80 5794 114
rect 6126 80 6142 114
rect 6176 80 6192 114
rect 6816 104 6850 164
rect 7664 18 7698 1462
rect 8386 1352 8420 1402
rect 8008 1318 9002 1352
rect 9808 1328 9842 1406
rect 7912 1237 7946 1256
rect 7912 1165 7946 1177
rect 7912 1093 7946 1109
rect 7912 1021 7946 1041
rect 7912 949 7946 973
rect 7912 877 7946 905
rect 7912 805 7946 837
rect 7912 735 7946 769
rect 7912 667 7946 699
rect 7912 599 7946 627
rect 7912 531 7946 555
rect 7912 463 7946 483
rect 7912 395 7946 411
rect 7912 327 7946 339
rect 7912 200 7946 267
rect 8008 1237 8042 1318
rect 8008 1165 8042 1177
rect 8008 1093 8042 1109
rect 8008 1021 8042 1041
rect 8008 949 8042 973
rect 8008 877 8042 905
rect 8008 805 8042 837
rect 8008 735 8042 769
rect 8008 667 8042 699
rect 8008 599 8042 627
rect 8008 531 8042 555
rect 8008 463 8042 483
rect 8008 395 8042 411
rect 8008 327 8042 339
rect 8008 248 8042 267
rect 8104 1237 8138 1256
rect 8104 1165 8138 1177
rect 8104 1093 8138 1109
rect 8104 1021 8138 1041
rect 8104 949 8138 973
rect 8104 877 8138 905
rect 8104 805 8138 837
rect 8104 735 8138 769
rect 8104 667 8138 699
rect 8104 599 8138 627
rect 8104 531 8138 555
rect 8104 463 8138 483
rect 8104 395 8138 411
rect 8104 327 8138 339
rect 8104 200 8138 267
rect 8200 1237 8234 1318
rect 8200 1165 8234 1177
rect 8200 1093 8234 1109
rect 8200 1021 8234 1041
rect 8200 949 8234 973
rect 8200 877 8234 905
rect 8200 805 8234 837
rect 8200 735 8234 769
rect 8200 667 8234 699
rect 8200 599 8234 627
rect 8200 531 8234 555
rect 8200 463 8234 483
rect 8200 395 8234 411
rect 8200 327 8234 339
rect 8200 248 8234 267
rect 8296 1237 8330 1256
rect 8296 1165 8330 1177
rect 8296 1093 8330 1109
rect 8296 1021 8330 1041
rect 8296 949 8330 973
rect 8296 877 8330 905
rect 8296 805 8330 837
rect 8296 735 8330 769
rect 8296 667 8330 699
rect 8296 599 8330 627
rect 8296 531 8330 555
rect 8296 463 8330 483
rect 8296 395 8330 411
rect 8296 327 8330 339
rect 8296 200 8330 267
rect 8392 1237 8426 1318
rect 8392 1165 8426 1177
rect 8392 1093 8426 1109
rect 8392 1021 8426 1041
rect 8392 949 8426 973
rect 8392 877 8426 905
rect 8392 805 8426 837
rect 8392 735 8426 769
rect 8392 667 8426 699
rect 8392 599 8426 627
rect 8392 531 8426 555
rect 8392 463 8426 483
rect 8392 395 8426 411
rect 8392 327 8426 339
rect 8392 248 8426 267
rect 8488 1237 8522 1256
rect 8488 1165 8522 1177
rect 8488 1093 8522 1109
rect 8488 1021 8522 1041
rect 8488 949 8522 973
rect 8488 877 8522 905
rect 8488 805 8522 837
rect 8488 735 8522 769
rect 8488 667 8522 699
rect 8488 599 8522 627
rect 8488 531 8522 555
rect 8488 463 8522 483
rect 8488 395 8522 411
rect 8488 327 8522 339
rect 8488 200 8522 267
rect 8584 1237 8618 1318
rect 8584 1165 8618 1177
rect 8584 1093 8618 1109
rect 8584 1021 8618 1041
rect 8584 949 8618 973
rect 8584 877 8618 905
rect 8584 805 8618 837
rect 8584 735 8618 769
rect 8584 667 8618 699
rect 8584 599 8618 627
rect 8584 531 8618 555
rect 8584 463 8618 483
rect 8584 395 8618 411
rect 8584 327 8618 339
rect 8584 250 8618 267
rect 8680 1237 8714 1256
rect 8680 1165 8714 1177
rect 8680 1093 8714 1109
rect 8680 1021 8714 1041
rect 8680 949 8714 973
rect 8680 877 8714 905
rect 8680 805 8714 837
rect 8680 735 8714 769
rect 8680 667 8714 699
rect 8680 599 8714 627
rect 8680 531 8714 555
rect 8680 463 8714 483
rect 8680 395 8714 411
rect 8680 327 8714 339
rect 8680 200 8714 267
rect 8776 1237 8810 1318
rect 8776 1165 8810 1177
rect 8776 1093 8810 1109
rect 8776 1021 8810 1041
rect 8776 949 8810 973
rect 8776 877 8810 905
rect 8776 805 8810 837
rect 8776 735 8810 769
rect 8776 667 8810 699
rect 8776 599 8810 627
rect 8776 531 8810 555
rect 8776 463 8810 483
rect 8776 395 8810 411
rect 8776 327 8810 339
rect 8776 250 8810 267
rect 8872 1237 8906 1256
rect 8872 1165 8906 1177
rect 8872 1093 8906 1109
rect 8872 1021 8906 1041
rect 8872 949 8906 973
rect 8872 877 8906 905
rect 8872 805 8906 837
rect 8872 735 8906 769
rect 8872 667 8906 699
rect 8872 599 8906 627
rect 8872 531 8906 555
rect 8872 463 8906 483
rect 8872 395 8906 411
rect 8872 327 8906 339
rect 8872 200 8906 267
rect 8968 1237 9002 1318
rect 9326 1294 10322 1328
rect 8968 1165 9002 1177
rect 8968 1093 9002 1109
rect 8968 1021 9002 1041
rect 8968 949 9002 973
rect 8968 877 9002 905
rect 8968 805 9002 837
rect 8968 735 9002 769
rect 8968 667 9002 699
rect 8968 599 9002 627
rect 8968 531 9002 555
rect 8968 463 9002 483
rect 8968 395 9002 411
rect 8968 327 9002 339
rect 8968 250 9002 267
rect 9232 1235 9266 1254
rect 9232 1163 9266 1175
rect 9232 1091 9266 1107
rect 9232 1019 9266 1039
rect 9232 947 9266 971
rect 9232 875 9266 903
rect 9232 803 9266 835
rect 9232 733 9266 767
rect 9232 665 9266 697
rect 9232 597 9266 625
rect 9232 529 9266 553
rect 9232 461 9266 481
rect 9232 393 9266 409
rect 9232 325 9266 337
rect 7912 166 8906 200
rect 9232 196 9266 265
rect 9328 1235 9362 1294
rect 9328 1163 9362 1175
rect 9328 1091 9362 1107
rect 9328 1019 9362 1039
rect 9328 947 9362 971
rect 9328 875 9362 903
rect 9328 803 9362 835
rect 9328 733 9362 767
rect 9328 665 9362 697
rect 9328 597 9362 625
rect 9328 529 9362 553
rect 9328 461 9362 481
rect 9328 393 9362 409
rect 9328 325 9362 337
rect 9328 246 9362 265
rect 9424 1235 9458 1252
rect 9424 1163 9458 1175
rect 9424 1091 9458 1107
rect 9424 1019 9458 1039
rect 9424 947 9458 971
rect 9424 875 9458 903
rect 9424 803 9458 835
rect 9424 733 9458 767
rect 9424 665 9458 697
rect 9424 597 9458 625
rect 9424 529 9458 553
rect 9424 461 9458 481
rect 9424 393 9458 409
rect 9424 325 9458 337
rect 9424 196 9458 265
rect 9520 1235 9554 1294
rect 9520 1163 9554 1175
rect 9520 1091 9554 1107
rect 9520 1019 9554 1039
rect 9520 947 9554 971
rect 9520 875 9554 903
rect 9520 803 9554 835
rect 9520 733 9554 767
rect 9520 665 9554 697
rect 9520 597 9554 625
rect 9520 529 9554 553
rect 9520 461 9554 481
rect 9520 393 9554 409
rect 9520 325 9554 337
rect 9520 246 9554 265
rect 9616 1235 9650 1252
rect 9616 1163 9650 1175
rect 9616 1091 9650 1107
rect 9616 1019 9650 1039
rect 9616 947 9650 971
rect 9616 875 9650 903
rect 9616 803 9650 835
rect 9616 733 9650 767
rect 9616 665 9650 697
rect 9616 597 9650 625
rect 9616 529 9650 553
rect 9616 461 9650 481
rect 9616 393 9650 409
rect 9616 325 9650 337
rect 9616 196 9650 265
rect 9712 1235 9746 1294
rect 9712 1163 9746 1175
rect 9712 1091 9746 1107
rect 9712 1019 9746 1039
rect 9712 947 9746 971
rect 9712 875 9746 903
rect 9712 803 9746 835
rect 9712 733 9746 767
rect 9712 665 9746 697
rect 9712 597 9746 625
rect 9712 529 9746 553
rect 9712 461 9746 481
rect 9712 393 9746 409
rect 9712 325 9746 337
rect 9712 246 9746 265
rect 9808 1235 9842 1252
rect 9808 1163 9842 1175
rect 9808 1091 9842 1107
rect 9808 1019 9842 1039
rect 9808 947 9842 971
rect 9808 875 9842 903
rect 9808 803 9842 835
rect 9808 733 9842 767
rect 9808 665 9842 697
rect 9808 597 9842 625
rect 9808 529 9842 553
rect 9808 461 9842 481
rect 9808 393 9842 409
rect 9808 325 9842 337
rect 9808 196 9842 265
rect 9904 1235 9938 1294
rect 9904 1163 9938 1175
rect 9904 1091 9938 1107
rect 9904 1019 9938 1039
rect 9904 947 9938 971
rect 9904 875 9938 903
rect 9904 803 9938 835
rect 9904 733 9938 767
rect 9904 665 9938 697
rect 9904 597 9938 625
rect 9904 529 9938 553
rect 9904 461 9938 481
rect 9904 393 9938 409
rect 9904 325 9938 337
rect 9904 246 9938 265
rect 10000 1235 10034 1252
rect 10000 1163 10034 1175
rect 10000 1091 10034 1107
rect 10000 1019 10034 1039
rect 10000 947 10034 971
rect 10000 875 10034 903
rect 10000 803 10034 835
rect 10000 733 10034 767
rect 10000 665 10034 697
rect 10000 597 10034 625
rect 10000 529 10034 553
rect 10000 461 10034 481
rect 10000 393 10034 409
rect 10000 325 10034 337
rect 10000 196 10034 265
rect 10096 1235 10130 1294
rect 10096 1163 10130 1175
rect 10096 1091 10130 1107
rect 10096 1019 10130 1039
rect 10096 947 10130 971
rect 10096 875 10130 903
rect 10096 803 10130 835
rect 10096 733 10130 767
rect 10096 665 10130 697
rect 10096 597 10130 625
rect 10096 529 10130 553
rect 10096 461 10130 481
rect 10096 393 10130 409
rect 10096 325 10130 337
rect 10096 246 10130 265
rect 10192 1235 10226 1252
rect 10192 1163 10226 1175
rect 10192 1091 10226 1107
rect 10192 1019 10226 1039
rect 10192 947 10226 971
rect 10192 875 10226 903
rect 10192 803 10226 835
rect 10192 733 10226 767
rect 10192 665 10226 697
rect 10192 597 10226 625
rect 10192 529 10226 553
rect 10192 461 10226 481
rect 10192 393 10226 409
rect 10192 325 10226 337
rect 10192 196 10226 265
rect 10288 1235 10322 1294
rect 10288 1163 10322 1175
rect 10288 1091 10322 1107
rect 10288 1019 10322 1039
rect 10288 947 10322 971
rect 10288 875 10322 903
rect 10288 803 10322 835
rect 10288 733 10322 767
rect 10288 665 10322 697
rect 10288 597 10322 625
rect 10288 529 10322 553
rect 10288 461 10322 481
rect 10288 393 10322 409
rect 10288 325 10322 337
rect 10288 248 10322 265
rect 10384 1235 10418 1252
rect 10384 1163 10418 1175
rect 10384 1091 10418 1107
rect 10384 1019 10418 1039
rect 10384 947 10418 971
rect 10384 875 10418 903
rect 10384 803 10418 835
rect 10384 733 10418 767
rect 10384 665 10418 697
rect 10384 597 10418 625
rect 10384 529 10418 553
rect 10384 461 10418 481
rect 10384 393 10418 409
rect 10384 325 10418 337
rect 10384 196 10418 265
rect 8480 130 8514 166
rect 9232 162 10418 196
rect 8758 80 8774 114
rect 8808 80 8824 114
rect 9214 78 9230 112
rect 9264 78 9280 112
rect 9904 102 9938 162
rect 4656 13 4708 16
rect -2026 -106 722 -18
rect 4656 -21 4665 13
rect 4699 -21 4708 13
rect 4656 -24 4708 -21
rect 7656 15 7708 18
rect 7656 -19 7665 15
rect 7699 -19 7708 15
rect 10664 14 10698 1464
rect 14152 1448 14186 1604
rect 15450 1458 15466 1492
rect 15500 1458 15516 1492
rect 13964 1414 14186 1448
rect 11474 1350 11508 1400
rect 11096 1316 12090 1350
rect 11000 1235 11034 1254
rect 11000 1163 11034 1175
rect 11000 1091 11034 1107
rect 11000 1019 11034 1039
rect 11000 947 11034 971
rect 11000 875 11034 903
rect 11000 803 11034 835
rect 11000 733 11034 767
rect 11000 665 11034 697
rect 11000 597 11034 625
rect 11000 529 11034 553
rect 11000 461 11034 481
rect 11000 393 11034 409
rect 11000 325 11034 337
rect 11000 198 11034 265
rect 11096 1235 11130 1316
rect 11096 1163 11130 1175
rect 11096 1091 11130 1107
rect 11096 1019 11130 1039
rect 11096 947 11130 971
rect 11096 875 11130 903
rect 11096 803 11130 835
rect 11096 733 11130 767
rect 11096 665 11130 697
rect 11096 597 11130 625
rect 11096 529 11130 553
rect 11096 461 11130 481
rect 11096 393 11130 409
rect 11096 325 11130 337
rect 11096 246 11130 265
rect 11192 1235 11226 1254
rect 11192 1163 11226 1175
rect 11192 1091 11226 1107
rect 11192 1019 11226 1039
rect 11192 947 11226 971
rect 11192 875 11226 903
rect 11192 803 11226 835
rect 11192 733 11226 767
rect 11192 665 11226 697
rect 11192 597 11226 625
rect 11192 529 11226 553
rect 11192 461 11226 481
rect 11192 393 11226 409
rect 11192 325 11226 337
rect 11192 198 11226 265
rect 11288 1235 11322 1316
rect 11288 1163 11322 1175
rect 11288 1091 11322 1107
rect 11288 1019 11322 1039
rect 11288 947 11322 971
rect 11288 875 11322 903
rect 11288 803 11322 835
rect 11288 733 11322 767
rect 11288 665 11322 697
rect 11288 597 11322 625
rect 11288 529 11322 553
rect 11288 461 11322 481
rect 11288 393 11322 409
rect 11288 325 11322 337
rect 11288 246 11322 265
rect 11384 1235 11418 1254
rect 11384 1163 11418 1175
rect 11384 1091 11418 1107
rect 11384 1019 11418 1039
rect 11384 947 11418 971
rect 11384 875 11418 903
rect 11384 803 11418 835
rect 11384 733 11418 767
rect 11384 665 11418 697
rect 11384 597 11418 625
rect 11384 529 11418 553
rect 11384 461 11418 481
rect 11384 393 11418 409
rect 11384 325 11418 337
rect 11384 198 11418 265
rect 11480 1235 11514 1316
rect 11480 1163 11514 1175
rect 11480 1091 11514 1107
rect 11480 1019 11514 1039
rect 11480 947 11514 971
rect 11480 875 11514 903
rect 11480 803 11514 835
rect 11480 733 11514 767
rect 11480 665 11514 697
rect 11480 597 11514 625
rect 11480 529 11514 553
rect 11480 461 11514 481
rect 11480 393 11514 409
rect 11480 325 11514 337
rect 11480 246 11514 265
rect 11576 1235 11610 1254
rect 11576 1163 11610 1175
rect 11576 1091 11610 1107
rect 11576 1019 11610 1039
rect 11576 947 11610 971
rect 11576 875 11610 903
rect 11576 803 11610 835
rect 11576 733 11610 767
rect 11576 665 11610 697
rect 11576 597 11610 625
rect 11576 529 11610 553
rect 11576 461 11610 481
rect 11576 393 11610 409
rect 11576 325 11610 337
rect 11576 198 11610 265
rect 11672 1235 11706 1316
rect 11672 1163 11706 1175
rect 11672 1091 11706 1107
rect 11672 1019 11706 1039
rect 11672 947 11706 971
rect 11672 875 11706 903
rect 11672 803 11706 835
rect 11672 733 11706 767
rect 11672 665 11706 697
rect 11672 597 11706 625
rect 11672 529 11706 553
rect 11672 461 11706 481
rect 11672 393 11706 409
rect 11672 325 11706 337
rect 11672 248 11706 265
rect 11768 1235 11802 1254
rect 11768 1163 11802 1175
rect 11768 1091 11802 1107
rect 11768 1019 11802 1039
rect 11768 947 11802 971
rect 11768 875 11802 903
rect 11768 803 11802 835
rect 11768 733 11802 767
rect 11768 665 11802 697
rect 11768 597 11802 625
rect 11768 529 11802 553
rect 11768 461 11802 481
rect 11768 393 11802 409
rect 11768 325 11802 337
rect 11768 198 11802 265
rect 11864 1235 11898 1316
rect 11864 1163 11898 1175
rect 11864 1091 11898 1107
rect 11864 1019 11898 1039
rect 11864 947 11898 971
rect 11864 875 11898 903
rect 11864 803 11898 835
rect 11864 733 11898 767
rect 11864 665 11898 697
rect 11864 597 11898 625
rect 11864 529 11898 553
rect 11864 461 11898 481
rect 11864 393 11898 409
rect 11864 325 11898 337
rect 11864 248 11898 265
rect 11960 1235 11994 1254
rect 11960 1163 11994 1175
rect 11960 1091 11994 1107
rect 11960 1019 11994 1039
rect 11960 947 11994 971
rect 11960 875 11994 903
rect 11960 803 11994 835
rect 11960 733 11994 767
rect 11960 665 11994 697
rect 11960 597 11994 625
rect 11960 529 11994 553
rect 11960 461 11994 481
rect 11960 393 11994 409
rect 11960 325 11994 337
rect 11960 198 11994 265
rect 12056 1235 12090 1316
rect 12964 1302 12998 1380
rect 12482 1268 13478 1302
rect 12056 1163 12090 1175
rect 12056 1091 12090 1107
rect 12056 1019 12090 1039
rect 12056 947 12090 971
rect 12056 875 12090 903
rect 12056 803 12090 835
rect 12056 733 12090 767
rect 12056 665 12090 697
rect 12056 597 12090 625
rect 12056 529 12090 553
rect 12056 461 12090 481
rect 12056 393 12090 409
rect 12056 325 12090 337
rect 12056 248 12090 265
rect 12388 1209 12422 1228
rect 12388 1137 12422 1149
rect 12388 1065 12422 1081
rect 12388 993 12422 1013
rect 12388 921 12422 945
rect 12388 849 12422 877
rect 12388 777 12422 809
rect 12388 707 12422 741
rect 12388 639 12422 671
rect 12388 571 12422 599
rect 12388 503 12422 527
rect 12388 435 12422 455
rect 12388 367 12422 383
rect 12388 299 12422 311
rect 11000 164 11994 198
rect 12388 170 12422 239
rect 12484 1209 12518 1268
rect 12484 1137 12518 1149
rect 12484 1065 12518 1081
rect 12484 993 12518 1013
rect 12484 921 12518 945
rect 12484 849 12518 877
rect 12484 777 12518 809
rect 12484 707 12518 741
rect 12484 639 12518 671
rect 12484 571 12518 599
rect 12484 503 12518 527
rect 12484 435 12518 455
rect 12484 367 12518 383
rect 12484 299 12518 311
rect 12484 220 12518 239
rect 12580 1209 12614 1226
rect 12580 1137 12614 1149
rect 12580 1065 12614 1081
rect 12580 993 12614 1013
rect 12580 921 12614 945
rect 12580 849 12614 877
rect 12580 777 12614 809
rect 12580 707 12614 741
rect 12580 639 12614 671
rect 12580 571 12614 599
rect 12580 503 12614 527
rect 12580 435 12614 455
rect 12580 367 12614 383
rect 12580 299 12614 311
rect 12580 170 12614 239
rect 12676 1209 12710 1268
rect 12676 1137 12710 1149
rect 12676 1065 12710 1081
rect 12676 993 12710 1013
rect 12676 921 12710 945
rect 12676 849 12710 877
rect 12676 777 12710 809
rect 12676 707 12710 741
rect 12676 639 12710 671
rect 12676 571 12710 599
rect 12676 503 12710 527
rect 12676 435 12710 455
rect 12676 367 12710 383
rect 12676 299 12710 311
rect 12676 220 12710 239
rect 12772 1209 12806 1226
rect 12772 1137 12806 1149
rect 12772 1065 12806 1081
rect 12772 993 12806 1013
rect 12772 921 12806 945
rect 12772 849 12806 877
rect 12772 777 12806 809
rect 12772 707 12806 741
rect 12772 639 12806 671
rect 12772 571 12806 599
rect 12772 503 12806 527
rect 12772 435 12806 455
rect 12772 367 12806 383
rect 12772 299 12806 311
rect 12772 170 12806 239
rect 12868 1209 12902 1268
rect 12868 1137 12902 1149
rect 12868 1065 12902 1081
rect 12868 993 12902 1013
rect 12868 921 12902 945
rect 12868 849 12902 877
rect 12868 777 12902 809
rect 12868 707 12902 741
rect 12868 639 12902 671
rect 12868 571 12902 599
rect 12868 503 12902 527
rect 12868 435 12902 455
rect 12868 367 12902 383
rect 12868 299 12902 311
rect 12868 220 12902 239
rect 12964 1209 12998 1226
rect 12964 1137 12998 1149
rect 12964 1065 12998 1081
rect 12964 993 12998 1013
rect 12964 921 12998 945
rect 12964 849 12998 877
rect 12964 777 12998 809
rect 12964 707 12998 741
rect 12964 639 12998 671
rect 12964 571 12998 599
rect 12964 503 12998 527
rect 12964 435 12998 455
rect 12964 367 12998 383
rect 12964 299 12998 311
rect 12964 170 12998 239
rect 13060 1209 13094 1268
rect 13060 1137 13094 1149
rect 13060 1065 13094 1081
rect 13060 993 13094 1013
rect 13060 921 13094 945
rect 13060 849 13094 877
rect 13060 777 13094 809
rect 13060 707 13094 741
rect 13060 639 13094 671
rect 13060 571 13094 599
rect 13060 503 13094 527
rect 13060 435 13094 455
rect 13060 367 13094 383
rect 13060 299 13094 311
rect 13060 220 13094 239
rect 13156 1209 13190 1226
rect 13156 1137 13190 1149
rect 13156 1065 13190 1081
rect 13156 993 13190 1013
rect 13156 921 13190 945
rect 13156 849 13190 877
rect 13156 777 13190 809
rect 13156 707 13190 741
rect 13156 639 13190 671
rect 13156 571 13190 599
rect 13156 503 13190 527
rect 13156 435 13190 455
rect 13156 367 13190 383
rect 13156 299 13190 311
rect 13156 170 13190 239
rect 13252 1209 13286 1268
rect 13252 1137 13286 1149
rect 13252 1065 13286 1081
rect 13252 993 13286 1013
rect 13252 921 13286 945
rect 13252 849 13286 877
rect 13252 777 13286 809
rect 13252 707 13286 741
rect 13252 639 13286 671
rect 13252 571 13286 599
rect 13252 503 13286 527
rect 13252 435 13286 455
rect 13252 367 13286 383
rect 13252 299 13286 311
rect 13252 220 13286 239
rect 13348 1209 13382 1226
rect 13348 1137 13382 1149
rect 13348 1065 13382 1081
rect 13348 993 13382 1013
rect 13348 921 13382 945
rect 13348 849 13382 877
rect 13348 777 13382 809
rect 13348 707 13382 741
rect 13348 639 13382 671
rect 13348 571 13382 599
rect 13348 503 13382 527
rect 13348 435 13382 455
rect 13348 367 13382 383
rect 13348 299 13382 311
rect 13348 170 13382 239
rect 13444 1209 13478 1268
rect 13444 1137 13478 1149
rect 13444 1065 13478 1081
rect 13444 993 13478 1013
rect 13444 921 13478 945
rect 13444 849 13478 877
rect 13444 777 13478 809
rect 13444 707 13478 741
rect 13444 639 13478 671
rect 13444 571 13478 599
rect 13444 503 13478 527
rect 13444 435 13478 455
rect 13444 367 13478 383
rect 13444 299 13478 311
rect 13444 222 13478 239
rect 13540 1209 13574 1226
rect 13540 1137 13574 1149
rect 13540 1065 13574 1081
rect 13540 993 13574 1013
rect 13540 921 13574 945
rect 13540 849 13574 877
rect 13540 777 13574 809
rect 13540 707 13574 741
rect 13540 639 13574 671
rect 13540 571 13574 599
rect 13540 503 13574 527
rect 13540 435 13574 455
rect 13540 367 13574 383
rect 13540 299 13574 311
rect 13540 170 13574 239
rect 11568 128 11602 164
rect 12388 136 13574 170
rect 11846 78 11862 112
rect 11896 78 11912 112
rect 12370 52 12386 86
rect 12420 52 12436 86
rect 13060 76 13094 136
rect 7656 -22 7708 -19
rect 10654 11 10706 14
rect 10654 -23 10663 11
rect 10697 -23 10706 11
rect 13964 -12 13998 1414
rect 14630 1324 14664 1374
rect 14252 1290 15246 1324
rect 14156 1209 14190 1228
rect 14156 1137 14190 1149
rect 14156 1065 14190 1081
rect 14156 993 14190 1013
rect 14156 921 14190 945
rect 14156 849 14190 877
rect 14156 777 14190 809
rect 14156 707 14190 741
rect 14156 639 14190 671
rect 14156 571 14190 599
rect 14156 503 14190 527
rect 14156 435 14190 455
rect 14156 367 14190 383
rect 14156 299 14190 311
rect 14156 172 14190 239
rect 14252 1209 14286 1290
rect 14252 1137 14286 1149
rect 14252 1065 14286 1081
rect 14252 993 14286 1013
rect 14252 921 14286 945
rect 14252 849 14286 877
rect 14252 777 14286 809
rect 14252 707 14286 741
rect 14252 639 14286 671
rect 14252 571 14286 599
rect 14252 503 14286 527
rect 14252 435 14286 455
rect 14252 367 14286 383
rect 14252 299 14286 311
rect 14252 220 14286 239
rect 14348 1209 14382 1228
rect 14348 1137 14382 1149
rect 14348 1065 14382 1081
rect 14348 993 14382 1013
rect 14348 921 14382 945
rect 14348 849 14382 877
rect 14348 777 14382 809
rect 14348 707 14382 741
rect 14348 639 14382 671
rect 14348 571 14382 599
rect 14348 503 14382 527
rect 14348 435 14382 455
rect 14348 367 14382 383
rect 14348 299 14382 311
rect 14348 172 14382 239
rect 14444 1209 14478 1290
rect 14444 1137 14478 1149
rect 14444 1065 14478 1081
rect 14444 993 14478 1013
rect 14444 921 14478 945
rect 14444 849 14478 877
rect 14444 777 14478 809
rect 14444 707 14478 741
rect 14444 639 14478 671
rect 14444 571 14478 599
rect 14444 503 14478 527
rect 14444 435 14478 455
rect 14444 367 14478 383
rect 14444 299 14478 311
rect 14444 220 14478 239
rect 14540 1209 14574 1228
rect 14540 1137 14574 1149
rect 14540 1065 14574 1081
rect 14540 993 14574 1013
rect 14540 921 14574 945
rect 14540 849 14574 877
rect 14540 777 14574 809
rect 14540 707 14574 741
rect 14540 639 14574 671
rect 14540 571 14574 599
rect 14540 503 14574 527
rect 14540 435 14574 455
rect 14540 367 14574 383
rect 14540 299 14574 311
rect 14540 172 14574 239
rect 14636 1209 14670 1290
rect 14636 1137 14670 1149
rect 14636 1065 14670 1081
rect 14636 993 14670 1013
rect 14636 921 14670 945
rect 14636 849 14670 877
rect 14636 777 14670 809
rect 14636 707 14670 741
rect 14636 639 14670 671
rect 14636 571 14670 599
rect 14636 503 14670 527
rect 14636 435 14670 455
rect 14636 367 14670 383
rect 14636 299 14670 311
rect 14636 220 14670 239
rect 14732 1209 14766 1228
rect 14732 1137 14766 1149
rect 14732 1065 14766 1081
rect 14732 993 14766 1013
rect 14732 921 14766 945
rect 14732 849 14766 877
rect 14732 777 14766 809
rect 14732 707 14766 741
rect 14732 639 14766 671
rect 14732 571 14766 599
rect 14732 503 14766 527
rect 14732 435 14766 455
rect 14732 367 14766 383
rect 14732 299 14766 311
rect 14732 172 14766 239
rect 14828 1209 14862 1290
rect 14828 1137 14862 1149
rect 14828 1065 14862 1081
rect 14828 993 14862 1013
rect 14828 921 14862 945
rect 14828 849 14862 877
rect 14828 777 14862 809
rect 14828 707 14862 741
rect 14828 639 14862 671
rect 14828 571 14862 599
rect 14828 503 14862 527
rect 14828 435 14862 455
rect 14828 367 14862 383
rect 14828 299 14862 311
rect 14828 222 14862 239
rect 14924 1209 14958 1228
rect 14924 1137 14958 1149
rect 14924 1065 14958 1081
rect 14924 993 14958 1013
rect 14924 921 14958 945
rect 14924 849 14958 877
rect 14924 777 14958 809
rect 14924 707 14958 741
rect 14924 639 14958 671
rect 14924 571 14958 599
rect 14924 503 14958 527
rect 14924 435 14958 455
rect 14924 367 14958 383
rect 14924 299 14958 311
rect 14924 172 14958 239
rect 15020 1209 15054 1290
rect 15020 1137 15054 1149
rect 15020 1065 15054 1081
rect 15020 993 15054 1013
rect 15020 921 15054 945
rect 15020 849 15054 877
rect 15020 777 15054 809
rect 15020 707 15054 741
rect 15020 639 15054 671
rect 15020 571 15054 599
rect 15020 503 15054 527
rect 15020 435 15054 455
rect 15020 367 15054 383
rect 15020 299 15054 311
rect 15020 222 15054 239
rect 15116 1209 15150 1228
rect 15116 1137 15150 1149
rect 15116 1065 15150 1081
rect 15116 993 15150 1013
rect 15116 921 15150 945
rect 15116 849 15150 877
rect 15116 777 15150 809
rect 15116 707 15150 741
rect 15116 639 15150 671
rect 15116 571 15150 599
rect 15116 503 15150 527
rect 15116 435 15150 455
rect 15116 367 15150 383
rect 15116 299 15150 311
rect 15116 172 15150 239
rect 15212 1209 15246 1290
rect 15212 1137 15246 1149
rect 15212 1065 15246 1081
rect 15212 993 15246 1013
rect 15212 921 15246 945
rect 15212 849 15246 877
rect 15212 777 15246 809
rect 15212 707 15246 741
rect 15212 639 15246 671
rect 15212 571 15246 599
rect 15212 503 15246 527
rect 15212 435 15246 455
rect 15212 367 15246 383
rect 15212 299 15246 311
rect 15212 222 15246 239
rect 15422 1261 15456 1336
rect 15422 1193 15456 1223
rect 15422 1125 15456 1151
rect 15422 1057 15456 1079
rect 15422 989 15456 1007
rect 15422 921 15456 935
rect 15422 853 15456 863
rect 15422 785 15456 791
rect 15422 717 15456 719
rect 15422 681 15456 683
rect 15422 609 15456 615
rect 15422 537 15456 547
rect 15422 465 15456 479
rect 15422 393 15456 411
rect 15422 321 15456 343
rect 15422 249 15456 275
rect 14156 138 15150 172
rect 15422 177 15456 207
rect 14724 102 14758 138
rect 15422 96 15456 139
rect 15510 1261 15544 1304
rect 15510 1193 15544 1223
rect 15510 1125 15544 1151
rect 15510 1057 15544 1079
rect 15510 989 15544 1007
rect 15510 921 15544 935
rect 15510 853 15544 863
rect 15510 785 15544 791
rect 15510 717 15544 719
rect 15510 681 15544 683
rect 15510 609 15544 615
rect 15510 537 15544 547
rect 15510 465 15544 479
rect 15510 393 15544 411
rect 15510 321 15544 343
rect 15510 249 15544 275
rect 15510 177 15544 207
rect 15002 52 15018 86
rect 15052 52 15068 86
rect 15510 52 15544 139
rect 15510 16 15544 18
rect 10654 -26 10706 -23
rect 13956 -15 14008 -12
rect 13956 -49 13965 -15
rect 13999 -49 14008 -15
rect 13956 -52 14008 -49
rect 13964 -56 13998 -52
<< viali >>
rect 764 6858 798 6892
rect 288 6773 322 6807
rect 3720 6842 3754 6876
rect 2440 6754 2474 6788
rect 2728 6769 2762 6803
rect 3244 6757 3278 6791
rect 6750 6842 6784 6876
rect 5396 6738 5430 6772
rect 5684 6753 5718 6787
rect 6274 6757 6308 6791
rect 194 6565 228 6591
rect 194 6557 228 6565
rect 194 6497 228 6519
rect 194 6485 228 6497
rect 194 6429 228 6447
rect 194 6413 228 6429
rect 194 6361 228 6375
rect 194 6341 228 6361
rect 194 6293 228 6303
rect 194 6269 228 6293
rect 194 6225 228 6231
rect 194 6197 228 6225
rect 194 6157 228 6159
rect 194 6125 228 6157
rect 194 6055 228 6087
rect 194 6053 228 6055
rect -1652 5895 -1618 5921
rect -1652 5887 -1618 5895
rect -1652 5827 -1618 5849
rect -1652 5815 -1618 5827
rect -1652 5759 -1618 5777
rect -1652 5743 -1618 5759
rect -1652 5691 -1618 5705
rect -1652 5671 -1618 5691
rect -1652 5623 -1618 5633
rect -1652 5599 -1618 5623
rect -1652 5555 -1618 5561
rect -1652 5527 -1618 5555
rect -1652 5487 -1618 5489
rect -1652 5455 -1618 5487
rect -1652 5385 -1618 5417
rect -1652 5383 -1618 5385
rect -1652 5317 -1618 5345
rect -1652 5311 -1618 5317
rect -1652 5249 -1618 5273
rect -1652 5239 -1618 5249
rect -1652 5181 -1618 5201
rect -1652 5167 -1618 5181
rect -1652 5113 -1618 5129
rect -1652 5095 -1618 5113
rect -1652 5045 -1618 5057
rect -1652 5023 -1618 5045
rect -1652 4977 -1618 4985
rect -1652 4951 -1618 4977
rect -1554 5895 -1520 5921
rect -1554 5887 -1520 5895
rect -1554 5827 -1520 5849
rect -1554 5815 -1520 5827
rect -1554 5759 -1520 5777
rect -1554 5743 -1520 5759
rect -1554 5691 -1520 5705
rect -1554 5671 -1520 5691
rect -1554 5623 -1520 5633
rect -1554 5599 -1520 5623
rect -1554 5555 -1520 5561
rect -1554 5527 -1520 5555
rect -1554 5487 -1520 5489
rect -1554 5455 -1520 5487
rect -1554 5385 -1520 5417
rect -1554 5383 -1520 5385
rect -1554 5317 -1520 5345
rect -1554 5311 -1520 5317
rect -1554 5249 -1520 5273
rect -1554 5239 -1520 5249
rect -1554 5181 -1520 5201
rect -1554 5167 -1520 5181
rect -1554 5113 -1520 5129
rect -1554 5095 -1520 5113
rect -1554 5045 -1520 5057
rect -1554 5023 -1520 5045
rect -1554 4977 -1520 4985
rect -1554 4951 -1520 4977
rect -1456 5895 -1422 5921
rect -1456 5887 -1422 5895
rect -1456 5827 -1422 5849
rect -1456 5815 -1422 5827
rect -1456 5759 -1422 5777
rect -1456 5743 -1422 5759
rect -1456 5691 -1422 5705
rect -1456 5671 -1422 5691
rect -1456 5623 -1422 5633
rect -1456 5599 -1422 5623
rect -1456 5555 -1422 5561
rect -1456 5527 -1422 5555
rect -1456 5487 -1422 5489
rect -1456 5455 -1422 5487
rect -1456 5385 -1422 5417
rect -1456 5383 -1422 5385
rect -1456 5317 -1422 5345
rect -1456 5311 -1422 5317
rect -1456 5249 -1422 5273
rect -1456 5239 -1422 5249
rect -1456 5181 -1422 5201
rect -1456 5167 -1422 5181
rect -1456 5113 -1422 5129
rect -1456 5095 -1422 5113
rect -1456 5045 -1422 5057
rect -1456 5023 -1422 5045
rect -1456 4977 -1422 4985
rect -1456 4951 -1422 4977
rect -1358 5895 -1324 5921
rect -1358 5887 -1324 5895
rect -1358 5827 -1324 5849
rect -1358 5815 -1324 5827
rect -1358 5759 -1324 5777
rect -1358 5743 -1324 5759
rect -1358 5691 -1324 5705
rect -1358 5671 -1324 5691
rect -1358 5623 -1324 5633
rect -1358 5599 -1324 5623
rect -1358 5555 -1324 5561
rect -1358 5527 -1324 5555
rect -1358 5487 -1324 5489
rect -1358 5455 -1324 5487
rect -1358 5385 -1324 5417
rect -1358 5383 -1324 5385
rect -1358 5317 -1324 5345
rect -1358 5311 -1324 5317
rect -1358 5249 -1324 5273
rect -1358 5239 -1324 5249
rect -1358 5181 -1324 5201
rect -1358 5167 -1324 5181
rect -1358 5113 -1324 5129
rect -1358 5095 -1324 5113
rect -1358 5045 -1324 5057
rect -1358 5023 -1324 5045
rect -1358 4977 -1324 4985
rect -1358 4951 -1324 4977
rect -1260 5895 -1226 5921
rect -1260 5887 -1226 5895
rect -1260 5827 -1226 5849
rect -1260 5815 -1226 5827
rect -1260 5759 -1226 5777
rect -1260 5743 -1226 5759
rect -1260 5691 -1226 5705
rect -1260 5671 -1226 5691
rect -1260 5623 -1226 5633
rect -1260 5599 -1226 5623
rect -1260 5555 -1226 5561
rect -1260 5527 -1226 5555
rect -1260 5487 -1226 5489
rect -1260 5455 -1226 5487
rect -1260 5385 -1226 5417
rect -1260 5383 -1226 5385
rect -1260 5317 -1226 5345
rect -1260 5311 -1226 5317
rect -1260 5249 -1226 5273
rect -1260 5239 -1226 5249
rect -1260 5181 -1226 5201
rect -1260 5167 -1226 5181
rect -1260 5113 -1226 5129
rect -1260 5095 -1226 5113
rect -1260 5045 -1226 5057
rect -1260 5023 -1226 5045
rect -1260 4977 -1226 4985
rect -1260 4951 -1226 4977
rect -1162 5895 -1128 5921
rect -1162 5887 -1128 5895
rect -1162 5827 -1128 5849
rect -1162 5815 -1128 5827
rect -1162 5759 -1128 5777
rect -1162 5743 -1128 5759
rect -1162 5691 -1128 5705
rect -1162 5671 -1128 5691
rect -1162 5623 -1128 5633
rect -1162 5599 -1128 5623
rect -1162 5555 -1128 5561
rect -1162 5527 -1128 5555
rect -1162 5487 -1128 5489
rect -1162 5455 -1128 5487
rect -1162 5385 -1128 5417
rect -1162 5383 -1128 5385
rect -1162 5317 -1128 5345
rect -1162 5311 -1128 5317
rect -1162 5249 -1128 5273
rect -1162 5239 -1128 5249
rect -1162 5181 -1128 5201
rect -1162 5167 -1128 5181
rect -1162 5113 -1128 5129
rect -1162 5095 -1128 5113
rect -1162 5045 -1128 5057
rect -1162 5023 -1128 5045
rect -1162 4977 -1128 4985
rect -1162 4951 -1128 4977
rect -1064 5895 -1030 5921
rect -1064 5887 -1030 5895
rect -1064 5827 -1030 5849
rect -1064 5815 -1030 5827
rect -1064 5759 -1030 5777
rect -1064 5743 -1030 5759
rect -1064 5691 -1030 5705
rect -1064 5671 -1030 5691
rect -1064 5623 -1030 5633
rect -1064 5599 -1030 5623
rect -1064 5555 -1030 5561
rect -1064 5527 -1030 5555
rect -1064 5487 -1030 5489
rect -1064 5455 -1030 5487
rect -1064 5385 -1030 5417
rect -1064 5383 -1030 5385
rect -1064 5317 -1030 5345
rect -1064 5311 -1030 5317
rect -1064 5249 -1030 5273
rect -1064 5239 -1030 5249
rect -1064 5181 -1030 5201
rect -1064 5167 -1030 5181
rect -1064 5113 -1030 5129
rect -1064 5095 -1030 5113
rect -1064 5045 -1030 5057
rect -1064 5023 -1030 5045
rect -1064 4977 -1030 4985
rect -1064 4951 -1030 4977
rect -966 5895 -932 5921
rect -966 5887 -932 5895
rect -966 5827 -932 5849
rect -966 5815 -932 5827
rect -966 5759 -932 5777
rect -966 5743 -932 5759
rect -966 5691 -932 5705
rect -966 5671 -932 5691
rect -966 5623 -932 5633
rect -966 5599 -932 5623
rect -966 5555 -932 5561
rect -966 5527 -932 5555
rect -966 5487 -932 5489
rect -966 5455 -932 5487
rect -966 5385 -932 5417
rect -966 5383 -932 5385
rect -966 5317 -932 5345
rect -966 5311 -932 5317
rect -966 5249 -932 5273
rect -966 5239 -932 5249
rect -966 5181 -932 5201
rect -966 5167 -932 5181
rect -966 5113 -932 5129
rect -966 5095 -932 5113
rect -966 5045 -932 5057
rect -966 5023 -932 5045
rect -966 4977 -932 4985
rect -966 4951 -932 4977
rect -868 5895 -834 5921
rect -868 5887 -834 5895
rect -868 5827 -834 5849
rect -868 5815 -834 5827
rect -868 5759 -834 5777
rect -868 5743 -834 5759
rect -868 5691 -834 5705
rect -868 5671 -834 5691
rect -868 5623 -834 5633
rect -868 5599 -834 5623
rect 194 5987 228 6015
rect 194 5981 228 5987
rect 194 5919 228 5943
rect 194 5909 228 5919
rect 194 5851 228 5871
rect 194 5837 228 5851
rect 194 5783 228 5799
rect 194 5765 228 5783
rect 194 5715 228 5727
rect 194 5693 228 5715
rect 194 5647 228 5655
rect 194 5621 228 5647
rect 290 6565 324 6591
rect 290 6557 324 6565
rect 290 6497 324 6519
rect 290 6485 324 6497
rect 290 6429 324 6447
rect 290 6413 324 6429
rect 290 6361 324 6375
rect 290 6341 324 6361
rect 290 6293 324 6303
rect 290 6269 324 6293
rect 290 6225 324 6231
rect 290 6197 324 6225
rect 290 6157 324 6159
rect 290 6125 324 6157
rect 290 6055 324 6087
rect 290 6053 324 6055
rect 290 5987 324 6015
rect 290 5981 324 5987
rect 290 5919 324 5943
rect 290 5909 324 5919
rect 290 5851 324 5871
rect 290 5837 324 5851
rect 290 5783 324 5799
rect 290 5765 324 5783
rect 290 5715 324 5727
rect 290 5693 324 5715
rect 290 5647 324 5655
rect 290 5621 324 5647
rect -868 5555 -834 5561
rect -868 5527 -834 5555
rect 386 6565 420 6591
rect 386 6557 420 6565
rect 386 6497 420 6519
rect 386 6485 420 6497
rect 386 6429 420 6447
rect 386 6413 420 6429
rect 386 6361 420 6375
rect 386 6341 420 6361
rect 386 6293 420 6303
rect 386 6269 420 6293
rect 386 6225 420 6231
rect 386 6197 420 6225
rect 386 6157 420 6159
rect 386 6125 420 6157
rect 386 6055 420 6087
rect 386 6053 420 6055
rect 386 5987 420 6015
rect 386 5981 420 5987
rect 386 5919 420 5943
rect 386 5909 420 5919
rect 386 5851 420 5871
rect 386 5837 420 5851
rect 386 5783 420 5799
rect 386 5765 420 5783
rect 386 5715 420 5727
rect 386 5693 420 5715
rect 386 5647 420 5655
rect 386 5621 420 5647
rect 482 6565 516 6591
rect 482 6557 516 6565
rect 482 6497 516 6519
rect 482 6485 516 6497
rect 482 6429 516 6447
rect 482 6413 516 6429
rect 482 6361 516 6375
rect 482 6341 516 6361
rect 482 6293 516 6303
rect 482 6269 516 6293
rect 482 6225 516 6231
rect 482 6197 516 6225
rect 482 6157 516 6159
rect 482 6125 516 6157
rect 482 6055 516 6087
rect 482 6053 516 6055
rect 482 5987 516 6015
rect 482 5981 516 5987
rect 482 5919 516 5943
rect 482 5909 516 5919
rect 482 5851 516 5871
rect 482 5837 516 5851
rect 482 5783 516 5799
rect 482 5765 516 5783
rect 482 5715 516 5727
rect 482 5693 516 5715
rect 482 5647 516 5655
rect 482 5621 516 5647
rect 578 6565 612 6591
rect 578 6557 612 6565
rect 578 6497 612 6519
rect 578 6485 612 6497
rect 578 6429 612 6447
rect 578 6413 612 6429
rect 578 6361 612 6375
rect 578 6341 612 6361
rect 578 6293 612 6303
rect 578 6269 612 6293
rect 578 6225 612 6231
rect 578 6197 612 6225
rect 578 6157 612 6159
rect 578 6125 612 6157
rect 578 6055 612 6087
rect 578 6053 612 6055
rect 578 5987 612 6015
rect 578 5981 612 5987
rect 578 5919 612 5943
rect 578 5909 612 5919
rect 578 5851 612 5871
rect 578 5837 612 5851
rect 578 5783 612 5799
rect 578 5765 612 5783
rect 578 5715 612 5727
rect 578 5693 612 5715
rect 578 5647 612 5655
rect 578 5621 612 5647
rect 674 6565 708 6591
rect 674 6557 708 6565
rect 674 6497 708 6519
rect 674 6485 708 6497
rect 674 6429 708 6447
rect 674 6413 708 6429
rect 674 6361 708 6375
rect 674 6341 708 6361
rect 674 6293 708 6303
rect 674 6269 708 6293
rect 674 6225 708 6231
rect 674 6197 708 6225
rect 674 6157 708 6159
rect 674 6125 708 6157
rect 674 6055 708 6087
rect 674 6053 708 6055
rect 674 5987 708 6015
rect 674 5981 708 5987
rect 674 5919 708 5943
rect 674 5909 708 5919
rect 674 5851 708 5871
rect 674 5837 708 5851
rect 674 5783 708 5799
rect 674 5765 708 5783
rect 674 5715 708 5727
rect 674 5693 708 5715
rect 674 5647 708 5655
rect 674 5621 708 5647
rect 770 6565 804 6591
rect 770 6557 804 6565
rect 770 6497 804 6519
rect 770 6485 804 6497
rect 770 6429 804 6447
rect 770 6413 804 6429
rect 770 6361 804 6375
rect 770 6341 804 6361
rect 770 6293 804 6303
rect 770 6269 804 6293
rect 770 6225 804 6231
rect 770 6197 804 6225
rect 770 6157 804 6159
rect 770 6125 804 6157
rect 770 6055 804 6087
rect 770 6053 804 6055
rect 770 5987 804 6015
rect 770 5981 804 5987
rect 770 5919 804 5943
rect 770 5909 804 5919
rect 770 5851 804 5871
rect 770 5837 804 5851
rect 770 5783 804 5799
rect 770 5765 804 5783
rect 770 5715 804 5727
rect 770 5693 804 5715
rect 770 5647 804 5655
rect 770 5621 804 5647
rect 866 6565 900 6591
rect 866 6557 900 6565
rect 866 6497 900 6519
rect 866 6485 900 6497
rect 866 6429 900 6447
rect 866 6413 900 6429
rect 866 6361 900 6375
rect 866 6341 900 6361
rect 866 6293 900 6303
rect 866 6269 900 6293
rect 866 6225 900 6231
rect 866 6197 900 6225
rect 866 6157 900 6159
rect 866 6125 900 6157
rect 866 6055 900 6087
rect 866 6053 900 6055
rect 866 5987 900 6015
rect 866 5981 900 5987
rect 866 5919 900 5943
rect 866 5909 900 5919
rect 866 5851 900 5871
rect 866 5837 900 5851
rect 866 5783 900 5799
rect 866 5765 900 5783
rect 866 5715 900 5727
rect 866 5693 900 5715
rect 866 5647 900 5655
rect 866 5621 900 5647
rect 962 6565 996 6591
rect 962 6557 996 6565
rect 962 6497 996 6519
rect 962 6485 996 6497
rect 962 6429 996 6447
rect 962 6413 996 6429
rect 962 6361 996 6375
rect 962 6341 996 6361
rect 962 6293 996 6303
rect 962 6269 996 6293
rect 962 6225 996 6231
rect 962 6197 996 6225
rect 962 6157 996 6159
rect 962 6125 996 6157
rect 962 6055 996 6087
rect 962 6053 996 6055
rect 962 5987 996 6015
rect 962 5981 996 5987
rect 962 5919 996 5943
rect 962 5909 996 5919
rect 962 5851 996 5871
rect 962 5837 996 5851
rect 962 5783 996 5799
rect 962 5765 996 5783
rect 962 5715 996 5727
rect 962 5693 996 5715
rect 962 5647 996 5655
rect 962 5621 996 5647
rect 1058 6565 1092 6591
rect 1058 6557 1092 6565
rect 1058 6497 1092 6519
rect 1058 6485 1092 6497
rect 1058 6429 1092 6447
rect 1058 6413 1092 6429
rect 1058 6361 1092 6375
rect 1058 6341 1092 6361
rect 1058 6293 1092 6303
rect 1058 6269 1092 6293
rect 1058 6225 1092 6231
rect 1058 6197 1092 6225
rect 1058 6157 1092 6159
rect 1058 6125 1092 6157
rect 1058 6055 1092 6087
rect 1058 6053 1092 6055
rect 1058 5987 1092 6015
rect 1058 5981 1092 5987
rect 1058 5919 1092 5943
rect 1058 5909 1092 5919
rect 1058 5851 1092 5871
rect 1058 5837 1092 5851
rect 1058 5783 1092 5799
rect 1058 5765 1092 5783
rect 1058 5715 1092 5727
rect 1058 5693 1092 5715
rect 1058 5647 1092 5655
rect 1058 5621 1092 5647
rect 1154 6565 1188 6591
rect 1154 6557 1188 6565
rect 1154 6497 1188 6519
rect 1154 6485 1188 6497
rect 1154 6429 1188 6447
rect 1154 6413 1188 6429
rect 1154 6361 1188 6375
rect 1154 6341 1188 6361
rect 1154 6293 1188 6303
rect 1154 6269 1188 6293
rect 1154 6225 1188 6231
rect 1154 6197 1188 6225
rect 1154 6157 1188 6159
rect 1154 6125 1188 6157
rect 1154 6055 1188 6087
rect 1154 6053 1188 6055
rect 1154 5987 1188 6015
rect 1154 5981 1188 5987
rect 1154 5919 1188 5943
rect 1154 5909 1188 5919
rect 1154 5851 1188 5871
rect 1154 5837 1188 5851
rect 1154 5783 1188 5799
rect 1154 5765 1188 5783
rect 1154 5715 1188 5727
rect 1154 5693 1188 5715
rect 1154 5647 1188 5655
rect 1154 5621 1188 5647
rect 1250 6565 1284 6591
rect 1250 6557 1284 6565
rect 1250 6497 1284 6519
rect 1250 6485 1284 6497
rect 1250 6429 1284 6447
rect 1250 6413 1284 6429
rect 1250 6361 1284 6375
rect 1250 6341 1284 6361
rect 1250 6293 1284 6303
rect 1250 6269 1284 6293
rect 1250 6225 1284 6231
rect 1250 6197 1284 6225
rect 1250 6157 1284 6159
rect 1250 6125 1284 6157
rect 1250 6055 1284 6087
rect 1250 6053 1284 6055
rect 1250 5987 1284 6015
rect 1250 5981 1284 5987
rect 1250 5919 1284 5943
rect 1250 5909 1284 5919
rect 1250 5851 1284 5871
rect 1250 5837 1284 5851
rect 1250 5783 1284 5799
rect 1250 5765 1284 5783
rect 1250 5715 1284 5727
rect 1250 5693 1284 5715
rect 1250 5647 1284 5655
rect 1250 5621 1284 5647
rect 1346 6565 1380 6591
rect 1346 6557 1380 6565
rect 1346 6497 1380 6519
rect 1346 6485 1380 6497
rect 1346 6429 1380 6447
rect 1346 6413 1380 6429
rect 1346 6361 1380 6375
rect 1346 6341 1380 6361
rect 1346 6293 1380 6303
rect 1346 6269 1380 6293
rect 1346 6225 1380 6231
rect 1346 6197 1380 6225
rect 1346 6157 1380 6159
rect 1346 6125 1380 6157
rect 1346 6055 1380 6087
rect 1346 6053 1380 6055
rect 1346 5987 1380 6015
rect 1346 5981 1380 5987
rect 1346 5919 1380 5943
rect 1346 5909 1380 5919
rect 1346 5851 1380 5871
rect 1346 5837 1380 5851
rect 1346 5783 1380 5799
rect 1346 5765 1380 5783
rect 1346 5715 1380 5727
rect 1346 5693 1380 5715
rect 1346 5647 1380 5655
rect 1346 5621 1380 5647
rect 1960 6561 1994 6587
rect 1960 6553 1994 6561
rect 1960 6493 1994 6515
rect 1960 6481 1994 6493
rect 1960 6425 1994 6443
rect 1960 6409 1994 6425
rect 1960 6357 1994 6371
rect 1960 6337 1994 6357
rect 1960 6289 1994 6299
rect 1960 6265 1994 6289
rect 1960 6221 1994 6227
rect 1960 6193 1994 6221
rect 1960 6153 1994 6155
rect 1960 6121 1994 6153
rect 1960 6051 1994 6083
rect 1960 6049 1994 6051
rect 1960 5983 1994 6011
rect 1960 5977 1994 5983
rect 1960 5915 1994 5939
rect 1960 5905 1994 5915
rect 1960 5847 1994 5867
rect 1960 5833 1994 5847
rect 1960 5779 1994 5795
rect 1960 5761 1994 5779
rect 1960 5711 1994 5723
rect 1960 5689 1994 5711
rect 1960 5643 1994 5651
rect 1960 5617 1994 5643
rect 2056 6561 2090 6587
rect 2056 6553 2090 6561
rect 2056 6493 2090 6515
rect 2056 6481 2090 6493
rect 2056 6425 2090 6443
rect 2056 6409 2090 6425
rect 2056 6357 2090 6371
rect 2056 6337 2090 6357
rect 2056 6289 2090 6299
rect 2056 6265 2090 6289
rect 2056 6221 2090 6227
rect 2056 6193 2090 6221
rect 2056 6153 2090 6155
rect 2056 6121 2090 6153
rect 2056 6051 2090 6083
rect 2056 6049 2090 6051
rect 2056 5983 2090 6011
rect 2056 5977 2090 5983
rect 2056 5915 2090 5939
rect 2056 5905 2090 5915
rect 2056 5847 2090 5867
rect 2056 5833 2090 5847
rect 2056 5779 2090 5795
rect 2056 5761 2090 5779
rect 2056 5711 2090 5723
rect 2056 5689 2090 5711
rect 2056 5643 2090 5651
rect 2056 5617 2090 5643
rect 2152 6561 2186 6587
rect 2152 6553 2186 6561
rect 2152 6493 2186 6515
rect 2152 6481 2186 6493
rect 2152 6425 2186 6443
rect 2152 6409 2186 6425
rect 2152 6357 2186 6371
rect 2152 6337 2186 6357
rect 2152 6289 2186 6299
rect 2152 6265 2186 6289
rect 2152 6221 2186 6227
rect 2152 6193 2186 6221
rect 2152 6153 2186 6155
rect 2152 6121 2186 6153
rect 2152 6051 2186 6083
rect 2152 6049 2186 6051
rect 2152 5983 2186 6011
rect 2152 5977 2186 5983
rect 2152 5915 2186 5939
rect 2152 5905 2186 5915
rect 2152 5847 2186 5867
rect 2152 5833 2186 5847
rect 2152 5779 2186 5795
rect 2152 5761 2186 5779
rect 2152 5711 2186 5723
rect 2152 5689 2186 5711
rect 2152 5643 2186 5651
rect 2152 5617 2186 5643
rect 2248 6561 2282 6587
rect 2248 6553 2282 6561
rect 2248 6493 2282 6515
rect 2248 6481 2282 6493
rect 2248 6425 2282 6443
rect 2248 6409 2282 6425
rect 2248 6357 2282 6371
rect 2248 6337 2282 6357
rect 2248 6289 2282 6299
rect 2248 6265 2282 6289
rect 2248 6221 2282 6227
rect 2248 6193 2282 6221
rect 2248 6153 2282 6155
rect 2248 6121 2282 6153
rect 2248 6051 2282 6083
rect 2248 6049 2282 6051
rect 2248 5983 2282 6011
rect 2248 5977 2282 5983
rect 2248 5915 2282 5939
rect 2248 5905 2282 5915
rect 2248 5847 2282 5867
rect 2248 5833 2282 5847
rect 2248 5779 2282 5795
rect 2248 5761 2282 5779
rect 2248 5711 2282 5723
rect 2248 5689 2282 5711
rect 2248 5643 2282 5651
rect 2248 5617 2282 5643
rect 2344 6561 2378 6587
rect 2344 6553 2378 6561
rect 2344 6493 2378 6515
rect 2344 6481 2378 6493
rect 2344 6425 2378 6443
rect 2344 6409 2378 6425
rect 2344 6357 2378 6371
rect 2344 6337 2378 6357
rect 2344 6289 2378 6299
rect 2344 6265 2378 6289
rect 2344 6221 2378 6227
rect 2344 6193 2378 6221
rect 2344 6153 2378 6155
rect 2344 6121 2378 6153
rect 2344 6051 2378 6083
rect 2344 6049 2378 6051
rect 2344 5983 2378 6011
rect 2344 5977 2378 5983
rect 2344 5915 2378 5939
rect 2344 5905 2378 5915
rect 2344 5847 2378 5867
rect 2344 5833 2378 5847
rect 2344 5779 2378 5795
rect 2344 5761 2378 5779
rect 2344 5711 2378 5723
rect 2344 5689 2378 5711
rect 2344 5643 2378 5651
rect 2344 5617 2378 5643
rect 2440 6561 2474 6587
rect 2440 6553 2474 6561
rect 2440 6493 2474 6515
rect 2440 6481 2474 6493
rect 2440 6425 2474 6443
rect 2440 6409 2474 6425
rect 2440 6357 2474 6371
rect 2440 6337 2474 6357
rect 2440 6289 2474 6299
rect 2440 6265 2474 6289
rect 2440 6221 2474 6227
rect 2440 6193 2474 6221
rect 2440 6153 2474 6155
rect 2440 6121 2474 6153
rect 2440 6051 2474 6083
rect 2440 6049 2474 6051
rect 2440 5983 2474 6011
rect 2440 5977 2474 5983
rect 2440 5915 2474 5939
rect 2440 5905 2474 5915
rect 2440 5847 2474 5867
rect 2440 5833 2474 5847
rect 2440 5779 2474 5795
rect 2440 5761 2474 5779
rect 2440 5711 2474 5723
rect 2440 5689 2474 5711
rect 2440 5643 2474 5651
rect 2440 5617 2474 5643
rect 2536 6561 2570 6587
rect 2536 6553 2570 6561
rect 2536 6493 2570 6515
rect 2536 6481 2570 6493
rect 2536 6425 2570 6443
rect 2536 6409 2570 6425
rect 2536 6357 2570 6371
rect 2536 6337 2570 6357
rect 2536 6289 2570 6299
rect 2536 6265 2570 6289
rect 2536 6221 2570 6227
rect 2536 6193 2570 6221
rect 2536 6153 2570 6155
rect 2536 6121 2570 6153
rect 2536 6051 2570 6083
rect 2536 6049 2570 6051
rect 2536 5983 2570 6011
rect 2536 5977 2570 5983
rect 2536 5915 2570 5939
rect 2536 5905 2570 5915
rect 2536 5847 2570 5867
rect 2536 5833 2570 5847
rect 2536 5779 2570 5795
rect 2536 5761 2570 5779
rect 2536 5711 2570 5723
rect 2536 5689 2570 5711
rect 2536 5643 2570 5651
rect 2536 5617 2570 5643
rect 2632 6561 2666 6587
rect 2632 6553 2666 6561
rect 2632 6493 2666 6515
rect 2632 6481 2666 6493
rect 2632 6425 2666 6443
rect 2632 6409 2666 6425
rect 2632 6357 2666 6371
rect 2632 6337 2666 6357
rect 2632 6289 2666 6299
rect 2632 6265 2666 6289
rect 2632 6221 2666 6227
rect 2632 6193 2666 6221
rect 2632 6153 2666 6155
rect 2632 6121 2666 6153
rect 2632 6051 2666 6083
rect 2632 6049 2666 6051
rect 2632 5983 2666 6011
rect 2632 5977 2666 5983
rect 2632 5915 2666 5939
rect 2632 5905 2666 5915
rect 2632 5847 2666 5867
rect 2632 5833 2666 5847
rect 2632 5779 2666 5795
rect 2632 5761 2666 5779
rect 2632 5711 2666 5723
rect 2632 5689 2666 5711
rect 2632 5643 2666 5651
rect 2632 5617 2666 5643
rect 2728 6561 2762 6587
rect 2728 6553 2762 6561
rect 2728 6493 2762 6515
rect 2728 6481 2762 6493
rect 2728 6425 2762 6443
rect 2728 6409 2762 6425
rect 2728 6357 2762 6371
rect 2728 6337 2762 6357
rect 2728 6289 2762 6299
rect 2728 6265 2762 6289
rect 2728 6221 2762 6227
rect 2728 6193 2762 6221
rect 2728 6153 2762 6155
rect 2728 6121 2762 6153
rect 2728 6051 2762 6083
rect 2728 6049 2762 6051
rect 2728 5983 2762 6011
rect 2728 5977 2762 5983
rect 2728 5915 2762 5939
rect 2728 5905 2762 5915
rect 2728 5847 2762 5867
rect 2728 5833 2762 5847
rect 2728 5779 2762 5795
rect 2728 5761 2762 5779
rect 2728 5711 2762 5723
rect 2728 5689 2762 5711
rect 2728 5643 2762 5651
rect 2728 5617 2762 5643
rect 9838 6840 9872 6874
rect 8426 6738 8460 6772
rect 8714 6753 8748 6787
rect 9362 6755 9396 6789
rect 3150 6549 3184 6575
rect 3150 6541 3184 6549
rect 3150 6481 3184 6503
rect 3150 6469 3184 6481
rect 3150 6413 3184 6431
rect 3150 6397 3184 6413
rect 3150 6345 3184 6359
rect 3150 6325 3184 6345
rect 3150 6277 3184 6287
rect 3150 6253 3184 6277
rect 3150 6209 3184 6215
rect 3150 6181 3184 6209
rect 3150 6141 3184 6143
rect 3150 6109 3184 6141
rect 3150 6039 3184 6071
rect 3150 6037 3184 6039
rect 3150 5971 3184 5999
rect 3150 5965 3184 5971
rect 3150 5903 3184 5927
rect 3150 5893 3184 5903
rect 3150 5835 3184 5855
rect 3150 5821 3184 5835
rect 3150 5767 3184 5783
rect 3150 5749 3184 5767
rect 3150 5699 3184 5711
rect 3150 5677 3184 5699
rect 3150 5631 3184 5639
rect 3150 5605 3184 5631
rect 3246 6549 3280 6575
rect 3246 6541 3280 6549
rect 3246 6481 3280 6503
rect 3246 6469 3280 6481
rect 3246 6413 3280 6431
rect 3246 6397 3280 6413
rect 3246 6345 3280 6359
rect 3246 6325 3280 6345
rect 3246 6277 3280 6287
rect 3246 6253 3280 6277
rect 3246 6209 3280 6215
rect 3246 6181 3280 6209
rect 3246 6141 3280 6143
rect 3246 6109 3280 6141
rect 3246 6039 3280 6071
rect 3246 6037 3280 6039
rect 3246 5971 3280 5999
rect 3246 5965 3280 5971
rect 3246 5903 3280 5927
rect 3246 5893 3280 5903
rect 3246 5835 3280 5855
rect 3246 5821 3280 5835
rect 3246 5767 3280 5783
rect 3246 5749 3280 5767
rect 3246 5699 3280 5711
rect 3246 5677 3280 5699
rect 3246 5631 3280 5639
rect 3246 5605 3280 5631
rect -868 5487 -834 5489
rect -868 5455 -834 5487
rect -868 5385 -834 5417
rect -868 5383 -834 5385
rect 3342 6549 3376 6575
rect 3342 6541 3376 6549
rect 3342 6481 3376 6503
rect 3342 6469 3376 6481
rect 3342 6413 3376 6431
rect 3342 6397 3376 6413
rect 3342 6345 3376 6359
rect 3342 6325 3376 6345
rect 3342 6277 3376 6287
rect 3342 6253 3376 6277
rect 3342 6209 3376 6215
rect 3342 6181 3376 6209
rect 3342 6141 3376 6143
rect 3342 6109 3376 6141
rect 3342 6039 3376 6071
rect 3342 6037 3376 6039
rect 3342 5971 3376 5999
rect 3342 5965 3376 5971
rect 3342 5903 3376 5927
rect 3342 5893 3376 5903
rect 3342 5835 3376 5855
rect 3342 5821 3376 5835
rect 3342 5767 3376 5783
rect 3342 5749 3376 5767
rect 3342 5699 3376 5711
rect 3342 5677 3376 5699
rect 3342 5631 3376 5639
rect 3342 5605 3376 5631
rect 3438 6549 3472 6575
rect 3438 6541 3472 6549
rect 3438 6481 3472 6503
rect 3438 6469 3472 6481
rect 3438 6413 3472 6431
rect 3438 6397 3472 6413
rect 3438 6345 3472 6359
rect 3438 6325 3472 6345
rect 3438 6277 3472 6287
rect 3438 6253 3472 6277
rect 3438 6209 3472 6215
rect 3438 6181 3472 6209
rect 3438 6141 3472 6143
rect 3438 6109 3472 6141
rect 3438 6039 3472 6071
rect 3438 6037 3472 6039
rect 3438 5971 3472 5999
rect 3438 5965 3472 5971
rect 3438 5903 3472 5927
rect 3438 5893 3472 5903
rect 3438 5835 3472 5855
rect 3438 5821 3472 5835
rect 3438 5767 3472 5783
rect 3438 5749 3472 5767
rect 3438 5699 3472 5711
rect 3438 5677 3472 5699
rect 3438 5631 3472 5639
rect 3438 5605 3472 5631
rect 3534 6549 3568 6575
rect 3534 6541 3568 6549
rect 3534 6481 3568 6503
rect 3534 6469 3568 6481
rect 3534 6413 3568 6431
rect 3534 6397 3568 6413
rect 3534 6345 3568 6359
rect 3534 6325 3568 6345
rect 3534 6277 3568 6287
rect 3534 6253 3568 6277
rect 3534 6209 3568 6215
rect 3534 6181 3568 6209
rect 3534 6141 3568 6143
rect 3534 6109 3568 6141
rect 3534 6039 3568 6071
rect 3534 6037 3568 6039
rect 3534 5971 3568 5999
rect 3534 5965 3568 5971
rect 3534 5903 3568 5927
rect 3534 5893 3568 5903
rect 3534 5835 3568 5855
rect 3534 5821 3568 5835
rect 3534 5767 3568 5783
rect 3534 5749 3568 5767
rect 3534 5699 3568 5711
rect 3534 5677 3568 5699
rect 3534 5631 3568 5639
rect 3534 5605 3568 5631
rect 3630 6549 3664 6575
rect 3630 6541 3664 6549
rect 3630 6481 3664 6503
rect 3630 6469 3664 6481
rect 3630 6413 3664 6431
rect 3630 6397 3664 6413
rect 3630 6345 3664 6359
rect 3630 6325 3664 6345
rect 3630 6277 3664 6287
rect 3630 6253 3664 6277
rect 3630 6209 3664 6215
rect 3630 6181 3664 6209
rect 3630 6141 3664 6143
rect 3630 6109 3664 6141
rect 3630 6039 3664 6071
rect 3630 6037 3664 6039
rect 3630 5971 3664 5999
rect 3630 5965 3664 5971
rect 3630 5903 3664 5927
rect 3630 5893 3664 5903
rect 3630 5835 3664 5855
rect 3630 5821 3664 5835
rect 3630 5767 3664 5783
rect 3630 5749 3664 5767
rect 3630 5699 3664 5711
rect 3630 5677 3664 5699
rect 3630 5631 3664 5639
rect 3630 5605 3664 5631
rect 3726 6549 3760 6575
rect 3726 6541 3760 6549
rect 3726 6481 3760 6503
rect 3726 6469 3760 6481
rect 3726 6413 3760 6431
rect 3726 6397 3760 6413
rect 3726 6345 3760 6359
rect 3726 6325 3760 6345
rect 3726 6277 3760 6287
rect 3726 6253 3760 6277
rect 3726 6209 3760 6215
rect 3726 6181 3760 6209
rect 3726 6141 3760 6143
rect 3726 6109 3760 6141
rect 3726 6039 3760 6071
rect 3726 6037 3760 6039
rect 3726 5971 3760 5999
rect 3726 5965 3760 5971
rect 3726 5903 3760 5927
rect 3726 5893 3760 5903
rect 3726 5835 3760 5855
rect 3726 5821 3760 5835
rect 3726 5767 3760 5783
rect 3726 5749 3760 5767
rect 3726 5699 3760 5711
rect 3726 5677 3760 5699
rect 3726 5631 3760 5639
rect 3726 5605 3760 5631
rect 3822 6549 3856 6575
rect 3822 6541 3856 6549
rect 3822 6481 3856 6503
rect 3822 6469 3856 6481
rect 3822 6413 3856 6431
rect 3822 6397 3856 6413
rect 3822 6345 3856 6359
rect 3822 6325 3856 6345
rect 3822 6277 3856 6287
rect 3822 6253 3856 6277
rect 3822 6209 3856 6215
rect 3822 6181 3856 6209
rect 3822 6141 3856 6143
rect 3822 6109 3856 6141
rect 3822 6039 3856 6071
rect 3822 6037 3856 6039
rect 3822 5971 3856 5999
rect 3822 5965 3856 5971
rect 3822 5903 3856 5927
rect 3822 5893 3856 5903
rect 3822 5835 3856 5855
rect 3822 5821 3856 5835
rect 3822 5767 3856 5783
rect 3822 5749 3856 5767
rect 3822 5699 3856 5711
rect 3822 5677 3856 5699
rect 3822 5631 3856 5639
rect 3822 5605 3856 5631
rect 3918 6549 3952 6575
rect 3918 6541 3952 6549
rect 3918 6481 3952 6503
rect 3918 6469 3952 6481
rect 3918 6413 3952 6431
rect 3918 6397 3952 6413
rect 3918 6345 3952 6359
rect 3918 6325 3952 6345
rect 3918 6277 3952 6287
rect 3918 6253 3952 6277
rect 3918 6209 3952 6215
rect 3918 6181 3952 6209
rect 3918 6141 3952 6143
rect 3918 6109 3952 6141
rect 3918 6039 3952 6071
rect 3918 6037 3952 6039
rect 3918 5971 3952 5999
rect 3918 5965 3952 5971
rect 3918 5903 3952 5927
rect 3918 5893 3952 5903
rect 3918 5835 3952 5855
rect 3918 5821 3952 5835
rect 3918 5767 3952 5783
rect 3918 5749 3952 5767
rect 3918 5699 3952 5711
rect 3918 5677 3952 5699
rect 3918 5631 3952 5639
rect 3918 5605 3952 5631
rect 4014 6549 4048 6575
rect 4014 6541 4048 6549
rect 4014 6481 4048 6503
rect 4014 6469 4048 6481
rect 4014 6413 4048 6431
rect 4014 6397 4048 6413
rect 4014 6345 4048 6359
rect 4014 6325 4048 6345
rect 4014 6277 4048 6287
rect 4014 6253 4048 6277
rect 4014 6209 4048 6215
rect 4014 6181 4048 6209
rect 4014 6141 4048 6143
rect 4014 6109 4048 6141
rect 4014 6039 4048 6071
rect 4014 6037 4048 6039
rect 4014 5971 4048 5999
rect 4014 5965 4048 5971
rect 4014 5903 4048 5927
rect 4014 5893 4048 5903
rect 4014 5835 4048 5855
rect 4014 5821 4048 5835
rect 4014 5767 4048 5783
rect 4014 5749 4048 5767
rect 4014 5699 4048 5711
rect 4014 5677 4048 5699
rect 4014 5631 4048 5639
rect 4014 5605 4048 5631
rect 4110 6549 4144 6575
rect 4110 6541 4144 6549
rect 4110 6481 4144 6503
rect 4110 6469 4144 6481
rect 4110 6413 4144 6431
rect 4110 6397 4144 6413
rect 4110 6345 4144 6359
rect 4110 6325 4144 6345
rect 4110 6277 4144 6287
rect 4110 6253 4144 6277
rect 4110 6209 4144 6215
rect 4110 6181 4144 6209
rect 4110 6141 4144 6143
rect 4110 6109 4144 6141
rect 4110 6039 4144 6071
rect 4110 6037 4144 6039
rect 4110 5971 4144 5999
rect 4110 5965 4144 5971
rect 4110 5903 4144 5927
rect 4110 5893 4144 5903
rect 4110 5835 4144 5855
rect 4110 5821 4144 5835
rect 4110 5767 4144 5783
rect 4110 5749 4144 5767
rect 4110 5699 4144 5711
rect 4110 5677 4144 5699
rect 4110 5631 4144 5639
rect 4110 5605 4144 5631
rect 4206 6549 4240 6575
rect 4206 6541 4240 6549
rect 4206 6481 4240 6503
rect 4206 6469 4240 6481
rect 4206 6413 4240 6431
rect 4206 6397 4240 6413
rect 4206 6345 4240 6359
rect 4206 6325 4240 6345
rect 4206 6277 4240 6287
rect 4206 6253 4240 6277
rect 4206 6209 4240 6215
rect 4206 6181 4240 6209
rect 4206 6141 4240 6143
rect 4206 6109 4240 6141
rect 4206 6039 4240 6071
rect 4206 6037 4240 6039
rect 4206 5971 4240 5999
rect 4206 5965 4240 5971
rect 4206 5903 4240 5927
rect 4206 5893 4240 5903
rect 4206 5835 4240 5855
rect 4206 5821 4240 5835
rect 4206 5767 4240 5783
rect 4206 5749 4240 5767
rect 4206 5699 4240 5711
rect 4206 5677 4240 5699
rect 4206 5631 4240 5639
rect 4206 5605 4240 5631
rect 4302 6549 4336 6575
rect 4302 6541 4336 6549
rect 4302 6481 4336 6503
rect 4302 6469 4336 6481
rect 4302 6413 4336 6431
rect 4302 6397 4336 6413
rect 4302 6345 4336 6359
rect 4302 6325 4336 6345
rect 4302 6277 4336 6287
rect 4302 6253 4336 6277
rect 4302 6209 4336 6215
rect 4302 6181 4336 6209
rect 4302 6141 4336 6143
rect 4302 6109 4336 6141
rect 4302 6039 4336 6071
rect 4302 6037 4336 6039
rect 4302 5971 4336 5999
rect 4302 5965 4336 5971
rect 4302 5903 4336 5927
rect 4302 5893 4336 5903
rect 4302 5835 4336 5855
rect 4302 5821 4336 5835
rect 4302 5767 4336 5783
rect 4302 5749 4336 5767
rect 4302 5699 4336 5711
rect 4302 5677 4336 5699
rect 4302 5631 4336 5639
rect 4302 5605 4336 5631
rect 4916 6545 4950 6571
rect 4916 6537 4950 6545
rect 4916 6477 4950 6499
rect 4916 6465 4950 6477
rect 4916 6409 4950 6427
rect 4916 6393 4950 6409
rect 4916 6341 4950 6355
rect 4916 6321 4950 6341
rect 4916 6273 4950 6283
rect 4916 6249 4950 6273
rect 4916 6205 4950 6211
rect 4916 6177 4950 6205
rect 4916 6137 4950 6139
rect 4916 6105 4950 6137
rect 4916 6035 4950 6067
rect 4916 6033 4950 6035
rect 4916 5967 4950 5995
rect 4916 5961 4950 5967
rect 4916 5899 4950 5923
rect 4916 5889 4950 5899
rect 4916 5831 4950 5851
rect 4916 5817 4950 5831
rect 4916 5763 4950 5779
rect 4916 5745 4950 5763
rect 4916 5695 4950 5707
rect 4916 5673 4950 5695
rect 4916 5627 4950 5635
rect 4916 5601 4950 5627
rect 5012 6545 5046 6571
rect 5012 6537 5046 6545
rect 5012 6477 5046 6499
rect 5012 6465 5046 6477
rect 5012 6409 5046 6427
rect 5012 6393 5046 6409
rect 5012 6341 5046 6355
rect 5012 6321 5046 6341
rect 5012 6273 5046 6283
rect 5012 6249 5046 6273
rect 5012 6205 5046 6211
rect 5012 6177 5046 6205
rect 5012 6137 5046 6139
rect 5012 6105 5046 6137
rect 5012 6035 5046 6067
rect 5012 6033 5046 6035
rect 5012 5967 5046 5995
rect 5012 5961 5046 5967
rect 5012 5899 5046 5923
rect 5012 5889 5046 5899
rect 5012 5831 5046 5851
rect 5012 5817 5046 5831
rect 5012 5763 5046 5779
rect 5012 5745 5046 5763
rect 5012 5695 5046 5707
rect 5012 5673 5046 5695
rect 5012 5627 5046 5635
rect 5012 5601 5046 5627
rect 880 5372 914 5406
rect 5108 6545 5142 6571
rect 5108 6537 5142 6545
rect 5108 6477 5142 6499
rect 5108 6465 5142 6477
rect 5108 6409 5142 6427
rect 5108 6393 5142 6409
rect 5108 6341 5142 6355
rect 5108 6321 5142 6341
rect 5108 6273 5142 6283
rect 5108 6249 5142 6273
rect 5108 6205 5142 6211
rect 5108 6177 5142 6205
rect 5108 6137 5142 6139
rect 5108 6105 5142 6137
rect 5108 6035 5142 6067
rect 5108 6033 5142 6035
rect 5108 5967 5142 5995
rect 5108 5961 5142 5967
rect 5108 5899 5142 5923
rect 5108 5889 5142 5899
rect 5108 5831 5142 5851
rect 5108 5817 5142 5831
rect 5108 5763 5142 5779
rect 5108 5745 5142 5763
rect 5108 5695 5142 5707
rect 5108 5673 5142 5695
rect 5108 5627 5142 5635
rect 5108 5601 5142 5627
rect 5204 6545 5238 6571
rect 5204 6537 5238 6545
rect 5204 6477 5238 6499
rect 5204 6465 5238 6477
rect 5204 6409 5238 6427
rect 5204 6393 5238 6409
rect 5204 6341 5238 6355
rect 5204 6321 5238 6341
rect 5204 6273 5238 6283
rect 5204 6249 5238 6273
rect 5204 6205 5238 6211
rect 5204 6177 5238 6205
rect 5204 6137 5238 6139
rect 5204 6105 5238 6137
rect 5204 6035 5238 6067
rect 5204 6033 5238 6035
rect 5204 5967 5238 5995
rect 5204 5961 5238 5967
rect 5204 5899 5238 5923
rect 5204 5889 5238 5899
rect 5204 5831 5238 5851
rect 5204 5817 5238 5831
rect 5204 5763 5238 5779
rect 5204 5745 5238 5763
rect 5204 5695 5238 5707
rect 5204 5673 5238 5695
rect 5204 5627 5238 5635
rect 5204 5601 5238 5627
rect 5300 6545 5334 6571
rect 5300 6537 5334 6545
rect 5300 6477 5334 6499
rect 5300 6465 5334 6477
rect 5300 6409 5334 6427
rect 5300 6393 5334 6409
rect 5300 6341 5334 6355
rect 5300 6321 5334 6341
rect 5300 6273 5334 6283
rect 5300 6249 5334 6273
rect 5300 6205 5334 6211
rect 5300 6177 5334 6205
rect 5300 6137 5334 6139
rect 5300 6105 5334 6137
rect 5300 6035 5334 6067
rect 5300 6033 5334 6035
rect 5300 5967 5334 5995
rect 5300 5961 5334 5967
rect 5300 5899 5334 5923
rect 5300 5889 5334 5899
rect 5300 5831 5334 5851
rect 5300 5817 5334 5831
rect 5300 5763 5334 5779
rect 5300 5745 5334 5763
rect 5300 5695 5334 5707
rect 5300 5673 5334 5695
rect 5300 5627 5334 5635
rect 5300 5601 5334 5627
rect 5396 6545 5430 6571
rect 5396 6537 5430 6545
rect 5396 6477 5430 6499
rect 5396 6465 5430 6477
rect 5396 6409 5430 6427
rect 5396 6393 5430 6409
rect 5396 6341 5430 6355
rect 5396 6321 5430 6341
rect 5396 6273 5430 6283
rect 5396 6249 5430 6273
rect 5396 6205 5430 6211
rect 5396 6177 5430 6205
rect 5396 6137 5430 6139
rect 5396 6105 5430 6137
rect 5396 6035 5430 6067
rect 5396 6033 5430 6035
rect 5396 5967 5430 5995
rect 5396 5961 5430 5967
rect 5396 5899 5430 5923
rect 5396 5889 5430 5899
rect 5396 5831 5430 5851
rect 5396 5817 5430 5831
rect 5396 5763 5430 5779
rect 5396 5745 5430 5763
rect 5396 5695 5430 5707
rect 5396 5673 5430 5695
rect 5396 5627 5430 5635
rect 5396 5601 5430 5627
rect 5492 6545 5526 6571
rect 5492 6537 5526 6545
rect 5492 6477 5526 6499
rect 5492 6465 5526 6477
rect 5492 6409 5526 6427
rect 5492 6393 5526 6409
rect 5492 6341 5526 6355
rect 5492 6321 5526 6341
rect 5492 6273 5526 6283
rect 5492 6249 5526 6273
rect 5492 6205 5526 6211
rect 5492 6177 5526 6205
rect 5492 6137 5526 6139
rect 5492 6105 5526 6137
rect 5492 6035 5526 6067
rect 5492 6033 5526 6035
rect 5492 5967 5526 5995
rect 5492 5961 5526 5967
rect 5492 5899 5526 5923
rect 5492 5889 5526 5899
rect 5492 5831 5526 5851
rect 5492 5817 5526 5831
rect 5492 5763 5526 5779
rect 5492 5745 5526 5763
rect 5492 5695 5526 5707
rect 5492 5673 5526 5695
rect 5492 5627 5526 5635
rect 5492 5601 5526 5627
rect 5588 6545 5622 6571
rect 5588 6537 5622 6545
rect 5588 6477 5622 6499
rect 5588 6465 5622 6477
rect 5588 6409 5622 6427
rect 5588 6393 5622 6409
rect 5588 6341 5622 6355
rect 5588 6321 5622 6341
rect 5588 6273 5622 6283
rect 5588 6249 5622 6273
rect 5588 6205 5622 6211
rect 5588 6177 5622 6205
rect 5588 6137 5622 6139
rect 5588 6105 5622 6137
rect 5588 6035 5622 6067
rect 5588 6033 5622 6035
rect 5588 5967 5622 5995
rect 5588 5961 5622 5967
rect 5588 5899 5622 5923
rect 5588 5889 5622 5899
rect 5588 5831 5622 5851
rect 5588 5817 5622 5831
rect 5588 5763 5622 5779
rect 5588 5745 5622 5763
rect 5588 5695 5622 5707
rect 5588 5673 5622 5695
rect 5588 5627 5622 5635
rect 5588 5601 5622 5627
rect 5684 6545 5718 6571
rect 5684 6537 5718 6545
rect 5684 6477 5718 6499
rect 5684 6465 5718 6477
rect 5684 6409 5718 6427
rect 5684 6393 5718 6409
rect 5684 6341 5718 6355
rect 5684 6321 5718 6341
rect 5684 6273 5718 6283
rect 5684 6249 5718 6273
rect 5684 6205 5718 6211
rect 5684 6177 5718 6205
rect 5684 6137 5718 6139
rect 5684 6105 5718 6137
rect 5684 6035 5718 6067
rect 5684 6033 5718 6035
rect 5684 5967 5718 5995
rect 5684 5961 5718 5967
rect 5684 5899 5718 5923
rect 5684 5889 5718 5899
rect 5684 5831 5718 5851
rect 5684 5817 5718 5831
rect 5684 5763 5718 5779
rect 5684 5745 5718 5763
rect 5684 5695 5718 5707
rect 5684 5673 5718 5695
rect 5684 5627 5718 5635
rect 5684 5601 5718 5627
rect 12994 6814 13028 6848
rect 11514 6736 11548 6770
rect 11802 6751 11836 6785
rect 12518 6729 12552 6763
rect 6180 6549 6214 6575
rect 6180 6541 6214 6549
rect 6180 6481 6214 6503
rect 6180 6469 6214 6481
rect 6180 6413 6214 6431
rect 6180 6397 6214 6413
rect 6180 6345 6214 6359
rect 6180 6325 6214 6345
rect 6180 6277 6214 6287
rect 6180 6253 6214 6277
rect 6180 6209 6214 6215
rect 6180 6181 6214 6209
rect 6180 6141 6214 6143
rect 6180 6109 6214 6141
rect 6180 6039 6214 6071
rect 6180 6037 6214 6039
rect 6180 5971 6214 5999
rect 6180 5965 6214 5971
rect 6180 5903 6214 5927
rect 6180 5893 6214 5903
rect 6180 5835 6214 5855
rect 6180 5821 6214 5835
rect 6180 5767 6214 5783
rect 6180 5749 6214 5767
rect 6180 5699 6214 5711
rect 6180 5677 6214 5699
rect 6180 5631 6214 5639
rect 6180 5605 6214 5631
rect 6276 6549 6310 6575
rect 6276 6541 6310 6549
rect 6276 6481 6310 6503
rect 6276 6469 6310 6481
rect 6276 6413 6310 6431
rect 6276 6397 6310 6413
rect 6276 6345 6310 6359
rect 6276 6325 6310 6345
rect 6276 6277 6310 6287
rect 6276 6253 6310 6277
rect 6276 6209 6310 6215
rect 6276 6181 6310 6209
rect 6276 6141 6310 6143
rect 6276 6109 6310 6141
rect 6276 6039 6310 6071
rect 6276 6037 6310 6039
rect 6276 5971 6310 5999
rect 6276 5965 6310 5971
rect 6276 5903 6310 5927
rect 6276 5893 6310 5903
rect 6276 5835 6310 5855
rect 6276 5821 6310 5835
rect 6276 5767 6310 5783
rect 6276 5749 6310 5767
rect 6276 5699 6310 5711
rect 6276 5677 6310 5699
rect 6276 5631 6310 5639
rect 6276 5605 6310 5631
rect 2344 5376 2378 5410
rect 6372 6549 6406 6575
rect 6372 6541 6406 6549
rect 6372 6481 6406 6503
rect 6372 6469 6406 6481
rect 6372 6413 6406 6431
rect 6372 6397 6406 6413
rect 6372 6345 6406 6359
rect 6372 6325 6406 6345
rect 6372 6277 6406 6287
rect 6372 6253 6406 6277
rect 6372 6209 6406 6215
rect 6372 6181 6406 6209
rect 6372 6141 6406 6143
rect 6372 6109 6406 6141
rect 6372 6039 6406 6071
rect 6372 6037 6406 6039
rect 6372 5971 6406 5999
rect 6372 5965 6406 5971
rect 6372 5903 6406 5927
rect 6372 5893 6406 5903
rect 6372 5835 6406 5855
rect 6372 5821 6406 5835
rect 6372 5767 6406 5783
rect 6372 5749 6406 5767
rect 6372 5699 6406 5711
rect 6372 5677 6406 5699
rect 6372 5631 6406 5639
rect 6372 5605 6406 5631
rect 6468 6549 6502 6575
rect 6468 6541 6502 6549
rect 6468 6481 6502 6503
rect 6468 6469 6502 6481
rect 6468 6413 6502 6431
rect 6468 6397 6502 6413
rect 6468 6345 6502 6359
rect 6468 6325 6502 6345
rect 6468 6277 6502 6287
rect 6468 6253 6502 6277
rect 6468 6209 6502 6215
rect 6468 6181 6502 6209
rect 6468 6141 6502 6143
rect 6468 6109 6502 6141
rect 6468 6039 6502 6071
rect 6468 6037 6502 6039
rect 6468 5971 6502 5999
rect 6468 5965 6502 5971
rect 6468 5903 6502 5927
rect 6468 5893 6502 5903
rect 6468 5835 6502 5855
rect 6468 5821 6502 5835
rect 6468 5767 6502 5783
rect 6468 5749 6502 5767
rect 6468 5699 6502 5711
rect 6468 5677 6502 5699
rect 6468 5631 6502 5639
rect 6468 5605 6502 5631
rect 6564 6549 6598 6575
rect 6564 6541 6598 6549
rect 6564 6481 6598 6503
rect 6564 6469 6598 6481
rect 6564 6413 6598 6431
rect 6564 6397 6598 6413
rect 6564 6345 6598 6359
rect 6564 6325 6598 6345
rect 6564 6277 6598 6287
rect 6564 6253 6598 6277
rect 6564 6209 6598 6215
rect 6564 6181 6598 6209
rect 6564 6141 6598 6143
rect 6564 6109 6598 6141
rect 6564 6039 6598 6071
rect 6564 6037 6598 6039
rect 6564 5971 6598 5999
rect 6564 5965 6598 5971
rect 6564 5903 6598 5927
rect 6564 5893 6598 5903
rect 6564 5835 6598 5855
rect 6564 5821 6598 5835
rect 6564 5767 6598 5783
rect 6564 5749 6598 5767
rect 6564 5699 6598 5711
rect 6564 5677 6598 5699
rect 6564 5631 6598 5639
rect 6564 5605 6598 5631
rect 6660 6549 6694 6575
rect 6660 6541 6694 6549
rect 6660 6481 6694 6503
rect 6660 6469 6694 6481
rect 6660 6413 6694 6431
rect 6660 6397 6694 6413
rect 6660 6345 6694 6359
rect 6660 6325 6694 6345
rect 6660 6277 6694 6287
rect 6660 6253 6694 6277
rect 6660 6209 6694 6215
rect 6660 6181 6694 6209
rect 6660 6141 6694 6143
rect 6660 6109 6694 6141
rect 6660 6039 6694 6071
rect 6660 6037 6694 6039
rect 6660 5971 6694 5999
rect 6660 5965 6694 5971
rect 6660 5903 6694 5927
rect 6660 5893 6694 5903
rect 6660 5835 6694 5855
rect 6660 5821 6694 5835
rect 6660 5767 6694 5783
rect 6660 5749 6694 5767
rect 6660 5699 6694 5711
rect 6660 5677 6694 5699
rect 6660 5631 6694 5639
rect 6660 5605 6694 5631
rect 6756 6549 6790 6575
rect 6756 6541 6790 6549
rect 6756 6481 6790 6503
rect 6756 6469 6790 6481
rect 6756 6413 6790 6431
rect 6756 6397 6790 6413
rect 6756 6345 6790 6359
rect 6756 6325 6790 6345
rect 6756 6277 6790 6287
rect 6756 6253 6790 6277
rect 6756 6209 6790 6215
rect 6756 6181 6790 6209
rect 6756 6141 6790 6143
rect 6756 6109 6790 6141
rect 6756 6039 6790 6071
rect 6756 6037 6790 6039
rect 6756 5971 6790 5999
rect 6756 5965 6790 5971
rect 6756 5903 6790 5927
rect 6756 5893 6790 5903
rect 6756 5835 6790 5855
rect 6756 5821 6790 5835
rect 6756 5767 6790 5783
rect 6756 5749 6790 5767
rect 6756 5699 6790 5711
rect 6756 5677 6790 5699
rect 6756 5631 6790 5639
rect 6756 5605 6790 5631
rect 6852 6549 6886 6575
rect 6852 6541 6886 6549
rect 6852 6481 6886 6503
rect 6852 6469 6886 6481
rect 6852 6413 6886 6431
rect 6852 6397 6886 6413
rect 6852 6345 6886 6359
rect 6852 6325 6886 6345
rect 6852 6277 6886 6287
rect 6852 6253 6886 6277
rect 6852 6209 6886 6215
rect 6852 6181 6886 6209
rect 6852 6141 6886 6143
rect 6852 6109 6886 6141
rect 6852 6039 6886 6071
rect 6852 6037 6886 6039
rect 6852 5971 6886 5999
rect 6852 5965 6886 5971
rect 6852 5903 6886 5927
rect 6852 5893 6886 5903
rect 6852 5835 6886 5855
rect 6852 5821 6886 5835
rect 6852 5767 6886 5783
rect 6852 5749 6886 5767
rect 6852 5699 6886 5711
rect 6852 5677 6886 5699
rect 6852 5631 6886 5639
rect 6852 5605 6886 5631
rect 6948 6549 6982 6575
rect 6948 6541 6982 6549
rect 6948 6481 6982 6503
rect 6948 6469 6982 6481
rect 6948 6413 6982 6431
rect 6948 6397 6982 6413
rect 6948 6345 6982 6359
rect 6948 6325 6982 6345
rect 6948 6277 6982 6287
rect 6948 6253 6982 6277
rect 6948 6209 6982 6215
rect 6948 6181 6982 6209
rect 6948 6141 6982 6143
rect 6948 6109 6982 6141
rect 6948 6039 6982 6071
rect 6948 6037 6982 6039
rect 6948 5971 6982 5999
rect 6948 5965 6982 5971
rect 6948 5903 6982 5927
rect 6948 5893 6982 5903
rect 6948 5835 6982 5855
rect 6948 5821 6982 5835
rect 6948 5767 6982 5783
rect 6948 5749 6982 5767
rect 6948 5699 6982 5711
rect 6948 5677 6982 5699
rect 6948 5631 6982 5639
rect 6948 5605 6982 5631
rect 7044 6549 7078 6575
rect 7044 6541 7078 6549
rect 7044 6481 7078 6503
rect 7044 6469 7078 6481
rect 7044 6413 7078 6431
rect 7044 6397 7078 6413
rect 7044 6345 7078 6359
rect 7044 6325 7078 6345
rect 7044 6277 7078 6287
rect 7044 6253 7078 6277
rect 7044 6209 7078 6215
rect 7044 6181 7078 6209
rect 7044 6141 7078 6143
rect 7044 6109 7078 6141
rect 7044 6039 7078 6071
rect 7044 6037 7078 6039
rect 7044 5971 7078 5999
rect 7044 5965 7078 5971
rect 7044 5903 7078 5927
rect 7044 5893 7078 5903
rect 7044 5835 7078 5855
rect 7044 5821 7078 5835
rect 7044 5767 7078 5783
rect 7044 5749 7078 5767
rect 7044 5699 7078 5711
rect 7044 5677 7078 5699
rect 7044 5631 7078 5639
rect 7044 5605 7078 5631
rect 7140 6549 7174 6575
rect 7140 6541 7174 6549
rect 7140 6481 7174 6503
rect 7140 6469 7174 6481
rect 7140 6413 7174 6431
rect 7140 6397 7174 6413
rect 7140 6345 7174 6359
rect 7140 6325 7174 6345
rect 7140 6277 7174 6287
rect 7140 6253 7174 6277
rect 7140 6209 7174 6215
rect 7140 6181 7174 6209
rect 7140 6141 7174 6143
rect 7140 6109 7174 6141
rect 7140 6039 7174 6071
rect 7140 6037 7174 6039
rect 7140 5971 7174 5999
rect 7140 5965 7174 5971
rect 7140 5903 7174 5927
rect 7140 5893 7174 5903
rect 7140 5835 7174 5855
rect 7140 5821 7174 5835
rect 7140 5767 7174 5783
rect 7140 5749 7174 5767
rect 7140 5699 7174 5711
rect 7140 5677 7174 5699
rect 7140 5631 7174 5639
rect 7140 5605 7174 5631
rect 7236 6549 7270 6575
rect 7236 6541 7270 6549
rect 7236 6481 7270 6503
rect 7236 6469 7270 6481
rect 7236 6413 7270 6431
rect 7236 6397 7270 6413
rect 7236 6345 7270 6359
rect 7236 6325 7270 6345
rect 7236 6277 7270 6287
rect 7236 6253 7270 6277
rect 7236 6209 7270 6215
rect 7236 6181 7270 6209
rect 7236 6141 7270 6143
rect 7236 6109 7270 6141
rect 7236 6039 7270 6071
rect 7236 6037 7270 6039
rect 7236 5971 7270 5999
rect 7236 5965 7270 5971
rect 7236 5903 7270 5927
rect 7236 5893 7270 5903
rect 7236 5835 7270 5855
rect 7236 5821 7270 5835
rect 7236 5767 7270 5783
rect 7236 5749 7270 5767
rect 7236 5699 7270 5711
rect 7236 5677 7270 5699
rect 7236 5631 7270 5639
rect 7236 5605 7270 5631
rect 7332 6549 7366 6575
rect 7332 6541 7366 6549
rect 7332 6481 7366 6503
rect 7332 6469 7366 6481
rect 7332 6413 7366 6431
rect 7332 6397 7366 6413
rect 7332 6345 7366 6359
rect 7332 6325 7366 6345
rect 7332 6277 7366 6287
rect 7332 6253 7366 6277
rect 7332 6209 7366 6215
rect 7332 6181 7366 6209
rect 7332 6141 7366 6143
rect 7332 6109 7366 6141
rect 7332 6039 7366 6071
rect 7332 6037 7366 6039
rect 7332 5971 7366 5999
rect 7332 5965 7366 5971
rect 7332 5903 7366 5927
rect 7332 5893 7366 5903
rect 7332 5835 7366 5855
rect 7332 5821 7366 5835
rect 7332 5767 7366 5783
rect 7332 5749 7366 5767
rect 7332 5699 7366 5711
rect 7332 5677 7366 5699
rect 7332 5631 7366 5639
rect 7332 5605 7366 5631
rect 7946 6545 7980 6571
rect 7946 6537 7980 6545
rect 7946 6477 7980 6499
rect 7946 6465 7980 6477
rect 7946 6409 7980 6427
rect 7946 6393 7980 6409
rect 7946 6341 7980 6355
rect 7946 6321 7980 6341
rect 7946 6273 7980 6283
rect 7946 6249 7980 6273
rect 7946 6205 7980 6211
rect 7946 6177 7980 6205
rect 7946 6137 7980 6139
rect 7946 6105 7980 6137
rect 7946 6035 7980 6067
rect 7946 6033 7980 6035
rect 7946 5967 7980 5995
rect 7946 5961 7980 5967
rect 7946 5899 7980 5923
rect 7946 5889 7980 5899
rect 7946 5831 7980 5851
rect 7946 5817 7980 5831
rect 7946 5763 7980 5779
rect 7946 5745 7980 5763
rect 7946 5695 7980 5707
rect 7946 5673 7980 5695
rect 7946 5627 7980 5635
rect 7946 5601 7980 5627
rect 8042 6545 8076 6571
rect 8042 6537 8076 6545
rect 8042 6477 8076 6499
rect 8042 6465 8076 6477
rect 8042 6409 8076 6427
rect 8042 6393 8076 6409
rect 8042 6341 8076 6355
rect 8042 6321 8076 6341
rect 8042 6273 8076 6283
rect 8042 6249 8076 6273
rect 8042 6205 8076 6211
rect 8042 6177 8076 6205
rect 8042 6137 8076 6139
rect 8042 6105 8076 6137
rect 8042 6035 8076 6067
rect 8042 6033 8076 6035
rect 8042 5967 8076 5995
rect 8042 5961 8076 5967
rect 8042 5899 8076 5923
rect 8042 5889 8076 5899
rect 8042 5831 8076 5851
rect 8042 5817 8076 5831
rect 8042 5763 8076 5779
rect 8042 5745 8076 5763
rect 8042 5695 8076 5707
rect 8042 5673 8076 5695
rect 8042 5627 8076 5635
rect 8042 5601 8076 5627
rect 8138 6545 8172 6571
rect 8138 6537 8172 6545
rect 8138 6477 8172 6499
rect 8138 6465 8172 6477
rect 8138 6409 8172 6427
rect 8138 6393 8172 6409
rect 8138 6341 8172 6355
rect 8138 6321 8172 6341
rect 8138 6273 8172 6283
rect 8138 6249 8172 6273
rect 8138 6205 8172 6211
rect 8138 6177 8172 6205
rect 8138 6137 8172 6139
rect 8138 6105 8172 6137
rect 8138 6035 8172 6067
rect 8138 6033 8172 6035
rect 8138 5967 8172 5995
rect 8138 5961 8172 5967
rect 8138 5899 8172 5923
rect 8138 5889 8172 5899
rect 8138 5831 8172 5851
rect 8138 5817 8172 5831
rect 8138 5763 8172 5779
rect 8138 5745 8172 5763
rect 8138 5695 8172 5707
rect 8138 5673 8172 5695
rect 8138 5627 8172 5635
rect 8138 5601 8172 5627
rect 8234 6545 8268 6571
rect 8234 6537 8268 6545
rect 8234 6477 8268 6499
rect 8234 6465 8268 6477
rect 8234 6409 8268 6427
rect 8234 6393 8268 6409
rect 8234 6341 8268 6355
rect 8234 6321 8268 6341
rect 8234 6273 8268 6283
rect 8234 6249 8268 6273
rect 8234 6205 8268 6211
rect 8234 6177 8268 6205
rect 8234 6137 8268 6139
rect 8234 6105 8268 6137
rect 8234 6035 8268 6067
rect 8234 6033 8268 6035
rect 8234 5967 8268 5995
rect 8234 5961 8268 5967
rect 8234 5899 8268 5923
rect 8234 5889 8268 5899
rect 8234 5831 8268 5851
rect 8234 5817 8268 5831
rect 8234 5763 8268 5779
rect 8234 5745 8268 5763
rect 8234 5695 8268 5707
rect 8234 5673 8268 5695
rect 8234 5627 8268 5635
rect 8234 5601 8268 5627
rect 8330 6545 8364 6571
rect 8330 6537 8364 6545
rect 8330 6477 8364 6499
rect 8330 6465 8364 6477
rect 8330 6409 8364 6427
rect 8330 6393 8364 6409
rect 8330 6341 8364 6355
rect 8330 6321 8364 6341
rect 8330 6273 8364 6283
rect 8330 6249 8364 6273
rect 8330 6205 8364 6211
rect 8330 6177 8364 6205
rect 8330 6137 8364 6139
rect 8330 6105 8364 6137
rect 8330 6035 8364 6067
rect 8330 6033 8364 6035
rect 8330 5967 8364 5995
rect 8330 5961 8364 5967
rect 8330 5899 8364 5923
rect 8330 5889 8364 5899
rect 8330 5831 8364 5851
rect 8330 5817 8364 5831
rect 8330 5763 8364 5779
rect 8330 5745 8364 5763
rect 8330 5695 8364 5707
rect 8330 5673 8364 5695
rect 8330 5627 8364 5635
rect 8330 5601 8364 5627
rect 8426 6545 8460 6571
rect 8426 6537 8460 6545
rect 8426 6477 8460 6499
rect 8426 6465 8460 6477
rect 8426 6409 8460 6427
rect 8426 6393 8460 6409
rect 8426 6341 8460 6355
rect 8426 6321 8460 6341
rect 8426 6273 8460 6283
rect 8426 6249 8460 6273
rect 8426 6205 8460 6211
rect 8426 6177 8460 6205
rect 8426 6137 8460 6139
rect 8426 6105 8460 6137
rect 8426 6035 8460 6067
rect 8426 6033 8460 6035
rect 8426 5967 8460 5995
rect 8426 5961 8460 5967
rect 8426 5899 8460 5923
rect 8426 5889 8460 5899
rect 8426 5831 8460 5851
rect 8426 5817 8460 5831
rect 8426 5763 8460 5779
rect 8426 5745 8460 5763
rect 8426 5695 8460 5707
rect 8426 5673 8460 5695
rect 8426 5627 8460 5635
rect 8426 5601 8460 5627
rect 8522 6545 8556 6571
rect 8522 6537 8556 6545
rect 8522 6477 8556 6499
rect 8522 6465 8556 6477
rect 8522 6409 8556 6427
rect 8522 6393 8556 6409
rect 8522 6341 8556 6355
rect 8522 6321 8556 6341
rect 8522 6273 8556 6283
rect 8522 6249 8556 6273
rect 8522 6205 8556 6211
rect 8522 6177 8556 6205
rect 8522 6137 8556 6139
rect 8522 6105 8556 6137
rect 8522 6035 8556 6067
rect 8522 6033 8556 6035
rect 8522 5967 8556 5995
rect 8522 5961 8556 5967
rect 8522 5899 8556 5923
rect 8522 5889 8556 5899
rect 8522 5831 8556 5851
rect 8522 5817 8556 5831
rect 8522 5763 8556 5779
rect 8522 5745 8556 5763
rect 8522 5695 8556 5707
rect 8522 5673 8556 5695
rect 8522 5627 8556 5635
rect 8522 5601 8556 5627
rect 8618 6545 8652 6571
rect 8618 6537 8652 6545
rect 8618 6477 8652 6499
rect 8618 6465 8652 6477
rect 8618 6409 8652 6427
rect 8618 6393 8652 6409
rect 8618 6341 8652 6355
rect 8618 6321 8652 6341
rect 8618 6273 8652 6283
rect 8618 6249 8652 6273
rect 8618 6205 8652 6211
rect 8618 6177 8652 6205
rect 8618 6137 8652 6139
rect 8618 6105 8652 6137
rect 8618 6035 8652 6067
rect 8618 6033 8652 6035
rect 8618 5967 8652 5995
rect 8618 5961 8652 5967
rect 8618 5899 8652 5923
rect 8618 5889 8652 5899
rect 8618 5831 8652 5851
rect 8618 5817 8652 5831
rect 8618 5763 8652 5779
rect 8618 5745 8652 5763
rect 8618 5695 8652 5707
rect 8618 5673 8652 5695
rect 8618 5627 8652 5635
rect 8618 5601 8652 5627
rect 8714 6545 8748 6571
rect 8714 6537 8748 6545
rect 8714 6477 8748 6499
rect 8714 6465 8748 6477
rect 8714 6409 8748 6427
rect 8714 6393 8748 6409
rect 8714 6341 8748 6355
rect 8714 6321 8748 6341
rect 8714 6273 8748 6283
rect 8714 6249 8748 6273
rect 8714 6205 8748 6211
rect 8714 6177 8748 6205
rect 8714 6137 8748 6139
rect 8714 6105 8748 6137
rect 8714 6035 8748 6067
rect 8714 6033 8748 6035
rect 8714 5967 8748 5995
rect 8714 5961 8748 5967
rect 8714 5899 8748 5923
rect 8714 5889 8748 5899
rect 8714 5831 8748 5851
rect 8714 5817 8748 5831
rect 8714 5763 8748 5779
rect 8714 5745 8748 5763
rect 8714 5695 8748 5707
rect 8714 5673 8748 5695
rect 8714 5627 8748 5635
rect 8714 5601 8748 5627
rect 14670 6710 14704 6744
rect 14958 6725 14992 6759
rect 9268 6547 9302 6573
rect 9268 6539 9302 6547
rect 9268 6479 9302 6501
rect 9268 6467 9302 6479
rect 9268 6411 9302 6429
rect 9268 6395 9302 6411
rect 9268 6343 9302 6357
rect 9268 6323 9302 6343
rect 9268 6275 9302 6285
rect 9268 6251 9302 6275
rect 9268 6207 9302 6213
rect 9268 6179 9302 6207
rect 9268 6139 9302 6141
rect 9268 6107 9302 6139
rect 9268 6037 9302 6069
rect 9268 6035 9302 6037
rect 9268 5969 9302 5997
rect 9268 5963 9302 5969
rect 9268 5901 9302 5925
rect 9268 5891 9302 5901
rect 9268 5833 9302 5853
rect 9268 5819 9302 5833
rect 9268 5765 9302 5781
rect 9268 5747 9302 5765
rect 9268 5697 9302 5709
rect 9268 5675 9302 5697
rect 9268 5629 9302 5637
rect 9268 5603 9302 5629
rect 9364 6547 9398 6573
rect 9364 6539 9398 6547
rect 9364 6479 9398 6501
rect 9364 6467 9398 6479
rect 9364 6411 9398 6429
rect 9364 6395 9398 6411
rect 9364 6343 9398 6357
rect 9364 6323 9398 6343
rect 9364 6275 9398 6285
rect 9364 6251 9398 6275
rect 9364 6207 9398 6213
rect 9364 6179 9398 6207
rect 9364 6139 9398 6141
rect 9364 6107 9398 6139
rect 9364 6037 9398 6069
rect 9364 6035 9398 6037
rect 9364 5969 9398 5997
rect 9364 5963 9398 5969
rect 9364 5901 9398 5925
rect 9364 5891 9398 5901
rect 9364 5833 9398 5853
rect 9364 5819 9398 5833
rect 9364 5765 9398 5781
rect 9364 5747 9398 5765
rect 9364 5697 9398 5709
rect 9364 5675 9398 5697
rect 9364 5629 9398 5637
rect 9364 5603 9398 5629
rect 3836 5356 3870 5390
rect 5300 5360 5334 5394
rect 9460 6547 9494 6573
rect 9460 6539 9494 6547
rect 9460 6479 9494 6501
rect 9460 6467 9494 6479
rect 9460 6411 9494 6429
rect 9460 6395 9494 6411
rect 9460 6343 9494 6357
rect 9460 6323 9494 6343
rect 9460 6275 9494 6285
rect 9460 6251 9494 6275
rect 9460 6207 9494 6213
rect 9460 6179 9494 6207
rect 9460 6139 9494 6141
rect 9460 6107 9494 6139
rect 9460 6037 9494 6069
rect 9460 6035 9494 6037
rect 9460 5969 9494 5997
rect 9460 5963 9494 5969
rect 9460 5901 9494 5925
rect 9460 5891 9494 5901
rect 9460 5833 9494 5853
rect 9460 5819 9494 5833
rect 9460 5765 9494 5781
rect 9460 5747 9494 5765
rect 9460 5697 9494 5709
rect 9460 5675 9494 5697
rect 9460 5629 9494 5637
rect 9460 5603 9494 5629
rect 9556 6547 9590 6573
rect 9556 6539 9590 6547
rect 9556 6479 9590 6501
rect 9556 6467 9590 6479
rect 9556 6411 9590 6429
rect 9556 6395 9590 6411
rect 9556 6343 9590 6357
rect 9556 6323 9590 6343
rect 9556 6275 9590 6285
rect 9556 6251 9590 6275
rect 9556 6207 9590 6213
rect 9556 6179 9590 6207
rect 9556 6139 9590 6141
rect 9556 6107 9590 6139
rect 9556 6037 9590 6069
rect 9556 6035 9590 6037
rect 9556 5969 9590 5997
rect 9556 5963 9590 5969
rect 9556 5901 9590 5925
rect 9556 5891 9590 5901
rect 9556 5833 9590 5853
rect 9556 5819 9590 5833
rect 9556 5765 9590 5781
rect 9556 5747 9590 5765
rect 9556 5697 9590 5709
rect 9556 5675 9590 5697
rect 9556 5629 9590 5637
rect 9556 5603 9590 5629
rect 9652 6547 9686 6573
rect 9652 6539 9686 6547
rect 9652 6479 9686 6501
rect 9652 6467 9686 6479
rect 9652 6411 9686 6429
rect 9652 6395 9686 6411
rect 9652 6343 9686 6357
rect 9652 6323 9686 6343
rect 9652 6275 9686 6285
rect 9652 6251 9686 6275
rect 9652 6207 9686 6213
rect 9652 6179 9686 6207
rect 9652 6139 9686 6141
rect 9652 6107 9686 6139
rect 9652 6037 9686 6069
rect 9652 6035 9686 6037
rect 9652 5969 9686 5997
rect 9652 5963 9686 5969
rect 9652 5901 9686 5925
rect 9652 5891 9686 5901
rect 9652 5833 9686 5853
rect 9652 5819 9686 5833
rect 9652 5765 9686 5781
rect 9652 5747 9686 5765
rect 9652 5697 9686 5709
rect 9652 5675 9686 5697
rect 9652 5629 9686 5637
rect 9652 5603 9686 5629
rect 9748 6547 9782 6573
rect 9748 6539 9782 6547
rect 9748 6479 9782 6501
rect 9748 6467 9782 6479
rect 9748 6411 9782 6429
rect 9748 6395 9782 6411
rect 9748 6343 9782 6357
rect 9748 6323 9782 6343
rect 9748 6275 9782 6285
rect 9748 6251 9782 6275
rect 9748 6207 9782 6213
rect 9748 6179 9782 6207
rect 9748 6139 9782 6141
rect 9748 6107 9782 6139
rect 9748 6037 9782 6069
rect 9748 6035 9782 6037
rect 9748 5969 9782 5997
rect 9748 5963 9782 5969
rect 9748 5901 9782 5925
rect 9748 5891 9782 5901
rect 9748 5833 9782 5853
rect 9748 5819 9782 5833
rect 9748 5765 9782 5781
rect 9748 5747 9782 5765
rect 9748 5697 9782 5709
rect 9748 5675 9782 5697
rect 9748 5629 9782 5637
rect 9748 5603 9782 5629
rect 9844 6547 9878 6573
rect 9844 6539 9878 6547
rect 9844 6479 9878 6501
rect 9844 6467 9878 6479
rect 9844 6411 9878 6429
rect 9844 6395 9878 6411
rect 9844 6343 9878 6357
rect 9844 6323 9878 6343
rect 9844 6275 9878 6285
rect 9844 6251 9878 6275
rect 9844 6207 9878 6213
rect 9844 6179 9878 6207
rect 9844 6139 9878 6141
rect 9844 6107 9878 6139
rect 9844 6037 9878 6069
rect 9844 6035 9878 6037
rect 9844 5969 9878 5997
rect 9844 5963 9878 5969
rect 9844 5901 9878 5925
rect 9844 5891 9878 5901
rect 9844 5833 9878 5853
rect 9844 5819 9878 5833
rect 9844 5765 9878 5781
rect 9844 5747 9878 5765
rect 9844 5697 9878 5709
rect 9844 5675 9878 5697
rect 9844 5629 9878 5637
rect 9844 5603 9878 5629
rect 9940 6547 9974 6573
rect 9940 6539 9974 6547
rect 9940 6479 9974 6501
rect 9940 6467 9974 6479
rect 9940 6411 9974 6429
rect 9940 6395 9974 6411
rect 9940 6343 9974 6357
rect 9940 6323 9974 6343
rect 9940 6275 9974 6285
rect 9940 6251 9974 6275
rect 9940 6207 9974 6213
rect 9940 6179 9974 6207
rect 9940 6139 9974 6141
rect 9940 6107 9974 6139
rect 9940 6037 9974 6069
rect 9940 6035 9974 6037
rect 9940 5969 9974 5997
rect 9940 5963 9974 5969
rect 9940 5901 9974 5925
rect 9940 5891 9974 5901
rect 9940 5833 9974 5853
rect 9940 5819 9974 5833
rect 9940 5765 9974 5781
rect 9940 5747 9974 5765
rect 9940 5697 9974 5709
rect 9940 5675 9974 5697
rect 9940 5629 9974 5637
rect 9940 5603 9974 5629
rect 10036 6547 10070 6573
rect 10036 6539 10070 6547
rect 10036 6479 10070 6501
rect 10036 6467 10070 6479
rect 10036 6411 10070 6429
rect 10036 6395 10070 6411
rect 10036 6343 10070 6357
rect 10036 6323 10070 6343
rect 10036 6275 10070 6285
rect 10036 6251 10070 6275
rect 10036 6207 10070 6213
rect 10036 6179 10070 6207
rect 10036 6139 10070 6141
rect 10036 6107 10070 6139
rect 10036 6037 10070 6069
rect 10036 6035 10070 6037
rect 10036 5969 10070 5997
rect 10036 5963 10070 5969
rect 10036 5901 10070 5925
rect 10036 5891 10070 5901
rect 10036 5833 10070 5853
rect 10036 5819 10070 5833
rect 10036 5765 10070 5781
rect 10036 5747 10070 5765
rect 10036 5697 10070 5709
rect 10036 5675 10070 5697
rect 10036 5629 10070 5637
rect 10036 5603 10070 5629
rect 10132 6547 10166 6573
rect 10132 6539 10166 6547
rect 10132 6479 10166 6501
rect 10132 6467 10166 6479
rect 10132 6411 10166 6429
rect 10132 6395 10166 6411
rect 10132 6343 10166 6357
rect 10132 6323 10166 6343
rect 10132 6275 10166 6285
rect 10132 6251 10166 6275
rect 10132 6207 10166 6213
rect 10132 6179 10166 6207
rect 10132 6139 10166 6141
rect 10132 6107 10166 6139
rect 10132 6037 10166 6069
rect 10132 6035 10166 6037
rect 10132 5969 10166 5997
rect 10132 5963 10166 5969
rect 10132 5901 10166 5925
rect 10132 5891 10166 5901
rect 10132 5833 10166 5853
rect 10132 5819 10166 5833
rect 10132 5765 10166 5781
rect 10132 5747 10166 5765
rect 10132 5697 10166 5709
rect 10132 5675 10166 5697
rect 10132 5629 10166 5637
rect 10132 5603 10166 5629
rect 10228 6547 10262 6573
rect 10228 6539 10262 6547
rect 10228 6479 10262 6501
rect 10228 6467 10262 6479
rect 10228 6411 10262 6429
rect 10228 6395 10262 6411
rect 10228 6343 10262 6357
rect 10228 6323 10262 6343
rect 10228 6275 10262 6285
rect 10228 6251 10262 6275
rect 10228 6207 10262 6213
rect 10228 6179 10262 6207
rect 10228 6139 10262 6141
rect 10228 6107 10262 6139
rect 10228 6037 10262 6069
rect 10228 6035 10262 6037
rect 10228 5969 10262 5997
rect 10228 5963 10262 5969
rect 10228 5901 10262 5925
rect 10228 5891 10262 5901
rect 10228 5833 10262 5853
rect 10228 5819 10262 5833
rect 10228 5765 10262 5781
rect 10228 5747 10262 5765
rect 10228 5697 10262 5709
rect 10228 5675 10262 5697
rect 10228 5629 10262 5637
rect 10228 5603 10262 5629
rect 10324 6547 10358 6573
rect 10324 6539 10358 6547
rect 10324 6479 10358 6501
rect 10324 6467 10358 6479
rect 10324 6411 10358 6429
rect 10324 6395 10358 6411
rect 10324 6343 10358 6357
rect 10324 6323 10358 6343
rect 10324 6275 10358 6285
rect 10324 6251 10358 6275
rect 10324 6207 10358 6213
rect 10324 6179 10358 6207
rect 10324 6139 10358 6141
rect 10324 6107 10358 6139
rect 10324 6037 10358 6069
rect 10324 6035 10358 6037
rect 10324 5969 10358 5997
rect 10324 5963 10358 5969
rect 10324 5901 10358 5925
rect 10324 5891 10358 5901
rect 10324 5833 10358 5853
rect 10324 5819 10358 5833
rect 10324 5765 10358 5781
rect 10324 5747 10358 5765
rect 10324 5697 10358 5709
rect 10324 5675 10358 5697
rect 10324 5629 10358 5637
rect 10324 5603 10358 5629
rect 10420 6547 10454 6573
rect 10420 6539 10454 6547
rect 10420 6479 10454 6501
rect 10420 6467 10454 6479
rect 10420 6411 10454 6429
rect 10420 6395 10454 6411
rect 10420 6343 10454 6357
rect 10420 6323 10454 6343
rect 10420 6275 10454 6285
rect 10420 6251 10454 6275
rect 10420 6207 10454 6213
rect 10420 6179 10454 6207
rect 10420 6139 10454 6141
rect 10420 6107 10454 6139
rect 10420 6037 10454 6069
rect 10420 6035 10454 6037
rect 10420 5969 10454 5997
rect 10420 5963 10454 5969
rect 10420 5901 10454 5925
rect 10420 5891 10454 5901
rect 10420 5833 10454 5853
rect 10420 5819 10454 5833
rect 10420 5765 10454 5781
rect 10420 5747 10454 5765
rect 10420 5697 10454 5709
rect 10420 5675 10454 5697
rect 10420 5629 10454 5637
rect 10420 5603 10454 5629
rect 11034 6543 11068 6569
rect 11034 6535 11068 6543
rect 11034 6475 11068 6497
rect 11034 6463 11068 6475
rect 11034 6407 11068 6425
rect 11034 6391 11068 6407
rect 11034 6339 11068 6353
rect 11034 6319 11068 6339
rect 11034 6271 11068 6281
rect 11034 6247 11068 6271
rect 11034 6203 11068 6209
rect 11034 6175 11068 6203
rect 11034 6135 11068 6137
rect 11034 6103 11068 6135
rect 11034 6033 11068 6065
rect 11034 6031 11068 6033
rect 11034 5965 11068 5993
rect 11034 5959 11068 5965
rect 11034 5897 11068 5921
rect 11034 5887 11068 5897
rect 11034 5829 11068 5849
rect 11034 5815 11068 5829
rect 11034 5761 11068 5777
rect 11034 5743 11068 5761
rect 11034 5693 11068 5705
rect 11034 5671 11068 5693
rect 11034 5625 11068 5633
rect 11034 5599 11068 5625
rect 11130 6543 11164 6569
rect 11130 6535 11164 6543
rect 11130 6475 11164 6497
rect 11130 6463 11164 6475
rect 11130 6407 11164 6425
rect 11130 6391 11164 6407
rect 11130 6339 11164 6353
rect 11130 6319 11164 6339
rect 11130 6271 11164 6281
rect 11130 6247 11164 6271
rect 11130 6203 11164 6209
rect 11130 6175 11164 6203
rect 11130 6135 11164 6137
rect 11130 6103 11164 6135
rect 11130 6033 11164 6065
rect 11130 6031 11164 6033
rect 11130 5965 11164 5993
rect 11130 5959 11164 5965
rect 11130 5897 11164 5921
rect 11130 5887 11164 5897
rect 11130 5829 11164 5849
rect 11130 5815 11164 5829
rect 11130 5761 11164 5777
rect 11130 5743 11164 5761
rect 11130 5693 11164 5705
rect 11130 5671 11164 5693
rect 11130 5625 11164 5633
rect 11130 5599 11164 5625
rect 11226 6543 11260 6569
rect 11226 6535 11260 6543
rect 11226 6475 11260 6497
rect 11226 6463 11260 6475
rect 11226 6407 11260 6425
rect 11226 6391 11260 6407
rect 11226 6339 11260 6353
rect 11226 6319 11260 6339
rect 11226 6271 11260 6281
rect 11226 6247 11260 6271
rect 11226 6203 11260 6209
rect 11226 6175 11260 6203
rect 11226 6135 11260 6137
rect 11226 6103 11260 6135
rect 11226 6033 11260 6065
rect 11226 6031 11260 6033
rect 11226 5965 11260 5993
rect 11226 5959 11260 5965
rect 11226 5897 11260 5921
rect 11226 5887 11260 5897
rect 11226 5829 11260 5849
rect 11226 5815 11260 5829
rect 11226 5761 11260 5777
rect 11226 5743 11260 5761
rect 11226 5693 11260 5705
rect 11226 5671 11260 5693
rect 11226 5625 11260 5633
rect 11226 5599 11260 5625
rect 11322 6543 11356 6569
rect 11322 6535 11356 6543
rect 11322 6475 11356 6497
rect 11322 6463 11356 6475
rect 11322 6407 11356 6425
rect 11322 6391 11356 6407
rect 11322 6339 11356 6353
rect 11322 6319 11356 6339
rect 11322 6271 11356 6281
rect 11322 6247 11356 6271
rect 11322 6203 11356 6209
rect 11322 6175 11356 6203
rect 11322 6135 11356 6137
rect 11322 6103 11356 6135
rect 11322 6033 11356 6065
rect 11322 6031 11356 6033
rect 11322 5965 11356 5993
rect 11322 5959 11356 5965
rect 11322 5897 11356 5921
rect 11322 5887 11356 5897
rect 11322 5829 11356 5849
rect 11322 5815 11356 5829
rect 11322 5761 11356 5777
rect 11322 5743 11356 5761
rect 11322 5693 11356 5705
rect 11322 5671 11356 5693
rect 11322 5625 11356 5633
rect 11322 5599 11356 5625
rect 11418 6543 11452 6569
rect 11418 6535 11452 6543
rect 11418 6475 11452 6497
rect 11418 6463 11452 6475
rect 11418 6407 11452 6425
rect 11418 6391 11452 6407
rect 11418 6339 11452 6353
rect 11418 6319 11452 6339
rect 11418 6271 11452 6281
rect 11418 6247 11452 6271
rect 11418 6203 11452 6209
rect 11418 6175 11452 6203
rect 11418 6135 11452 6137
rect 11418 6103 11452 6135
rect 11418 6033 11452 6065
rect 11418 6031 11452 6033
rect 11418 5965 11452 5993
rect 11418 5959 11452 5965
rect 11418 5897 11452 5921
rect 11418 5887 11452 5897
rect 11418 5829 11452 5849
rect 11418 5815 11452 5829
rect 11418 5761 11452 5777
rect 11418 5743 11452 5761
rect 11418 5693 11452 5705
rect 11418 5671 11452 5693
rect 11418 5625 11452 5633
rect 11418 5599 11452 5625
rect 11514 6543 11548 6569
rect 11514 6535 11548 6543
rect 11514 6475 11548 6497
rect 11514 6463 11548 6475
rect 11514 6407 11548 6425
rect 11514 6391 11548 6407
rect 11514 6339 11548 6353
rect 11514 6319 11548 6339
rect 11514 6271 11548 6281
rect 11514 6247 11548 6271
rect 11514 6203 11548 6209
rect 11514 6175 11548 6203
rect 11514 6135 11548 6137
rect 11514 6103 11548 6135
rect 11514 6033 11548 6065
rect 11514 6031 11548 6033
rect 11514 5965 11548 5993
rect 11514 5959 11548 5965
rect 11514 5897 11548 5921
rect 11514 5887 11548 5897
rect 11514 5829 11548 5849
rect 11514 5815 11548 5829
rect 11514 5761 11548 5777
rect 11514 5743 11548 5761
rect 11514 5693 11548 5705
rect 11514 5671 11548 5693
rect 11514 5625 11548 5633
rect 11514 5599 11548 5625
rect 11610 6543 11644 6569
rect 11610 6535 11644 6543
rect 11610 6475 11644 6497
rect 11610 6463 11644 6475
rect 11610 6407 11644 6425
rect 11610 6391 11644 6407
rect 11610 6339 11644 6353
rect 11610 6319 11644 6339
rect 11610 6271 11644 6281
rect 11610 6247 11644 6271
rect 11610 6203 11644 6209
rect 11610 6175 11644 6203
rect 11610 6135 11644 6137
rect 11610 6103 11644 6135
rect 11610 6033 11644 6065
rect 11610 6031 11644 6033
rect 11610 5965 11644 5993
rect 11610 5959 11644 5965
rect 11610 5897 11644 5921
rect 11610 5887 11644 5897
rect 11610 5829 11644 5849
rect 11610 5815 11644 5829
rect 11610 5761 11644 5777
rect 11610 5743 11644 5761
rect 11610 5693 11644 5705
rect 11610 5671 11644 5693
rect 11610 5625 11644 5633
rect 11610 5599 11644 5625
rect 11706 6543 11740 6569
rect 11706 6535 11740 6543
rect 11706 6475 11740 6497
rect 11706 6463 11740 6475
rect 11706 6407 11740 6425
rect 11706 6391 11740 6407
rect 11706 6339 11740 6353
rect 11706 6319 11740 6339
rect 11706 6271 11740 6281
rect 11706 6247 11740 6271
rect 11706 6203 11740 6209
rect 11706 6175 11740 6203
rect 11706 6135 11740 6137
rect 11706 6103 11740 6135
rect 11706 6033 11740 6065
rect 11706 6031 11740 6033
rect 11706 5965 11740 5993
rect 11706 5959 11740 5965
rect 11706 5897 11740 5921
rect 11706 5887 11740 5897
rect 11706 5829 11740 5849
rect 11706 5815 11740 5829
rect 11706 5761 11740 5777
rect 11706 5743 11740 5761
rect 11706 5693 11740 5705
rect 11706 5671 11740 5693
rect 11706 5625 11740 5633
rect 11706 5599 11740 5625
rect 11802 6543 11836 6569
rect 11802 6535 11836 6543
rect 11802 6475 11836 6497
rect 11802 6463 11836 6475
rect 11802 6407 11836 6425
rect 11802 6391 11836 6407
rect 11802 6339 11836 6353
rect 11802 6319 11836 6339
rect 11802 6271 11836 6281
rect 11802 6247 11836 6271
rect 11802 6203 11836 6209
rect 11802 6175 11836 6203
rect 11802 6135 11836 6137
rect 11802 6103 11836 6135
rect 11802 6033 11836 6065
rect 11802 6031 11836 6033
rect 11802 5965 11836 5993
rect 11802 5959 11836 5965
rect 11802 5897 11836 5921
rect 11802 5887 11836 5897
rect 11802 5829 11836 5849
rect 11802 5815 11836 5829
rect 11802 5761 11836 5777
rect 11802 5743 11836 5761
rect 11802 5693 11836 5705
rect 11802 5671 11836 5693
rect 11802 5625 11836 5633
rect 11802 5599 11836 5625
rect 12424 6521 12458 6547
rect 12424 6513 12458 6521
rect 12424 6453 12458 6475
rect 12424 6441 12458 6453
rect 12424 6385 12458 6403
rect 12424 6369 12458 6385
rect 12424 6317 12458 6331
rect 12424 6297 12458 6317
rect 12424 6249 12458 6259
rect 12424 6225 12458 6249
rect 12424 6181 12458 6187
rect 12424 6153 12458 6181
rect 12424 6113 12458 6115
rect 12424 6081 12458 6113
rect 12424 6011 12458 6043
rect 12424 6009 12458 6011
rect 12424 5943 12458 5971
rect 12424 5937 12458 5943
rect 12424 5875 12458 5899
rect 12424 5865 12458 5875
rect 12424 5807 12458 5827
rect 12424 5793 12458 5807
rect 12424 5739 12458 5755
rect 12424 5721 12458 5739
rect 12424 5671 12458 5683
rect 12424 5649 12458 5671
rect 12424 5603 12458 5611
rect 12424 5577 12458 5603
rect 12520 6521 12554 6547
rect 12520 6513 12554 6521
rect 12520 6453 12554 6475
rect 12520 6441 12554 6453
rect 12520 6385 12554 6403
rect 12520 6369 12554 6385
rect 12520 6317 12554 6331
rect 12520 6297 12554 6317
rect 12520 6249 12554 6259
rect 12520 6225 12554 6249
rect 12520 6181 12554 6187
rect 12520 6153 12554 6181
rect 12520 6113 12554 6115
rect 12520 6081 12554 6113
rect 12520 6011 12554 6043
rect 12520 6009 12554 6011
rect 12520 5943 12554 5971
rect 12520 5937 12554 5943
rect 12520 5875 12554 5899
rect 12520 5865 12554 5875
rect 12520 5807 12554 5827
rect 12520 5793 12554 5807
rect 12520 5739 12554 5755
rect 12520 5721 12554 5739
rect 12520 5671 12554 5683
rect 12520 5649 12554 5671
rect 12520 5603 12554 5611
rect 12520 5577 12554 5603
rect 6866 5356 6900 5390
rect 8330 5360 8364 5394
rect 12616 6521 12650 6547
rect 12616 6513 12650 6521
rect 12616 6453 12650 6475
rect 12616 6441 12650 6453
rect 12616 6385 12650 6403
rect 12616 6369 12650 6385
rect 12616 6317 12650 6331
rect 12616 6297 12650 6317
rect 12616 6249 12650 6259
rect 12616 6225 12650 6249
rect 12616 6181 12650 6187
rect 12616 6153 12650 6181
rect 12616 6113 12650 6115
rect 12616 6081 12650 6113
rect 12616 6011 12650 6043
rect 12616 6009 12650 6011
rect 12616 5943 12650 5971
rect 12616 5937 12650 5943
rect 12616 5875 12650 5899
rect 12616 5865 12650 5875
rect 12616 5807 12650 5827
rect 12616 5793 12650 5807
rect 12616 5739 12650 5755
rect 12616 5721 12650 5739
rect 12616 5671 12650 5683
rect 12616 5649 12650 5671
rect 12616 5603 12650 5611
rect 12616 5577 12650 5603
rect 12712 6521 12746 6547
rect 12712 6513 12746 6521
rect 12712 6453 12746 6475
rect 12712 6441 12746 6453
rect 12712 6385 12746 6403
rect 12712 6369 12746 6385
rect 12712 6317 12746 6331
rect 12712 6297 12746 6317
rect 12712 6249 12746 6259
rect 12712 6225 12746 6249
rect 12712 6181 12746 6187
rect 12712 6153 12746 6181
rect 12712 6113 12746 6115
rect 12712 6081 12746 6113
rect 12712 6011 12746 6043
rect 12712 6009 12746 6011
rect 12712 5943 12746 5971
rect 12712 5937 12746 5943
rect 12712 5875 12746 5899
rect 12712 5865 12746 5875
rect 12712 5807 12746 5827
rect 12712 5793 12746 5807
rect 12712 5739 12746 5755
rect 12712 5721 12746 5739
rect 12712 5671 12746 5683
rect 12712 5649 12746 5671
rect 12712 5603 12746 5611
rect 12712 5577 12746 5603
rect 12808 6521 12842 6547
rect 12808 6513 12842 6521
rect 12808 6453 12842 6475
rect 12808 6441 12842 6453
rect 12808 6385 12842 6403
rect 12808 6369 12842 6385
rect 12808 6317 12842 6331
rect 12808 6297 12842 6317
rect 12808 6249 12842 6259
rect 12808 6225 12842 6249
rect 12808 6181 12842 6187
rect 12808 6153 12842 6181
rect 12808 6113 12842 6115
rect 12808 6081 12842 6113
rect 12808 6011 12842 6043
rect 12808 6009 12842 6011
rect 12808 5943 12842 5971
rect 12808 5937 12842 5943
rect 12808 5875 12842 5899
rect 12808 5865 12842 5875
rect 12808 5807 12842 5827
rect 12808 5793 12842 5807
rect 12808 5739 12842 5755
rect 12808 5721 12842 5739
rect 12808 5671 12842 5683
rect 12808 5649 12842 5671
rect 12808 5603 12842 5611
rect 12808 5577 12842 5603
rect 12904 6521 12938 6547
rect 12904 6513 12938 6521
rect 12904 6453 12938 6475
rect 12904 6441 12938 6453
rect 12904 6385 12938 6403
rect 12904 6369 12938 6385
rect 12904 6317 12938 6331
rect 12904 6297 12938 6317
rect 12904 6249 12938 6259
rect 12904 6225 12938 6249
rect 12904 6181 12938 6187
rect 12904 6153 12938 6181
rect 12904 6113 12938 6115
rect 12904 6081 12938 6113
rect 12904 6011 12938 6043
rect 12904 6009 12938 6011
rect 12904 5943 12938 5971
rect 12904 5937 12938 5943
rect 12904 5875 12938 5899
rect 12904 5865 12938 5875
rect 12904 5807 12938 5827
rect 12904 5793 12938 5807
rect 12904 5739 12938 5755
rect 12904 5721 12938 5739
rect 12904 5671 12938 5683
rect 12904 5649 12938 5671
rect 12904 5603 12938 5611
rect 12904 5577 12938 5603
rect 13000 6521 13034 6547
rect 13000 6513 13034 6521
rect 13000 6453 13034 6475
rect 13000 6441 13034 6453
rect 13000 6385 13034 6403
rect 13000 6369 13034 6385
rect 13000 6317 13034 6331
rect 13000 6297 13034 6317
rect 13000 6249 13034 6259
rect 13000 6225 13034 6249
rect 13000 6181 13034 6187
rect 13000 6153 13034 6181
rect 13000 6113 13034 6115
rect 13000 6081 13034 6113
rect 13000 6011 13034 6043
rect 13000 6009 13034 6011
rect 13000 5943 13034 5971
rect 13000 5937 13034 5943
rect 13000 5875 13034 5899
rect 13000 5865 13034 5875
rect 13000 5807 13034 5827
rect 13000 5793 13034 5807
rect 13000 5739 13034 5755
rect 13000 5721 13034 5739
rect 13000 5671 13034 5683
rect 13000 5649 13034 5671
rect 13000 5603 13034 5611
rect 13000 5577 13034 5603
rect 13096 6521 13130 6547
rect 13096 6513 13130 6521
rect 13096 6453 13130 6475
rect 13096 6441 13130 6453
rect 13096 6385 13130 6403
rect 13096 6369 13130 6385
rect 13096 6317 13130 6331
rect 13096 6297 13130 6317
rect 13096 6249 13130 6259
rect 13096 6225 13130 6249
rect 13096 6181 13130 6187
rect 13096 6153 13130 6181
rect 13096 6113 13130 6115
rect 13096 6081 13130 6113
rect 13096 6011 13130 6043
rect 13096 6009 13130 6011
rect 13096 5943 13130 5971
rect 13096 5937 13130 5943
rect 13096 5875 13130 5899
rect 13096 5865 13130 5875
rect 13096 5807 13130 5827
rect 13096 5793 13130 5807
rect 13096 5739 13130 5755
rect 13096 5721 13130 5739
rect 13096 5671 13130 5683
rect 13096 5649 13130 5671
rect 13096 5603 13130 5611
rect 13096 5577 13130 5603
rect 13192 6521 13226 6547
rect 13192 6513 13226 6521
rect 13192 6453 13226 6475
rect 13192 6441 13226 6453
rect 13192 6385 13226 6403
rect 13192 6369 13226 6385
rect 13192 6317 13226 6331
rect 13192 6297 13226 6317
rect 13192 6249 13226 6259
rect 13192 6225 13226 6249
rect 13192 6181 13226 6187
rect 13192 6153 13226 6181
rect 13192 6113 13226 6115
rect 13192 6081 13226 6113
rect 13192 6011 13226 6043
rect 13192 6009 13226 6011
rect 13192 5943 13226 5971
rect 13192 5937 13226 5943
rect 13192 5875 13226 5899
rect 13192 5865 13226 5875
rect 13192 5807 13226 5827
rect 13192 5793 13226 5807
rect 13192 5739 13226 5755
rect 13192 5721 13226 5739
rect 13192 5671 13226 5683
rect 13192 5649 13226 5671
rect 13192 5603 13226 5611
rect 13192 5577 13226 5603
rect 13288 6521 13322 6547
rect 13288 6513 13322 6521
rect 13288 6453 13322 6475
rect 13288 6441 13322 6453
rect 13288 6385 13322 6403
rect 13288 6369 13322 6385
rect 13288 6317 13322 6331
rect 13288 6297 13322 6317
rect 13288 6249 13322 6259
rect 13288 6225 13322 6249
rect 13288 6181 13322 6187
rect 13288 6153 13322 6181
rect 13288 6113 13322 6115
rect 13288 6081 13322 6113
rect 13288 6011 13322 6043
rect 13288 6009 13322 6011
rect 13288 5943 13322 5971
rect 13288 5937 13322 5943
rect 13288 5875 13322 5899
rect 13288 5865 13322 5875
rect 13288 5807 13322 5827
rect 13288 5793 13322 5807
rect 13288 5739 13322 5755
rect 13288 5721 13322 5739
rect 13288 5671 13322 5683
rect 13288 5649 13322 5671
rect 13288 5603 13322 5611
rect 13288 5577 13322 5603
rect 13384 6521 13418 6547
rect 13384 6513 13418 6521
rect 13384 6453 13418 6475
rect 13384 6441 13418 6453
rect 13384 6385 13418 6403
rect 13384 6369 13418 6385
rect 13384 6317 13418 6331
rect 13384 6297 13418 6317
rect 13384 6249 13418 6259
rect 13384 6225 13418 6249
rect 13384 6181 13418 6187
rect 13384 6153 13418 6181
rect 13384 6113 13418 6115
rect 13384 6081 13418 6113
rect 13384 6011 13418 6043
rect 13384 6009 13418 6011
rect 13384 5943 13418 5971
rect 13384 5937 13418 5943
rect 13384 5875 13418 5899
rect 13384 5865 13418 5875
rect 13384 5807 13418 5827
rect 13384 5793 13418 5807
rect 13384 5739 13418 5755
rect 13384 5721 13418 5739
rect 13384 5671 13418 5683
rect 13384 5649 13418 5671
rect 13384 5603 13418 5611
rect 13384 5577 13418 5603
rect 13480 6521 13514 6547
rect 13480 6513 13514 6521
rect 13480 6453 13514 6475
rect 13480 6441 13514 6453
rect 13480 6385 13514 6403
rect 13480 6369 13514 6385
rect 13480 6317 13514 6331
rect 13480 6297 13514 6317
rect 13480 6249 13514 6259
rect 13480 6225 13514 6249
rect 13480 6181 13514 6187
rect 13480 6153 13514 6181
rect 13480 6113 13514 6115
rect 13480 6081 13514 6113
rect 13480 6011 13514 6043
rect 13480 6009 13514 6011
rect 13480 5943 13514 5971
rect 13480 5937 13514 5943
rect 13480 5875 13514 5899
rect 13480 5865 13514 5875
rect 13480 5807 13514 5827
rect 13480 5793 13514 5807
rect 13480 5739 13514 5755
rect 13480 5721 13514 5739
rect 13480 5671 13514 5683
rect 13480 5649 13514 5671
rect 13480 5603 13514 5611
rect 13480 5577 13514 5603
rect 13576 6521 13610 6547
rect 13576 6513 13610 6521
rect 13576 6453 13610 6475
rect 13576 6441 13610 6453
rect 13576 6385 13610 6403
rect 13576 6369 13610 6385
rect 13576 6317 13610 6331
rect 13576 6297 13610 6317
rect 13576 6249 13610 6259
rect 13576 6225 13610 6249
rect 13576 6181 13610 6187
rect 13576 6153 13610 6181
rect 13576 6113 13610 6115
rect 13576 6081 13610 6113
rect 13576 6011 13610 6043
rect 13576 6009 13610 6011
rect 13576 5943 13610 5971
rect 13576 5937 13610 5943
rect 13576 5875 13610 5899
rect 13576 5865 13610 5875
rect 13576 5807 13610 5827
rect 13576 5793 13610 5807
rect 13576 5739 13610 5755
rect 13576 5721 13610 5739
rect 13576 5671 13610 5683
rect 13576 5649 13610 5671
rect 13576 5603 13610 5611
rect 13576 5577 13610 5603
rect 14190 6517 14224 6543
rect 14190 6509 14224 6517
rect 14190 6449 14224 6471
rect 14190 6437 14224 6449
rect 14190 6381 14224 6399
rect 14190 6365 14224 6381
rect 14190 6313 14224 6327
rect 14190 6293 14224 6313
rect 14190 6245 14224 6255
rect 14190 6221 14224 6245
rect 14190 6177 14224 6183
rect 14190 6149 14224 6177
rect 14190 6109 14224 6111
rect 14190 6077 14224 6109
rect 14190 6007 14224 6039
rect 14190 6005 14224 6007
rect 14190 5939 14224 5967
rect 14190 5933 14224 5939
rect 14190 5871 14224 5895
rect 14190 5861 14224 5871
rect 14190 5803 14224 5823
rect 14190 5789 14224 5803
rect 14190 5735 14224 5751
rect 14190 5717 14224 5735
rect 14190 5667 14224 5679
rect 14190 5645 14224 5667
rect 14190 5599 14224 5607
rect 14190 5573 14224 5599
rect 14286 6517 14320 6543
rect 14286 6509 14320 6517
rect 14286 6449 14320 6471
rect 14286 6437 14320 6449
rect 14286 6381 14320 6399
rect 14286 6365 14320 6381
rect 14286 6313 14320 6327
rect 14286 6293 14320 6313
rect 14286 6245 14320 6255
rect 14286 6221 14320 6245
rect 14286 6177 14320 6183
rect 14286 6149 14320 6177
rect 14286 6109 14320 6111
rect 14286 6077 14320 6109
rect 14286 6007 14320 6039
rect 14286 6005 14320 6007
rect 14286 5939 14320 5967
rect 14286 5933 14320 5939
rect 14286 5871 14320 5895
rect 14286 5861 14320 5871
rect 14286 5803 14320 5823
rect 14286 5789 14320 5803
rect 14286 5735 14320 5751
rect 14286 5717 14320 5735
rect 14286 5667 14320 5679
rect 14286 5645 14320 5667
rect 14286 5599 14320 5607
rect 14286 5573 14320 5599
rect 9954 5354 9988 5388
rect 14382 6517 14416 6543
rect 14382 6509 14416 6517
rect 14382 6449 14416 6471
rect 14382 6437 14416 6449
rect 14382 6381 14416 6399
rect 14382 6365 14416 6381
rect 14382 6313 14416 6327
rect 14382 6293 14416 6313
rect 14382 6245 14416 6255
rect 14382 6221 14416 6245
rect 14382 6177 14416 6183
rect 14382 6149 14416 6177
rect 14382 6109 14416 6111
rect 14382 6077 14416 6109
rect 14382 6007 14416 6039
rect 14382 6005 14416 6007
rect 14382 5939 14416 5967
rect 14382 5933 14416 5939
rect 14382 5871 14416 5895
rect 14382 5861 14416 5871
rect 14382 5803 14416 5823
rect 14382 5789 14416 5803
rect 14382 5735 14416 5751
rect 14382 5717 14416 5735
rect 14382 5667 14416 5679
rect 14382 5645 14416 5667
rect 14382 5599 14416 5607
rect 14382 5573 14416 5599
rect 14478 6517 14512 6543
rect 14478 6509 14512 6517
rect 14478 6449 14512 6471
rect 14478 6437 14512 6449
rect 14478 6381 14512 6399
rect 14478 6365 14512 6381
rect 14478 6313 14512 6327
rect 14478 6293 14512 6313
rect 14478 6245 14512 6255
rect 14478 6221 14512 6245
rect 14478 6177 14512 6183
rect 14478 6149 14512 6177
rect 14478 6109 14512 6111
rect 14478 6077 14512 6109
rect 14478 6007 14512 6039
rect 14478 6005 14512 6007
rect 14478 5939 14512 5967
rect 14478 5933 14512 5939
rect 14478 5871 14512 5895
rect 14478 5861 14512 5871
rect 14478 5803 14512 5823
rect 14478 5789 14512 5803
rect 14478 5735 14512 5751
rect 14478 5717 14512 5735
rect 14478 5667 14512 5679
rect 14478 5645 14512 5667
rect 14478 5599 14512 5607
rect 14478 5573 14512 5599
rect 14574 6517 14608 6543
rect 14574 6509 14608 6517
rect 14574 6449 14608 6471
rect 14574 6437 14608 6449
rect 14574 6381 14608 6399
rect 14574 6365 14608 6381
rect 14574 6313 14608 6327
rect 14574 6293 14608 6313
rect 14574 6245 14608 6255
rect 14574 6221 14608 6245
rect 14574 6177 14608 6183
rect 14574 6149 14608 6177
rect 14574 6109 14608 6111
rect 14574 6077 14608 6109
rect 14574 6007 14608 6039
rect 14574 6005 14608 6007
rect 14574 5939 14608 5967
rect 14574 5933 14608 5939
rect 14574 5871 14608 5895
rect 14574 5861 14608 5871
rect 14574 5803 14608 5823
rect 14574 5789 14608 5803
rect 14574 5735 14608 5751
rect 14574 5717 14608 5735
rect 14574 5667 14608 5679
rect 14574 5645 14608 5667
rect 14574 5599 14608 5607
rect 14574 5573 14608 5599
rect 14670 6517 14704 6543
rect 14670 6509 14704 6517
rect 14670 6449 14704 6471
rect 14670 6437 14704 6449
rect 14670 6381 14704 6399
rect 14670 6365 14704 6381
rect 14670 6313 14704 6327
rect 14670 6293 14704 6313
rect 14670 6245 14704 6255
rect 14670 6221 14704 6245
rect 14670 6177 14704 6183
rect 14670 6149 14704 6177
rect 14670 6109 14704 6111
rect 14670 6077 14704 6109
rect 14670 6007 14704 6039
rect 14670 6005 14704 6007
rect 14670 5939 14704 5967
rect 14670 5933 14704 5939
rect 14670 5871 14704 5895
rect 14670 5861 14704 5871
rect 14670 5803 14704 5823
rect 14670 5789 14704 5803
rect 14670 5735 14704 5751
rect 14670 5717 14704 5735
rect 14670 5667 14704 5679
rect 14670 5645 14704 5667
rect 14670 5599 14704 5607
rect 14670 5573 14704 5599
rect 14766 6517 14800 6543
rect 14766 6509 14800 6517
rect 14766 6449 14800 6471
rect 14766 6437 14800 6449
rect 14766 6381 14800 6399
rect 14766 6365 14800 6381
rect 14766 6313 14800 6327
rect 14766 6293 14800 6313
rect 14766 6245 14800 6255
rect 14766 6221 14800 6245
rect 14766 6177 14800 6183
rect 14766 6149 14800 6177
rect 14766 6109 14800 6111
rect 14766 6077 14800 6109
rect 14766 6007 14800 6039
rect 14766 6005 14800 6007
rect 14766 5939 14800 5967
rect 14766 5933 14800 5939
rect 14766 5871 14800 5895
rect 14766 5861 14800 5871
rect 14766 5803 14800 5823
rect 14766 5789 14800 5803
rect 14766 5735 14800 5751
rect 14766 5717 14800 5735
rect 14766 5667 14800 5679
rect 14766 5645 14800 5667
rect 14766 5599 14800 5607
rect 14766 5573 14800 5599
rect 14862 6517 14896 6543
rect 14862 6509 14896 6517
rect 14862 6449 14896 6471
rect 14862 6437 14896 6449
rect 14862 6381 14896 6399
rect 14862 6365 14896 6381
rect 14862 6313 14896 6327
rect 14862 6293 14896 6313
rect 14862 6245 14896 6255
rect 14862 6221 14896 6245
rect 14862 6177 14896 6183
rect 14862 6149 14896 6177
rect 14862 6109 14896 6111
rect 14862 6077 14896 6109
rect 14862 6007 14896 6039
rect 14862 6005 14896 6007
rect 14862 5939 14896 5967
rect 14862 5933 14896 5939
rect 14862 5871 14896 5895
rect 14862 5861 14896 5871
rect 14862 5803 14896 5823
rect 14862 5789 14896 5803
rect 14862 5735 14896 5751
rect 14862 5717 14896 5735
rect 14862 5667 14896 5679
rect 14862 5645 14896 5667
rect 14862 5599 14896 5607
rect 14862 5573 14896 5599
rect 14958 6517 14992 6543
rect 14958 6509 14992 6517
rect 14958 6449 14992 6471
rect 14958 6437 14992 6449
rect 14958 6381 14992 6399
rect 14958 6365 14992 6381
rect 14958 6313 14992 6327
rect 14958 6293 14992 6313
rect 14958 6245 14992 6255
rect 14958 6221 14992 6245
rect 14958 6177 14992 6183
rect 14958 6149 14992 6177
rect 14958 6109 14992 6111
rect 14958 6077 14992 6109
rect 14958 6007 14992 6039
rect 15614 6148 15648 6182
rect 14958 6005 14992 6007
rect 14958 5939 14992 5967
rect 14958 5933 14992 5939
rect 14958 5871 14992 5895
rect 14958 5861 14992 5871
rect 14958 5803 14992 5823
rect 14958 5789 14992 5803
rect 14958 5735 14992 5751
rect 14958 5717 14992 5735
rect 14958 5667 14992 5679
rect 14958 5645 14992 5667
rect 14958 5599 14992 5607
rect 14958 5573 14992 5599
rect 15518 5861 15552 5879
rect 15518 5845 15552 5861
rect 15518 5793 15552 5807
rect 15518 5773 15552 5793
rect 15518 5725 15552 5735
rect 15518 5701 15552 5725
rect 15518 5657 15552 5663
rect 15518 5629 15552 5657
rect 15518 5589 15552 5591
rect 15518 5557 15552 5589
rect 11418 5358 11452 5392
rect 15518 5487 15552 5519
rect 15518 5485 15552 5487
rect -868 5317 -834 5345
rect 13110 5328 13144 5362
rect 14574 5332 14608 5366
rect 15518 5419 15552 5447
rect 15518 5413 15552 5419
rect 15518 5351 15552 5375
rect 15518 5341 15552 5351
rect -868 5311 -834 5317
rect -868 5249 -834 5273
rect -868 5239 -834 5249
rect -868 5181 -834 5201
rect -868 5167 -834 5181
rect -868 5113 -834 5129
rect 15518 5283 15552 5303
rect 15518 5269 15552 5283
rect 15518 5215 15552 5231
rect 15518 5197 15552 5215
rect 15518 5147 15552 5159
rect 15518 5125 15552 5147
rect -868 5095 -834 5113
rect -868 5045 -834 5057
rect -868 5023 -834 5045
rect 1580 5090 1614 5124
rect 4536 5074 4570 5108
rect 7566 5074 7600 5108
rect 10654 5072 10688 5106
rect -868 4977 -834 4985
rect -868 4951 -834 4977
rect 1484 4903 1518 4929
rect 1484 4895 1518 4903
rect 1484 4835 1518 4857
rect 1484 4823 1518 4835
rect -1067 4735 -1033 4769
rect 1484 4767 1518 4785
rect 1484 4751 1518 4767
rect 1484 4699 1518 4713
rect 1484 4679 1518 4699
rect 1484 4631 1518 4641
rect 1484 4607 1518 4631
rect 1484 4563 1518 4569
rect 1484 4535 1518 4563
rect 1484 4495 1518 4497
rect 1484 4463 1518 4495
rect 1484 4393 1518 4425
rect 1484 4391 1518 4393
rect 1484 4325 1518 4353
rect 1484 4319 1518 4325
rect 1484 4257 1518 4281
rect 1484 4247 1518 4257
rect 1484 4189 1518 4209
rect 1484 4175 1518 4189
rect 1484 4121 1518 4137
rect 1484 4103 1518 4121
rect 1484 4053 1518 4065
rect 1484 4031 1518 4053
rect 1484 3985 1518 3993
rect 1484 3959 1518 3985
rect 1580 4903 1614 4929
rect 1580 4895 1614 4903
rect 1580 4835 1614 4857
rect 1580 4823 1614 4835
rect 1580 4767 1614 4785
rect 1580 4751 1614 4767
rect 1580 4699 1614 4713
rect 1580 4679 1614 4699
rect 1580 4631 1614 4641
rect 1580 4607 1614 4631
rect 1580 4563 1614 4569
rect 1580 4535 1614 4563
rect 1580 4495 1614 4497
rect 1580 4463 1614 4495
rect 1580 4393 1614 4425
rect 1580 4391 1614 4393
rect 1580 4325 1614 4353
rect 1580 4319 1614 4325
rect 1580 4257 1614 4281
rect 1580 4247 1614 4257
rect 1580 4189 1614 4209
rect 1580 4175 1614 4189
rect 1580 4121 1614 4137
rect 1580 4103 1614 4121
rect 1580 4053 1614 4065
rect 1580 4031 1614 4053
rect 1580 3985 1614 3993
rect 1580 3959 1614 3985
rect 1676 4903 1710 4929
rect 1676 4895 1710 4903
rect 1676 4835 1710 4857
rect 1676 4823 1710 4835
rect 1676 4767 1710 4785
rect 1676 4751 1710 4767
rect 1676 4699 1710 4713
rect 1676 4679 1710 4699
rect 1676 4631 1710 4641
rect 1676 4607 1710 4631
rect 1676 4563 1710 4569
rect 1676 4535 1710 4563
rect 1676 4495 1710 4497
rect 1676 4463 1710 4495
rect 1676 4393 1710 4425
rect 1676 4391 1710 4393
rect 1676 4325 1710 4353
rect 1676 4319 1710 4325
rect 1676 4257 1710 4281
rect 1676 4247 1710 4257
rect 1676 4189 1710 4209
rect 1676 4175 1710 4189
rect 1676 4121 1710 4137
rect 1676 4103 1710 4121
rect 1676 4053 1710 4065
rect 1676 4031 1710 4053
rect 1676 3985 1710 3993
rect 1676 3959 1710 3985
rect 1772 4903 1806 4929
rect 1772 4895 1806 4903
rect 1772 4835 1806 4857
rect 1772 4823 1806 4835
rect 1772 4767 1806 4785
rect 1772 4751 1806 4767
rect 1772 4699 1806 4713
rect 1772 4679 1806 4699
rect 1772 4631 1806 4641
rect 1772 4607 1806 4631
rect 1772 4563 1806 4569
rect 1772 4535 1806 4563
rect 1772 4495 1806 4497
rect 1772 4463 1806 4495
rect 1772 4393 1806 4425
rect 1772 4391 1806 4393
rect 1772 4325 1806 4353
rect 1772 4319 1806 4325
rect 1772 4257 1806 4281
rect 1772 4247 1806 4257
rect 1772 4189 1806 4209
rect 1772 4175 1806 4189
rect 1772 4121 1806 4137
rect 1772 4103 1806 4121
rect 1772 4053 1806 4065
rect 1772 4031 1806 4053
rect 1772 3985 1806 3993
rect 1772 3959 1806 3985
rect 13810 5046 13844 5080
rect 1868 4903 1902 4929
rect 1868 4895 1902 4903
rect 1868 4835 1902 4857
rect 1868 4823 1902 4835
rect 1868 4767 1902 4785
rect 1868 4751 1902 4767
rect 1868 4699 1902 4713
rect 1868 4679 1902 4699
rect 1868 4631 1902 4641
rect 1868 4607 1902 4631
rect 1868 4563 1902 4569
rect 1868 4535 1902 4563
rect 1868 4495 1902 4497
rect 1868 4463 1902 4495
rect 1868 4393 1902 4425
rect 1868 4391 1902 4393
rect 1868 4325 1902 4353
rect 1868 4319 1902 4325
rect 1868 4257 1902 4281
rect 1868 4247 1902 4257
rect 1868 4189 1902 4209
rect 1868 4175 1902 4189
rect 1868 4121 1902 4137
rect 1868 4103 1902 4121
rect 1868 4053 1902 4065
rect 1868 4031 1902 4053
rect 1868 3985 1902 3993
rect 1868 3959 1902 3985
rect 4440 4887 4474 4913
rect 4440 4879 4474 4887
rect 4440 4819 4474 4841
rect 4440 4807 4474 4819
rect 4440 4751 4474 4769
rect 4440 4735 4474 4751
rect 4440 4683 4474 4697
rect 4440 4663 4474 4683
rect 4440 4615 4474 4625
rect 4440 4591 4474 4615
rect 4440 4547 4474 4553
rect 4440 4519 4474 4547
rect 4440 4479 4474 4481
rect 4440 4447 4474 4479
rect 4440 4377 4474 4409
rect 4440 4375 4474 4377
rect 4440 4309 4474 4337
rect 4440 4303 4474 4309
rect 4440 4241 4474 4265
rect 4440 4231 4474 4241
rect 4440 4173 4474 4193
rect 4440 4159 4474 4173
rect 4440 4105 4474 4121
rect 4440 4087 4474 4105
rect 4440 4037 4474 4049
rect 4440 4015 4474 4037
rect 4440 3969 4474 3977
rect 4440 3943 4474 3969
rect 4536 4887 4570 4913
rect 4536 4879 4570 4887
rect 4536 4819 4570 4841
rect 4536 4807 4570 4819
rect 4536 4751 4570 4769
rect 4536 4735 4570 4751
rect 4536 4683 4570 4697
rect 4536 4663 4570 4683
rect 4536 4615 4570 4625
rect 4536 4591 4570 4615
rect 4536 4547 4570 4553
rect 4536 4519 4570 4547
rect 4536 4479 4570 4481
rect 4536 4447 4570 4479
rect 4536 4377 4570 4409
rect 4536 4375 4570 4377
rect 4536 4309 4570 4337
rect 4536 4303 4570 4309
rect 4536 4241 4570 4265
rect 4536 4231 4570 4241
rect 4536 4173 4570 4193
rect 4536 4159 4570 4173
rect 4536 4105 4570 4121
rect 4536 4087 4570 4105
rect 4536 4037 4570 4049
rect 4536 4015 4570 4037
rect 4536 3969 4570 3977
rect 4536 3943 4570 3969
rect 4632 4887 4666 4913
rect 4632 4879 4666 4887
rect 4632 4819 4666 4841
rect 4632 4807 4666 4819
rect 4632 4751 4666 4769
rect 4632 4735 4666 4751
rect 4632 4683 4666 4697
rect 4632 4663 4666 4683
rect 4632 4615 4666 4625
rect 4632 4591 4666 4615
rect 4632 4547 4666 4553
rect 4632 4519 4666 4547
rect 4632 4479 4666 4481
rect 4632 4447 4666 4479
rect 4632 4377 4666 4409
rect 4632 4375 4666 4377
rect 4632 4309 4666 4337
rect 4632 4303 4666 4309
rect 4632 4241 4666 4265
rect 4632 4231 4666 4241
rect 4632 4173 4666 4193
rect 4632 4159 4666 4173
rect 4632 4105 4666 4121
rect 4632 4087 4666 4105
rect 4632 4037 4666 4049
rect 4632 4015 4666 4037
rect 4632 3969 4666 3977
rect 4632 3943 4666 3969
rect 4728 4887 4762 4913
rect 4728 4879 4762 4887
rect 4728 4819 4762 4841
rect 4728 4807 4762 4819
rect 4728 4751 4762 4769
rect 4728 4735 4762 4751
rect 4728 4683 4762 4697
rect 4728 4663 4762 4683
rect 4728 4615 4762 4625
rect 4728 4591 4762 4615
rect 4728 4547 4762 4553
rect 4728 4519 4762 4547
rect 4728 4479 4762 4481
rect 4728 4447 4762 4479
rect 4728 4377 4762 4409
rect 4728 4375 4762 4377
rect 4728 4309 4762 4337
rect 4728 4303 4762 4309
rect 4728 4241 4762 4265
rect 4728 4231 4762 4241
rect 4728 4173 4762 4193
rect 4728 4159 4762 4173
rect 4728 4105 4762 4121
rect 4728 4087 4762 4105
rect 4728 4037 4762 4049
rect 4728 4015 4762 4037
rect 4728 3969 4762 3977
rect 4728 3943 4762 3969
rect 4824 4887 4858 4913
rect 4824 4879 4858 4887
rect 4824 4819 4858 4841
rect 4824 4807 4858 4819
rect 4824 4751 4858 4769
rect 4824 4735 4858 4751
rect 4824 4683 4858 4697
rect 4824 4663 4858 4683
rect 4824 4615 4858 4625
rect 4824 4591 4858 4615
rect 4824 4547 4858 4553
rect 4824 4519 4858 4547
rect 4824 4479 4858 4481
rect 4824 4447 4858 4479
rect 4824 4377 4858 4409
rect 4824 4375 4858 4377
rect 4824 4309 4858 4337
rect 4824 4303 4858 4309
rect 4824 4241 4858 4265
rect 4824 4231 4858 4241
rect 4824 4173 4858 4193
rect 4824 4159 4858 4173
rect 4824 4105 4858 4121
rect 4824 4087 4858 4105
rect 4824 4037 4858 4049
rect 4824 4015 4858 4037
rect 4824 3969 4858 3977
rect 4824 3943 4858 3969
rect 7470 4887 7504 4913
rect 7470 4879 7504 4887
rect 7470 4819 7504 4841
rect 7470 4807 7504 4819
rect 7470 4751 7504 4769
rect 7470 4735 7504 4751
rect 7470 4683 7504 4697
rect 7470 4663 7504 4683
rect 7470 4615 7504 4625
rect 7470 4591 7504 4615
rect 7470 4547 7504 4553
rect 7470 4519 7504 4547
rect 7470 4479 7504 4481
rect 7470 4447 7504 4479
rect 7470 4377 7504 4409
rect 7470 4375 7504 4377
rect 7470 4309 7504 4337
rect 7470 4303 7504 4309
rect 7470 4241 7504 4265
rect 7470 4231 7504 4241
rect 7470 4173 7504 4193
rect 7470 4159 7504 4173
rect 7470 4105 7504 4121
rect 7470 4087 7504 4105
rect 7470 4037 7504 4049
rect 7470 4015 7504 4037
rect 7470 3969 7504 3977
rect 7470 3943 7504 3969
rect 7566 4887 7600 4913
rect 7566 4879 7600 4887
rect 7566 4819 7600 4841
rect 7566 4807 7600 4819
rect 7566 4751 7600 4769
rect 7566 4735 7600 4751
rect 7566 4683 7600 4697
rect 7566 4663 7600 4683
rect 7566 4615 7600 4625
rect 7566 4591 7600 4615
rect 7566 4547 7600 4553
rect 7566 4519 7600 4547
rect 7566 4479 7600 4481
rect 7566 4447 7600 4479
rect 7566 4377 7600 4409
rect 7566 4375 7600 4377
rect 7566 4309 7600 4337
rect 7566 4303 7600 4309
rect 7566 4241 7600 4265
rect 7566 4231 7600 4241
rect 7566 4173 7600 4193
rect 7566 4159 7600 4173
rect 7566 4105 7600 4121
rect 7566 4087 7600 4105
rect 7566 4037 7600 4049
rect 7566 4015 7600 4037
rect 7566 3969 7600 3977
rect 7566 3943 7600 3969
rect 1580 3743 1614 3777
rect 7662 4887 7696 4913
rect 7662 4879 7696 4887
rect 7662 4819 7696 4841
rect 7662 4807 7696 4819
rect 7662 4751 7696 4769
rect 7662 4735 7696 4751
rect 7662 4683 7696 4697
rect 7662 4663 7696 4683
rect 7662 4615 7696 4625
rect 7662 4591 7696 4615
rect 7662 4547 7696 4553
rect 7662 4519 7696 4547
rect 7662 4479 7696 4481
rect 7662 4447 7696 4479
rect 7662 4377 7696 4409
rect 7662 4375 7696 4377
rect 7662 4309 7696 4337
rect 7662 4303 7696 4309
rect 7662 4241 7696 4265
rect 7662 4231 7696 4241
rect 7662 4173 7696 4193
rect 7662 4159 7696 4173
rect 7662 4105 7696 4121
rect 7662 4087 7696 4105
rect 7662 4037 7696 4049
rect 7662 4015 7696 4037
rect 7662 3969 7696 3977
rect 7662 3943 7696 3969
rect 7758 4887 7792 4913
rect 7758 4879 7792 4887
rect 7758 4819 7792 4841
rect 7758 4807 7792 4819
rect 7758 4751 7792 4769
rect 7758 4735 7792 4751
rect 7758 4683 7792 4697
rect 7758 4663 7792 4683
rect 7758 4615 7792 4625
rect 7758 4591 7792 4615
rect 7758 4547 7792 4553
rect 7758 4519 7792 4547
rect 7758 4479 7792 4481
rect 7758 4447 7792 4479
rect 7758 4377 7792 4409
rect 7758 4375 7792 4377
rect 7758 4309 7792 4337
rect 7758 4303 7792 4309
rect 7758 4241 7792 4265
rect 7758 4231 7792 4241
rect 7758 4173 7792 4193
rect 7758 4159 7792 4173
rect 7758 4105 7792 4121
rect 7758 4087 7792 4105
rect 7758 4037 7792 4049
rect 7758 4015 7792 4037
rect 7758 3969 7792 3977
rect 7758 3943 7792 3969
rect 15518 5079 15552 5087
rect 15518 5053 15552 5079
rect 15518 5011 15552 5015
rect 7854 4887 7888 4913
rect 7854 4879 7888 4887
rect 7854 4819 7888 4841
rect 7854 4807 7888 4819
rect 7854 4751 7888 4769
rect 7854 4735 7888 4751
rect 7854 4683 7888 4697
rect 7854 4663 7888 4683
rect 7854 4615 7888 4625
rect 7854 4591 7888 4615
rect 7854 4547 7888 4553
rect 7854 4519 7888 4547
rect 7854 4479 7888 4481
rect 7854 4447 7888 4479
rect 7854 4377 7888 4409
rect 7854 4375 7888 4377
rect 7854 4309 7888 4337
rect 7854 4303 7888 4309
rect 7854 4241 7888 4265
rect 7854 4231 7888 4241
rect 7854 4173 7888 4193
rect 7854 4159 7888 4173
rect 7854 4105 7888 4121
rect 7854 4087 7888 4105
rect 7854 4037 7888 4049
rect 7854 4015 7888 4037
rect 7854 3969 7888 3977
rect 7854 3943 7888 3969
rect 10558 4885 10592 4911
rect 10558 4877 10592 4885
rect 10558 4817 10592 4839
rect 10558 4805 10592 4817
rect 10558 4749 10592 4767
rect 10558 4733 10592 4749
rect 10558 4681 10592 4695
rect 10558 4661 10592 4681
rect 10558 4613 10592 4623
rect 10558 4589 10592 4613
rect 10558 4545 10592 4551
rect 10558 4517 10592 4545
rect 10558 4477 10592 4479
rect 10558 4445 10592 4477
rect 10558 4375 10592 4407
rect 10558 4373 10592 4375
rect 10558 4307 10592 4335
rect 10558 4301 10592 4307
rect 10558 4239 10592 4263
rect 10558 4229 10592 4239
rect 10558 4171 10592 4191
rect 10558 4157 10592 4171
rect 10558 4103 10592 4119
rect 10558 4085 10592 4103
rect 10558 4035 10592 4047
rect 10558 4013 10592 4035
rect 10558 3967 10592 3975
rect 10558 3941 10592 3967
rect 10654 4885 10688 4911
rect 10654 4877 10688 4885
rect 10654 4817 10688 4839
rect 10654 4805 10688 4817
rect 10654 4749 10688 4767
rect 10654 4733 10688 4749
rect 10654 4681 10688 4695
rect 10654 4661 10688 4681
rect 10654 4613 10688 4623
rect 10654 4589 10688 4613
rect 10654 4545 10688 4551
rect 10654 4517 10688 4545
rect 10654 4477 10688 4479
rect 10654 4445 10688 4477
rect 10654 4375 10688 4407
rect 10654 4373 10688 4375
rect 10654 4307 10688 4335
rect 10654 4301 10688 4307
rect 10654 4239 10688 4263
rect 10654 4229 10688 4239
rect 10654 4171 10688 4191
rect 10654 4157 10688 4171
rect 10654 4103 10688 4119
rect 10654 4085 10688 4103
rect 10654 4035 10688 4047
rect 10654 4013 10688 4035
rect 10654 3967 10688 3975
rect 10654 3941 10688 3967
rect 10750 4885 10784 4911
rect 10750 4877 10784 4885
rect 10750 4817 10784 4839
rect 10750 4805 10784 4817
rect 10750 4749 10784 4767
rect 10750 4733 10784 4749
rect 10750 4681 10784 4695
rect 10750 4661 10784 4681
rect 10750 4613 10784 4623
rect 10750 4589 10784 4613
rect 10750 4545 10784 4551
rect 10750 4517 10784 4545
rect 10750 4477 10784 4479
rect 10750 4445 10784 4477
rect 10750 4375 10784 4407
rect 10750 4373 10784 4375
rect 10750 4307 10784 4335
rect 10750 4301 10784 4307
rect 10750 4239 10784 4263
rect 10750 4229 10784 4239
rect 10750 4171 10784 4191
rect 10750 4157 10784 4171
rect 10750 4103 10784 4119
rect 10750 4085 10784 4103
rect 10750 4035 10784 4047
rect 10750 4013 10784 4035
rect 10750 3967 10784 3975
rect 10750 3941 10784 3967
rect 10846 4885 10880 4911
rect 10846 4877 10880 4885
rect 10846 4817 10880 4839
rect 10846 4805 10880 4817
rect 10846 4749 10880 4767
rect 10846 4733 10880 4749
rect 10846 4681 10880 4695
rect 10846 4661 10880 4681
rect 10846 4613 10880 4623
rect 10846 4589 10880 4613
rect 10846 4545 10880 4551
rect 10846 4517 10880 4545
rect 10846 4477 10880 4479
rect 10846 4445 10880 4477
rect 10846 4375 10880 4407
rect 10846 4373 10880 4375
rect 10846 4307 10880 4335
rect 10846 4301 10880 4307
rect 10846 4239 10880 4263
rect 10846 4229 10880 4239
rect 10846 4171 10880 4191
rect 10846 4157 10880 4171
rect 10846 4103 10880 4119
rect 10846 4085 10880 4103
rect 10846 4035 10880 4047
rect 10846 4013 10880 4035
rect 10846 3967 10880 3975
rect 10846 3941 10880 3967
rect 15518 4981 15552 5011
rect 10942 4885 10976 4911
rect 10942 4877 10976 4885
rect 10942 4817 10976 4839
rect 10942 4805 10976 4817
rect 10942 4749 10976 4767
rect 10942 4733 10976 4749
rect 10942 4681 10976 4695
rect 10942 4661 10976 4681
rect 10942 4613 10976 4623
rect 10942 4589 10976 4613
rect 10942 4545 10976 4551
rect 10942 4517 10976 4545
rect 10942 4477 10976 4479
rect 10942 4445 10976 4477
rect 10942 4375 10976 4407
rect 10942 4373 10976 4375
rect 10942 4307 10976 4335
rect 10942 4301 10976 4307
rect 10942 4239 10976 4263
rect 10942 4229 10976 4239
rect 10942 4171 10976 4191
rect 10942 4157 10976 4171
rect 10942 4103 10976 4119
rect 10942 4085 10976 4103
rect 10942 4035 10976 4047
rect 10942 4013 10976 4035
rect 10942 3967 10976 3975
rect 10942 3941 10976 3967
rect 13714 4859 13748 4885
rect 13714 4851 13748 4859
rect 13714 4791 13748 4813
rect 13714 4779 13748 4791
rect 13714 4723 13748 4741
rect 13714 4707 13748 4723
rect 13714 4655 13748 4669
rect 13714 4635 13748 4655
rect 13714 4587 13748 4597
rect 13714 4563 13748 4587
rect 13714 4519 13748 4525
rect 13714 4491 13748 4519
rect 13714 4451 13748 4453
rect 13714 4419 13748 4451
rect 13714 4349 13748 4381
rect 13714 4347 13748 4349
rect 13714 4281 13748 4309
rect 13714 4275 13748 4281
rect 13714 4213 13748 4237
rect 13714 4203 13748 4213
rect 13714 4145 13748 4165
rect 13714 4131 13748 4145
rect 13714 4077 13748 4093
rect 13714 4059 13748 4077
rect 13714 4009 13748 4021
rect 13714 3987 13748 4009
rect 13714 3941 13748 3949
rect 13714 3915 13748 3941
rect 13810 4859 13844 4885
rect 13810 4851 13844 4859
rect 13810 4791 13844 4813
rect 13810 4779 13844 4791
rect 13810 4723 13844 4741
rect 13810 4707 13844 4723
rect 13810 4655 13844 4669
rect 13810 4635 13844 4655
rect 13810 4587 13844 4597
rect 13810 4563 13844 4587
rect 13810 4519 13844 4525
rect 13810 4491 13844 4519
rect 13810 4451 13844 4453
rect 13810 4419 13844 4451
rect 13810 4349 13844 4381
rect 13810 4347 13844 4349
rect 13810 4281 13844 4309
rect 13810 4275 13844 4281
rect 13810 4213 13844 4237
rect 13810 4203 13844 4213
rect 13810 4145 13844 4165
rect 13810 4131 13844 4145
rect 13810 4077 13844 4093
rect 13810 4059 13844 4077
rect 13810 4009 13844 4021
rect 13810 3987 13844 4009
rect 13810 3941 13844 3949
rect 13810 3915 13844 3941
rect 1676 3720 1710 3754
rect 1772 3743 1806 3777
rect 4536 3727 4570 3761
rect 4632 3704 4666 3738
rect 4728 3727 4762 3761
rect 7566 3727 7600 3761
rect 13906 4859 13940 4885
rect 13906 4851 13940 4859
rect 13906 4791 13940 4813
rect 13906 4779 13940 4791
rect 13906 4723 13940 4741
rect 13906 4707 13940 4723
rect 13906 4655 13940 4669
rect 13906 4635 13940 4655
rect 13906 4587 13940 4597
rect 13906 4563 13940 4587
rect 13906 4519 13940 4525
rect 13906 4491 13940 4519
rect 13906 4451 13940 4453
rect 13906 4419 13940 4451
rect 13906 4349 13940 4381
rect 13906 4347 13940 4349
rect 13906 4281 13940 4309
rect 13906 4275 13940 4281
rect 13906 4213 13940 4237
rect 13906 4203 13940 4213
rect 13906 4145 13940 4165
rect 13906 4131 13940 4145
rect 13906 4077 13940 4093
rect 13906 4059 13940 4077
rect 13906 4009 13940 4021
rect 13906 3987 13940 4009
rect 13906 3941 13940 3949
rect 13906 3915 13940 3941
rect 14002 4859 14036 4885
rect 14002 4851 14036 4859
rect 14002 4791 14036 4813
rect 14002 4779 14036 4791
rect 14002 4723 14036 4741
rect 14002 4707 14036 4723
rect 14002 4655 14036 4669
rect 14002 4635 14036 4655
rect 14002 4587 14036 4597
rect 14002 4563 14036 4587
rect 14002 4519 14036 4525
rect 14002 4491 14036 4519
rect 14002 4451 14036 4453
rect 14002 4419 14036 4451
rect 14002 4349 14036 4381
rect 14002 4347 14036 4349
rect 14002 4281 14036 4309
rect 14002 4275 14036 4281
rect 14002 4213 14036 4237
rect 14002 4203 14036 4213
rect 14002 4145 14036 4165
rect 14002 4131 14036 4145
rect 14002 4077 14036 4093
rect 14002 4059 14036 4077
rect 14002 4009 14036 4021
rect 14002 3987 14036 4009
rect 14002 3941 14036 3949
rect 14002 3915 14036 3941
rect 14098 4859 14132 4885
rect 14098 4851 14132 4859
rect 14098 4791 14132 4813
rect 14098 4779 14132 4791
rect 14098 4723 14132 4741
rect 14098 4707 14132 4723
rect 14098 4655 14132 4669
rect 14098 4635 14132 4655
rect 14098 4587 14132 4597
rect 14098 4563 14132 4587
rect 14098 4519 14132 4525
rect 14098 4491 14132 4519
rect 14098 4451 14132 4453
rect 14098 4419 14132 4451
rect 14098 4349 14132 4381
rect 14098 4347 14132 4349
rect 14098 4281 14132 4309
rect 14098 4275 14132 4281
rect 14098 4213 14132 4237
rect 14098 4203 14132 4213
rect 14098 4145 14132 4165
rect 14098 4131 14132 4145
rect 14098 4077 14132 4093
rect 14098 4059 14132 4077
rect 14098 4009 14132 4021
rect 14098 3987 14132 4009
rect 14098 3941 14132 3949
rect 14098 3915 14132 3941
rect 15518 4909 15552 4943
rect 15518 4841 15552 4871
rect 15518 4837 15552 4841
rect 15518 4773 15552 4799
rect 15518 4765 15552 4773
rect 15518 4705 15552 4727
rect 15518 4693 15552 4705
rect 15518 4637 15552 4655
rect 15518 4621 15552 4637
rect 15518 4569 15552 4583
rect 15518 4549 15552 4569
rect 15518 4501 15552 4511
rect 15518 4477 15552 4501
rect 15518 4433 15552 4439
rect 15518 4405 15552 4433
rect 15518 4365 15552 4367
rect 15518 4333 15552 4365
rect 15518 4263 15552 4295
rect 15518 4261 15552 4263
rect 15518 4195 15552 4223
rect 15518 4189 15552 4195
rect 15518 4127 15552 4151
rect 15518 4117 15552 4127
rect 15518 4059 15552 4079
rect 15518 4045 15552 4059
rect 15518 3991 15552 4007
rect 15518 3973 15552 3991
rect 15614 5861 15648 5879
rect 15614 5845 15648 5861
rect 15614 5793 15648 5807
rect 15614 5773 15648 5793
rect 15614 5725 15648 5735
rect 15614 5701 15648 5725
rect 15614 5657 15648 5663
rect 15614 5629 15648 5657
rect 15614 5589 15648 5591
rect 15614 5557 15648 5589
rect 15614 5487 15648 5519
rect 15614 5485 15648 5487
rect 15614 5419 15648 5447
rect 15614 5413 15648 5419
rect 15614 5351 15648 5375
rect 15614 5341 15648 5351
rect 15614 5283 15648 5303
rect 15614 5269 15648 5283
rect 15614 5215 15648 5231
rect 15614 5197 15648 5215
rect 15614 5147 15648 5159
rect 15614 5125 15648 5147
rect 15614 5079 15648 5087
rect 15614 5053 15648 5079
rect 15614 5011 15648 5015
rect 15614 4981 15648 5011
rect 15614 4909 15648 4943
rect 15614 4841 15648 4871
rect 15614 4837 15648 4841
rect 15614 4773 15648 4799
rect 15614 4765 15648 4773
rect 15614 4705 15648 4727
rect 15614 4693 15648 4705
rect 15614 4637 15648 4655
rect 15614 4621 15648 4637
rect 15614 4569 15648 4583
rect 15614 4549 15648 4569
rect 15614 4501 15648 4511
rect 15614 4477 15648 4501
rect 15614 4433 15648 4439
rect 15614 4405 15648 4433
rect 15614 4365 15648 4367
rect 15614 4333 15648 4365
rect 15614 4263 15648 4295
rect 15614 4261 15648 4263
rect 15614 4195 15648 4223
rect 15614 4189 15648 4195
rect 15614 4127 15648 4151
rect 15614 4117 15648 4127
rect 15614 4059 15648 4079
rect 15614 4045 15648 4059
rect 15614 3991 15648 4007
rect 15614 3973 15648 3991
rect 15710 5861 15744 5879
rect 15710 5845 15744 5861
rect 15710 5793 15744 5807
rect 15710 5773 15744 5793
rect 15710 5725 15744 5735
rect 15710 5701 15744 5725
rect 15710 5657 15744 5663
rect 15710 5629 15744 5657
rect 15710 5589 15744 5591
rect 15710 5557 15744 5589
rect 15710 5487 15744 5519
rect 15710 5485 15744 5487
rect 15710 5419 15744 5447
rect 15710 5413 15744 5419
rect 15710 5351 15744 5375
rect 15710 5341 15744 5351
rect 15710 5283 15744 5303
rect 15710 5269 15744 5283
rect 15710 5215 15744 5231
rect 15710 5197 15744 5215
rect 15710 5147 15744 5159
rect 15710 5125 15744 5147
rect 15710 5079 15744 5087
rect 15710 5053 15744 5079
rect 15710 5011 15744 5015
rect 15710 4981 15744 5011
rect 15710 4909 15744 4943
rect 15710 4841 15744 4871
rect 15710 4837 15744 4841
rect 15710 4773 15744 4799
rect 15710 4765 15744 4773
rect 15710 4705 15744 4727
rect 15710 4693 15744 4705
rect 15710 4637 15744 4655
rect 15710 4621 15744 4637
rect 15710 4569 15744 4583
rect 15710 4549 15744 4569
rect 15710 4501 15744 4511
rect 15710 4477 15744 4501
rect 15710 4433 15744 4439
rect 15710 4405 15744 4433
rect 15710 4365 15744 4367
rect 15710 4333 15744 4365
rect 15710 4263 15744 4295
rect 15710 4261 15744 4263
rect 15710 4195 15744 4223
rect 15710 4189 15744 4195
rect 15710 4127 15744 4151
rect 15710 4117 15744 4127
rect 15710 4059 15744 4079
rect 15710 4045 15744 4059
rect 15710 3991 15744 4007
rect 15710 3973 15744 3991
rect 7662 3704 7696 3738
rect 7758 3727 7792 3761
rect 10654 3725 10688 3759
rect 10750 3702 10784 3736
rect 10846 3725 10880 3759
rect 13810 3699 13844 3733
rect 15566 3745 15600 3779
rect 13906 3676 13940 3710
rect 14002 3699 14036 3733
rect 15710 3726 15744 3760
rect -1590 3394 -1556 3428
rect -1110 3290 -1076 3324
rect -1686 3195 -1652 3221
rect -1686 3187 -1652 3195
rect -1686 3127 -1652 3149
rect -1686 3115 -1652 3127
rect -1686 3059 -1652 3077
rect -1686 3043 -1652 3059
rect -1686 2991 -1652 3005
rect -1686 2971 -1652 2991
rect -1686 2923 -1652 2933
rect -1686 2899 -1652 2923
rect -1686 2855 -1652 2861
rect -1686 2827 -1652 2855
rect -1686 2787 -1652 2789
rect -1686 2755 -1652 2787
rect -1686 2685 -1652 2717
rect -1686 2683 -1652 2685
rect -1686 2617 -1652 2645
rect -1686 2611 -1652 2617
rect -1686 2549 -1652 2573
rect -1686 2539 -1652 2549
rect -1686 2481 -1652 2501
rect -1686 2467 -1652 2481
rect -1686 2413 -1652 2429
rect -1686 2395 -1652 2413
rect -1686 2345 -1652 2357
rect -1686 2323 -1652 2345
rect -1686 2277 -1652 2285
rect -1686 2251 -1652 2277
rect -1590 3195 -1556 3221
rect -1590 3187 -1556 3195
rect -1590 3127 -1556 3149
rect -1590 3115 -1556 3127
rect -1590 3059 -1556 3077
rect -1590 3043 -1556 3059
rect -1590 2991 -1556 3005
rect -1590 2971 -1556 2991
rect -1590 2923 -1556 2933
rect -1590 2899 -1556 2923
rect -1590 2855 -1556 2861
rect -1590 2827 -1556 2855
rect -1590 2787 -1556 2789
rect -1590 2755 -1556 2787
rect -1590 2685 -1556 2717
rect -1590 2683 -1556 2685
rect -1590 2617 -1556 2645
rect -1590 2611 -1556 2617
rect -1590 2549 -1556 2573
rect -1590 2539 -1556 2549
rect -1590 2481 -1556 2501
rect -1590 2467 -1556 2481
rect -1590 2413 -1556 2429
rect -1590 2395 -1556 2413
rect -1590 2345 -1556 2357
rect -1590 2323 -1556 2345
rect -1590 2277 -1556 2285
rect -1590 2251 -1556 2277
rect -1494 3195 -1460 3221
rect -1494 3187 -1460 3195
rect -1494 3127 -1460 3149
rect -1494 3115 -1460 3127
rect -1494 3059 -1460 3077
rect -1494 3043 -1460 3059
rect -1494 2991 -1460 3005
rect -1494 2971 -1460 2991
rect -1494 2923 -1460 2933
rect -1494 2899 -1460 2923
rect -1494 2855 -1460 2861
rect -1494 2827 -1460 2855
rect -1494 2787 -1460 2789
rect -1494 2755 -1460 2787
rect -1494 2685 -1460 2717
rect -1494 2683 -1460 2685
rect -1494 2617 -1460 2645
rect -1494 2611 -1460 2617
rect -1494 2549 -1460 2573
rect -1494 2539 -1460 2549
rect -1494 2481 -1460 2501
rect -1494 2467 -1460 2481
rect -1494 2413 -1460 2429
rect -1494 2395 -1460 2413
rect -1494 2345 -1460 2357
rect -1494 2323 -1460 2345
rect -1494 2277 -1460 2285
rect -1494 2251 -1460 2277
rect -1398 3195 -1364 3221
rect -1398 3187 -1364 3195
rect -1398 3127 -1364 3149
rect -1398 3115 -1364 3127
rect -1398 3059 -1364 3077
rect -1398 3043 -1364 3059
rect -1398 2991 -1364 3005
rect -1398 2971 -1364 2991
rect -1398 2923 -1364 2933
rect -1398 2899 -1364 2923
rect -1398 2855 -1364 2861
rect -1398 2827 -1364 2855
rect -1398 2787 -1364 2789
rect -1398 2755 -1364 2787
rect -1398 2685 -1364 2717
rect -1398 2683 -1364 2685
rect -1398 2617 -1364 2645
rect -1398 2611 -1364 2617
rect -1398 2549 -1364 2573
rect -1398 2539 -1364 2549
rect -1398 2481 -1364 2501
rect -1398 2467 -1364 2481
rect -1398 2413 -1364 2429
rect -1398 2395 -1364 2413
rect -1398 2345 -1364 2357
rect -1398 2323 -1364 2345
rect -1398 2277 -1364 2285
rect -1398 2251 -1364 2277
rect -1302 3195 -1268 3221
rect -1302 3187 -1268 3195
rect -1302 3127 -1268 3149
rect -1302 3115 -1268 3127
rect -1302 3059 -1268 3077
rect -1302 3043 -1268 3059
rect -1302 2991 -1268 3005
rect -1302 2971 -1268 2991
rect -1302 2923 -1268 2933
rect -1302 2899 -1268 2923
rect -1302 2855 -1268 2861
rect -1302 2827 -1268 2855
rect -1302 2787 -1268 2789
rect -1302 2755 -1268 2787
rect -1302 2685 -1268 2717
rect -1302 2683 -1268 2685
rect -1302 2617 -1268 2645
rect -1302 2611 -1268 2617
rect -1302 2549 -1268 2573
rect -1302 2539 -1268 2549
rect -1302 2481 -1268 2501
rect -1302 2467 -1268 2481
rect -1302 2413 -1268 2429
rect -1302 2395 -1268 2413
rect -1302 2345 -1268 2357
rect -1302 2323 -1268 2345
rect -1302 2277 -1268 2285
rect -1302 2251 -1268 2277
rect -1206 3195 -1172 3221
rect -1206 3187 -1172 3195
rect -1206 3127 -1172 3149
rect -1206 3115 -1172 3127
rect -1206 3059 -1172 3077
rect -1206 3043 -1172 3059
rect -1206 2991 -1172 3005
rect -1206 2971 -1172 2991
rect -1206 2923 -1172 2933
rect -1206 2899 -1172 2923
rect -1206 2855 -1172 2861
rect -1206 2827 -1172 2855
rect -1206 2787 -1172 2789
rect -1206 2755 -1172 2787
rect -1206 2685 -1172 2717
rect -1206 2683 -1172 2685
rect -1206 2617 -1172 2645
rect -1206 2611 -1172 2617
rect -1206 2549 -1172 2573
rect -1206 2539 -1172 2549
rect -1206 2481 -1172 2501
rect -1206 2467 -1172 2481
rect -1206 2413 -1172 2429
rect -1206 2395 -1172 2413
rect -1206 2345 -1172 2357
rect -1206 2323 -1172 2345
rect -1206 2277 -1172 2285
rect -1206 2251 -1172 2277
rect -1110 3195 -1076 3221
rect -1110 3187 -1076 3195
rect -1110 3127 -1076 3149
rect -1110 3115 -1076 3127
rect -1110 3059 -1076 3077
rect -1110 3043 -1076 3059
rect -1110 2991 -1076 3005
rect -1110 2971 -1076 2991
rect -1110 2923 -1076 2933
rect -1110 2899 -1076 2923
rect -1110 2855 -1076 2861
rect -1110 2827 -1076 2855
rect -1110 2787 -1076 2789
rect -1110 2755 -1076 2787
rect -1110 2685 -1076 2717
rect -1110 2683 -1076 2685
rect -1110 2617 -1076 2645
rect -1110 2611 -1076 2617
rect -1110 2549 -1076 2573
rect -1110 2539 -1076 2549
rect -1110 2481 -1076 2501
rect -1110 2467 -1076 2481
rect -1110 2413 -1076 2429
rect -1110 2395 -1076 2413
rect -1110 2345 -1076 2357
rect -1110 2323 -1076 2345
rect -1110 2277 -1076 2285
rect -1110 2251 -1076 2277
rect -1014 3195 -980 3221
rect -1014 3187 -980 3195
rect -1014 3127 -980 3149
rect -1014 3115 -980 3127
rect -1014 3059 -980 3077
rect -1014 3043 -980 3059
rect -1014 2991 -980 3005
rect -1014 2971 -980 2991
rect -1014 2923 -980 2933
rect -1014 2899 -980 2923
rect -1014 2855 -980 2861
rect -1014 2827 -980 2855
rect -1014 2787 -980 2789
rect -1014 2755 -980 2787
rect -1014 2685 -980 2717
rect -1014 2683 -980 2685
rect -1014 2617 -980 2645
rect -1014 2611 -980 2617
rect -1014 2549 -980 2573
rect -1014 2539 -980 2549
rect -1014 2481 -980 2501
rect -1014 2467 -980 2481
rect -1014 2413 -980 2429
rect -1014 2395 -980 2413
rect -1014 2345 -980 2357
rect -1014 2323 -980 2345
rect -1014 2277 -980 2285
rect -1014 2251 -980 2277
rect -918 3195 -884 3221
rect -918 3187 -884 3195
rect -918 3127 -884 3149
rect -918 3115 -884 3127
rect -918 3059 -884 3077
rect -918 3043 -884 3059
rect -918 2991 -884 3005
rect -918 2971 -884 2991
rect 1578 2968 1612 3002
rect -918 2923 -884 2933
rect -918 2899 -884 2923
rect 1674 2960 1708 2994
rect 4534 2952 4568 2986
rect 4630 2944 4664 2978
rect 7564 2952 7598 2986
rect -918 2855 -884 2861
rect -918 2827 -884 2855
rect 7660 2944 7694 2978
rect 10652 2950 10686 2984
rect 10748 2942 10782 2976
rect -918 2787 -884 2789
rect -918 2755 -884 2787
rect -918 2685 -884 2717
rect -918 2683 -884 2685
rect -918 2617 -884 2645
rect -918 2611 -884 2617
rect -918 2549 -884 2573
rect -918 2539 -884 2549
rect -918 2481 -884 2501
rect -918 2467 -884 2481
rect -918 2413 -884 2429
rect -918 2395 -884 2413
rect -918 2345 -884 2357
rect -918 2323 -884 2345
rect -918 2277 -884 2285
rect -918 2251 -884 2277
rect -1097 2138 -1063 2172
rect 1482 2789 1516 2815
rect 1482 2781 1516 2789
rect 1482 2721 1516 2743
rect 1482 2709 1516 2721
rect 1482 2653 1516 2671
rect 1482 2637 1516 2653
rect 1482 2585 1516 2599
rect 1482 2565 1516 2585
rect 1482 2517 1516 2527
rect 1482 2493 1516 2517
rect 1482 2449 1516 2455
rect 1482 2421 1516 2449
rect 1482 2381 1516 2383
rect 1482 2349 1516 2381
rect 1482 2279 1516 2311
rect 1482 2277 1516 2279
rect 1482 2211 1516 2239
rect 1482 2205 1516 2211
rect 1482 2143 1516 2167
rect 1482 2133 1516 2143
rect 1482 2075 1516 2095
rect 1482 2061 1516 2075
rect 1482 2007 1516 2023
rect 1482 1989 1516 2007
rect 1482 1939 1516 1951
rect 1482 1917 1516 1939
rect 1482 1871 1516 1879
rect 1482 1845 1516 1871
rect 1578 2789 1612 2815
rect 1578 2781 1612 2789
rect 1578 2721 1612 2743
rect 1578 2709 1612 2721
rect 1578 2653 1612 2671
rect 1578 2637 1612 2653
rect 1578 2585 1612 2599
rect 1578 2565 1612 2585
rect 1578 2517 1612 2527
rect 1578 2493 1612 2517
rect 1578 2449 1612 2455
rect 1578 2421 1612 2449
rect 1578 2381 1612 2383
rect 1578 2349 1612 2381
rect 1578 2279 1612 2311
rect 1578 2277 1612 2279
rect 1578 2211 1612 2239
rect 1578 2205 1612 2211
rect 1578 2143 1612 2167
rect 1578 2133 1612 2143
rect 1578 2075 1612 2095
rect 1578 2061 1612 2075
rect 1578 2007 1612 2023
rect 1578 1989 1612 2007
rect 1578 1939 1612 1951
rect 1578 1917 1612 1939
rect 1578 1871 1612 1879
rect 1578 1845 1612 1871
rect 1674 2789 1708 2815
rect 1674 2781 1708 2789
rect 1674 2721 1708 2743
rect 1674 2709 1708 2721
rect 1674 2653 1708 2671
rect 1674 2637 1708 2653
rect 1674 2585 1708 2599
rect 1674 2565 1708 2585
rect 1674 2517 1708 2527
rect 1674 2493 1708 2517
rect 1674 2449 1708 2455
rect 1674 2421 1708 2449
rect 1674 2381 1708 2383
rect 1674 2349 1708 2381
rect 1674 2279 1708 2311
rect 1674 2277 1708 2279
rect 1674 2211 1708 2239
rect 1674 2205 1708 2211
rect 1674 2143 1708 2167
rect 1674 2133 1708 2143
rect 1674 2075 1708 2095
rect 1674 2061 1708 2075
rect 1674 2007 1708 2023
rect 1674 1989 1708 2007
rect 1674 1939 1708 1951
rect 1674 1917 1708 1939
rect 1674 1871 1708 1879
rect 1674 1845 1708 1871
rect 1770 2789 1804 2815
rect 1770 2781 1804 2789
rect 1770 2721 1804 2743
rect 1770 2709 1804 2721
rect 1770 2653 1804 2671
rect 1770 2637 1804 2653
rect 1770 2585 1804 2599
rect 1770 2565 1804 2585
rect 1770 2517 1804 2527
rect 1770 2493 1804 2517
rect 1770 2449 1804 2455
rect 1770 2421 1804 2449
rect 1770 2381 1804 2383
rect 1770 2349 1804 2381
rect 1770 2279 1804 2311
rect 1770 2277 1804 2279
rect 1770 2211 1804 2239
rect 1770 2205 1804 2211
rect 1770 2143 1804 2167
rect 1770 2133 1804 2143
rect 1770 2075 1804 2095
rect 1770 2061 1804 2075
rect 1770 2007 1804 2023
rect 1770 1989 1804 2007
rect 1770 1939 1804 1951
rect 1770 1917 1804 1939
rect 1770 1871 1804 1879
rect 1770 1845 1804 1871
rect 1866 2789 1900 2815
rect 1866 2781 1900 2789
rect 1866 2721 1900 2743
rect 1866 2709 1900 2721
rect 1866 2653 1900 2671
rect 1866 2637 1900 2653
rect 1866 2585 1900 2599
rect 1866 2565 1900 2585
rect 1866 2517 1900 2527
rect 1866 2493 1900 2517
rect 1866 2449 1900 2455
rect 1866 2421 1900 2449
rect 4438 2773 4472 2799
rect 4438 2765 4472 2773
rect 4438 2705 4472 2727
rect 4438 2693 4472 2705
rect 4438 2637 4472 2655
rect 4438 2621 4472 2637
rect 4438 2569 4472 2583
rect 4438 2549 4472 2569
rect 4438 2501 4472 2511
rect 4438 2477 4472 2501
rect 4438 2433 4472 2439
rect 2579 2394 2613 2428
rect 4438 2405 4472 2433
rect 1866 2381 1900 2383
rect 1866 2349 1900 2381
rect 4438 2365 4472 2367
rect 2392 2316 2426 2350
rect 1866 2279 1900 2311
rect 1866 2277 1900 2279
rect 1866 2211 1900 2239
rect 1866 2205 1900 2211
rect 1866 2143 1900 2167
rect 1866 2133 1900 2143
rect 1866 2075 1900 2095
rect 1866 2061 1900 2075
rect 1866 2007 1900 2023
rect 1866 1989 1900 2007
rect 1866 1939 1900 1951
rect 1866 1917 1900 1939
rect 2500 2227 2534 2229
rect 2500 2195 2534 2227
rect 2500 2125 2534 2157
rect 2500 2123 2534 2125
rect 2658 2227 2692 2229
rect 2658 2195 2692 2227
rect 2658 2125 2692 2157
rect 2658 2123 2692 2125
rect 4438 2333 4472 2365
rect 4438 2263 4472 2295
rect 4438 2261 4472 2263
rect 4438 2195 4472 2223
rect 4438 2189 4472 2195
rect 4438 2127 4472 2151
rect 4438 2117 4472 2127
rect 1866 1871 1900 1879
rect 1866 1845 1900 1871
rect 4438 2059 4472 2079
rect 4438 2045 4472 2059
rect 4438 1991 4472 2007
rect 4438 1973 4472 1991
rect 4438 1923 4472 1935
rect 4438 1901 4472 1923
rect 1578 1662 1612 1696
rect 4438 1855 4472 1863
rect 4438 1829 4472 1855
rect 4534 2773 4568 2799
rect 4534 2765 4568 2773
rect 4534 2705 4568 2727
rect 4534 2693 4568 2705
rect 4534 2637 4568 2655
rect 4534 2621 4568 2637
rect 4534 2569 4568 2583
rect 4534 2549 4568 2569
rect 4534 2501 4568 2511
rect 4534 2477 4568 2501
rect 4534 2433 4568 2439
rect 4534 2405 4568 2433
rect 4534 2365 4568 2367
rect 4534 2333 4568 2365
rect 4534 2263 4568 2295
rect 4534 2261 4568 2263
rect 4534 2195 4568 2223
rect 4534 2189 4568 2195
rect 4534 2127 4568 2151
rect 4534 2117 4568 2127
rect 4534 2059 4568 2079
rect 4534 2045 4568 2059
rect 4534 1991 4568 2007
rect 4534 1973 4568 1991
rect 4534 1923 4568 1935
rect 4534 1901 4568 1923
rect 4534 1855 4568 1863
rect 4534 1829 4568 1855
rect 4630 2773 4664 2799
rect 4630 2765 4664 2773
rect 4630 2705 4664 2727
rect 4630 2693 4664 2705
rect 4630 2637 4664 2655
rect 4630 2621 4664 2637
rect 4630 2569 4664 2583
rect 4630 2549 4664 2569
rect 4630 2501 4664 2511
rect 4630 2477 4664 2501
rect 4630 2433 4664 2439
rect 4630 2405 4664 2433
rect 4630 2365 4664 2367
rect 4630 2333 4664 2365
rect 4630 2263 4664 2295
rect 4630 2261 4664 2263
rect 4630 2195 4664 2223
rect 4630 2189 4664 2195
rect 4630 2127 4664 2151
rect 4630 2117 4664 2127
rect 4630 2059 4664 2079
rect 4630 2045 4664 2059
rect 4630 1991 4664 2007
rect 4630 1973 4664 1991
rect 4630 1923 4664 1935
rect 4630 1901 4664 1923
rect 4630 1855 4664 1863
rect 4630 1829 4664 1855
rect 13808 2924 13842 2958
rect 13904 2916 13938 2950
rect 4726 2773 4760 2799
rect 4726 2765 4760 2773
rect 4726 2705 4760 2727
rect 4726 2693 4760 2705
rect 4726 2637 4760 2655
rect 4726 2621 4760 2637
rect 4726 2569 4760 2583
rect 4726 2549 4760 2569
rect 4726 2501 4760 2511
rect 4726 2477 4760 2501
rect 4726 2433 4760 2439
rect 4726 2405 4760 2433
rect 4726 2365 4760 2367
rect 4726 2333 4760 2365
rect 4726 2263 4760 2295
rect 4726 2261 4760 2263
rect 4726 2195 4760 2223
rect 4726 2189 4760 2195
rect 4726 2127 4760 2151
rect 4726 2117 4760 2127
rect 4726 2059 4760 2079
rect 4726 2045 4760 2059
rect 4726 1991 4760 2007
rect 4726 1973 4760 1991
rect 4726 1923 4760 1935
rect 4726 1901 4760 1923
rect 4726 1855 4760 1863
rect 4726 1829 4760 1855
rect 4822 2773 4856 2799
rect 4822 2765 4856 2773
rect 4822 2705 4856 2727
rect 4822 2693 4856 2705
rect 4822 2637 4856 2655
rect 4822 2621 4856 2637
rect 4822 2569 4856 2583
rect 4822 2549 4856 2569
rect 4822 2501 4856 2511
rect 4822 2477 4856 2501
rect 4822 2433 4856 2439
rect 4822 2405 4856 2433
rect 7468 2773 7502 2799
rect 7468 2765 7502 2773
rect 7468 2705 7502 2727
rect 7468 2693 7502 2705
rect 7468 2637 7502 2655
rect 7468 2621 7502 2637
rect 7468 2569 7502 2583
rect 7468 2549 7502 2569
rect 7468 2501 7502 2511
rect 7468 2477 7502 2501
rect 7468 2433 7502 2439
rect 5579 2394 5613 2428
rect 7468 2405 7502 2433
rect 4822 2365 4856 2367
rect 4822 2333 4856 2365
rect 7468 2365 7502 2367
rect 5392 2316 5426 2350
rect 4822 2263 4856 2295
rect 4822 2261 4856 2263
rect 4822 2195 4856 2223
rect 4822 2189 4856 2195
rect 4822 2127 4856 2151
rect 4822 2117 4856 2127
rect 4822 2059 4856 2079
rect 4822 2045 4856 2059
rect 4822 1991 4856 2007
rect 4822 1973 4856 1991
rect 4822 1923 4856 1935
rect 4822 1901 4856 1923
rect 4822 1855 4856 1863
rect 4822 1829 4856 1855
rect 5500 2227 5534 2229
rect 5500 2195 5534 2227
rect 5500 2125 5534 2157
rect 5500 2123 5534 2125
rect 5658 2227 5692 2229
rect 5658 2195 5692 2227
rect 5658 2125 5692 2157
rect 5658 2123 5692 2125
rect 7468 2333 7502 2365
rect 7468 2263 7502 2295
rect 7468 2261 7502 2263
rect 7468 2195 7502 2223
rect 7468 2189 7502 2195
rect 7468 2127 7502 2151
rect 7468 2117 7502 2127
rect 7468 2059 7502 2079
rect 7468 2045 7502 2059
rect 7468 1991 7502 2007
rect 7468 1973 7502 1991
rect 7468 1923 7502 1935
rect 7468 1901 7502 1923
rect 7468 1855 7502 1863
rect 7468 1829 7502 1855
rect 7564 2773 7598 2799
rect 7564 2765 7598 2773
rect 7564 2705 7598 2727
rect 7564 2693 7598 2705
rect 7564 2637 7598 2655
rect 7564 2621 7598 2637
rect 7564 2569 7598 2583
rect 7564 2549 7598 2569
rect 7564 2501 7598 2511
rect 7564 2477 7598 2501
rect 7564 2433 7598 2439
rect 7564 2405 7598 2433
rect 7564 2365 7598 2367
rect 7564 2333 7598 2365
rect 7564 2263 7598 2295
rect 7564 2261 7598 2263
rect 7564 2195 7598 2223
rect 7564 2189 7598 2195
rect 7564 2127 7598 2151
rect 7564 2117 7598 2127
rect 7564 2059 7598 2079
rect 7564 2045 7598 2059
rect 7564 1991 7598 2007
rect 7564 1973 7598 1991
rect 7564 1923 7598 1935
rect 7564 1901 7598 1923
rect 7564 1855 7598 1863
rect 7564 1829 7598 1855
rect 7660 2773 7694 2799
rect 7660 2765 7694 2773
rect 7660 2705 7694 2727
rect 7660 2693 7694 2705
rect 7660 2637 7694 2655
rect 7660 2621 7694 2637
rect 7660 2569 7694 2583
rect 7660 2549 7694 2569
rect 7660 2501 7694 2511
rect 7660 2477 7694 2501
rect 7660 2433 7694 2439
rect 7660 2405 7694 2433
rect 7660 2365 7694 2367
rect 7660 2333 7694 2365
rect 7660 2263 7694 2295
rect 7660 2261 7694 2263
rect 7660 2195 7694 2223
rect 7660 2189 7694 2195
rect 7660 2127 7694 2151
rect 7660 2117 7694 2127
rect 7660 2059 7694 2079
rect 7660 2045 7694 2059
rect 7660 1991 7694 2007
rect 7660 1973 7694 1991
rect 7660 1923 7694 1935
rect 7660 1901 7694 1923
rect 7660 1855 7694 1863
rect 7660 1829 7694 1855
rect 7756 2773 7790 2799
rect 7756 2765 7790 2773
rect 7756 2705 7790 2727
rect 7756 2693 7790 2705
rect 7756 2637 7790 2655
rect 7756 2621 7790 2637
rect 7756 2569 7790 2583
rect 7756 2549 7790 2569
rect 7756 2501 7790 2511
rect 7756 2477 7790 2501
rect 7756 2433 7790 2439
rect 7756 2405 7790 2433
rect 7756 2365 7790 2367
rect 7756 2333 7790 2365
rect 7756 2263 7790 2295
rect 7756 2261 7790 2263
rect 7756 2195 7790 2223
rect 7756 2189 7790 2195
rect 7756 2127 7790 2151
rect 7756 2117 7790 2127
rect 7756 2059 7790 2079
rect 7756 2045 7790 2059
rect 7756 1991 7790 2007
rect 7756 1973 7790 1991
rect 7756 1923 7790 1935
rect 7756 1901 7790 1923
rect 7756 1855 7790 1863
rect 7756 1829 7790 1855
rect 7852 2773 7886 2799
rect 7852 2765 7886 2773
rect 7852 2705 7886 2727
rect 7852 2693 7886 2705
rect 7852 2637 7886 2655
rect 7852 2621 7886 2637
rect 7852 2569 7886 2583
rect 7852 2549 7886 2569
rect 7852 2501 7886 2511
rect 7852 2477 7886 2501
rect 7852 2433 7886 2439
rect 7852 2405 7886 2433
rect 10556 2771 10590 2797
rect 10556 2763 10590 2771
rect 10556 2703 10590 2725
rect 10556 2691 10590 2703
rect 10556 2635 10590 2653
rect 10556 2619 10590 2635
rect 10556 2567 10590 2581
rect 10556 2547 10590 2567
rect 10556 2499 10590 2509
rect 10556 2475 10590 2499
rect 10556 2431 10590 2437
rect 8579 2394 8613 2428
rect 10556 2403 10590 2431
rect 7852 2365 7886 2367
rect 7852 2333 7886 2365
rect 10556 2363 10590 2365
rect 8392 2316 8426 2350
rect 7852 2263 7886 2295
rect 7852 2261 7886 2263
rect 7852 2195 7886 2223
rect 7852 2189 7886 2195
rect 7852 2127 7886 2151
rect 7852 2117 7886 2127
rect 7852 2059 7886 2079
rect 7852 2045 7886 2059
rect 7852 1991 7886 2007
rect 7852 1973 7886 1991
rect 7852 1923 7886 1935
rect 7852 1901 7886 1923
rect 7852 1855 7886 1863
rect 7852 1829 7886 1855
rect 8500 2227 8534 2229
rect 8500 2195 8534 2227
rect 8500 2125 8534 2157
rect 8500 2123 8534 2125
rect 8658 2227 8692 2229
rect 8658 2195 8692 2227
rect 8658 2125 8692 2157
rect 8658 2123 8692 2125
rect 10556 2331 10590 2363
rect 10556 2261 10590 2293
rect 10556 2259 10590 2261
rect 10556 2193 10590 2221
rect 10556 2187 10590 2193
rect 10556 2125 10590 2149
rect 10556 2115 10590 2125
rect 4534 1646 4568 1680
rect 10556 2057 10590 2077
rect 10556 2043 10590 2057
rect 10556 1989 10590 2005
rect 10556 1971 10590 1989
rect 10556 1921 10590 1933
rect 10556 1899 10590 1921
rect 10556 1853 10590 1861
rect 10556 1827 10590 1853
rect 7564 1646 7598 1680
rect 10652 2771 10686 2797
rect 10652 2763 10686 2771
rect 10652 2703 10686 2725
rect 10652 2691 10686 2703
rect 10652 2635 10686 2653
rect 10652 2619 10686 2635
rect 10652 2567 10686 2581
rect 10652 2547 10686 2567
rect 10652 2499 10686 2509
rect 10652 2475 10686 2499
rect 10652 2431 10686 2437
rect 10652 2403 10686 2431
rect 10652 2363 10686 2365
rect 10652 2331 10686 2363
rect 10652 2261 10686 2293
rect 10652 2259 10686 2261
rect 10652 2193 10686 2221
rect 10652 2187 10686 2193
rect 10652 2125 10686 2149
rect 10652 2115 10686 2125
rect 10652 2057 10686 2077
rect 10652 2043 10686 2057
rect 10652 1989 10686 2005
rect 10652 1971 10686 1989
rect 10652 1921 10686 1933
rect 10652 1899 10686 1921
rect 10652 1853 10686 1861
rect 10652 1827 10686 1853
rect 10748 2771 10782 2797
rect 10748 2763 10782 2771
rect 10748 2703 10782 2725
rect 10748 2691 10782 2703
rect 10748 2635 10782 2653
rect 10748 2619 10782 2635
rect 10748 2567 10782 2581
rect 10748 2547 10782 2567
rect 10748 2499 10782 2509
rect 10748 2475 10782 2499
rect 10748 2431 10782 2437
rect 10748 2403 10782 2431
rect 10748 2363 10782 2365
rect 10748 2331 10782 2363
rect 10748 2261 10782 2293
rect 10748 2259 10782 2261
rect 10748 2193 10782 2221
rect 10748 2187 10782 2193
rect 10748 2125 10782 2149
rect 10748 2115 10782 2125
rect 10748 2057 10782 2077
rect 10748 2043 10782 2057
rect 10748 1989 10782 2005
rect 10748 1971 10782 1989
rect 10748 1921 10782 1933
rect 10748 1899 10782 1921
rect 10748 1853 10782 1861
rect 10748 1827 10782 1853
rect 10844 2771 10878 2797
rect 10844 2763 10878 2771
rect 10844 2703 10878 2725
rect 10844 2691 10878 2703
rect 10844 2635 10878 2653
rect 10844 2619 10878 2635
rect 10844 2567 10878 2581
rect 10844 2547 10878 2567
rect 10844 2499 10878 2509
rect 10844 2475 10878 2499
rect 10844 2431 10878 2437
rect 10844 2403 10878 2431
rect 10844 2363 10878 2365
rect 10844 2331 10878 2363
rect 10844 2261 10878 2293
rect 10844 2259 10878 2261
rect 10844 2193 10878 2221
rect 10844 2187 10878 2193
rect 10844 2125 10878 2149
rect 10844 2115 10878 2125
rect 10844 2057 10878 2077
rect 10844 2043 10878 2057
rect 10844 1989 10878 2005
rect 10844 1971 10878 1989
rect 10844 1921 10878 1933
rect 10844 1899 10878 1921
rect 10844 1853 10878 1861
rect 10844 1827 10878 1853
rect 10940 2771 10974 2797
rect 10940 2763 10974 2771
rect 10940 2703 10974 2725
rect 10940 2691 10974 2703
rect 10940 2635 10974 2653
rect 10940 2619 10974 2635
rect 10940 2567 10974 2581
rect 10940 2547 10974 2567
rect 10940 2499 10974 2509
rect 10940 2475 10974 2499
rect 10940 2431 10974 2437
rect 10940 2403 10974 2431
rect 13712 2745 13746 2771
rect 13712 2737 13746 2745
rect 13712 2677 13746 2699
rect 13712 2665 13746 2677
rect 13712 2609 13746 2627
rect 13712 2593 13746 2609
rect 13712 2541 13746 2555
rect 13712 2521 13746 2541
rect 13712 2473 13746 2483
rect 13712 2449 13746 2473
rect 11579 2394 11613 2428
rect 13712 2405 13746 2411
rect 10940 2363 10974 2365
rect 10940 2331 10974 2363
rect 13712 2377 13746 2405
rect 11392 2316 11426 2350
rect 10940 2261 10974 2293
rect 10940 2259 10974 2261
rect 10940 2193 10974 2221
rect 10940 2187 10974 2193
rect 10940 2125 10974 2149
rect 10940 2115 10974 2125
rect 10940 2057 10974 2077
rect 10940 2043 10974 2057
rect 10940 1989 10974 2005
rect 10940 1971 10974 1989
rect 10940 1921 10974 1933
rect 10940 1899 10974 1921
rect 10940 1853 10974 1861
rect 10940 1827 10974 1853
rect 11500 2227 11534 2229
rect 11500 2195 11534 2227
rect 11500 2125 11534 2157
rect 11500 2123 11534 2125
rect 11658 2227 11692 2229
rect 11658 2195 11692 2227
rect 11658 2125 11692 2157
rect 11658 2123 11692 2125
rect 13712 2337 13746 2339
rect 13712 2305 13746 2337
rect 13712 2235 13746 2267
rect 13712 2233 13746 2235
rect 13712 2167 13746 2195
rect 13712 2161 13746 2167
rect 13712 2099 13746 2123
rect 13712 2089 13746 2099
rect 13712 2031 13746 2051
rect 13712 2017 13746 2031
rect 13712 1963 13746 1979
rect 13712 1945 13746 1963
rect 13712 1895 13746 1907
rect 13712 1873 13746 1895
rect 13712 1827 13746 1835
rect 13712 1801 13746 1827
rect 13808 2745 13842 2771
rect 13808 2737 13842 2745
rect 13808 2677 13842 2699
rect 13808 2665 13842 2677
rect 13808 2609 13842 2627
rect 13808 2593 13842 2609
rect 13808 2541 13842 2555
rect 13808 2521 13842 2541
rect 13808 2473 13842 2483
rect 13808 2449 13842 2473
rect 13808 2405 13842 2411
rect 13808 2377 13842 2405
rect 13808 2337 13842 2339
rect 13808 2305 13842 2337
rect 13808 2235 13842 2267
rect 13808 2233 13842 2235
rect 13808 2167 13842 2195
rect 13808 2161 13842 2167
rect 13808 2099 13842 2123
rect 13808 2089 13842 2099
rect 13808 2031 13842 2051
rect 13808 2017 13842 2031
rect 13808 1963 13842 1979
rect 13808 1945 13842 1963
rect 13808 1895 13842 1907
rect 13808 1873 13842 1895
rect 13808 1827 13842 1835
rect 13808 1801 13842 1827
rect 13904 2745 13938 2771
rect 13904 2737 13938 2745
rect 13904 2677 13938 2699
rect 13904 2665 13938 2677
rect 13904 2609 13938 2627
rect 13904 2593 13938 2609
rect 13904 2541 13938 2555
rect 13904 2521 13938 2541
rect 13904 2473 13938 2483
rect 13904 2449 13938 2473
rect 13904 2405 13938 2411
rect 13904 2377 13938 2405
rect 13904 2337 13938 2339
rect 13904 2305 13938 2337
rect 13904 2235 13938 2267
rect 13904 2233 13938 2235
rect 13904 2167 13938 2195
rect 13904 2161 13938 2167
rect 13904 2099 13938 2123
rect 13904 2089 13938 2099
rect 13904 2031 13938 2051
rect 13904 2017 13938 2031
rect 13904 1963 13938 1979
rect 13904 1945 13938 1963
rect 13904 1895 13938 1907
rect 13904 1873 13938 1895
rect 13904 1827 13938 1835
rect 13904 1801 13938 1827
rect 14000 2745 14034 2771
rect 14000 2737 14034 2745
rect 14000 2677 14034 2699
rect 14000 2665 14034 2677
rect 14000 2609 14034 2627
rect 14000 2593 14034 2609
rect 14000 2541 14034 2555
rect 14000 2521 14034 2541
rect 14000 2473 14034 2483
rect 14000 2449 14034 2473
rect 14000 2405 14034 2411
rect 14000 2377 14034 2405
rect 14000 2337 14034 2339
rect 14000 2305 14034 2337
rect 14000 2235 14034 2267
rect 14000 2233 14034 2235
rect 14000 2167 14034 2195
rect 14000 2161 14034 2167
rect 14000 2099 14034 2123
rect 14000 2089 14034 2099
rect 14000 2031 14034 2051
rect 14000 2017 14034 2031
rect 14000 1963 14034 1979
rect 14000 1945 14034 1963
rect 14000 1895 14034 1907
rect 14000 1873 14034 1895
rect 14000 1827 14034 1835
rect 14000 1801 14034 1827
rect 14096 2745 14130 2771
rect 14096 2737 14130 2745
rect 14096 2677 14130 2699
rect 14096 2665 14130 2677
rect 14096 2609 14130 2627
rect 14096 2593 14130 2609
rect 14096 2541 14130 2555
rect 14096 2521 14130 2541
rect 14096 2473 14130 2483
rect 14096 2449 14130 2473
rect 14096 2405 14130 2411
rect 14096 2377 14130 2405
rect 14579 2394 14613 2428
rect 14096 2337 14130 2339
rect 14096 2305 14130 2337
rect 14392 2316 14426 2350
rect 14096 2235 14130 2267
rect 14096 2233 14130 2235
rect 14096 2167 14130 2195
rect 14096 2161 14130 2167
rect 14096 2099 14130 2123
rect 14096 2089 14130 2099
rect 14096 2031 14130 2051
rect 14096 2017 14130 2031
rect 14096 1963 14130 1979
rect 14096 1945 14130 1963
rect 14096 1895 14130 1907
rect 14096 1873 14130 1895
rect 14096 1827 14130 1835
rect 14096 1801 14130 1827
rect 14500 2227 14534 2229
rect 14500 2195 14534 2227
rect 14500 2125 14534 2157
rect 14500 2123 14534 2125
rect 10652 1644 10686 1678
rect 13808 1618 13842 1652
rect 14658 2227 14692 2229
rect 14658 2195 14692 2227
rect 14658 2125 14692 2157
rect 14658 2123 14692 2125
rect 734 1424 768 1458
rect -1095 1264 -1061 1298
rect -899 1264 -865 1298
rect 158 1227 192 1253
rect 158 1219 192 1227
rect -1686 1025 -1652 1051
rect -1686 1017 -1652 1025
rect -1686 957 -1652 979
rect -1686 945 -1652 957
rect -1686 889 -1652 907
rect -1686 873 -1652 889
rect -1686 821 -1652 835
rect -1686 801 -1652 821
rect -1686 753 -1652 763
rect -1686 729 -1652 753
rect -1686 685 -1652 691
rect -1686 657 -1652 685
rect -1686 617 -1652 619
rect -1686 585 -1652 617
rect -1686 515 -1652 547
rect -1686 513 -1652 515
rect -1686 447 -1652 475
rect -1686 441 -1652 447
rect -1686 379 -1652 403
rect -1686 369 -1652 379
rect -1686 311 -1652 331
rect -1686 297 -1652 311
rect -1686 243 -1652 259
rect -1686 225 -1652 243
rect -1686 175 -1652 187
rect -1686 153 -1652 175
rect -1686 107 -1652 115
rect -1686 81 -1652 107
rect -1588 1025 -1554 1051
rect -1588 1017 -1554 1025
rect -1588 957 -1554 979
rect -1588 945 -1554 957
rect -1588 889 -1554 907
rect -1588 873 -1554 889
rect -1588 821 -1554 835
rect -1588 801 -1554 821
rect -1588 753 -1554 763
rect -1588 729 -1554 753
rect -1588 685 -1554 691
rect -1588 657 -1554 685
rect -1588 617 -1554 619
rect -1588 585 -1554 617
rect -1588 515 -1554 547
rect -1588 513 -1554 515
rect -1588 447 -1554 475
rect -1588 441 -1554 447
rect -1588 379 -1554 403
rect -1588 369 -1554 379
rect -1588 311 -1554 331
rect -1588 297 -1554 311
rect -1588 243 -1554 259
rect -1588 225 -1554 243
rect -1588 175 -1554 187
rect -1588 153 -1554 175
rect -1588 107 -1554 115
rect -1588 81 -1554 107
rect -1490 1025 -1456 1051
rect -1490 1017 -1456 1025
rect -1490 957 -1456 979
rect -1490 945 -1456 957
rect -1490 889 -1456 907
rect -1490 873 -1456 889
rect -1490 821 -1456 835
rect -1490 801 -1456 821
rect -1490 753 -1456 763
rect -1490 729 -1456 753
rect -1490 685 -1456 691
rect -1490 657 -1456 685
rect -1490 617 -1456 619
rect -1490 585 -1456 617
rect -1490 515 -1456 547
rect -1490 513 -1456 515
rect -1490 447 -1456 475
rect -1490 441 -1456 447
rect -1490 379 -1456 403
rect -1490 369 -1456 379
rect -1490 311 -1456 331
rect -1490 297 -1456 311
rect -1490 243 -1456 259
rect -1490 225 -1456 243
rect -1490 175 -1456 187
rect -1490 153 -1456 175
rect -1490 107 -1456 115
rect -1490 81 -1456 107
rect -1392 1025 -1358 1051
rect -1392 1017 -1358 1025
rect -1392 957 -1358 979
rect -1392 945 -1358 957
rect -1392 889 -1358 907
rect -1392 873 -1358 889
rect -1392 821 -1358 835
rect -1392 801 -1358 821
rect -1392 753 -1358 763
rect -1392 729 -1358 753
rect -1392 685 -1358 691
rect -1392 657 -1358 685
rect -1392 617 -1358 619
rect -1392 585 -1358 617
rect -1392 515 -1358 547
rect -1392 513 -1358 515
rect -1392 447 -1358 475
rect -1392 441 -1358 447
rect -1392 379 -1358 403
rect -1392 369 -1358 379
rect -1392 311 -1358 331
rect -1392 297 -1358 311
rect -1392 243 -1358 259
rect -1392 225 -1358 243
rect -1392 175 -1358 187
rect -1392 153 -1358 175
rect -1392 107 -1358 115
rect -1392 81 -1358 107
rect -1294 1025 -1260 1051
rect -1294 1017 -1260 1025
rect -1294 957 -1260 979
rect -1294 945 -1260 957
rect -1294 889 -1260 907
rect -1294 873 -1260 889
rect -1294 821 -1260 835
rect -1294 801 -1260 821
rect -1294 753 -1260 763
rect -1294 729 -1260 753
rect -1294 685 -1260 691
rect -1294 657 -1260 685
rect -1294 617 -1260 619
rect -1294 585 -1260 617
rect -1294 515 -1260 547
rect -1294 513 -1260 515
rect -1294 447 -1260 475
rect -1294 441 -1260 447
rect -1294 379 -1260 403
rect -1294 369 -1260 379
rect -1294 311 -1260 331
rect -1294 297 -1260 311
rect -1294 243 -1260 259
rect -1294 225 -1260 243
rect -1294 175 -1260 187
rect -1294 153 -1260 175
rect -1294 107 -1260 115
rect -1294 81 -1260 107
rect -1196 1025 -1162 1051
rect -1196 1017 -1162 1025
rect -1196 957 -1162 979
rect -1196 945 -1162 957
rect -1196 889 -1162 907
rect -1196 873 -1162 889
rect -1196 821 -1162 835
rect -1196 801 -1162 821
rect -1196 753 -1162 763
rect -1196 729 -1162 753
rect -1196 685 -1162 691
rect -1196 657 -1162 685
rect -1196 617 -1162 619
rect -1196 585 -1162 617
rect -1196 515 -1162 547
rect -1196 513 -1162 515
rect -1196 447 -1162 475
rect -1196 441 -1162 447
rect -1196 379 -1162 403
rect -1196 369 -1162 379
rect -1196 311 -1162 331
rect -1196 297 -1162 311
rect -1196 243 -1162 259
rect -1196 225 -1162 243
rect -1196 175 -1162 187
rect -1196 153 -1162 175
rect -1196 107 -1162 115
rect -1196 81 -1162 107
rect -1098 1025 -1064 1051
rect -1098 1017 -1064 1025
rect -1098 957 -1064 979
rect -1098 945 -1064 957
rect -1098 889 -1064 907
rect -1098 873 -1064 889
rect -1098 821 -1064 835
rect -1098 801 -1064 821
rect -1098 753 -1064 763
rect -1098 729 -1064 753
rect -1098 685 -1064 691
rect -1098 657 -1064 685
rect -1098 617 -1064 619
rect -1098 585 -1064 617
rect -1098 515 -1064 547
rect -1098 513 -1064 515
rect -1098 447 -1064 475
rect -1098 441 -1064 447
rect -1098 379 -1064 403
rect -1098 369 -1064 379
rect -1098 311 -1064 331
rect -1098 297 -1064 311
rect -1098 243 -1064 259
rect -1098 225 -1064 243
rect -1098 175 -1064 187
rect -1098 153 -1064 175
rect -1098 107 -1064 115
rect -1098 81 -1064 107
rect 158 1159 192 1181
rect 158 1147 192 1159
rect 158 1091 192 1109
rect 158 1075 192 1091
rect -1000 1025 -966 1051
rect -1000 1017 -966 1025
rect -1000 957 -966 979
rect -1000 945 -966 957
rect -1000 889 -966 907
rect -1000 873 -966 889
rect -1000 821 -966 835
rect -1000 801 -966 821
rect -1000 753 -966 763
rect -1000 729 -966 753
rect -1000 685 -966 691
rect -1000 657 -966 685
rect -1000 617 -966 619
rect -1000 585 -966 617
rect -1000 515 -966 547
rect -1000 513 -966 515
rect -1000 447 -966 475
rect -1000 441 -966 447
rect -1000 379 -966 403
rect -1000 369 -966 379
rect -1000 311 -966 331
rect -1000 297 -966 311
rect -1000 243 -966 259
rect -1000 225 -966 243
rect -1000 175 -966 187
rect -1000 153 -966 175
rect -1000 107 -966 115
rect -1000 81 -966 107
rect -902 1025 -868 1051
rect -902 1017 -868 1025
rect -902 957 -868 979
rect -902 945 -868 957
rect -902 889 -868 907
rect -902 873 -868 889
rect -902 821 -868 835
rect -902 801 -868 821
rect -902 753 -868 763
rect -902 729 -868 753
rect -902 685 -868 691
rect -902 657 -868 685
rect -902 617 -868 619
rect -902 585 -868 617
rect -902 515 -868 547
rect -902 513 -868 515
rect -902 447 -868 475
rect -902 441 -868 447
rect -902 379 -868 403
rect -902 369 -868 379
rect -902 311 -868 331
rect -902 297 -868 311
rect -902 243 -868 259
rect -902 225 -868 243
rect -902 175 -868 187
rect 158 1023 192 1037
rect 158 1003 192 1023
rect 158 955 192 965
rect 158 931 192 955
rect 158 887 192 893
rect 158 859 192 887
rect 158 819 192 821
rect 158 787 192 819
rect 158 717 192 749
rect 158 715 192 717
rect 158 649 192 677
rect 158 643 192 649
rect 158 581 192 605
rect 158 571 192 581
rect 158 513 192 533
rect 158 499 192 513
rect 158 445 192 461
rect 158 427 192 445
rect 158 377 192 389
rect 158 355 192 377
rect 158 309 192 317
rect 158 283 192 309
rect 254 1227 288 1253
rect 254 1219 288 1227
rect 254 1159 288 1181
rect 254 1147 288 1159
rect 254 1091 288 1109
rect 254 1075 288 1091
rect 254 1023 288 1037
rect 254 1003 288 1023
rect 254 955 288 965
rect 254 931 288 955
rect 254 887 288 893
rect 254 859 288 887
rect 254 819 288 821
rect 254 787 288 819
rect 254 717 288 749
rect 254 715 288 717
rect 254 649 288 677
rect 254 643 288 649
rect 254 581 288 605
rect 254 571 288 581
rect 254 513 288 533
rect 254 499 288 513
rect 254 445 288 461
rect 254 427 288 445
rect 254 377 288 389
rect 254 355 288 377
rect 254 309 288 317
rect 254 283 288 309
rect 350 1227 384 1253
rect 350 1219 384 1227
rect 350 1159 384 1181
rect 350 1147 384 1159
rect 350 1091 384 1109
rect 350 1075 384 1091
rect 350 1023 384 1037
rect 350 1003 384 1023
rect 350 955 384 965
rect 350 931 384 955
rect 350 887 384 893
rect 350 859 384 887
rect 350 819 384 821
rect 350 787 384 819
rect 350 717 384 749
rect 350 715 384 717
rect 350 649 384 677
rect 350 643 384 649
rect 350 581 384 605
rect 350 571 384 581
rect 350 513 384 533
rect 350 499 384 513
rect 350 445 384 461
rect 350 427 384 445
rect 350 377 384 389
rect 350 355 384 377
rect 350 309 384 317
rect 350 283 384 309
rect 446 1227 480 1253
rect 446 1219 480 1227
rect 446 1159 480 1181
rect 446 1147 480 1159
rect 446 1091 480 1109
rect 446 1075 480 1091
rect 446 1023 480 1037
rect 446 1003 480 1023
rect 446 955 480 965
rect 446 931 480 955
rect 446 887 480 893
rect 446 859 480 887
rect 446 819 480 821
rect 446 787 480 819
rect 446 717 480 749
rect 446 715 480 717
rect 446 649 480 677
rect 446 643 480 649
rect 446 581 480 605
rect 446 571 480 581
rect 446 513 480 533
rect 446 499 480 513
rect 446 445 480 461
rect 446 427 480 445
rect 446 377 480 389
rect 446 355 480 377
rect 446 309 480 317
rect 446 283 480 309
rect 542 1227 576 1253
rect 542 1219 576 1227
rect 542 1159 576 1181
rect 542 1147 576 1159
rect 542 1091 576 1109
rect 542 1075 576 1091
rect 542 1023 576 1037
rect 542 1003 576 1023
rect 542 955 576 965
rect 542 931 576 955
rect 542 887 576 893
rect 542 859 576 887
rect 542 819 576 821
rect 542 787 576 819
rect 542 717 576 749
rect 542 715 576 717
rect 542 649 576 677
rect 542 643 576 649
rect 542 581 576 605
rect 542 571 576 581
rect 542 513 576 533
rect 542 499 576 513
rect 542 445 576 461
rect 542 427 576 445
rect 542 377 576 389
rect 542 355 576 377
rect 542 309 576 317
rect 542 283 576 309
rect 638 1227 672 1253
rect 638 1219 672 1227
rect 638 1159 672 1181
rect 638 1147 672 1159
rect 638 1091 672 1109
rect 638 1075 672 1091
rect 638 1023 672 1037
rect 638 1003 672 1023
rect 638 955 672 965
rect 638 931 672 955
rect 638 887 672 893
rect 638 859 672 887
rect 638 819 672 821
rect 638 787 672 819
rect 638 717 672 749
rect 638 715 672 717
rect 638 649 672 677
rect 638 643 672 649
rect 638 581 672 605
rect 638 571 672 581
rect 638 513 672 533
rect 638 499 672 513
rect 638 445 672 461
rect 638 427 672 445
rect 638 377 672 389
rect 638 355 672 377
rect 638 309 672 317
rect 638 283 672 309
rect 734 1227 768 1253
rect 734 1219 768 1227
rect 734 1159 768 1181
rect 734 1147 768 1159
rect 734 1091 768 1109
rect 734 1075 768 1091
rect 734 1023 768 1037
rect 734 1003 768 1023
rect 734 955 768 965
rect 734 931 768 955
rect 734 887 768 893
rect 734 859 768 887
rect 734 819 768 821
rect 734 787 768 819
rect 734 717 768 749
rect 734 715 768 717
rect 734 649 768 677
rect 734 643 768 649
rect 734 581 768 605
rect 734 571 768 581
rect 734 513 768 533
rect 734 499 768 513
rect 734 445 768 461
rect 734 427 768 445
rect 734 377 768 389
rect 734 355 768 377
rect 734 309 768 317
rect 734 283 768 309
rect 830 1227 864 1253
rect 830 1219 864 1227
rect 830 1159 864 1181
rect 830 1147 864 1159
rect 830 1091 864 1109
rect 830 1075 864 1091
rect 830 1023 864 1037
rect 830 1003 864 1023
rect 830 955 864 965
rect 830 931 864 955
rect 830 887 864 893
rect 830 859 864 887
rect 830 819 864 821
rect 830 787 864 819
rect 830 717 864 749
rect 830 715 864 717
rect 830 649 864 677
rect 830 643 864 649
rect 830 581 864 605
rect 830 571 864 581
rect 830 513 864 533
rect 830 499 864 513
rect 830 445 864 461
rect 830 427 864 445
rect 830 377 864 389
rect 830 355 864 377
rect 830 309 864 317
rect 830 283 864 309
rect 926 1227 960 1253
rect 926 1219 960 1227
rect 926 1159 960 1181
rect 926 1147 960 1159
rect 926 1091 960 1109
rect 926 1075 960 1091
rect 926 1023 960 1037
rect 926 1003 960 1023
rect 926 955 960 965
rect 926 931 960 955
rect 926 887 960 893
rect 926 859 960 887
rect 926 819 960 821
rect 926 787 960 819
rect 926 717 960 749
rect 926 715 960 717
rect 926 649 960 677
rect 926 643 960 649
rect 926 581 960 605
rect 926 571 960 581
rect 926 513 960 533
rect 926 499 960 513
rect 926 445 960 461
rect 926 427 960 445
rect 926 377 960 389
rect 926 355 960 377
rect 926 309 960 317
rect 926 283 960 309
rect 1022 1227 1056 1253
rect 1022 1219 1056 1227
rect 1022 1159 1056 1181
rect 1022 1147 1056 1159
rect 1022 1091 1056 1109
rect 1022 1075 1056 1091
rect 1022 1023 1056 1037
rect 1022 1003 1056 1023
rect 1022 955 1056 965
rect 1022 931 1056 955
rect 1022 887 1056 893
rect 1022 859 1056 887
rect 1022 819 1056 821
rect 1022 787 1056 819
rect 1022 717 1056 749
rect 1022 715 1056 717
rect 1022 649 1056 677
rect 1022 643 1056 649
rect 1022 581 1056 605
rect 1022 571 1056 581
rect 1022 513 1056 533
rect 1022 499 1056 513
rect 1022 445 1056 461
rect 1022 427 1056 445
rect 1022 377 1056 389
rect 1022 355 1056 377
rect 1022 309 1056 317
rect 1022 283 1056 309
rect 1118 1227 1152 1253
rect 1118 1219 1152 1227
rect 1118 1159 1152 1181
rect 1118 1147 1152 1159
rect 1118 1091 1152 1109
rect 1118 1075 1152 1091
rect 1118 1023 1152 1037
rect 1118 1003 1152 1023
rect 1118 955 1152 965
rect 1118 931 1152 955
rect 1118 887 1152 893
rect 1118 859 1152 887
rect 1118 819 1152 821
rect 1118 787 1152 819
rect 1118 717 1152 749
rect 1118 715 1152 717
rect 1118 649 1152 677
rect 1118 643 1152 649
rect 1118 581 1152 605
rect 1118 571 1152 581
rect 1118 513 1152 533
rect 1118 499 1152 513
rect 1118 445 1152 461
rect 1118 427 1152 445
rect 1118 377 1152 389
rect 1118 355 1152 377
rect 1118 309 1152 317
rect 1118 283 1152 309
rect 1214 1227 1248 1253
rect 1214 1219 1248 1227
rect 1214 1159 1248 1181
rect 1214 1147 1248 1159
rect 1214 1091 1248 1109
rect 1214 1075 1248 1091
rect 1214 1023 1248 1037
rect 1214 1003 1248 1023
rect 1214 955 1248 965
rect 1214 931 1248 955
rect 1214 887 1248 893
rect 1214 859 1248 887
rect 1214 819 1248 821
rect 1214 787 1248 819
rect 1214 717 1248 749
rect 1214 715 1248 717
rect 1214 649 1248 677
rect 1214 643 1248 649
rect 1214 581 1248 605
rect 1214 571 1248 581
rect 1214 513 1248 533
rect 1214 499 1248 513
rect 1214 445 1248 461
rect 1214 427 1248 445
rect 1214 377 1248 389
rect 1214 355 1248 377
rect 1214 309 1248 317
rect 1214 283 1248 309
rect 1310 1227 1344 1253
rect 1310 1219 1344 1227
rect 1310 1159 1344 1181
rect 1310 1147 1344 1159
rect 1310 1091 1344 1109
rect 1310 1075 1344 1091
rect 1310 1023 1344 1037
rect 1310 1003 1344 1023
rect 1310 955 1344 965
rect 1310 931 1344 955
rect 1310 887 1344 893
rect 1310 859 1344 887
rect 1310 819 1344 821
rect 1310 787 1344 819
rect 1310 717 1344 749
rect 1310 715 1344 717
rect 1310 649 1344 677
rect 1310 643 1344 649
rect 1310 581 1344 605
rect 1310 571 1344 581
rect 1310 513 1344 533
rect 1310 499 1344 513
rect 1310 445 1344 461
rect 1310 427 1344 445
rect 1310 377 1344 389
rect 1310 355 1344 377
rect 1310 309 1344 317
rect 1310 283 1344 309
rect -902 153 -868 175
rect -902 107 -868 115
rect -902 81 -868 107
rect 156 96 190 130
rect 830 86 864 120
rect 2400 1418 2434 1452
rect 3690 1408 3724 1442
rect 1926 1227 1960 1253
rect 1926 1219 1960 1227
rect 1926 1159 1960 1181
rect 1926 1147 1960 1159
rect 1926 1091 1960 1109
rect 1926 1075 1960 1091
rect 1926 1023 1960 1037
rect 1926 1003 1960 1023
rect 1926 955 1960 965
rect 1926 931 1960 955
rect 1926 887 1960 893
rect 1926 859 1960 887
rect 1926 819 1960 821
rect 1926 787 1960 819
rect 1926 717 1960 749
rect 1926 715 1960 717
rect 1926 649 1960 677
rect 1926 643 1960 649
rect 1926 581 1960 605
rect 1926 571 1960 581
rect 1926 513 1960 533
rect 1926 499 1960 513
rect 1926 445 1960 461
rect 1926 427 1960 445
rect 1926 377 1960 389
rect 1926 355 1960 377
rect 1926 309 1960 317
rect 1926 283 1960 309
rect 2022 1227 2056 1253
rect 2022 1219 2056 1227
rect 2022 1159 2056 1181
rect 2022 1147 2056 1159
rect 2022 1091 2056 1109
rect 2022 1075 2056 1091
rect 2022 1023 2056 1037
rect 2022 1003 2056 1023
rect 2022 955 2056 965
rect 2022 931 2056 955
rect 2022 887 2056 893
rect 2022 859 2056 887
rect 2022 819 2056 821
rect 2022 787 2056 819
rect 2022 717 2056 749
rect 2022 715 2056 717
rect 2022 649 2056 677
rect 2022 643 2056 649
rect 2022 581 2056 605
rect 2022 571 2056 581
rect 2022 513 2056 533
rect 2022 499 2056 513
rect 2022 445 2056 461
rect 2022 427 2056 445
rect 2022 377 2056 389
rect 2022 355 2056 377
rect 2022 309 2056 317
rect 2022 283 2056 309
rect 2118 1227 2152 1253
rect 2118 1219 2152 1227
rect 2118 1159 2152 1181
rect 2118 1147 2152 1159
rect 2118 1091 2152 1109
rect 2118 1075 2152 1091
rect 2118 1023 2152 1037
rect 2118 1003 2152 1023
rect 2118 955 2152 965
rect 2118 931 2152 955
rect 2118 887 2152 893
rect 2118 859 2152 887
rect 2118 819 2152 821
rect 2118 787 2152 819
rect 2118 717 2152 749
rect 2118 715 2152 717
rect 2118 649 2152 677
rect 2118 643 2152 649
rect 2118 581 2152 605
rect 2118 571 2152 581
rect 2118 513 2152 533
rect 2118 499 2152 513
rect 2118 445 2152 461
rect 2118 427 2152 445
rect 2118 377 2152 389
rect 2118 355 2152 377
rect 2118 309 2152 317
rect 2118 283 2152 309
rect 2214 1227 2248 1253
rect 2214 1219 2248 1227
rect 2214 1159 2248 1181
rect 2214 1147 2248 1159
rect 2214 1091 2248 1109
rect 2214 1075 2248 1091
rect 2214 1023 2248 1037
rect 2214 1003 2248 1023
rect 2214 955 2248 965
rect 2214 931 2248 955
rect 2214 887 2248 893
rect 2214 859 2248 887
rect 2214 819 2248 821
rect 2214 787 2248 819
rect 2214 717 2248 749
rect 2214 715 2248 717
rect 2214 649 2248 677
rect 2214 643 2248 649
rect 2214 581 2248 605
rect 2214 571 2248 581
rect 2214 513 2248 533
rect 2214 499 2248 513
rect 2214 445 2248 461
rect 2214 427 2248 445
rect 2214 377 2248 389
rect 2214 355 2248 377
rect 2214 309 2248 317
rect 2214 283 2248 309
rect 2310 1227 2344 1253
rect 2310 1219 2344 1227
rect 2310 1159 2344 1181
rect 2310 1147 2344 1159
rect 2310 1091 2344 1109
rect 2310 1075 2344 1091
rect 2310 1023 2344 1037
rect 2310 1003 2344 1023
rect 2310 955 2344 965
rect 2310 931 2344 955
rect 2310 887 2344 893
rect 2310 859 2344 887
rect 2310 819 2344 821
rect 2310 787 2344 819
rect 2310 717 2344 749
rect 2310 715 2344 717
rect 2310 649 2344 677
rect 2310 643 2344 649
rect 2310 581 2344 605
rect 2310 571 2344 581
rect 2310 513 2344 533
rect 2310 499 2344 513
rect 2310 445 2344 461
rect 2310 427 2344 445
rect 2310 377 2344 389
rect 2310 355 2344 377
rect 2310 309 2344 317
rect 2310 283 2344 309
rect 2406 1227 2440 1253
rect 2406 1219 2440 1227
rect 2406 1159 2440 1181
rect 2406 1147 2440 1159
rect 2406 1091 2440 1109
rect 2406 1075 2440 1091
rect 2406 1023 2440 1037
rect 2406 1003 2440 1023
rect 2406 955 2440 965
rect 2406 931 2440 955
rect 2406 887 2440 893
rect 2406 859 2440 887
rect 2406 819 2440 821
rect 2406 787 2440 819
rect 2406 717 2440 749
rect 2406 715 2440 717
rect 2406 649 2440 677
rect 2406 643 2440 649
rect 2406 581 2440 605
rect 2406 571 2440 581
rect 2406 513 2440 533
rect 2406 499 2440 513
rect 2406 445 2440 461
rect 2406 427 2440 445
rect 2406 377 2440 389
rect 2406 355 2440 377
rect 2406 309 2440 317
rect 2406 283 2440 309
rect 2502 1227 2536 1253
rect 2502 1219 2536 1227
rect 2502 1159 2536 1181
rect 2502 1147 2536 1159
rect 2502 1091 2536 1109
rect 2502 1075 2536 1091
rect 2502 1023 2536 1037
rect 2502 1003 2536 1023
rect 2502 955 2536 965
rect 2502 931 2536 955
rect 2502 887 2536 893
rect 2502 859 2536 887
rect 2502 819 2536 821
rect 2502 787 2536 819
rect 2502 717 2536 749
rect 2502 715 2536 717
rect 2502 649 2536 677
rect 2502 643 2536 649
rect 2502 581 2536 605
rect 2502 571 2536 581
rect 2502 513 2536 533
rect 2502 499 2536 513
rect 2502 445 2536 461
rect 2502 427 2536 445
rect 2502 377 2536 389
rect 2502 355 2536 377
rect 2502 309 2536 317
rect 2502 283 2536 309
rect 2598 1227 2632 1253
rect 2598 1219 2632 1227
rect 2598 1159 2632 1181
rect 2598 1147 2632 1159
rect 2598 1091 2632 1109
rect 2598 1075 2632 1091
rect 2598 1023 2632 1037
rect 2598 1003 2632 1023
rect 2598 955 2632 965
rect 2598 931 2632 955
rect 2598 887 2632 893
rect 2598 859 2632 887
rect 2598 819 2632 821
rect 2598 787 2632 819
rect 2598 717 2632 749
rect 2598 715 2632 717
rect 2598 649 2632 677
rect 2598 643 2632 649
rect 2598 581 2632 605
rect 2598 571 2632 581
rect 2598 513 2632 533
rect 2598 499 2632 513
rect 2598 445 2632 461
rect 2598 427 2632 445
rect 2598 377 2632 389
rect 2598 355 2632 377
rect 2598 309 2632 317
rect 2598 283 2632 309
rect 2694 1227 2728 1253
rect 2694 1219 2728 1227
rect 2694 1159 2728 1181
rect 2694 1147 2728 1159
rect 2694 1091 2728 1109
rect 2694 1075 2728 1091
rect 2694 1023 2728 1037
rect 2694 1003 2728 1023
rect 2694 955 2728 965
rect 2694 931 2728 955
rect 2694 887 2728 893
rect 2694 859 2728 887
rect 2694 819 2728 821
rect 2694 787 2728 819
rect 2694 717 2728 749
rect 2694 715 2728 717
rect 2694 649 2728 677
rect 2694 643 2728 649
rect 2694 581 2728 605
rect 2694 571 2728 581
rect 2694 513 2728 533
rect 2694 499 2728 513
rect 2694 445 2728 461
rect 2694 427 2728 445
rect 2694 377 2728 389
rect 2694 355 2728 377
rect 2694 309 2728 317
rect 2694 283 2728 309
rect 2790 1227 2824 1253
rect 2790 1219 2824 1227
rect 2790 1159 2824 1181
rect 2790 1147 2824 1159
rect 2790 1091 2824 1109
rect 2790 1075 2824 1091
rect 2790 1023 2824 1037
rect 2790 1003 2824 1023
rect 2790 955 2824 965
rect 2790 931 2824 955
rect 2790 887 2824 893
rect 2790 859 2824 887
rect 2790 819 2824 821
rect 2790 787 2824 819
rect 2790 717 2824 749
rect 2790 715 2824 717
rect 2790 649 2824 677
rect 2790 643 2824 649
rect 2790 581 2824 605
rect 2790 571 2824 581
rect 2790 513 2824 533
rect 2790 499 2824 513
rect 2790 445 2824 461
rect 2790 427 2824 445
rect 2790 377 2824 389
rect 2790 355 2824 377
rect 2790 309 2824 317
rect 2790 283 2824 309
rect 2886 1227 2920 1253
rect 2886 1219 2920 1227
rect 2886 1159 2920 1181
rect 2886 1147 2920 1159
rect 2886 1091 2920 1109
rect 2886 1075 2920 1091
rect 2886 1023 2920 1037
rect 2886 1003 2920 1023
rect 2886 955 2920 965
rect 2886 931 2920 955
rect 2886 887 2920 893
rect 2886 859 2920 887
rect 2886 819 2920 821
rect 2886 787 2920 819
rect 2886 717 2920 749
rect 2886 715 2920 717
rect 2886 649 2920 677
rect 2886 643 2920 649
rect 2886 581 2920 605
rect 2886 571 2920 581
rect 2886 513 2920 533
rect 2886 499 2920 513
rect 2886 445 2920 461
rect 2886 427 2920 445
rect 2886 377 2920 389
rect 2886 355 2920 377
rect 2886 309 2920 317
rect 2886 283 2920 309
rect 2982 1227 3016 1253
rect 2982 1219 3016 1227
rect 2982 1159 3016 1181
rect 2982 1147 3016 1159
rect 2982 1091 3016 1109
rect 2982 1075 3016 1091
rect 2982 1023 3016 1037
rect 2982 1003 3016 1023
rect 2982 955 3016 965
rect 2982 931 3016 955
rect 2982 887 3016 893
rect 2982 859 3016 887
rect 2982 819 3016 821
rect 2982 787 3016 819
rect 2982 717 3016 749
rect 2982 715 3016 717
rect 2982 649 3016 677
rect 2982 643 3016 649
rect 2982 581 3016 605
rect 2982 571 3016 581
rect 2982 513 3016 533
rect 2982 499 3016 513
rect 2982 445 3016 461
rect 2982 427 3016 445
rect 2982 377 3016 389
rect 2982 355 3016 377
rect 2982 309 3016 317
rect 2982 283 3016 309
rect 3114 1211 3148 1237
rect 3114 1203 3148 1211
rect 3114 1143 3148 1165
rect 3114 1131 3148 1143
rect 3114 1075 3148 1093
rect 3114 1059 3148 1075
rect 3114 1007 3148 1021
rect 3114 987 3148 1007
rect 3114 939 3148 949
rect 3114 915 3148 939
rect 3114 871 3148 877
rect 3114 843 3148 871
rect 3114 803 3148 805
rect 3114 771 3148 803
rect 3114 701 3148 733
rect 3114 699 3148 701
rect 3114 633 3148 661
rect 3114 627 3148 633
rect 3114 565 3148 589
rect 3114 555 3148 565
rect 3114 497 3148 517
rect 3114 483 3148 497
rect 3114 429 3148 445
rect 3114 411 3148 429
rect 3114 361 3148 373
rect 3114 339 3148 361
rect 3114 293 3148 301
rect 3114 267 3148 293
rect 3210 1211 3244 1237
rect 3210 1203 3244 1211
rect 3210 1143 3244 1165
rect 3210 1131 3244 1143
rect 3210 1075 3244 1093
rect 3210 1059 3244 1075
rect 3210 1007 3244 1021
rect 3210 987 3244 1007
rect 3210 939 3244 949
rect 3210 915 3244 939
rect 3210 871 3244 877
rect 3210 843 3244 871
rect 3210 803 3244 805
rect 3210 771 3244 803
rect 3210 701 3244 733
rect 3210 699 3244 701
rect 3210 633 3244 661
rect 3210 627 3244 633
rect 3210 565 3244 589
rect 3210 555 3244 565
rect 3210 497 3244 517
rect 3210 483 3244 497
rect 3210 429 3244 445
rect 3210 411 3244 429
rect 3210 361 3244 373
rect 3210 339 3244 361
rect 3210 293 3244 301
rect 3210 267 3244 293
rect 3306 1211 3340 1237
rect 3306 1203 3340 1211
rect 3306 1143 3340 1165
rect 3306 1131 3340 1143
rect 3306 1075 3340 1093
rect 3306 1059 3340 1075
rect 3306 1007 3340 1021
rect 3306 987 3340 1007
rect 3306 939 3340 949
rect 3306 915 3340 939
rect 3306 871 3340 877
rect 3306 843 3340 871
rect 3306 803 3340 805
rect 3306 771 3340 803
rect 3306 701 3340 733
rect 3306 699 3340 701
rect 3306 633 3340 661
rect 3306 627 3340 633
rect 3306 565 3340 589
rect 3306 555 3340 565
rect 3306 497 3340 517
rect 3306 483 3340 497
rect 3306 429 3340 445
rect 3306 411 3340 429
rect 3306 361 3340 373
rect 3306 339 3340 361
rect 3306 293 3340 301
rect 3306 267 3340 293
rect 3402 1211 3436 1237
rect 3402 1203 3436 1211
rect 3402 1143 3436 1165
rect 3402 1131 3436 1143
rect 3402 1075 3436 1093
rect 3402 1059 3436 1075
rect 3402 1007 3436 1021
rect 3402 987 3436 1007
rect 3402 939 3436 949
rect 3402 915 3436 939
rect 3402 871 3436 877
rect 3402 843 3436 871
rect 3402 803 3436 805
rect 3402 771 3436 803
rect 3402 701 3436 733
rect 3402 699 3436 701
rect 3402 633 3436 661
rect 3402 627 3436 633
rect 3402 565 3436 589
rect 3402 555 3436 565
rect 3402 497 3436 517
rect 3402 483 3436 497
rect 3402 429 3436 445
rect 3402 411 3436 429
rect 3402 361 3436 373
rect 3402 339 3436 361
rect 3402 293 3436 301
rect 3402 267 3436 293
rect 3498 1211 3532 1237
rect 3498 1203 3532 1211
rect 3498 1143 3532 1165
rect 3498 1131 3532 1143
rect 3498 1075 3532 1093
rect 3498 1059 3532 1075
rect 3498 1007 3532 1021
rect 3498 987 3532 1007
rect 3498 939 3532 949
rect 3498 915 3532 939
rect 3498 871 3532 877
rect 3498 843 3532 871
rect 3498 803 3532 805
rect 3498 771 3532 803
rect 3498 701 3532 733
rect 3498 699 3532 701
rect 3498 633 3532 661
rect 3498 627 3532 633
rect 3498 565 3532 589
rect 3498 555 3532 565
rect 3498 497 3532 517
rect 3498 483 3532 497
rect 3498 429 3532 445
rect 3498 411 3532 429
rect 3498 361 3532 373
rect 3498 339 3532 361
rect 3498 293 3532 301
rect 3498 267 3532 293
rect 3594 1211 3628 1237
rect 3594 1203 3628 1211
rect 3594 1143 3628 1165
rect 3594 1131 3628 1143
rect 3594 1075 3628 1093
rect 3594 1059 3628 1075
rect 3594 1007 3628 1021
rect 3594 987 3628 1007
rect 3594 939 3628 949
rect 3594 915 3628 939
rect 3594 871 3628 877
rect 3594 843 3628 871
rect 3594 803 3628 805
rect 3594 771 3628 803
rect 3594 701 3628 733
rect 3594 699 3628 701
rect 3594 633 3628 661
rect 3594 627 3628 633
rect 3594 565 3628 589
rect 3594 555 3628 565
rect 3594 497 3628 517
rect 3594 483 3628 497
rect 3594 429 3628 445
rect 3594 411 3628 429
rect 3594 361 3628 373
rect 3594 339 3628 361
rect 3594 293 3628 301
rect 3594 267 3628 293
rect 3690 1211 3724 1237
rect 3690 1203 3724 1211
rect 3690 1143 3724 1165
rect 3690 1131 3724 1143
rect 3690 1075 3724 1093
rect 3690 1059 3724 1075
rect 3690 1007 3724 1021
rect 3690 987 3724 1007
rect 3690 939 3724 949
rect 3690 915 3724 939
rect 3690 871 3724 877
rect 3690 843 3724 871
rect 3690 803 3724 805
rect 3690 771 3724 803
rect 3690 701 3724 733
rect 3690 699 3724 701
rect 3690 633 3724 661
rect 3690 627 3724 633
rect 3690 565 3724 589
rect 3690 555 3724 565
rect 3690 497 3724 517
rect 3690 483 3724 497
rect 3690 429 3724 445
rect 3690 411 3724 429
rect 3690 361 3724 373
rect 3690 339 3724 361
rect 3690 293 3724 301
rect 3690 267 3724 293
rect 3786 1211 3820 1237
rect 3786 1203 3820 1211
rect 3786 1143 3820 1165
rect 3786 1131 3820 1143
rect 3786 1075 3820 1093
rect 3786 1059 3820 1075
rect 3786 1007 3820 1021
rect 3786 987 3820 1007
rect 3786 939 3820 949
rect 3786 915 3820 939
rect 3786 871 3820 877
rect 3786 843 3820 871
rect 3786 803 3820 805
rect 3786 771 3820 803
rect 3786 701 3820 733
rect 3786 699 3820 701
rect 3786 633 3820 661
rect 3786 627 3820 633
rect 3786 565 3820 589
rect 3786 555 3820 565
rect 3786 497 3820 517
rect 3786 483 3820 497
rect 3786 429 3820 445
rect 3786 411 3820 429
rect 3786 361 3820 373
rect 3786 339 3820 361
rect 3786 293 3820 301
rect 3786 267 3820 293
rect 3882 1211 3916 1237
rect 3882 1203 3916 1211
rect 3882 1143 3916 1165
rect 3882 1131 3916 1143
rect 3882 1075 3916 1093
rect 3882 1059 3916 1075
rect 3882 1007 3916 1021
rect 3882 987 3916 1007
rect 3882 939 3916 949
rect 3882 915 3916 939
rect 3882 871 3916 877
rect 3882 843 3916 871
rect 3882 803 3916 805
rect 3882 771 3916 803
rect 3882 701 3916 733
rect 3882 699 3916 701
rect 3882 633 3916 661
rect 3882 627 3916 633
rect 3882 565 3916 589
rect 3882 555 3916 565
rect 3882 497 3916 517
rect 3882 483 3916 497
rect 3882 429 3916 445
rect 3882 411 3916 429
rect 3882 361 3916 373
rect 3882 339 3916 361
rect 3882 293 3916 301
rect 3882 267 3916 293
rect 3978 1211 4012 1237
rect 3978 1203 4012 1211
rect 3978 1143 4012 1165
rect 3978 1131 4012 1143
rect 3978 1075 4012 1093
rect 3978 1059 4012 1075
rect 3978 1007 4012 1021
rect 3978 987 4012 1007
rect 3978 939 4012 949
rect 3978 915 4012 939
rect 3978 871 4012 877
rect 3978 843 4012 871
rect 3978 803 4012 805
rect 3978 771 4012 803
rect 3978 701 4012 733
rect 3978 699 4012 701
rect 3978 633 4012 661
rect 3978 627 4012 633
rect 3978 565 4012 589
rect 3978 555 4012 565
rect 3978 497 4012 517
rect 3978 483 4012 497
rect 3978 429 4012 445
rect 3978 411 4012 429
rect 3978 361 4012 373
rect 3978 339 4012 361
rect 3978 293 4012 301
rect 3978 267 4012 293
rect 4074 1211 4108 1237
rect 4074 1203 4108 1211
rect 4074 1143 4108 1165
rect 4074 1131 4108 1143
rect 4074 1075 4108 1093
rect 4074 1059 4108 1075
rect 4074 1007 4108 1021
rect 4074 987 4108 1007
rect 4074 939 4108 949
rect 4074 915 4108 939
rect 4074 871 4108 877
rect 4074 843 4108 871
rect 4074 803 4108 805
rect 4074 771 4108 803
rect 4074 701 4108 733
rect 4074 699 4108 701
rect 4074 633 4108 661
rect 4074 627 4108 633
rect 4074 565 4108 589
rect 4074 555 4108 565
rect 4074 497 4108 517
rect 4074 483 4108 497
rect 4074 429 4108 445
rect 4074 411 4108 429
rect 4074 361 4108 373
rect 4074 339 4108 361
rect 4074 293 4108 301
rect 4074 267 4108 293
rect 4170 1211 4204 1237
rect 4170 1203 4204 1211
rect 4170 1143 4204 1165
rect 4170 1131 4204 1143
rect 4170 1075 4204 1093
rect 4170 1059 4204 1075
rect 4170 1007 4204 1021
rect 4170 987 4204 1007
rect 4170 939 4204 949
rect 4170 915 4204 939
rect 4170 871 4204 877
rect 4170 843 4204 871
rect 4170 803 4204 805
rect 4170 771 4204 803
rect 4170 701 4204 733
rect 4170 699 4204 701
rect 4170 633 4204 661
rect 4170 627 4204 633
rect 4170 565 4204 589
rect 4170 555 4204 565
rect 4170 497 4204 517
rect 4170 483 4204 497
rect 4170 429 4204 445
rect 4170 411 4204 429
rect 4170 361 4204 373
rect 4170 339 4204 361
rect 4170 293 4204 301
rect 4170 267 4204 293
rect 4266 1211 4300 1237
rect 4266 1203 4300 1211
rect 4266 1143 4300 1165
rect 4266 1131 4300 1143
rect 4266 1075 4300 1093
rect 4266 1059 4300 1075
rect 4266 1007 4300 1021
rect 4266 987 4300 1007
rect 4266 939 4300 949
rect 4266 915 4300 939
rect 4266 871 4300 877
rect 4266 843 4300 871
rect 4266 803 4300 805
rect 4266 771 4300 803
rect 4266 701 4300 733
rect 4266 699 4300 701
rect 4266 633 4300 661
rect 4266 627 4300 633
rect 4266 565 4300 589
rect 4266 555 4300 565
rect 4266 497 4300 517
rect 4266 483 4300 497
rect 4266 429 4300 445
rect 4266 411 4300 429
rect 4266 361 4300 373
rect 4266 339 4300 361
rect 4266 293 4300 301
rect 4266 267 4300 293
rect 2494 112 2528 146
rect 2788 96 2822 130
rect 3112 80 3146 114
rect 3786 70 3820 104
rect 1664 -10 1698 24
rect 5356 1402 5390 1436
rect 6720 1408 6754 1442
rect 4882 1211 4916 1237
rect 4882 1203 4916 1211
rect 4882 1143 4916 1165
rect 4882 1131 4916 1143
rect 4882 1075 4916 1093
rect 4882 1059 4916 1075
rect 4882 1007 4916 1021
rect 4882 987 4916 1007
rect 4882 939 4916 949
rect 4882 915 4916 939
rect 4882 871 4916 877
rect 4882 843 4916 871
rect 4882 803 4916 805
rect 4882 771 4916 803
rect 4882 701 4916 733
rect 4882 699 4916 701
rect 4882 633 4916 661
rect 4882 627 4916 633
rect 4882 565 4916 589
rect 4882 555 4916 565
rect 4882 497 4916 517
rect 4882 483 4916 497
rect 4882 429 4916 445
rect 4882 411 4916 429
rect 4882 361 4916 373
rect 4882 339 4916 361
rect 4882 293 4916 301
rect 4882 267 4916 293
rect 4978 1211 5012 1237
rect 4978 1203 5012 1211
rect 4978 1143 5012 1165
rect 4978 1131 5012 1143
rect 4978 1075 5012 1093
rect 4978 1059 5012 1075
rect 4978 1007 5012 1021
rect 4978 987 5012 1007
rect 4978 939 5012 949
rect 4978 915 5012 939
rect 4978 871 5012 877
rect 4978 843 5012 871
rect 4978 803 5012 805
rect 4978 771 5012 803
rect 4978 701 5012 733
rect 4978 699 5012 701
rect 4978 633 5012 661
rect 4978 627 5012 633
rect 4978 565 5012 589
rect 4978 555 5012 565
rect 4978 497 5012 517
rect 4978 483 5012 497
rect 4978 429 5012 445
rect 4978 411 5012 429
rect 4978 361 5012 373
rect 4978 339 5012 361
rect 4978 293 5012 301
rect 4978 267 5012 293
rect 5074 1211 5108 1237
rect 5074 1203 5108 1211
rect 5074 1143 5108 1165
rect 5074 1131 5108 1143
rect 5074 1075 5108 1093
rect 5074 1059 5108 1075
rect 5074 1007 5108 1021
rect 5074 987 5108 1007
rect 5074 939 5108 949
rect 5074 915 5108 939
rect 5074 871 5108 877
rect 5074 843 5108 871
rect 5074 803 5108 805
rect 5074 771 5108 803
rect 5074 701 5108 733
rect 5074 699 5108 701
rect 5074 633 5108 661
rect 5074 627 5108 633
rect 5074 565 5108 589
rect 5074 555 5108 565
rect 5074 497 5108 517
rect 5074 483 5108 497
rect 5074 429 5108 445
rect 5074 411 5108 429
rect 5074 361 5108 373
rect 5074 339 5108 361
rect 5074 293 5108 301
rect 5074 267 5108 293
rect 5170 1211 5204 1237
rect 5170 1203 5204 1211
rect 5170 1143 5204 1165
rect 5170 1131 5204 1143
rect 5170 1075 5204 1093
rect 5170 1059 5204 1075
rect 5170 1007 5204 1021
rect 5170 987 5204 1007
rect 5170 939 5204 949
rect 5170 915 5204 939
rect 5170 871 5204 877
rect 5170 843 5204 871
rect 5170 803 5204 805
rect 5170 771 5204 803
rect 5170 701 5204 733
rect 5170 699 5204 701
rect 5170 633 5204 661
rect 5170 627 5204 633
rect 5170 565 5204 589
rect 5170 555 5204 565
rect 5170 497 5204 517
rect 5170 483 5204 497
rect 5170 429 5204 445
rect 5170 411 5204 429
rect 5170 361 5204 373
rect 5170 339 5204 361
rect 5170 293 5204 301
rect 5170 267 5204 293
rect 5266 1211 5300 1237
rect 5266 1203 5300 1211
rect 5266 1143 5300 1165
rect 5266 1131 5300 1143
rect 5266 1075 5300 1093
rect 5266 1059 5300 1075
rect 5266 1007 5300 1021
rect 5266 987 5300 1007
rect 5266 939 5300 949
rect 5266 915 5300 939
rect 5266 871 5300 877
rect 5266 843 5300 871
rect 5266 803 5300 805
rect 5266 771 5300 803
rect 5266 701 5300 733
rect 5266 699 5300 701
rect 5266 633 5300 661
rect 5266 627 5300 633
rect 5266 565 5300 589
rect 5266 555 5300 565
rect 5266 497 5300 517
rect 5266 483 5300 497
rect 5266 429 5300 445
rect 5266 411 5300 429
rect 5266 361 5300 373
rect 5266 339 5300 361
rect 5266 293 5300 301
rect 5266 267 5300 293
rect 5362 1211 5396 1237
rect 5362 1203 5396 1211
rect 5362 1143 5396 1165
rect 5362 1131 5396 1143
rect 5362 1075 5396 1093
rect 5362 1059 5396 1075
rect 5362 1007 5396 1021
rect 5362 987 5396 1007
rect 5362 939 5396 949
rect 5362 915 5396 939
rect 5362 871 5396 877
rect 5362 843 5396 871
rect 5362 803 5396 805
rect 5362 771 5396 803
rect 5362 701 5396 733
rect 5362 699 5396 701
rect 5362 633 5396 661
rect 5362 627 5396 633
rect 5362 565 5396 589
rect 5362 555 5396 565
rect 5362 497 5396 517
rect 5362 483 5396 497
rect 5362 429 5396 445
rect 5362 411 5396 429
rect 5362 361 5396 373
rect 5362 339 5396 361
rect 5362 293 5396 301
rect 5362 267 5396 293
rect 5458 1211 5492 1237
rect 5458 1203 5492 1211
rect 5458 1143 5492 1165
rect 5458 1131 5492 1143
rect 5458 1075 5492 1093
rect 5458 1059 5492 1075
rect 5458 1007 5492 1021
rect 5458 987 5492 1007
rect 5458 939 5492 949
rect 5458 915 5492 939
rect 5458 871 5492 877
rect 5458 843 5492 871
rect 5458 803 5492 805
rect 5458 771 5492 803
rect 5458 701 5492 733
rect 5458 699 5492 701
rect 5458 633 5492 661
rect 5458 627 5492 633
rect 5458 565 5492 589
rect 5458 555 5492 565
rect 5458 497 5492 517
rect 5458 483 5492 497
rect 5458 429 5492 445
rect 5458 411 5492 429
rect 5458 361 5492 373
rect 5458 339 5492 361
rect 5458 293 5492 301
rect 5458 267 5492 293
rect 5554 1211 5588 1237
rect 5554 1203 5588 1211
rect 5554 1143 5588 1165
rect 5554 1131 5588 1143
rect 5554 1075 5588 1093
rect 5554 1059 5588 1075
rect 5554 1007 5588 1021
rect 5554 987 5588 1007
rect 5554 939 5588 949
rect 5554 915 5588 939
rect 5554 871 5588 877
rect 5554 843 5588 871
rect 5554 803 5588 805
rect 5554 771 5588 803
rect 5554 701 5588 733
rect 5554 699 5588 701
rect 5554 633 5588 661
rect 5554 627 5588 633
rect 5554 565 5588 589
rect 5554 555 5588 565
rect 5554 497 5588 517
rect 5554 483 5588 497
rect 5554 429 5588 445
rect 5554 411 5588 429
rect 5554 361 5588 373
rect 5554 339 5588 361
rect 5554 293 5588 301
rect 5554 267 5588 293
rect 5650 1211 5684 1237
rect 5650 1203 5684 1211
rect 5650 1143 5684 1165
rect 5650 1131 5684 1143
rect 5650 1075 5684 1093
rect 5650 1059 5684 1075
rect 5650 1007 5684 1021
rect 5650 987 5684 1007
rect 5650 939 5684 949
rect 5650 915 5684 939
rect 5650 871 5684 877
rect 5650 843 5684 871
rect 5650 803 5684 805
rect 5650 771 5684 803
rect 5650 701 5684 733
rect 5650 699 5684 701
rect 5650 633 5684 661
rect 5650 627 5684 633
rect 5650 565 5684 589
rect 5650 555 5684 565
rect 5650 497 5684 517
rect 5650 483 5684 497
rect 5650 429 5684 445
rect 5650 411 5684 429
rect 5650 361 5684 373
rect 5650 339 5684 361
rect 5650 293 5684 301
rect 5650 267 5684 293
rect 5746 1211 5780 1237
rect 5746 1203 5780 1211
rect 5746 1143 5780 1165
rect 5746 1131 5780 1143
rect 5746 1075 5780 1093
rect 5746 1059 5780 1075
rect 5746 1007 5780 1021
rect 5746 987 5780 1007
rect 5746 939 5780 949
rect 5746 915 5780 939
rect 5746 871 5780 877
rect 5746 843 5780 871
rect 5746 803 5780 805
rect 5746 771 5780 803
rect 5746 701 5780 733
rect 5746 699 5780 701
rect 5746 633 5780 661
rect 5746 627 5780 633
rect 5746 565 5780 589
rect 5746 555 5780 565
rect 5746 497 5780 517
rect 5746 483 5780 497
rect 5746 429 5780 445
rect 5746 411 5780 429
rect 5746 361 5780 373
rect 5746 339 5780 361
rect 5746 293 5780 301
rect 5746 267 5780 293
rect 5842 1211 5876 1237
rect 5842 1203 5876 1211
rect 5842 1143 5876 1165
rect 5842 1131 5876 1143
rect 5842 1075 5876 1093
rect 5842 1059 5876 1075
rect 5842 1007 5876 1021
rect 5842 987 5876 1007
rect 5842 939 5876 949
rect 5842 915 5876 939
rect 5842 871 5876 877
rect 5842 843 5876 871
rect 5842 803 5876 805
rect 5842 771 5876 803
rect 5842 701 5876 733
rect 5842 699 5876 701
rect 5842 633 5876 661
rect 5842 627 5876 633
rect 5842 565 5876 589
rect 5842 555 5876 565
rect 5842 497 5876 517
rect 5842 483 5876 497
rect 5842 429 5876 445
rect 5842 411 5876 429
rect 5842 361 5876 373
rect 5842 339 5876 361
rect 5842 293 5876 301
rect 5842 267 5876 293
rect 5938 1211 5972 1237
rect 5938 1203 5972 1211
rect 5938 1143 5972 1165
rect 5938 1131 5972 1143
rect 5938 1075 5972 1093
rect 5938 1059 5972 1075
rect 5938 1007 5972 1021
rect 5938 987 5972 1007
rect 5938 939 5972 949
rect 5938 915 5972 939
rect 5938 871 5972 877
rect 5938 843 5972 871
rect 5938 803 5972 805
rect 5938 771 5972 803
rect 5938 701 5972 733
rect 5938 699 5972 701
rect 5938 633 5972 661
rect 5938 627 5972 633
rect 5938 565 5972 589
rect 5938 555 5972 565
rect 5938 497 5972 517
rect 5938 483 5972 497
rect 5938 429 5972 445
rect 5938 411 5972 429
rect 5938 361 5972 373
rect 5938 339 5972 361
rect 5938 293 5972 301
rect 5938 267 5972 293
rect 6144 1211 6178 1237
rect 6144 1203 6178 1211
rect 6144 1143 6178 1165
rect 6144 1131 6178 1143
rect 6144 1075 6178 1093
rect 6144 1059 6178 1075
rect 6144 1007 6178 1021
rect 6144 987 6178 1007
rect 6144 939 6178 949
rect 6144 915 6178 939
rect 6144 871 6178 877
rect 6144 843 6178 871
rect 6144 803 6178 805
rect 6144 771 6178 803
rect 6144 701 6178 733
rect 6144 699 6178 701
rect 6144 633 6178 661
rect 6144 627 6178 633
rect 6144 565 6178 589
rect 6144 555 6178 565
rect 6144 497 6178 517
rect 6144 483 6178 497
rect 6144 429 6178 445
rect 6144 411 6178 429
rect 6144 361 6178 373
rect 6144 339 6178 361
rect 6144 293 6178 301
rect 6144 267 6178 293
rect 6240 1211 6274 1237
rect 6240 1203 6274 1211
rect 6240 1143 6274 1165
rect 6240 1131 6274 1143
rect 6240 1075 6274 1093
rect 6240 1059 6274 1075
rect 6240 1007 6274 1021
rect 6240 987 6274 1007
rect 6240 939 6274 949
rect 6240 915 6274 939
rect 6240 871 6274 877
rect 6240 843 6274 871
rect 6240 803 6274 805
rect 6240 771 6274 803
rect 6240 701 6274 733
rect 6240 699 6274 701
rect 6240 633 6274 661
rect 6240 627 6274 633
rect 6240 565 6274 589
rect 6240 555 6274 565
rect 6240 497 6274 517
rect 6240 483 6274 497
rect 6240 429 6274 445
rect 6240 411 6274 429
rect 6240 361 6274 373
rect 6240 339 6274 361
rect 6240 293 6274 301
rect 6240 267 6274 293
rect 6336 1211 6370 1237
rect 6336 1203 6370 1211
rect 6336 1143 6370 1165
rect 6336 1131 6370 1143
rect 6336 1075 6370 1093
rect 6336 1059 6370 1075
rect 6336 1007 6370 1021
rect 6336 987 6370 1007
rect 6336 939 6370 949
rect 6336 915 6370 939
rect 6336 871 6370 877
rect 6336 843 6370 871
rect 6336 803 6370 805
rect 6336 771 6370 803
rect 6336 701 6370 733
rect 6336 699 6370 701
rect 6336 633 6370 661
rect 6336 627 6370 633
rect 6336 565 6370 589
rect 6336 555 6370 565
rect 6336 497 6370 517
rect 6336 483 6370 497
rect 6336 429 6370 445
rect 6336 411 6370 429
rect 6336 361 6370 373
rect 6336 339 6370 361
rect 6336 293 6370 301
rect 6336 267 6370 293
rect 6432 1211 6466 1237
rect 6432 1203 6466 1211
rect 6432 1143 6466 1165
rect 6432 1131 6466 1143
rect 6432 1075 6466 1093
rect 6432 1059 6466 1075
rect 6432 1007 6466 1021
rect 6432 987 6466 1007
rect 6432 939 6466 949
rect 6432 915 6466 939
rect 6432 871 6466 877
rect 6432 843 6466 871
rect 6432 803 6466 805
rect 6432 771 6466 803
rect 6432 701 6466 733
rect 6432 699 6466 701
rect 6432 633 6466 661
rect 6432 627 6466 633
rect 6432 565 6466 589
rect 6432 555 6466 565
rect 6432 497 6466 517
rect 6432 483 6466 497
rect 6432 429 6466 445
rect 6432 411 6466 429
rect 6432 361 6466 373
rect 6432 339 6466 361
rect 6432 293 6466 301
rect 6432 267 6466 293
rect 6528 1211 6562 1237
rect 6528 1203 6562 1211
rect 6528 1143 6562 1165
rect 6528 1131 6562 1143
rect 6528 1075 6562 1093
rect 6528 1059 6562 1075
rect 6528 1007 6562 1021
rect 6528 987 6562 1007
rect 6528 939 6562 949
rect 6528 915 6562 939
rect 6528 871 6562 877
rect 6528 843 6562 871
rect 6528 803 6562 805
rect 6528 771 6562 803
rect 6528 701 6562 733
rect 6528 699 6562 701
rect 6528 633 6562 661
rect 6528 627 6562 633
rect 6528 565 6562 589
rect 6528 555 6562 565
rect 6528 497 6562 517
rect 6528 483 6562 497
rect 6528 429 6562 445
rect 6528 411 6562 429
rect 6528 361 6562 373
rect 6528 339 6562 361
rect 6528 293 6562 301
rect 6528 267 6562 293
rect 6624 1211 6658 1237
rect 6624 1203 6658 1211
rect 6624 1143 6658 1165
rect 6624 1131 6658 1143
rect 6624 1075 6658 1093
rect 6624 1059 6658 1075
rect 6624 1007 6658 1021
rect 6624 987 6658 1007
rect 6624 939 6658 949
rect 6624 915 6658 939
rect 6624 871 6658 877
rect 6624 843 6658 871
rect 6624 803 6658 805
rect 6624 771 6658 803
rect 6624 701 6658 733
rect 6624 699 6658 701
rect 6624 633 6658 661
rect 6624 627 6658 633
rect 6624 565 6658 589
rect 6624 555 6658 565
rect 6624 497 6658 517
rect 6624 483 6658 497
rect 6624 429 6658 445
rect 6624 411 6658 429
rect 6624 361 6658 373
rect 6624 339 6658 361
rect 6624 293 6658 301
rect 6624 267 6658 293
rect 6720 1211 6754 1237
rect 6720 1203 6754 1211
rect 6720 1143 6754 1165
rect 6720 1131 6754 1143
rect 6720 1075 6754 1093
rect 6720 1059 6754 1075
rect 6720 1007 6754 1021
rect 6720 987 6754 1007
rect 6720 939 6754 949
rect 6720 915 6754 939
rect 6720 871 6754 877
rect 6720 843 6754 871
rect 6720 803 6754 805
rect 6720 771 6754 803
rect 6720 701 6754 733
rect 6720 699 6754 701
rect 6720 633 6754 661
rect 6720 627 6754 633
rect 6720 565 6754 589
rect 6720 555 6754 565
rect 6720 497 6754 517
rect 6720 483 6754 497
rect 6720 429 6754 445
rect 6720 411 6754 429
rect 6720 361 6754 373
rect 6720 339 6754 361
rect 6720 293 6754 301
rect 6720 267 6754 293
rect 6816 1211 6850 1237
rect 6816 1203 6850 1211
rect 6816 1143 6850 1165
rect 6816 1131 6850 1143
rect 6816 1075 6850 1093
rect 6816 1059 6850 1075
rect 6816 1007 6850 1021
rect 6816 987 6850 1007
rect 6816 939 6850 949
rect 6816 915 6850 939
rect 6816 871 6850 877
rect 6816 843 6850 871
rect 6816 803 6850 805
rect 6816 771 6850 803
rect 6816 701 6850 733
rect 6816 699 6850 701
rect 6816 633 6850 661
rect 6816 627 6850 633
rect 6816 565 6850 589
rect 6816 555 6850 565
rect 6816 497 6850 517
rect 6816 483 6850 497
rect 6816 429 6850 445
rect 6816 411 6850 429
rect 6816 361 6850 373
rect 6816 339 6850 361
rect 6816 293 6850 301
rect 6816 267 6850 293
rect 6912 1211 6946 1237
rect 6912 1203 6946 1211
rect 6912 1143 6946 1165
rect 6912 1131 6946 1143
rect 6912 1075 6946 1093
rect 6912 1059 6946 1075
rect 6912 1007 6946 1021
rect 6912 987 6946 1007
rect 6912 939 6946 949
rect 6912 915 6946 939
rect 6912 871 6946 877
rect 6912 843 6946 871
rect 6912 803 6946 805
rect 6912 771 6946 803
rect 6912 701 6946 733
rect 6912 699 6946 701
rect 6912 633 6946 661
rect 6912 627 6946 633
rect 6912 565 6946 589
rect 6912 555 6946 565
rect 6912 497 6946 517
rect 6912 483 6946 497
rect 6912 429 6946 445
rect 6912 411 6946 429
rect 6912 361 6946 373
rect 6912 339 6946 361
rect 6912 293 6946 301
rect 6912 267 6946 293
rect 7008 1211 7042 1237
rect 7008 1203 7042 1211
rect 7008 1143 7042 1165
rect 7008 1131 7042 1143
rect 7008 1075 7042 1093
rect 7008 1059 7042 1075
rect 7008 1007 7042 1021
rect 7008 987 7042 1007
rect 7008 939 7042 949
rect 7008 915 7042 939
rect 7008 871 7042 877
rect 7008 843 7042 871
rect 7008 803 7042 805
rect 7008 771 7042 803
rect 7008 701 7042 733
rect 7008 699 7042 701
rect 7008 633 7042 661
rect 7008 627 7042 633
rect 7008 565 7042 589
rect 7008 555 7042 565
rect 7008 497 7042 517
rect 7008 483 7042 497
rect 7008 429 7042 445
rect 7008 411 7042 429
rect 7008 361 7042 373
rect 7008 339 7042 361
rect 7008 293 7042 301
rect 7008 267 7042 293
rect 7104 1211 7138 1237
rect 7104 1203 7138 1211
rect 7104 1143 7138 1165
rect 7104 1131 7138 1143
rect 7104 1075 7138 1093
rect 7104 1059 7138 1075
rect 7104 1007 7138 1021
rect 7104 987 7138 1007
rect 7104 939 7138 949
rect 7104 915 7138 939
rect 7104 871 7138 877
rect 7104 843 7138 871
rect 7104 803 7138 805
rect 7104 771 7138 803
rect 7104 701 7138 733
rect 7104 699 7138 701
rect 7104 633 7138 661
rect 7104 627 7138 633
rect 7104 565 7138 589
rect 7104 555 7138 565
rect 7104 497 7138 517
rect 7104 483 7138 497
rect 7104 429 7138 445
rect 7104 411 7138 429
rect 7104 361 7138 373
rect 7104 339 7138 361
rect 7104 293 7138 301
rect 7104 267 7138 293
rect 7200 1211 7234 1237
rect 7200 1203 7234 1211
rect 7200 1143 7234 1165
rect 7200 1131 7234 1143
rect 7200 1075 7234 1093
rect 7200 1059 7234 1075
rect 7200 1007 7234 1021
rect 7200 987 7234 1007
rect 7200 939 7234 949
rect 7200 915 7234 939
rect 7200 871 7234 877
rect 7200 843 7234 871
rect 7200 803 7234 805
rect 7200 771 7234 803
rect 7200 701 7234 733
rect 7200 699 7234 701
rect 7200 633 7234 661
rect 7200 627 7234 633
rect 7200 565 7234 589
rect 7200 555 7234 565
rect 7200 497 7234 517
rect 7200 483 7234 497
rect 7200 429 7234 445
rect 7200 411 7234 429
rect 7200 361 7234 373
rect 7200 339 7234 361
rect 7200 293 7234 301
rect 7200 267 7234 293
rect 7296 1211 7330 1237
rect 7296 1203 7330 1211
rect 7296 1143 7330 1165
rect 7296 1131 7330 1143
rect 7296 1075 7330 1093
rect 7296 1059 7330 1075
rect 7296 1007 7330 1021
rect 7296 987 7330 1007
rect 7296 939 7330 949
rect 7296 915 7330 939
rect 7296 871 7330 877
rect 7296 843 7330 871
rect 7296 803 7330 805
rect 7296 771 7330 803
rect 7296 701 7330 733
rect 7296 699 7330 701
rect 7296 633 7330 661
rect 7296 627 7330 633
rect 7296 565 7330 589
rect 7296 555 7330 565
rect 7296 497 7330 517
rect 7296 483 7330 497
rect 7296 429 7330 445
rect 7296 411 7330 429
rect 7296 361 7330 373
rect 7296 339 7330 361
rect 7296 293 7330 301
rect 7296 267 7330 293
rect 5450 96 5484 130
rect 5744 80 5778 114
rect 6142 80 6176 114
rect 6816 70 6850 104
rect 8386 1402 8420 1436
rect 9808 1406 9842 1440
rect 7912 1211 7946 1237
rect 7912 1203 7946 1211
rect 7912 1143 7946 1165
rect 7912 1131 7946 1143
rect 7912 1075 7946 1093
rect 7912 1059 7946 1075
rect 7912 1007 7946 1021
rect 7912 987 7946 1007
rect 7912 939 7946 949
rect 7912 915 7946 939
rect 7912 871 7946 877
rect 7912 843 7946 871
rect 7912 803 7946 805
rect 7912 771 7946 803
rect 7912 701 7946 733
rect 7912 699 7946 701
rect 7912 633 7946 661
rect 7912 627 7946 633
rect 7912 565 7946 589
rect 7912 555 7946 565
rect 7912 497 7946 517
rect 7912 483 7946 497
rect 7912 429 7946 445
rect 7912 411 7946 429
rect 7912 361 7946 373
rect 7912 339 7946 361
rect 7912 293 7946 301
rect 7912 267 7946 293
rect 8008 1211 8042 1237
rect 8008 1203 8042 1211
rect 8008 1143 8042 1165
rect 8008 1131 8042 1143
rect 8008 1075 8042 1093
rect 8008 1059 8042 1075
rect 8008 1007 8042 1021
rect 8008 987 8042 1007
rect 8008 939 8042 949
rect 8008 915 8042 939
rect 8008 871 8042 877
rect 8008 843 8042 871
rect 8008 803 8042 805
rect 8008 771 8042 803
rect 8008 701 8042 733
rect 8008 699 8042 701
rect 8008 633 8042 661
rect 8008 627 8042 633
rect 8008 565 8042 589
rect 8008 555 8042 565
rect 8008 497 8042 517
rect 8008 483 8042 497
rect 8008 429 8042 445
rect 8008 411 8042 429
rect 8008 361 8042 373
rect 8008 339 8042 361
rect 8008 293 8042 301
rect 8008 267 8042 293
rect 8104 1211 8138 1237
rect 8104 1203 8138 1211
rect 8104 1143 8138 1165
rect 8104 1131 8138 1143
rect 8104 1075 8138 1093
rect 8104 1059 8138 1075
rect 8104 1007 8138 1021
rect 8104 987 8138 1007
rect 8104 939 8138 949
rect 8104 915 8138 939
rect 8104 871 8138 877
rect 8104 843 8138 871
rect 8104 803 8138 805
rect 8104 771 8138 803
rect 8104 701 8138 733
rect 8104 699 8138 701
rect 8104 633 8138 661
rect 8104 627 8138 633
rect 8104 565 8138 589
rect 8104 555 8138 565
rect 8104 497 8138 517
rect 8104 483 8138 497
rect 8104 429 8138 445
rect 8104 411 8138 429
rect 8104 361 8138 373
rect 8104 339 8138 361
rect 8104 293 8138 301
rect 8104 267 8138 293
rect 8200 1211 8234 1237
rect 8200 1203 8234 1211
rect 8200 1143 8234 1165
rect 8200 1131 8234 1143
rect 8200 1075 8234 1093
rect 8200 1059 8234 1075
rect 8200 1007 8234 1021
rect 8200 987 8234 1007
rect 8200 939 8234 949
rect 8200 915 8234 939
rect 8200 871 8234 877
rect 8200 843 8234 871
rect 8200 803 8234 805
rect 8200 771 8234 803
rect 8200 701 8234 733
rect 8200 699 8234 701
rect 8200 633 8234 661
rect 8200 627 8234 633
rect 8200 565 8234 589
rect 8200 555 8234 565
rect 8200 497 8234 517
rect 8200 483 8234 497
rect 8200 429 8234 445
rect 8200 411 8234 429
rect 8200 361 8234 373
rect 8200 339 8234 361
rect 8200 293 8234 301
rect 8200 267 8234 293
rect 8296 1211 8330 1237
rect 8296 1203 8330 1211
rect 8296 1143 8330 1165
rect 8296 1131 8330 1143
rect 8296 1075 8330 1093
rect 8296 1059 8330 1075
rect 8296 1007 8330 1021
rect 8296 987 8330 1007
rect 8296 939 8330 949
rect 8296 915 8330 939
rect 8296 871 8330 877
rect 8296 843 8330 871
rect 8296 803 8330 805
rect 8296 771 8330 803
rect 8296 701 8330 733
rect 8296 699 8330 701
rect 8296 633 8330 661
rect 8296 627 8330 633
rect 8296 565 8330 589
rect 8296 555 8330 565
rect 8296 497 8330 517
rect 8296 483 8330 497
rect 8296 429 8330 445
rect 8296 411 8330 429
rect 8296 361 8330 373
rect 8296 339 8330 361
rect 8296 293 8330 301
rect 8296 267 8330 293
rect 8392 1211 8426 1237
rect 8392 1203 8426 1211
rect 8392 1143 8426 1165
rect 8392 1131 8426 1143
rect 8392 1075 8426 1093
rect 8392 1059 8426 1075
rect 8392 1007 8426 1021
rect 8392 987 8426 1007
rect 8392 939 8426 949
rect 8392 915 8426 939
rect 8392 871 8426 877
rect 8392 843 8426 871
rect 8392 803 8426 805
rect 8392 771 8426 803
rect 8392 701 8426 733
rect 8392 699 8426 701
rect 8392 633 8426 661
rect 8392 627 8426 633
rect 8392 565 8426 589
rect 8392 555 8426 565
rect 8392 497 8426 517
rect 8392 483 8426 497
rect 8392 429 8426 445
rect 8392 411 8426 429
rect 8392 361 8426 373
rect 8392 339 8426 361
rect 8392 293 8426 301
rect 8392 267 8426 293
rect 8488 1211 8522 1237
rect 8488 1203 8522 1211
rect 8488 1143 8522 1165
rect 8488 1131 8522 1143
rect 8488 1075 8522 1093
rect 8488 1059 8522 1075
rect 8488 1007 8522 1021
rect 8488 987 8522 1007
rect 8488 939 8522 949
rect 8488 915 8522 939
rect 8488 871 8522 877
rect 8488 843 8522 871
rect 8488 803 8522 805
rect 8488 771 8522 803
rect 8488 701 8522 733
rect 8488 699 8522 701
rect 8488 633 8522 661
rect 8488 627 8522 633
rect 8488 565 8522 589
rect 8488 555 8522 565
rect 8488 497 8522 517
rect 8488 483 8522 497
rect 8488 429 8522 445
rect 8488 411 8522 429
rect 8488 361 8522 373
rect 8488 339 8522 361
rect 8488 293 8522 301
rect 8488 267 8522 293
rect 8584 1211 8618 1237
rect 8584 1203 8618 1211
rect 8584 1143 8618 1165
rect 8584 1131 8618 1143
rect 8584 1075 8618 1093
rect 8584 1059 8618 1075
rect 8584 1007 8618 1021
rect 8584 987 8618 1007
rect 8584 939 8618 949
rect 8584 915 8618 939
rect 8584 871 8618 877
rect 8584 843 8618 871
rect 8584 803 8618 805
rect 8584 771 8618 803
rect 8584 701 8618 733
rect 8584 699 8618 701
rect 8584 633 8618 661
rect 8584 627 8618 633
rect 8584 565 8618 589
rect 8584 555 8618 565
rect 8584 497 8618 517
rect 8584 483 8618 497
rect 8584 429 8618 445
rect 8584 411 8618 429
rect 8584 361 8618 373
rect 8584 339 8618 361
rect 8584 293 8618 301
rect 8584 267 8618 293
rect 8680 1211 8714 1237
rect 8680 1203 8714 1211
rect 8680 1143 8714 1165
rect 8680 1131 8714 1143
rect 8680 1075 8714 1093
rect 8680 1059 8714 1075
rect 8680 1007 8714 1021
rect 8680 987 8714 1007
rect 8680 939 8714 949
rect 8680 915 8714 939
rect 8680 871 8714 877
rect 8680 843 8714 871
rect 8680 803 8714 805
rect 8680 771 8714 803
rect 8680 701 8714 733
rect 8680 699 8714 701
rect 8680 633 8714 661
rect 8680 627 8714 633
rect 8680 565 8714 589
rect 8680 555 8714 565
rect 8680 497 8714 517
rect 8680 483 8714 497
rect 8680 429 8714 445
rect 8680 411 8714 429
rect 8680 361 8714 373
rect 8680 339 8714 361
rect 8680 293 8714 301
rect 8680 267 8714 293
rect 8776 1211 8810 1237
rect 8776 1203 8810 1211
rect 8776 1143 8810 1165
rect 8776 1131 8810 1143
rect 8776 1075 8810 1093
rect 8776 1059 8810 1075
rect 8776 1007 8810 1021
rect 8776 987 8810 1007
rect 8776 939 8810 949
rect 8776 915 8810 939
rect 8776 871 8810 877
rect 8776 843 8810 871
rect 8776 803 8810 805
rect 8776 771 8810 803
rect 8776 701 8810 733
rect 8776 699 8810 701
rect 8776 633 8810 661
rect 8776 627 8810 633
rect 8776 565 8810 589
rect 8776 555 8810 565
rect 8776 497 8810 517
rect 8776 483 8810 497
rect 8776 429 8810 445
rect 8776 411 8810 429
rect 8776 361 8810 373
rect 8776 339 8810 361
rect 8776 293 8810 301
rect 8776 267 8810 293
rect 8872 1211 8906 1237
rect 8872 1203 8906 1211
rect 8872 1143 8906 1165
rect 8872 1131 8906 1143
rect 8872 1075 8906 1093
rect 8872 1059 8906 1075
rect 8872 1007 8906 1021
rect 8872 987 8906 1007
rect 8872 939 8906 949
rect 8872 915 8906 939
rect 8872 871 8906 877
rect 8872 843 8906 871
rect 8872 803 8906 805
rect 8872 771 8906 803
rect 8872 701 8906 733
rect 8872 699 8906 701
rect 8872 633 8906 661
rect 8872 627 8906 633
rect 8872 565 8906 589
rect 8872 555 8906 565
rect 8872 497 8906 517
rect 8872 483 8906 497
rect 8872 429 8906 445
rect 8872 411 8906 429
rect 8872 361 8906 373
rect 8872 339 8906 361
rect 8872 293 8906 301
rect 8872 267 8906 293
rect 8968 1211 9002 1237
rect 8968 1203 9002 1211
rect 8968 1143 9002 1165
rect 8968 1131 9002 1143
rect 8968 1075 9002 1093
rect 8968 1059 9002 1075
rect 8968 1007 9002 1021
rect 8968 987 9002 1007
rect 8968 939 9002 949
rect 8968 915 9002 939
rect 8968 871 9002 877
rect 8968 843 9002 871
rect 8968 803 9002 805
rect 8968 771 9002 803
rect 8968 701 9002 733
rect 8968 699 9002 701
rect 8968 633 9002 661
rect 8968 627 9002 633
rect 8968 565 9002 589
rect 8968 555 9002 565
rect 8968 497 9002 517
rect 8968 483 9002 497
rect 8968 429 9002 445
rect 8968 411 9002 429
rect 8968 361 9002 373
rect 8968 339 9002 361
rect 8968 293 9002 301
rect 8968 267 9002 293
rect 9232 1209 9266 1235
rect 9232 1201 9266 1209
rect 9232 1141 9266 1163
rect 9232 1129 9266 1141
rect 9232 1073 9266 1091
rect 9232 1057 9266 1073
rect 9232 1005 9266 1019
rect 9232 985 9266 1005
rect 9232 937 9266 947
rect 9232 913 9266 937
rect 9232 869 9266 875
rect 9232 841 9266 869
rect 9232 801 9266 803
rect 9232 769 9266 801
rect 9232 699 9266 731
rect 9232 697 9266 699
rect 9232 631 9266 659
rect 9232 625 9266 631
rect 9232 563 9266 587
rect 9232 553 9266 563
rect 9232 495 9266 515
rect 9232 481 9266 495
rect 9232 427 9266 443
rect 9232 409 9266 427
rect 9232 359 9266 371
rect 9232 337 9266 359
rect 9232 291 9266 299
rect 9232 265 9266 291
rect 9328 1209 9362 1235
rect 9328 1201 9362 1209
rect 9328 1141 9362 1163
rect 9328 1129 9362 1141
rect 9328 1073 9362 1091
rect 9328 1057 9362 1073
rect 9328 1005 9362 1019
rect 9328 985 9362 1005
rect 9328 937 9362 947
rect 9328 913 9362 937
rect 9328 869 9362 875
rect 9328 841 9362 869
rect 9328 801 9362 803
rect 9328 769 9362 801
rect 9328 699 9362 731
rect 9328 697 9362 699
rect 9328 631 9362 659
rect 9328 625 9362 631
rect 9328 563 9362 587
rect 9328 553 9362 563
rect 9328 495 9362 515
rect 9328 481 9362 495
rect 9328 427 9362 443
rect 9328 409 9362 427
rect 9328 359 9362 371
rect 9328 337 9362 359
rect 9328 291 9362 299
rect 9328 265 9362 291
rect 9424 1209 9458 1235
rect 9424 1201 9458 1209
rect 9424 1141 9458 1163
rect 9424 1129 9458 1141
rect 9424 1073 9458 1091
rect 9424 1057 9458 1073
rect 9424 1005 9458 1019
rect 9424 985 9458 1005
rect 9424 937 9458 947
rect 9424 913 9458 937
rect 9424 869 9458 875
rect 9424 841 9458 869
rect 9424 801 9458 803
rect 9424 769 9458 801
rect 9424 699 9458 731
rect 9424 697 9458 699
rect 9424 631 9458 659
rect 9424 625 9458 631
rect 9424 563 9458 587
rect 9424 553 9458 563
rect 9424 495 9458 515
rect 9424 481 9458 495
rect 9424 427 9458 443
rect 9424 409 9458 427
rect 9424 359 9458 371
rect 9424 337 9458 359
rect 9424 291 9458 299
rect 9424 265 9458 291
rect 9520 1209 9554 1235
rect 9520 1201 9554 1209
rect 9520 1141 9554 1163
rect 9520 1129 9554 1141
rect 9520 1073 9554 1091
rect 9520 1057 9554 1073
rect 9520 1005 9554 1019
rect 9520 985 9554 1005
rect 9520 937 9554 947
rect 9520 913 9554 937
rect 9520 869 9554 875
rect 9520 841 9554 869
rect 9520 801 9554 803
rect 9520 769 9554 801
rect 9520 699 9554 731
rect 9520 697 9554 699
rect 9520 631 9554 659
rect 9520 625 9554 631
rect 9520 563 9554 587
rect 9520 553 9554 563
rect 9520 495 9554 515
rect 9520 481 9554 495
rect 9520 427 9554 443
rect 9520 409 9554 427
rect 9520 359 9554 371
rect 9520 337 9554 359
rect 9520 291 9554 299
rect 9520 265 9554 291
rect 9616 1209 9650 1235
rect 9616 1201 9650 1209
rect 9616 1141 9650 1163
rect 9616 1129 9650 1141
rect 9616 1073 9650 1091
rect 9616 1057 9650 1073
rect 9616 1005 9650 1019
rect 9616 985 9650 1005
rect 9616 937 9650 947
rect 9616 913 9650 937
rect 9616 869 9650 875
rect 9616 841 9650 869
rect 9616 801 9650 803
rect 9616 769 9650 801
rect 9616 699 9650 731
rect 9616 697 9650 699
rect 9616 631 9650 659
rect 9616 625 9650 631
rect 9616 563 9650 587
rect 9616 553 9650 563
rect 9616 495 9650 515
rect 9616 481 9650 495
rect 9616 427 9650 443
rect 9616 409 9650 427
rect 9616 359 9650 371
rect 9616 337 9650 359
rect 9616 291 9650 299
rect 9616 265 9650 291
rect 9712 1209 9746 1235
rect 9712 1201 9746 1209
rect 9712 1141 9746 1163
rect 9712 1129 9746 1141
rect 9712 1073 9746 1091
rect 9712 1057 9746 1073
rect 9712 1005 9746 1019
rect 9712 985 9746 1005
rect 9712 937 9746 947
rect 9712 913 9746 937
rect 9712 869 9746 875
rect 9712 841 9746 869
rect 9712 801 9746 803
rect 9712 769 9746 801
rect 9712 699 9746 731
rect 9712 697 9746 699
rect 9712 631 9746 659
rect 9712 625 9746 631
rect 9712 563 9746 587
rect 9712 553 9746 563
rect 9712 495 9746 515
rect 9712 481 9746 495
rect 9712 427 9746 443
rect 9712 409 9746 427
rect 9712 359 9746 371
rect 9712 337 9746 359
rect 9712 291 9746 299
rect 9712 265 9746 291
rect 9808 1209 9842 1235
rect 9808 1201 9842 1209
rect 9808 1141 9842 1163
rect 9808 1129 9842 1141
rect 9808 1073 9842 1091
rect 9808 1057 9842 1073
rect 9808 1005 9842 1019
rect 9808 985 9842 1005
rect 9808 937 9842 947
rect 9808 913 9842 937
rect 9808 869 9842 875
rect 9808 841 9842 869
rect 9808 801 9842 803
rect 9808 769 9842 801
rect 9808 699 9842 731
rect 9808 697 9842 699
rect 9808 631 9842 659
rect 9808 625 9842 631
rect 9808 563 9842 587
rect 9808 553 9842 563
rect 9808 495 9842 515
rect 9808 481 9842 495
rect 9808 427 9842 443
rect 9808 409 9842 427
rect 9808 359 9842 371
rect 9808 337 9842 359
rect 9808 291 9842 299
rect 9808 265 9842 291
rect 9904 1209 9938 1235
rect 9904 1201 9938 1209
rect 9904 1141 9938 1163
rect 9904 1129 9938 1141
rect 9904 1073 9938 1091
rect 9904 1057 9938 1073
rect 9904 1005 9938 1019
rect 9904 985 9938 1005
rect 9904 937 9938 947
rect 9904 913 9938 937
rect 9904 869 9938 875
rect 9904 841 9938 869
rect 9904 801 9938 803
rect 9904 769 9938 801
rect 9904 699 9938 731
rect 9904 697 9938 699
rect 9904 631 9938 659
rect 9904 625 9938 631
rect 9904 563 9938 587
rect 9904 553 9938 563
rect 9904 495 9938 515
rect 9904 481 9938 495
rect 9904 427 9938 443
rect 9904 409 9938 427
rect 9904 359 9938 371
rect 9904 337 9938 359
rect 9904 291 9938 299
rect 9904 265 9938 291
rect 10000 1209 10034 1235
rect 10000 1201 10034 1209
rect 10000 1141 10034 1163
rect 10000 1129 10034 1141
rect 10000 1073 10034 1091
rect 10000 1057 10034 1073
rect 10000 1005 10034 1019
rect 10000 985 10034 1005
rect 10000 937 10034 947
rect 10000 913 10034 937
rect 10000 869 10034 875
rect 10000 841 10034 869
rect 10000 801 10034 803
rect 10000 769 10034 801
rect 10000 699 10034 731
rect 10000 697 10034 699
rect 10000 631 10034 659
rect 10000 625 10034 631
rect 10000 563 10034 587
rect 10000 553 10034 563
rect 10000 495 10034 515
rect 10000 481 10034 495
rect 10000 427 10034 443
rect 10000 409 10034 427
rect 10000 359 10034 371
rect 10000 337 10034 359
rect 10000 291 10034 299
rect 10000 265 10034 291
rect 10096 1209 10130 1235
rect 10096 1201 10130 1209
rect 10096 1141 10130 1163
rect 10096 1129 10130 1141
rect 10096 1073 10130 1091
rect 10096 1057 10130 1073
rect 10096 1005 10130 1019
rect 10096 985 10130 1005
rect 10096 937 10130 947
rect 10096 913 10130 937
rect 10096 869 10130 875
rect 10096 841 10130 869
rect 10096 801 10130 803
rect 10096 769 10130 801
rect 10096 699 10130 731
rect 10096 697 10130 699
rect 10096 631 10130 659
rect 10096 625 10130 631
rect 10096 563 10130 587
rect 10096 553 10130 563
rect 10096 495 10130 515
rect 10096 481 10130 495
rect 10096 427 10130 443
rect 10096 409 10130 427
rect 10096 359 10130 371
rect 10096 337 10130 359
rect 10096 291 10130 299
rect 10096 265 10130 291
rect 10192 1209 10226 1235
rect 10192 1201 10226 1209
rect 10192 1141 10226 1163
rect 10192 1129 10226 1141
rect 10192 1073 10226 1091
rect 10192 1057 10226 1073
rect 10192 1005 10226 1019
rect 10192 985 10226 1005
rect 10192 937 10226 947
rect 10192 913 10226 937
rect 10192 869 10226 875
rect 10192 841 10226 869
rect 10192 801 10226 803
rect 10192 769 10226 801
rect 10192 699 10226 731
rect 10192 697 10226 699
rect 10192 631 10226 659
rect 10192 625 10226 631
rect 10192 563 10226 587
rect 10192 553 10226 563
rect 10192 495 10226 515
rect 10192 481 10226 495
rect 10192 427 10226 443
rect 10192 409 10226 427
rect 10192 359 10226 371
rect 10192 337 10226 359
rect 10192 291 10226 299
rect 10192 265 10226 291
rect 10288 1209 10322 1235
rect 10288 1201 10322 1209
rect 10288 1141 10322 1163
rect 10288 1129 10322 1141
rect 10288 1073 10322 1091
rect 10288 1057 10322 1073
rect 10288 1005 10322 1019
rect 10288 985 10322 1005
rect 10288 937 10322 947
rect 10288 913 10322 937
rect 10288 869 10322 875
rect 10288 841 10322 869
rect 10288 801 10322 803
rect 10288 769 10322 801
rect 10288 699 10322 731
rect 10288 697 10322 699
rect 10288 631 10322 659
rect 10288 625 10322 631
rect 10288 563 10322 587
rect 10288 553 10322 563
rect 10288 495 10322 515
rect 10288 481 10322 495
rect 10288 427 10322 443
rect 10288 409 10322 427
rect 10288 359 10322 371
rect 10288 337 10322 359
rect 10288 291 10322 299
rect 10288 265 10322 291
rect 10384 1209 10418 1235
rect 10384 1201 10418 1209
rect 10384 1141 10418 1163
rect 10384 1129 10418 1141
rect 10384 1073 10418 1091
rect 10384 1057 10418 1073
rect 10384 1005 10418 1019
rect 10384 985 10418 1005
rect 10384 937 10418 947
rect 10384 913 10418 937
rect 10384 869 10418 875
rect 10384 841 10418 869
rect 10384 801 10418 803
rect 10384 769 10418 801
rect 10384 699 10418 731
rect 10384 697 10418 699
rect 10384 631 10418 659
rect 10384 625 10418 631
rect 10384 563 10418 587
rect 10384 553 10418 563
rect 10384 495 10418 515
rect 10384 481 10418 495
rect 10384 427 10418 443
rect 10384 409 10418 427
rect 10384 359 10418 371
rect 10384 337 10418 359
rect 10384 291 10418 299
rect 10384 265 10418 291
rect 8480 96 8514 130
rect 8774 80 8808 114
rect 9230 78 9264 112
rect 9904 68 9938 102
rect 4665 -21 4699 13
rect 7665 -19 7699 15
rect 15466 1458 15500 1492
rect 11474 1400 11508 1434
rect 12964 1380 12998 1414
rect 11000 1209 11034 1235
rect 11000 1201 11034 1209
rect 11000 1141 11034 1163
rect 11000 1129 11034 1141
rect 11000 1073 11034 1091
rect 11000 1057 11034 1073
rect 11000 1005 11034 1019
rect 11000 985 11034 1005
rect 11000 937 11034 947
rect 11000 913 11034 937
rect 11000 869 11034 875
rect 11000 841 11034 869
rect 11000 801 11034 803
rect 11000 769 11034 801
rect 11000 699 11034 731
rect 11000 697 11034 699
rect 11000 631 11034 659
rect 11000 625 11034 631
rect 11000 563 11034 587
rect 11000 553 11034 563
rect 11000 495 11034 515
rect 11000 481 11034 495
rect 11000 427 11034 443
rect 11000 409 11034 427
rect 11000 359 11034 371
rect 11000 337 11034 359
rect 11000 291 11034 299
rect 11000 265 11034 291
rect 11096 1209 11130 1235
rect 11096 1201 11130 1209
rect 11096 1141 11130 1163
rect 11096 1129 11130 1141
rect 11096 1073 11130 1091
rect 11096 1057 11130 1073
rect 11096 1005 11130 1019
rect 11096 985 11130 1005
rect 11096 937 11130 947
rect 11096 913 11130 937
rect 11096 869 11130 875
rect 11096 841 11130 869
rect 11096 801 11130 803
rect 11096 769 11130 801
rect 11096 699 11130 731
rect 11096 697 11130 699
rect 11096 631 11130 659
rect 11096 625 11130 631
rect 11096 563 11130 587
rect 11096 553 11130 563
rect 11096 495 11130 515
rect 11096 481 11130 495
rect 11096 427 11130 443
rect 11096 409 11130 427
rect 11096 359 11130 371
rect 11096 337 11130 359
rect 11096 291 11130 299
rect 11096 265 11130 291
rect 11192 1209 11226 1235
rect 11192 1201 11226 1209
rect 11192 1141 11226 1163
rect 11192 1129 11226 1141
rect 11192 1073 11226 1091
rect 11192 1057 11226 1073
rect 11192 1005 11226 1019
rect 11192 985 11226 1005
rect 11192 937 11226 947
rect 11192 913 11226 937
rect 11192 869 11226 875
rect 11192 841 11226 869
rect 11192 801 11226 803
rect 11192 769 11226 801
rect 11192 699 11226 731
rect 11192 697 11226 699
rect 11192 631 11226 659
rect 11192 625 11226 631
rect 11192 563 11226 587
rect 11192 553 11226 563
rect 11192 495 11226 515
rect 11192 481 11226 495
rect 11192 427 11226 443
rect 11192 409 11226 427
rect 11192 359 11226 371
rect 11192 337 11226 359
rect 11192 291 11226 299
rect 11192 265 11226 291
rect 11288 1209 11322 1235
rect 11288 1201 11322 1209
rect 11288 1141 11322 1163
rect 11288 1129 11322 1141
rect 11288 1073 11322 1091
rect 11288 1057 11322 1073
rect 11288 1005 11322 1019
rect 11288 985 11322 1005
rect 11288 937 11322 947
rect 11288 913 11322 937
rect 11288 869 11322 875
rect 11288 841 11322 869
rect 11288 801 11322 803
rect 11288 769 11322 801
rect 11288 699 11322 731
rect 11288 697 11322 699
rect 11288 631 11322 659
rect 11288 625 11322 631
rect 11288 563 11322 587
rect 11288 553 11322 563
rect 11288 495 11322 515
rect 11288 481 11322 495
rect 11288 427 11322 443
rect 11288 409 11322 427
rect 11288 359 11322 371
rect 11288 337 11322 359
rect 11288 291 11322 299
rect 11288 265 11322 291
rect 11384 1209 11418 1235
rect 11384 1201 11418 1209
rect 11384 1141 11418 1163
rect 11384 1129 11418 1141
rect 11384 1073 11418 1091
rect 11384 1057 11418 1073
rect 11384 1005 11418 1019
rect 11384 985 11418 1005
rect 11384 937 11418 947
rect 11384 913 11418 937
rect 11384 869 11418 875
rect 11384 841 11418 869
rect 11384 801 11418 803
rect 11384 769 11418 801
rect 11384 699 11418 731
rect 11384 697 11418 699
rect 11384 631 11418 659
rect 11384 625 11418 631
rect 11384 563 11418 587
rect 11384 553 11418 563
rect 11384 495 11418 515
rect 11384 481 11418 495
rect 11384 427 11418 443
rect 11384 409 11418 427
rect 11384 359 11418 371
rect 11384 337 11418 359
rect 11384 291 11418 299
rect 11384 265 11418 291
rect 11480 1209 11514 1235
rect 11480 1201 11514 1209
rect 11480 1141 11514 1163
rect 11480 1129 11514 1141
rect 11480 1073 11514 1091
rect 11480 1057 11514 1073
rect 11480 1005 11514 1019
rect 11480 985 11514 1005
rect 11480 937 11514 947
rect 11480 913 11514 937
rect 11480 869 11514 875
rect 11480 841 11514 869
rect 11480 801 11514 803
rect 11480 769 11514 801
rect 11480 699 11514 731
rect 11480 697 11514 699
rect 11480 631 11514 659
rect 11480 625 11514 631
rect 11480 563 11514 587
rect 11480 553 11514 563
rect 11480 495 11514 515
rect 11480 481 11514 495
rect 11480 427 11514 443
rect 11480 409 11514 427
rect 11480 359 11514 371
rect 11480 337 11514 359
rect 11480 291 11514 299
rect 11480 265 11514 291
rect 11576 1209 11610 1235
rect 11576 1201 11610 1209
rect 11576 1141 11610 1163
rect 11576 1129 11610 1141
rect 11576 1073 11610 1091
rect 11576 1057 11610 1073
rect 11576 1005 11610 1019
rect 11576 985 11610 1005
rect 11576 937 11610 947
rect 11576 913 11610 937
rect 11576 869 11610 875
rect 11576 841 11610 869
rect 11576 801 11610 803
rect 11576 769 11610 801
rect 11576 699 11610 731
rect 11576 697 11610 699
rect 11576 631 11610 659
rect 11576 625 11610 631
rect 11576 563 11610 587
rect 11576 553 11610 563
rect 11576 495 11610 515
rect 11576 481 11610 495
rect 11576 427 11610 443
rect 11576 409 11610 427
rect 11576 359 11610 371
rect 11576 337 11610 359
rect 11576 291 11610 299
rect 11576 265 11610 291
rect 11672 1209 11706 1235
rect 11672 1201 11706 1209
rect 11672 1141 11706 1163
rect 11672 1129 11706 1141
rect 11672 1073 11706 1091
rect 11672 1057 11706 1073
rect 11672 1005 11706 1019
rect 11672 985 11706 1005
rect 11672 937 11706 947
rect 11672 913 11706 937
rect 11672 869 11706 875
rect 11672 841 11706 869
rect 11672 801 11706 803
rect 11672 769 11706 801
rect 11672 699 11706 731
rect 11672 697 11706 699
rect 11672 631 11706 659
rect 11672 625 11706 631
rect 11672 563 11706 587
rect 11672 553 11706 563
rect 11672 495 11706 515
rect 11672 481 11706 495
rect 11672 427 11706 443
rect 11672 409 11706 427
rect 11672 359 11706 371
rect 11672 337 11706 359
rect 11672 291 11706 299
rect 11672 265 11706 291
rect 11768 1209 11802 1235
rect 11768 1201 11802 1209
rect 11768 1141 11802 1163
rect 11768 1129 11802 1141
rect 11768 1073 11802 1091
rect 11768 1057 11802 1073
rect 11768 1005 11802 1019
rect 11768 985 11802 1005
rect 11768 937 11802 947
rect 11768 913 11802 937
rect 11768 869 11802 875
rect 11768 841 11802 869
rect 11768 801 11802 803
rect 11768 769 11802 801
rect 11768 699 11802 731
rect 11768 697 11802 699
rect 11768 631 11802 659
rect 11768 625 11802 631
rect 11768 563 11802 587
rect 11768 553 11802 563
rect 11768 495 11802 515
rect 11768 481 11802 495
rect 11768 427 11802 443
rect 11768 409 11802 427
rect 11768 359 11802 371
rect 11768 337 11802 359
rect 11768 291 11802 299
rect 11768 265 11802 291
rect 11864 1209 11898 1235
rect 11864 1201 11898 1209
rect 11864 1141 11898 1163
rect 11864 1129 11898 1141
rect 11864 1073 11898 1091
rect 11864 1057 11898 1073
rect 11864 1005 11898 1019
rect 11864 985 11898 1005
rect 11864 937 11898 947
rect 11864 913 11898 937
rect 11864 869 11898 875
rect 11864 841 11898 869
rect 11864 801 11898 803
rect 11864 769 11898 801
rect 11864 699 11898 731
rect 11864 697 11898 699
rect 11864 631 11898 659
rect 11864 625 11898 631
rect 11864 563 11898 587
rect 11864 553 11898 563
rect 11864 495 11898 515
rect 11864 481 11898 495
rect 11864 427 11898 443
rect 11864 409 11898 427
rect 11864 359 11898 371
rect 11864 337 11898 359
rect 11864 291 11898 299
rect 11864 265 11898 291
rect 11960 1209 11994 1235
rect 11960 1201 11994 1209
rect 11960 1141 11994 1163
rect 11960 1129 11994 1141
rect 11960 1073 11994 1091
rect 11960 1057 11994 1073
rect 11960 1005 11994 1019
rect 11960 985 11994 1005
rect 11960 937 11994 947
rect 11960 913 11994 937
rect 11960 869 11994 875
rect 11960 841 11994 869
rect 11960 801 11994 803
rect 11960 769 11994 801
rect 11960 699 11994 731
rect 11960 697 11994 699
rect 11960 631 11994 659
rect 11960 625 11994 631
rect 11960 563 11994 587
rect 11960 553 11994 563
rect 11960 495 11994 515
rect 11960 481 11994 495
rect 11960 427 11994 443
rect 11960 409 11994 427
rect 11960 359 11994 371
rect 11960 337 11994 359
rect 11960 291 11994 299
rect 11960 265 11994 291
rect 12056 1209 12090 1235
rect 12056 1201 12090 1209
rect 12056 1141 12090 1163
rect 12056 1129 12090 1141
rect 12056 1073 12090 1091
rect 12056 1057 12090 1073
rect 12056 1005 12090 1019
rect 12056 985 12090 1005
rect 12056 937 12090 947
rect 12056 913 12090 937
rect 12056 869 12090 875
rect 12056 841 12090 869
rect 12056 801 12090 803
rect 12056 769 12090 801
rect 12056 699 12090 731
rect 12056 697 12090 699
rect 12056 631 12090 659
rect 12056 625 12090 631
rect 12056 563 12090 587
rect 12056 553 12090 563
rect 12056 495 12090 515
rect 12056 481 12090 495
rect 12056 427 12090 443
rect 12056 409 12090 427
rect 12056 359 12090 371
rect 12056 337 12090 359
rect 12056 291 12090 299
rect 12056 265 12090 291
rect 12388 1183 12422 1209
rect 12388 1175 12422 1183
rect 12388 1115 12422 1137
rect 12388 1103 12422 1115
rect 12388 1047 12422 1065
rect 12388 1031 12422 1047
rect 12388 979 12422 993
rect 12388 959 12422 979
rect 12388 911 12422 921
rect 12388 887 12422 911
rect 12388 843 12422 849
rect 12388 815 12422 843
rect 12388 775 12422 777
rect 12388 743 12422 775
rect 12388 673 12422 705
rect 12388 671 12422 673
rect 12388 605 12422 633
rect 12388 599 12422 605
rect 12388 537 12422 561
rect 12388 527 12422 537
rect 12388 469 12422 489
rect 12388 455 12422 469
rect 12388 401 12422 417
rect 12388 383 12422 401
rect 12388 333 12422 345
rect 12388 311 12422 333
rect 12388 265 12422 273
rect 12388 239 12422 265
rect 12484 1183 12518 1209
rect 12484 1175 12518 1183
rect 12484 1115 12518 1137
rect 12484 1103 12518 1115
rect 12484 1047 12518 1065
rect 12484 1031 12518 1047
rect 12484 979 12518 993
rect 12484 959 12518 979
rect 12484 911 12518 921
rect 12484 887 12518 911
rect 12484 843 12518 849
rect 12484 815 12518 843
rect 12484 775 12518 777
rect 12484 743 12518 775
rect 12484 673 12518 705
rect 12484 671 12518 673
rect 12484 605 12518 633
rect 12484 599 12518 605
rect 12484 537 12518 561
rect 12484 527 12518 537
rect 12484 469 12518 489
rect 12484 455 12518 469
rect 12484 401 12518 417
rect 12484 383 12518 401
rect 12484 333 12518 345
rect 12484 311 12518 333
rect 12484 265 12518 273
rect 12484 239 12518 265
rect 12580 1183 12614 1209
rect 12580 1175 12614 1183
rect 12580 1115 12614 1137
rect 12580 1103 12614 1115
rect 12580 1047 12614 1065
rect 12580 1031 12614 1047
rect 12580 979 12614 993
rect 12580 959 12614 979
rect 12580 911 12614 921
rect 12580 887 12614 911
rect 12580 843 12614 849
rect 12580 815 12614 843
rect 12580 775 12614 777
rect 12580 743 12614 775
rect 12580 673 12614 705
rect 12580 671 12614 673
rect 12580 605 12614 633
rect 12580 599 12614 605
rect 12580 537 12614 561
rect 12580 527 12614 537
rect 12580 469 12614 489
rect 12580 455 12614 469
rect 12580 401 12614 417
rect 12580 383 12614 401
rect 12580 333 12614 345
rect 12580 311 12614 333
rect 12580 265 12614 273
rect 12580 239 12614 265
rect 12676 1183 12710 1209
rect 12676 1175 12710 1183
rect 12676 1115 12710 1137
rect 12676 1103 12710 1115
rect 12676 1047 12710 1065
rect 12676 1031 12710 1047
rect 12676 979 12710 993
rect 12676 959 12710 979
rect 12676 911 12710 921
rect 12676 887 12710 911
rect 12676 843 12710 849
rect 12676 815 12710 843
rect 12676 775 12710 777
rect 12676 743 12710 775
rect 12676 673 12710 705
rect 12676 671 12710 673
rect 12676 605 12710 633
rect 12676 599 12710 605
rect 12676 537 12710 561
rect 12676 527 12710 537
rect 12676 469 12710 489
rect 12676 455 12710 469
rect 12676 401 12710 417
rect 12676 383 12710 401
rect 12676 333 12710 345
rect 12676 311 12710 333
rect 12676 265 12710 273
rect 12676 239 12710 265
rect 12772 1183 12806 1209
rect 12772 1175 12806 1183
rect 12772 1115 12806 1137
rect 12772 1103 12806 1115
rect 12772 1047 12806 1065
rect 12772 1031 12806 1047
rect 12772 979 12806 993
rect 12772 959 12806 979
rect 12772 911 12806 921
rect 12772 887 12806 911
rect 12772 843 12806 849
rect 12772 815 12806 843
rect 12772 775 12806 777
rect 12772 743 12806 775
rect 12772 673 12806 705
rect 12772 671 12806 673
rect 12772 605 12806 633
rect 12772 599 12806 605
rect 12772 537 12806 561
rect 12772 527 12806 537
rect 12772 469 12806 489
rect 12772 455 12806 469
rect 12772 401 12806 417
rect 12772 383 12806 401
rect 12772 333 12806 345
rect 12772 311 12806 333
rect 12772 265 12806 273
rect 12772 239 12806 265
rect 12868 1183 12902 1209
rect 12868 1175 12902 1183
rect 12868 1115 12902 1137
rect 12868 1103 12902 1115
rect 12868 1047 12902 1065
rect 12868 1031 12902 1047
rect 12868 979 12902 993
rect 12868 959 12902 979
rect 12868 911 12902 921
rect 12868 887 12902 911
rect 12868 843 12902 849
rect 12868 815 12902 843
rect 12868 775 12902 777
rect 12868 743 12902 775
rect 12868 673 12902 705
rect 12868 671 12902 673
rect 12868 605 12902 633
rect 12868 599 12902 605
rect 12868 537 12902 561
rect 12868 527 12902 537
rect 12868 469 12902 489
rect 12868 455 12902 469
rect 12868 401 12902 417
rect 12868 383 12902 401
rect 12868 333 12902 345
rect 12868 311 12902 333
rect 12868 265 12902 273
rect 12868 239 12902 265
rect 12964 1183 12998 1209
rect 12964 1175 12998 1183
rect 12964 1115 12998 1137
rect 12964 1103 12998 1115
rect 12964 1047 12998 1065
rect 12964 1031 12998 1047
rect 12964 979 12998 993
rect 12964 959 12998 979
rect 12964 911 12998 921
rect 12964 887 12998 911
rect 12964 843 12998 849
rect 12964 815 12998 843
rect 12964 775 12998 777
rect 12964 743 12998 775
rect 12964 673 12998 705
rect 12964 671 12998 673
rect 12964 605 12998 633
rect 12964 599 12998 605
rect 12964 537 12998 561
rect 12964 527 12998 537
rect 12964 469 12998 489
rect 12964 455 12998 469
rect 12964 401 12998 417
rect 12964 383 12998 401
rect 12964 333 12998 345
rect 12964 311 12998 333
rect 12964 265 12998 273
rect 12964 239 12998 265
rect 13060 1183 13094 1209
rect 13060 1175 13094 1183
rect 13060 1115 13094 1137
rect 13060 1103 13094 1115
rect 13060 1047 13094 1065
rect 13060 1031 13094 1047
rect 13060 979 13094 993
rect 13060 959 13094 979
rect 13060 911 13094 921
rect 13060 887 13094 911
rect 13060 843 13094 849
rect 13060 815 13094 843
rect 13060 775 13094 777
rect 13060 743 13094 775
rect 13060 673 13094 705
rect 13060 671 13094 673
rect 13060 605 13094 633
rect 13060 599 13094 605
rect 13060 537 13094 561
rect 13060 527 13094 537
rect 13060 469 13094 489
rect 13060 455 13094 469
rect 13060 401 13094 417
rect 13060 383 13094 401
rect 13060 333 13094 345
rect 13060 311 13094 333
rect 13060 265 13094 273
rect 13060 239 13094 265
rect 13156 1183 13190 1209
rect 13156 1175 13190 1183
rect 13156 1115 13190 1137
rect 13156 1103 13190 1115
rect 13156 1047 13190 1065
rect 13156 1031 13190 1047
rect 13156 979 13190 993
rect 13156 959 13190 979
rect 13156 911 13190 921
rect 13156 887 13190 911
rect 13156 843 13190 849
rect 13156 815 13190 843
rect 13156 775 13190 777
rect 13156 743 13190 775
rect 13156 673 13190 705
rect 13156 671 13190 673
rect 13156 605 13190 633
rect 13156 599 13190 605
rect 13156 537 13190 561
rect 13156 527 13190 537
rect 13156 469 13190 489
rect 13156 455 13190 469
rect 13156 401 13190 417
rect 13156 383 13190 401
rect 13156 333 13190 345
rect 13156 311 13190 333
rect 13156 265 13190 273
rect 13156 239 13190 265
rect 13252 1183 13286 1209
rect 13252 1175 13286 1183
rect 13252 1115 13286 1137
rect 13252 1103 13286 1115
rect 13252 1047 13286 1065
rect 13252 1031 13286 1047
rect 13252 979 13286 993
rect 13252 959 13286 979
rect 13252 911 13286 921
rect 13252 887 13286 911
rect 13252 843 13286 849
rect 13252 815 13286 843
rect 13252 775 13286 777
rect 13252 743 13286 775
rect 13252 673 13286 705
rect 13252 671 13286 673
rect 13252 605 13286 633
rect 13252 599 13286 605
rect 13252 537 13286 561
rect 13252 527 13286 537
rect 13252 469 13286 489
rect 13252 455 13286 469
rect 13252 401 13286 417
rect 13252 383 13286 401
rect 13252 333 13286 345
rect 13252 311 13286 333
rect 13252 265 13286 273
rect 13252 239 13286 265
rect 13348 1183 13382 1209
rect 13348 1175 13382 1183
rect 13348 1115 13382 1137
rect 13348 1103 13382 1115
rect 13348 1047 13382 1065
rect 13348 1031 13382 1047
rect 13348 979 13382 993
rect 13348 959 13382 979
rect 13348 911 13382 921
rect 13348 887 13382 911
rect 13348 843 13382 849
rect 13348 815 13382 843
rect 13348 775 13382 777
rect 13348 743 13382 775
rect 13348 673 13382 705
rect 13348 671 13382 673
rect 13348 605 13382 633
rect 13348 599 13382 605
rect 13348 537 13382 561
rect 13348 527 13382 537
rect 13348 469 13382 489
rect 13348 455 13382 469
rect 13348 401 13382 417
rect 13348 383 13382 401
rect 13348 333 13382 345
rect 13348 311 13382 333
rect 13348 265 13382 273
rect 13348 239 13382 265
rect 13444 1183 13478 1209
rect 13444 1175 13478 1183
rect 13444 1115 13478 1137
rect 13444 1103 13478 1115
rect 13444 1047 13478 1065
rect 13444 1031 13478 1047
rect 13444 979 13478 993
rect 13444 959 13478 979
rect 13444 911 13478 921
rect 13444 887 13478 911
rect 13444 843 13478 849
rect 13444 815 13478 843
rect 13444 775 13478 777
rect 13444 743 13478 775
rect 13444 673 13478 705
rect 13444 671 13478 673
rect 13444 605 13478 633
rect 13444 599 13478 605
rect 13444 537 13478 561
rect 13444 527 13478 537
rect 13444 469 13478 489
rect 13444 455 13478 469
rect 13444 401 13478 417
rect 13444 383 13478 401
rect 13444 333 13478 345
rect 13444 311 13478 333
rect 13444 265 13478 273
rect 13444 239 13478 265
rect 13540 1183 13574 1209
rect 13540 1175 13574 1183
rect 13540 1115 13574 1137
rect 13540 1103 13574 1115
rect 13540 1047 13574 1065
rect 13540 1031 13574 1047
rect 13540 979 13574 993
rect 13540 959 13574 979
rect 13540 911 13574 921
rect 13540 887 13574 911
rect 13540 843 13574 849
rect 13540 815 13574 843
rect 13540 775 13574 777
rect 13540 743 13574 775
rect 13540 673 13574 705
rect 13540 671 13574 673
rect 13540 605 13574 633
rect 13540 599 13574 605
rect 13540 537 13574 561
rect 13540 527 13574 537
rect 13540 469 13574 489
rect 13540 455 13574 469
rect 13540 401 13574 417
rect 13540 383 13574 401
rect 13540 333 13574 345
rect 13540 311 13574 333
rect 13540 265 13574 273
rect 13540 239 13574 265
rect 11568 94 11602 128
rect 11862 78 11896 112
rect 12386 52 12420 86
rect 13060 42 13094 76
rect 10663 -23 10697 11
rect 14630 1374 14664 1408
rect 15422 1336 15456 1370
rect 14156 1183 14190 1209
rect 14156 1175 14190 1183
rect 14156 1115 14190 1137
rect 14156 1103 14190 1115
rect 14156 1047 14190 1065
rect 14156 1031 14190 1047
rect 14156 979 14190 993
rect 14156 959 14190 979
rect 14156 911 14190 921
rect 14156 887 14190 911
rect 14156 843 14190 849
rect 14156 815 14190 843
rect 14156 775 14190 777
rect 14156 743 14190 775
rect 14156 673 14190 705
rect 14156 671 14190 673
rect 14156 605 14190 633
rect 14156 599 14190 605
rect 14156 537 14190 561
rect 14156 527 14190 537
rect 14156 469 14190 489
rect 14156 455 14190 469
rect 14156 401 14190 417
rect 14156 383 14190 401
rect 14156 333 14190 345
rect 14156 311 14190 333
rect 14156 265 14190 273
rect 14156 239 14190 265
rect 14252 1183 14286 1209
rect 14252 1175 14286 1183
rect 14252 1115 14286 1137
rect 14252 1103 14286 1115
rect 14252 1047 14286 1065
rect 14252 1031 14286 1047
rect 14252 979 14286 993
rect 14252 959 14286 979
rect 14252 911 14286 921
rect 14252 887 14286 911
rect 14252 843 14286 849
rect 14252 815 14286 843
rect 14252 775 14286 777
rect 14252 743 14286 775
rect 14252 673 14286 705
rect 14252 671 14286 673
rect 14252 605 14286 633
rect 14252 599 14286 605
rect 14252 537 14286 561
rect 14252 527 14286 537
rect 14252 469 14286 489
rect 14252 455 14286 469
rect 14252 401 14286 417
rect 14252 383 14286 401
rect 14252 333 14286 345
rect 14252 311 14286 333
rect 14252 265 14286 273
rect 14252 239 14286 265
rect 14348 1183 14382 1209
rect 14348 1175 14382 1183
rect 14348 1115 14382 1137
rect 14348 1103 14382 1115
rect 14348 1047 14382 1065
rect 14348 1031 14382 1047
rect 14348 979 14382 993
rect 14348 959 14382 979
rect 14348 911 14382 921
rect 14348 887 14382 911
rect 14348 843 14382 849
rect 14348 815 14382 843
rect 14348 775 14382 777
rect 14348 743 14382 775
rect 14348 673 14382 705
rect 14348 671 14382 673
rect 14348 605 14382 633
rect 14348 599 14382 605
rect 14348 537 14382 561
rect 14348 527 14382 537
rect 14348 469 14382 489
rect 14348 455 14382 469
rect 14348 401 14382 417
rect 14348 383 14382 401
rect 14348 333 14382 345
rect 14348 311 14382 333
rect 14348 265 14382 273
rect 14348 239 14382 265
rect 14444 1183 14478 1209
rect 14444 1175 14478 1183
rect 14444 1115 14478 1137
rect 14444 1103 14478 1115
rect 14444 1047 14478 1065
rect 14444 1031 14478 1047
rect 14444 979 14478 993
rect 14444 959 14478 979
rect 14444 911 14478 921
rect 14444 887 14478 911
rect 14444 843 14478 849
rect 14444 815 14478 843
rect 14444 775 14478 777
rect 14444 743 14478 775
rect 14444 673 14478 705
rect 14444 671 14478 673
rect 14444 605 14478 633
rect 14444 599 14478 605
rect 14444 537 14478 561
rect 14444 527 14478 537
rect 14444 469 14478 489
rect 14444 455 14478 469
rect 14444 401 14478 417
rect 14444 383 14478 401
rect 14444 333 14478 345
rect 14444 311 14478 333
rect 14444 265 14478 273
rect 14444 239 14478 265
rect 14540 1183 14574 1209
rect 14540 1175 14574 1183
rect 14540 1115 14574 1137
rect 14540 1103 14574 1115
rect 14540 1047 14574 1065
rect 14540 1031 14574 1047
rect 14540 979 14574 993
rect 14540 959 14574 979
rect 14540 911 14574 921
rect 14540 887 14574 911
rect 14540 843 14574 849
rect 14540 815 14574 843
rect 14540 775 14574 777
rect 14540 743 14574 775
rect 14540 673 14574 705
rect 14540 671 14574 673
rect 14540 605 14574 633
rect 14540 599 14574 605
rect 14540 537 14574 561
rect 14540 527 14574 537
rect 14540 469 14574 489
rect 14540 455 14574 469
rect 14540 401 14574 417
rect 14540 383 14574 401
rect 14540 333 14574 345
rect 14540 311 14574 333
rect 14540 265 14574 273
rect 14540 239 14574 265
rect 14636 1183 14670 1209
rect 14636 1175 14670 1183
rect 14636 1115 14670 1137
rect 14636 1103 14670 1115
rect 14636 1047 14670 1065
rect 14636 1031 14670 1047
rect 14636 979 14670 993
rect 14636 959 14670 979
rect 14636 911 14670 921
rect 14636 887 14670 911
rect 14636 843 14670 849
rect 14636 815 14670 843
rect 14636 775 14670 777
rect 14636 743 14670 775
rect 14636 673 14670 705
rect 14636 671 14670 673
rect 14636 605 14670 633
rect 14636 599 14670 605
rect 14636 537 14670 561
rect 14636 527 14670 537
rect 14636 469 14670 489
rect 14636 455 14670 469
rect 14636 401 14670 417
rect 14636 383 14670 401
rect 14636 333 14670 345
rect 14636 311 14670 333
rect 14636 265 14670 273
rect 14636 239 14670 265
rect 14732 1183 14766 1209
rect 14732 1175 14766 1183
rect 14732 1115 14766 1137
rect 14732 1103 14766 1115
rect 14732 1047 14766 1065
rect 14732 1031 14766 1047
rect 14732 979 14766 993
rect 14732 959 14766 979
rect 14732 911 14766 921
rect 14732 887 14766 911
rect 14732 843 14766 849
rect 14732 815 14766 843
rect 14732 775 14766 777
rect 14732 743 14766 775
rect 14732 673 14766 705
rect 14732 671 14766 673
rect 14732 605 14766 633
rect 14732 599 14766 605
rect 14732 537 14766 561
rect 14732 527 14766 537
rect 14732 469 14766 489
rect 14732 455 14766 469
rect 14732 401 14766 417
rect 14732 383 14766 401
rect 14732 333 14766 345
rect 14732 311 14766 333
rect 14732 265 14766 273
rect 14732 239 14766 265
rect 14828 1183 14862 1209
rect 14828 1175 14862 1183
rect 14828 1115 14862 1137
rect 14828 1103 14862 1115
rect 14828 1047 14862 1065
rect 14828 1031 14862 1047
rect 14828 979 14862 993
rect 14828 959 14862 979
rect 14828 911 14862 921
rect 14828 887 14862 911
rect 14828 843 14862 849
rect 14828 815 14862 843
rect 14828 775 14862 777
rect 14828 743 14862 775
rect 14828 673 14862 705
rect 14828 671 14862 673
rect 14828 605 14862 633
rect 14828 599 14862 605
rect 14828 537 14862 561
rect 14828 527 14862 537
rect 14828 469 14862 489
rect 14828 455 14862 469
rect 14828 401 14862 417
rect 14828 383 14862 401
rect 14828 333 14862 345
rect 14828 311 14862 333
rect 14828 265 14862 273
rect 14828 239 14862 265
rect 14924 1183 14958 1209
rect 14924 1175 14958 1183
rect 14924 1115 14958 1137
rect 14924 1103 14958 1115
rect 14924 1047 14958 1065
rect 14924 1031 14958 1047
rect 14924 979 14958 993
rect 14924 959 14958 979
rect 14924 911 14958 921
rect 14924 887 14958 911
rect 14924 843 14958 849
rect 14924 815 14958 843
rect 14924 775 14958 777
rect 14924 743 14958 775
rect 14924 673 14958 705
rect 14924 671 14958 673
rect 14924 605 14958 633
rect 14924 599 14958 605
rect 14924 537 14958 561
rect 14924 527 14958 537
rect 14924 469 14958 489
rect 14924 455 14958 469
rect 14924 401 14958 417
rect 14924 383 14958 401
rect 14924 333 14958 345
rect 14924 311 14958 333
rect 14924 265 14958 273
rect 14924 239 14958 265
rect 15020 1183 15054 1209
rect 15020 1175 15054 1183
rect 15020 1115 15054 1137
rect 15020 1103 15054 1115
rect 15020 1047 15054 1065
rect 15020 1031 15054 1047
rect 15020 979 15054 993
rect 15020 959 15054 979
rect 15020 911 15054 921
rect 15020 887 15054 911
rect 15020 843 15054 849
rect 15020 815 15054 843
rect 15020 775 15054 777
rect 15020 743 15054 775
rect 15020 673 15054 705
rect 15020 671 15054 673
rect 15020 605 15054 633
rect 15020 599 15054 605
rect 15020 537 15054 561
rect 15020 527 15054 537
rect 15020 469 15054 489
rect 15020 455 15054 469
rect 15020 401 15054 417
rect 15020 383 15054 401
rect 15020 333 15054 345
rect 15020 311 15054 333
rect 15020 265 15054 273
rect 15020 239 15054 265
rect 15116 1183 15150 1209
rect 15116 1175 15150 1183
rect 15116 1115 15150 1137
rect 15116 1103 15150 1115
rect 15116 1047 15150 1065
rect 15116 1031 15150 1047
rect 15116 979 15150 993
rect 15116 959 15150 979
rect 15116 911 15150 921
rect 15116 887 15150 911
rect 15116 843 15150 849
rect 15116 815 15150 843
rect 15116 775 15150 777
rect 15116 743 15150 775
rect 15116 673 15150 705
rect 15116 671 15150 673
rect 15116 605 15150 633
rect 15116 599 15150 605
rect 15116 537 15150 561
rect 15116 527 15150 537
rect 15116 469 15150 489
rect 15116 455 15150 469
rect 15116 401 15150 417
rect 15116 383 15150 401
rect 15116 333 15150 345
rect 15116 311 15150 333
rect 15116 265 15150 273
rect 15116 239 15150 265
rect 15212 1183 15246 1209
rect 15212 1175 15246 1183
rect 15212 1115 15246 1137
rect 15212 1103 15246 1115
rect 15212 1047 15246 1065
rect 15212 1031 15246 1047
rect 15212 979 15246 993
rect 15212 959 15246 979
rect 15212 911 15246 921
rect 15212 887 15246 911
rect 15212 843 15246 849
rect 15212 815 15246 843
rect 15212 775 15246 777
rect 15212 743 15246 775
rect 15212 673 15246 705
rect 15212 671 15246 673
rect 15212 605 15246 633
rect 15212 599 15246 605
rect 15212 537 15246 561
rect 15212 527 15246 537
rect 15212 469 15246 489
rect 15212 455 15246 469
rect 15212 401 15246 417
rect 15212 383 15246 401
rect 15212 333 15246 345
rect 15212 311 15246 333
rect 15212 265 15246 273
rect 15212 239 15246 265
rect 15422 1227 15456 1257
rect 15422 1223 15456 1227
rect 15422 1159 15456 1185
rect 15422 1151 15456 1159
rect 15422 1091 15456 1113
rect 15422 1079 15456 1091
rect 15422 1023 15456 1041
rect 15422 1007 15456 1023
rect 15422 955 15456 969
rect 15422 935 15456 955
rect 15422 887 15456 897
rect 15422 863 15456 887
rect 15422 819 15456 825
rect 15422 791 15456 819
rect 15422 751 15456 753
rect 15422 719 15456 751
rect 15422 649 15456 681
rect 15422 647 15456 649
rect 15422 581 15456 609
rect 15422 575 15456 581
rect 15422 513 15456 537
rect 15422 503 15456 513
rect 15422 445 15456 465
rect 15422 431 15456 445
rect 15422 377 15456 393
rect 15422 359 15456 377
rect 15422 309 15456 321
rect 15422 287 15456 309
rect 15422 241 15456 249
rect 15422 215 15456 241
rect 15422 173 15456 177
rect 15422 143 15456 173
rect 14724 68 14758 102
rect 15510 1227 15544 1257
rect 15510 1223 15544 1227
rect 15510 1159 15544 1185
rect 15510 1151 15544 1159
rect 15510 1091 15544 1113
rect 15510 1079 15544 1091
rect 15510 1023 15544 1041
rect 15510 1007 15544 1023
rect 15510 955 15544 969
rect 15510 935 15544 955
rect 15510 887 15544 897
rect 15510 863 15544 887
rect 15510 819 15544 825
rect 15510 791 15544 819
rect 15510 751 15544 753
rect 15510 719 15544 751
rect 15510 649 15544 681
rect 15510 647 15544 649
rect 15510 581 15544 609
rect 15510 575 15544 581
rect 15510 513 15544 537
rect 15510 503 15544 513
rect 15510 445 15544 465
rect 15510 431 15544 445
rect 15510 377 15544 393
rect 15510 359 15544 377
rect 15510 309 15544 321
rect 15510 287 15544 309
rect 15510 241 15544 249
rect 15510 215 15544 241
rect 15510 173 15544 177
rect 15510 143 15544 173
rect 15018 52 15052 86
rect 15510 18 15544 52
rect 13965 -49 13999 -15
<< metal1 >>
rect 1738 7820 1748 7926
rect 1840 7820 1850 7926
rect -558 6998 12598 7210
rect -1658 5921 -1612 5936
rect -1658 5887 -1652 5921
rect -1618 5887 -1612 5921
rect -1658 5849 -1612 5887
rect -1658 5815 -1652 5849
rect -1618 5815 -1612 5849
rect -1658 5777 -1612 5815
rect -1658 5743 -1652 5777
rect -1618 5743 -1612 5777
rect -1658 5705 -1612 5743
rect -1658 5671 -1652 5705
rect -1618 5671 -1612 5705
rect -1658 5633 -1612 5671
rect -1658 5599 -1652 5633
rect -1618 5599 -1612 5633
rect -1658 5561 -1612 5599
rect -1658 5527 -1652 5561
rect -1618 5527 -1612 5561
rect -1658 5489 -1612 5527
rect -1658 5455 -1652 5489
rect -1618 5455 -1612 5489
rect -1658 5417 -1612 5455
rect -1658 5383 -1652 5417
rect -1618 5383 -1612 5417
rect -1658 5345 -1612 5383
rect -1658 5311 -1652 5345
rect -1618 5311 -1612 5345
rect -1658 5273 -1612 5311
rect -1658 5239 -1652 5273
rect -1618 5239 -1612 5273
rect -1658 5201 -1612 5239
rect -1658 5167 -1652 5201
rect -1618 5167 -1612 5201
rect -1658 5129 -1612 5167
rect -1658 5095 -1652 5129
rect -1618 5095 -1612 5129
rect -1658 5057 -1612 5095
rect -1658 5023 -1652 5057
rect -1618 5023 -1612 5057
rect -1658 4985 -1612 5023
rect -1658 4951 -1652 4985
rect -1618 4951 -1612 4985
rect -1658 4936 -1612 4951
rect -1560 5921 -1514 5936
rect -1560 5887 -1554 5921
rect -1520 5887 -1514 5921
rect -1560 5849 -1514 5887
rect -1560 5815 -1554 5849
rect -1520 5815 -1514 5849
rect -1560 5777 -1514 5815
rect -1560 5743 -1554 5777
rect -1520 5743 -1514 5777
rect -1560 5705 -1514 5743
rect -1560 5671 -1554 5705
rect -1520 5671 -1514 5705
rect -1560 5633 -1514 5671
rect -1560 5599 -1554 5633
rect -1520 5599 -1514 5633
rect -1560 5561 -1514 5599
rect -1560 5527 -1554 5561
rect -1520 5527 -1514 5561
rect -1560 5489 -1514 5527
rect -1560 5455 -1554 5489
rect -1520 5455 -1514 5489
rect -1560 5417 -1514 5455
rect -1560 5383 -1554 5417
rect -1520 5383 -1514 5417
rect -1560 5345 -1514 5383
rect -1560 5311 -1554 5345
rect -1520 5311 -1514 5345
rect -1560 5273 -1514 5311
rect -1560 5239 -1554 5273
rect -1520 5239 -1514 5273
rect -1560 5201 -1514 5239
rect -1560 5167 -1554 5201
rect -1520 5167 -1514 5201
rect -1560 5129 -1514 5167
rect -1560 5095 -1554 5129
rect -1520 5095 -1514 5129
rect -1560 5057 -1514 5095
rect -1560 5023 -1554 5057
rect -1520 5023 -1514 5057
rect -1560 4985 -1514 5023
rect -1560 4951 -1554 4985
rect -1520 4951 -1514 4985
rect -1560 4936 -1514 4951
rect -1462 5921 -1416 5936
rect -1462 5887 -1456 5921
rect -1422 5887 -1416 5921
rect -1462 5849 -1416 5887
rect -1462 5815 -1456 5849
rect -1422 5815 -1416 5849
rect -1462 5777 -1416 5815
rect -1462 5743 -1456 5777
rect -1422 5743 -1416 5777
rect -1462 5705 -1416 5743
rect -1462 5671 -1456 5705
rect -1422 5671 -1416 5705
rect -1462 5633 -1416 5671
rect -1462 5599 -1456 5633
rect -1422 5599 -1416 5633
rect -1462 5561 -1416 5599
rect -1462 5527 -1456 5561
rect -1422 5527 -1416 5561
rect -1462 5489 -1416 5527
rect -1462 5455 -1456 5489
rect -1422 5455 -1416 5489
rect -1462 5417 -1416 5455
rect -1462 5383 -1456 5417
rect -1422 5383 -1416 5417
rect -1462 5345 -1416 5383
rect -1462 5311 -1456 5345
rect -1422 5311 -1416 5345
rect -1462 5273 -1416 5311
rect -1462 5239 -1456 5273
rect -1422 5239 -1416 5273
rect -1462 5201 -1416 5239
rect -1462 5167 -1456 5201
rect -1422 5167 -1416 5201
rect -1462 5129 -1416 5167
rect -1462 5095 -1456 5129
rect -1422 5095 -1416 5129
rect -1462 5057 -1416 5095
rect -1462 5023 -1456 5057
rect -1422 5023 -1416 5057
rect -1462 4985 -1416 5023
rect -1462 4951 -1456 4985
rect -1422 4951 -1416 4985
rect -1462 4936 -1416 4951
rect -1364 5921 -1318 5936
rect -1364 5887 -1358 5921
rect -1324 5887 -1318 5921
rect -1364 5849 -1318 5887
rect -1364 5815 -1358 5849
rect -1324 5815 -1318 5849
rect -1364 5777 -1318 5815
rect -1364 5743 -1358 5777
rect -1324 5743 -1318 5777
rect -1364 5705 -1318 5743
rect -1364 5671 -1358 5705
rect -1324 5671 -1318 5705
rect -1364 5633 -1318 5671
rect -1364 5599 -1358 5633
rect -1324 5599 -1318 5633
rect -1364 5561 -1318 5599
rect -1364 5527 -1358 5561
rect -1324 5527 -1318 5561
rect -1364 5489 -1318 5527
rect -1364 5455 -1358 5489
rect -1324 5455 -1318 5489
rect -1364 5417 -1318 5455
rect -1364 5383 -1358 5417
rect -1324 5383 -1318 5417
rect -1364 5345 -1318 5383
rect -1364 5311 -1358 5345
rect -1324 5311 -1318 5345
rect -1364 5273 -1318 5311
rect -1364 5239 -1358 5273
rect -1324 5239 -1318 5273
rect -1364 5201 -1318 5239
rect -1364 5167 -1358 5201
rect -1324 5167 -1318 5201
rect -1364 5129 -1318 5167
rect -1364 5095 -1358 5129
rect -1324 5095 -1318 5129
rect -1364 5057 -1318 5095
rect -1364 5023 -1358 5057
rect -1324 5023 -1318 5057
rect -1364 4985 -1318 5023
rect -1364 4951 -1358 4985
rect -1324 4951 -1318 4985
rect -1364 4936 -1318 4951
rect -1266 5921 -1220 5936
rect -1266 5887 -1260 5921
rect -1226 5887 -1220 5921
rect -1266 5849 -1220 5887
rect -1266 5815 -1260 5849
rect -1226 5815 -1220 5849
rect -1266 5777 -1220 5815
rect -1266 5743 -1260 5777
rect -1226 5743 -1220 5777
rect -1266 5705 -1220 5743
rect -1266 5671 -1260 5705
rect -1226 5671 -1220 5705
rect -1266 5633 -1220 5671
rect -1266 5599 -1260 5633
rect -1226 5599 -1220 5633
rect -1266 5561 -1220 5599
rect -1266 5527 -1260 5561
rect -1226 5527 -1220 5561
rect -1266 5489 -1220 5527
rect -1266 5455 -1260 5489
rect -1226 5455 -1220 5489
rect -1266 5417 -1220 5455
rect -1266 5383 -1260 5417
rect -1226 5383 -1220 5417
rect -1266 5345 -1220 5383
rect -1266 5311 -1260 5345
rect -1226 5311 -1220 5345
rect -1266 5273 -1220 5311
rect -1266 5239 -1260 5273
rect -1226 5239 -1220 5273
rect -1266 5201 -1220 5239
rect -1266 5167 -1260 5201
rect -1226 5167 -1220 5201
rect -1266 5129 -1220 5167
rect -1266 5095 -1260 5129
rect -1226 5095 -1220 5129
rect -1266 5057 -1220 5095
rect -1266 5023 -1260 5057
rect -1226 5023 -1220 5057
rect -1266 4985 -1220 5023
rect -1266 4951 -1260 4985
rect -1226 4951 -1220 4985
rect -1266 4936 -1220 4951
rect -1168 5921 -1122 5936
rect -1168 5887 -1162 5921
rect -1128 5887 -1122 5921
rect -1168 5849 -1122 5887
rect -1168 5815 -1162 5849
rect -1128 5815 -1122 5849
rect -1168 5777 -1122 5815
rect -1168 5743 -1162 5777
rect -1128 5743 -1122 5777
rect -1168 5705 -1122 5743
rect -1168 5671 -1162 5705
rect -1128 5671 -1122 5705
rect -1168 5633 -1122 5671
rect -1168 5599 -1162 5633
rect -1128 5599 -1122 5633
rect -1168 5561 -1122 5599
rect -1168 5527 -1162 5561
rect -1128 5527 -1122 5561
rect -1168 5489 -1122 5527
rect -1168 5455 -1162 5489
rect -1128 5455 -1122 5489
rect -1168 5417 -1122 5455
rect -1168 5383 -1162 5417
rect -1128 5383 -1122 5417
rect -1168 5345 -1122 5383
rect -1168 5311 -1162 5345
rect -1128 5311 -1122 5345
rect -1168 5273 -1122 5311
rect -1168 5239 -1162 5273
rect -1128 5239 -1122 5273
rect -1168 5201 -1122 5239
rect -1168 5167 -1162 5201
rect -1128 5167 -1122 5201
rect -1168 5129 -1122 5167
rect -1168 5095 -1162 5129
rect -1128 5095 -1122 5129
rect -1168 5057 -1122 5095
rect -1168 5023 -1162 5057
rect -1128 5023 -1122 5057
rect -1168 4985 -1122 5023
rect -1168 4951 -1162 4985
rect -1128 4951 -1122 4985
rect -1168 4936 -1122 4951
rect -1070 5921 -1024 5936
rect -1070 5887 -1064 5921
rect -1030 5887 -1024 5921
rect -1070 5849 -1024 5887
rect -1070 5815 -1064 5849
rect -1030 5815 -1024 5849
rect -1070 5777 -1024 5815
rect -1070 5743 -1064 5777
rect -1030 5743 -1024 5777
rect -1070 5705 -1024 5743
rect -1070 5671 -1064 5705
rect -1030 5671 -1024 5705
rect -1070 5633 -1024 5671
rect -1070 5599 -1064 5633
rect -1030 5599 -1024 5633
rect -1070 5561 -1024 5599
rect -1070 5527 -1064 5561
rect -1030 5527 -1024 5561
rect -1070 5489 -1024 5527
rect -1070 5455 -1064 5489
rect -1030 5455 -1024 5489
rect -1070 5417 -1024 5455
rect -1070 5383 -1064 5417
rect -1030 5383 -1024 5417
rect -1070 5345 -1024 5383
rect -1070 5311 -1064 5345
rect -1030 5311 -1024 5345
rect -1070 5273 -1024 5311
rect -1070 5239 -1064 5273
rect -1030 5239 -1024 5273
rect -1070 5201 -1024 5239
rect -1070 5167 -1064 5201
rect -1030 5167 -1024 5201
rect -1070 5129 -1024 5167
rect -1070 5095 -1064 5129
rect -1030 5095 -1024 5129
rect -1070 5057 -1024 5095
rect -1070 5023 -1064 5057
rect -1030 5023 -1024 5057
rect -1070 4985 -1024 5023
rect -1070 4951 -1064 4985
rect -1030 4951 -1024 4985
rect -1070 4936 -1024 4951
rect -972 5921 -926 5936
rect -972 5887 -966 5921
rect -932 5887 -926 5921
rect -972 5849 -926 5887
rect -972 5815 -966 5849
rect -932 5815 -926 5849
rect -972 5777 -926 5815
rect -972 5743 -966 5777
rect -932 5743 -926 5777
rect -972 5705 -926 5743
rect -972 5671 -966 5705
rect -932 5671 -926 5705
rect -972 5633 -926 5671
rect -972 5599 -966 5633
rect -932 5599 -926 5633
rect -972 5561 -926 5599
rect -972 5527 -966 5561
rect -932 5527 -926 5561
rect -972 5489 -926 5527
rect -972 5455 -966 5489
rect -932 5455 -926 5489
rect -972 5417 -926 5455
rect -972 5383 -966 5417
rect -932 5383 -926 5417
rect -972 5345 -926 5383
rect -972 5311 -966 5345
rect -932 5311 -926 5345
rect -972 5273 -926 5311
rect -972 5239 -966 5273
rect -932 5239 -926 5273
rect -972 5201 -926 5239
rect -972 5167 -966 5201
rect -932 5167 -926 5201
rect -972 5129 -926 5167
rect -972 5095 -966 5129
rect -932 5095 -926 5129
rect -972 5057 -926 5095
rect -972 5023 -966 5057
rect -932 5023 -926 5057
rect -972 4985 -926 5023
rect -972 4951 -966 4985
rect -932 4951 -926 4985
rect -972 4936 -926 4951
rect -874 5921 -828 5936
rect -874 5887 -868 5921
rect -834 5887 -828 5921
rect -874 5849 -828 5887
rect -874 5815 -868 5849
rect -834 5815 -828 5849
rect -874 5777 -828 5815
rect -874 5743 -868 5777
rect -834 5743 -828 5777
rect -874 5705 -828 5743
rect -874 5671 -868 5705
rect -834 5671 -828 5705
rect -874 5633 -828 5671
rect -874 5599 -868 5633
rect -834 5599 -828 5633
rect -874 5561 -828 5599
rect -874 5527 -868 5561
rect -834 5527 -828 5561
rect -874 5489 -828 5527
rect -874 5455 -868 5489
rect -834 5455 -828 5489
rect -874 5417 -828 5455
rect -874 5383 -868 5417
rect -834 5383 -828 5417
rect -874 5345 -828 5383
rect -874 5311 -868 5345
rect -834 5311 -828 5345
rect -874 5273 -828 5311
rect -874 5239 -868 5273
rect -834 5239 -828 5273
rect -874 5201 -828 5239
rect -874 5167 -868 5201
rect -834 5167 -828 5201
rect -874 5129 -828 5167
rect -874 5095 -868 5129
rect -834 5095 -828 5129
rect -874 5057 -828 5095
rect -874 5023 -868 5057
rect -834 5023 -828 5057
rect -874 4985 -828 5023
rect -874 4951 -868 4985
rect -834 4951 -828 4985
rect -874 4936 -828 4951
rect -1126 4792 -1022 4794
rect -558 4792 -402 6998
rect 274 6807 336 6998
rect 1758 6947 1834 6950
rect 1758 6906 1770 6947
rect 752 6895 1770 6906
rect 1822 6906 1834 6947
rect 1822 6895 2488 6906
rect 752 6892 2488 6895
rect 752 6858 764 6892
rect 798 6858 2488 6892
rect 752 6848 2488 6858
rect 274 6773 288 6807
rect 322 6773 336 6807
rect 274 6762 336 6773
rect 2428 6788 2488 6848
rect 2758 6809 2960 6814
rect 2428 6754 2440 6788
rect 2474 6754 2488 6788
rect 2716 6803 2893 6809
rect 2716 6769 2728 6803
rect 2762 6769 2893 6803
rect 2716 6763 2893 6769
rect 2428 6744 2488 6754
rect 2758 6757 2893 6763
rect 2945 6757 2960 6809
rect 2758 6752 2960 6757
rect 3230 6791 3292 6998
rect 4668 6927 4760 6934
rect 4668 6890 4688 6927
rect 3708 6876 4688 6890
rect 3708 6842 3720 6876
rect 3754 6875 4688 6876
rect 4740 6890 4760 6927
rect 4740 6875 5444 6890
rect 3754 6842 5444 6875
rect 3708 6832 5444 6842
rect 3230 6757 3244 6791
rect 3278 6757 3292 6791
rect 3230 6742 3292 6757
rect 5384 6772 5444 6832
rect 5908 6803 5990 6806
rect 5908 6800 5923 6803
rect 5706 6793 5923 6800
rect 5384 6738 5396 6772
rect 5430 6738 5444 6772
rect 5672 6787 5923 6793
rect 5672 6753 5684 6787
rect 5718 6753 5923 6787
rect 5672 6751 5923 6753
rect 5975 6751 5990 6803
rect 5672 6748 5990 6751
rect 6260 6791 6322 6998
rect 7662 6934 7766 6952
rect 7662 6890 7688 6934
rect 6738 6882 7688 6890
rect 7740 6890 7766 6934
rect 7740 6882 8474 6890
rect 6738 6876 8474 6882
rect 6738 6842 6750 6876
rect 6784 6842 8474 6876
rect 6738 6832 8474 6842
rect 6260 6757 6274 6791
rect 6308 6757 6322 6791
rect 5672 6747 5950 6748
rect 5706 6742 5950 6747
rect 6260 6744 6322 6757
rect 8414 6772 8474 6832
rect 8740 6799 8972 6804
rect 8740 6793 8905 6799
rect 5384 6728 5444 6738
rect 8414 6738 8426 6772
rect 8460 6738 8474 6772
rect 8702 6787 8905 6793
rect 8702 6753 8714 6787
rect 8748 6753 8905 6787
rect 8702 6747 8905 6753
rect 8957 6747 8972 6799
rect 8740 6742 8972 6747
rect 9348 6789 9410 6998
rect 10730 6922 10838 6940
rect 10730 6888 10758 6922
rect 9826 6874 10758 6888
rect 9826 6840 9838 6874
rect 9872 6870 10758 6874
rect 10810 6888 10838 6922
rect 10810 6870 11562 6888
rect 9872 6840 11562 6870
rect 9826 6830 11562 6840
rect 9348 6755 9362 6789
rect 9396 6755 9410 6789
rect 9348 6742 9410 6755
rect 11502 6770 11562 6830
rect 11814 6801 12122 6806
rect 11814 6791 12055 6801
rect 8414 6728 8474 6738
rect 11502 6736 11514 6770
rect 11548 6736 11562 6770
rect 11790 6785 12055 6791
rect 11790 6751 11802 6785
rect 11836 6751 12055 6785
rect 11790 6749 12055 6751
rect 12107 6749 12122 6801
rect 11790 6745 12122 6749
rect 11814 6744 12122 6745
rect 12504 6763 12566 6998
rect 13922 6899 14036 6920
rect 13922 6862 13953 6899
rect 12982 6848 13953 6862
rect 12982 6814 12994 6848
rect 13028 6847 13953 6848
rect 14005 6862 14036 6899
rect 14005 6847 14718 6862
rect 13028 6814 14718 6847
rect 12982 6804 14718 6814
rect 11502 6726 11562 6736
rect 12504 6729 12518 6763
rect 12552 6729 12566 6763
rect 12504 6718 12566 6729
rect 14658 6744 14718 6804
rect 14658 6710 14670 6744
rect 14704 6710 14718 6744
rect 14844 6769 14978 6774
rect 14844 6717 14855 6769
rect 14907 6765 14978 6769
rect 14907 6759 15004 6765
rect 14907 6725 14958 6759
rect 14992 6725 15004 6759
rect 14907 6719 15004 6725
rect 14907 6717 14978 6719
rect 14844 6712 14978 6717
rect 14658 6700 14718 6710
rect 188 6591 234 6606
rect 188 6557 194 6591
rect 228 6557 234 6591
rect 188 6519 234 6557
rect 188 6485 194 6519
rect 228 6485 234 6519
rect 188 6447 234 6485
rect 188 6413 194 6447
rect 228 6413 234 6447
rect 188 6375 234 6413
rect 188 6341 194 6375
rect 228 6341 234 6375
rect 188 6303 234 6341
rect 188 6269 194 6303
rect 228 6269 234 6303
rect 188 6231 234 6269
rect 188 6197 194 6231
rect 228 6197 234 6231
rect 188 6159 234 6197
rect 188 6125 194 6159
rect 228 6125 234 6159
rect 188 6087 234 6125
rect 188 6053 194 6087
rect 228 6053 234 6087
rect 188 6015 234 6053
rect 188 5981 194 6015
rect 228 5981 234 6015
rect 188 5943 234 5981
rect 188 5909 194 5943
rect 228 5909 234 5943
rect 188 5871 234 5909
rect 188 5837 194 5871
rect 228 5837 234 5871
rect 188 5799 234 5837
rect 188 5765 194 5799
rect 228 5765 234 5799
rect 188 5727 234 5765
rect 188 5693 194 5727
rect 228 5693 234 5727
rect 188 5655 234 5693
rect 188 5621 194 5655
rect 228 5621 234 5655
rect 188 5606 234 5621
rect 284 6591 330 6606
rect 284 6557 290 6591
rect 324 6557 330 6591
rect 284 6519 330 6557
rect 284 6485 290 6519
rect 324 6485 330 6519
rect 284 6447 330 6485
rect 284 6413 290 6447
rect 324 6413 330 6447
rect 284 6375 330 6413
rect 284 6341 290 6375
rect 324 6341 330 6375
rect 284 6303 330 6341
rect 284 6269 290 6303
rect 324 6269 330 6303
rect 284 6231 330 6269
rect 284 6197 290 6231
rect 324 6197 330 6231
rect 284 6159 330 6197
rect 284 6125 290 6159
rect 324 6125 330 6159
rect 284 6087 330 6125
rect 284 6053 290 6087
rect 324 6053 330 6087
rect 284 6015 330 6053
rect 284 5981 290 6015
rect 324 5981 330 6015
rect 284 5943 330 5981
rect 284 5909 290 5943
rect 324 5909 330 5943
rect 284 5871 330 5909
rect 284 5837 290 5871
rect 324 5837 330 5871
rect 284 5799 330 5837
rect 284 5765 290 5799
rect 324 5765 330 5799
rect 284 5727 330 5765
rect 284 5693 290 5727
rect 324 5693 330 5727
rect 284 5655 330 5693
rect 284 5621 290 5655
rect 324 5621 330 5655
rect 284 5606 330 5621
rect 380 6591 426 6606
rect 380 6557 386 6591
rect 420 6557 426 6591
rect 380 6519 426 6557
rect 380 6485 386 6519
rect 420 6485 426 6519
rect 380 6447 426 6485
rect 380 6413 386 6447
rect 420 6413 426 6447
rect 380 6375 426 6413
rect 380 6341 386 6375
rect 420 6341 426 6375
rect 380 6303 426 6341
rect 380 6269 386 6303
rect 420 6269 426 6303
rect 380 6231 426 6269
rect 380 6197 386 6231
rect 420 6197 426 6231
rect 380 6159 426 6197
rect 380 6125 386 6159
rect 420 6125 426 6159
rect 380 6087 426 6125
rect 380 6053 386 6087
rect 420 6053 426 6087
rect 380 6015 426 6053
rect 380 5981 386 6015
rect 420 5981 426 6015
rect 380 5943 426 5981
rect 380 5909 386 5943
rect 420 5909 426 5943
rect 380 5871 426 5909
rect 380 5837 386 5871
rect 420 5837 426 5871
rect 380 5799 426 5837
rect 380 5765 386 5799
rect 420 5765 426 5799
rect 380 5727 426 5765
rect 380 5693 386 5727
rect 420 5693 426 5727
rect 380 5655 426 5693
rect 380 5621 386 5655
rect 420 5621 426 5655
rect 380 5606 426 5621
rect 476 6591 522 6606
rect 476 6557 482 6591
rect 516 6557 522 6591
rect 476 6519 522 6557
rect 476 6485 482 6519
rect 516 6485 522 6519
rect 476 6447 522 6485
rect 476 6413 482 6447
rect 516 6413 522 6447
rect 476 6375 522 6413
rect 476 6341 482 6375
rect 516 6341 522 6375
rect 476 6303 522 6341
rect 476 6269 482 6303
rect 516 6269 522 6303
rect 476 6231 522 6269
rect 476 6197 482 6231
rect 516 6197 522 6231
rect 476 6159 522 6197
rect 476 6125 482 6159
rect 516 6125 522 6159
rect 476 6087 522 6125
rect 476 6053 482 6087
rect 516 6053 522 6087
rect 476 6015 522 6053
rect 476 5981 482 6015
rect 516 5981 522 6015
rect 476 5943 522 5981
rect 476 5909 482 5943
rect 516 5909 522 5943
rect 476 5871 522 5909
rect 476 5837 482 5871
rect 516 5837 522 5871
rect 476 5799 522 5837
rect 476 5765 482 5799
rect 516 5765 522 5799
rect 476 5727 522 5765
rect 476 5693 482 5727
rect 516 5693 522 5727
rect 476 5655 522 5693
rect 476 5621 482 5655
rect 516 5621 522 5655
rect 476 5606 522 5621
rect 572 6591 618 6606
rect 572 6557 578 6591
rect 612 6557 618 6591
rect 572 6519 618 6557
rect 572 6485 578 6519
rect 612 6485 618 6519
rect 572 6447 618 6485
rect 572 6413 578 6447
rect 612 6413 618 6447
rect 572 6375 618 6413
rect 572 6341 578 6375
rect 612 6341 618 6375
rect 572 6303 618 6341
rect 572 6269 578 6303
rect 612 6269 618 6303
rect 572 6231 618 6269
rect 572 6197 578 6231
rect 612 6197 618 6231
rect 572 6159 618 6197
rect 572 6125 578 6159
rect 612 6125 618 6159
rect 572 6087 618 6125
rect 572 6053 578 6087
rect 612 6053 618 6087
rect 572 6015 618 6053
rect 572 5981 578 6015
rect 612 5981 618 6015
rect 572 5943 618 5981
rect 572 5909 578 5943
rect 612 5909 618 5943
rect 572 5871 618 5909
rect 572 5837 578 5871
rect 612 5837 618 5871
rect 572 5799 618 5837
rect 572 5765 578 5799
rect 612 5765 618 5799
rect 572 5727 618 5765
rect 572 5693 578 5727
rect 612 5693 618 5727
rect 572 5655 618 5693
rect 572 5621 578 5655
rect 612 5621 618 5655
rect 572 5606 618 5621
rect 668 6591 714 6606
rect 668 6557 674 6591
rect 708 6557 714 6591
rect 668 6519 714 6557
rect 668 6485 674 6519
rect 708 6485 714 6519
rect 668 6447 714 6485
rect 668 6413 674 6447
rect 708 6413 714 6447
rect 668 6375 714 6413
rect 668 6341 674 6375
rect 708 6341 714 6375
rect 668 6303 714 6341
rect 668 6269 674 6303
rect 708 6269 714 6303
rect 668 6231 714 6269
rect 668 6197 674 6231
rect 708 6197 714 6231
rect 668 6159 714 6197
rect 668 6125 674 6159
rect 708 6125 714 6159
rect 668 6087 714 6125
rect 668 6053 674 6087
rect 708 6053 714 6087
rect 668 6015 714 6053
rect 668 5981 674 6015
rect 708 5981 714 6015
rect 668 5943 714 5981
rect 668 5909 674 5943
rect 708 5909 714 5943
rect 668 5871 714 5909
rect 668 5837 674 5871
rect 708 5837 714 5871
rect 668 5799 714 5837
rect 668 5765 674 5799
rect 708 5765 714 5799
rect 668 5727 714 5765
rect 668 5693 674 5727
rect 708 5693 714 5727
rect 668 5655 714 5693
rect 668 5621 674 5655
rect 708 5621 714 5655
rect 668 5606 714 5621
rect 764 6591 810 6606
rect 764 6557 770 6591
rect 804 6557 810 6591
rect 764 6519 810 6557
rect 764 6485 770 6519
rect 804 6485 810 6519
rect 764 6447 810 6485
rect 764 6413 770 6447
rect 804 6413 810 6447
rect 764 6375 810 6413
rect 764 6341 770 6375
rect 804 6341 810 6375
rect 764 6303 810 6341
rect 764 6269 770 6303
rect 804 6269 810 6303
rect 764 6231 810 6269
rect 764 6197 770 6231
rect 804 6197 810 6231
rect 764 6159 810 6197
rect 764 6125 770 6159
rect 804 6125 810 6159
rect 764 6087 810 6125
rect 764 6053 770 6087
rect 804 6053 810 6087
rect 764 6015 810 6053
rect 764 5981 770 6015
rect 804 5981 810 6015
rect 764 5943 810 5981
rect 764 5909 770 5943
rect 804 5909 810 5943
rect 764 5871 810 5909
rect 764 5837 770 5871
rect 804 5837 810 5871
rect 764 5799 810 5837
rect 764 5765 770 5799
rect 804 5765 810 5799
rect 764 5727 810 5765
rect 764 5693 770 5727
rect 804 5693 810 5727
rect 764 5655 810 5693
rect 764 5621 770 5655
rect 804 5621 810 5655
rect 764 5606 810 5621
rect 860 6591 906 6606
rect 860 6557 866 6591
rect 900 6557 906 6591
rect 860 6519 906 6557
rect 860 6485 866 6519
rect 900 6485 906 6519
rect 860 6447 906 6485
rect 860 6413 866 6447
rect 900 6413 906 6447
rect 860 6375 906 6413
rect 860 6341 866 6375
rect 900 6341 906 6375
rect 860 6303 906 6341
rect 860 6269 866 6303
rect 900 6269 906 6303
rect 860 6231 906 6269
rect 860 6197 866 6231
rect 900 6197 906 6231
rect 860 6159 906 6197
rect 860 6125 866 6159
rect 900 6125 906 6159
rect 860 6087 906 6125
rect 860 6053 866 6087
rect 900 6053 906 6087
rect 860 6015 906 6053
rect 860 5981 866 6015
rect 900 5981 906 6015
rect 860 5943 906 5981
rect 860 5909 866 5943
rect 900 5909 906 5943
rect 860 5871 906 5909
rect 860 5837 866 5871
rect 900 5837 906 5871
rect 860 5799 906 5837
rect 860 5765 866 5799
rect 900 5765 906 5799
rect 860 5727 906 5765
rect 860 5693 866 5727
rect 900 5693 906 5727
rect 860 5655 906 5693
rect 860 5621 866 5655
rect 900 5621 906 5655
rect 860 5606 906 5621
rect 956 6591 1002 6606
rect 956 6557 962 6591
rect 996 6557 1002 6591
rect 956 6519 1002 6557
rect 956 6485 962 6519
rect 996 6485 1002 6519
rect 956 6447 1002 6485
rect 956 6413 962 6447
rect 996 6413 1002 6447
rect 956 6375 1002 6413
rect 956 6341 962 6375
rect 996 6341 1002 6375
rect 956 6303 1002 6341
rect 956 6269 962 6303
rect 996 6269 1002 6303
rect 956 6231 1002 6269
rect 956 6197 962 6231
rect 996 6197 1002 6231
rect 956 6159 1002 6197
rect 956 6125 962 6159
rect 996 6125 1002 6159
rect 956 6087 1002 6125
rect 956 6053 962 6087
rect 996 6053 1002 6087
rect 956 6015 1002 6053
rect 956 5981 962 6015
rect 996 5981 1002 6015
rect 956 5943 1002 5981
rect 956 5909 962 5943
rect 996 5909 1002 5943
rect 956 5871 1002 5909
rect 956 5837 962 5871
rect 996 5837 1002 5871
rect 956 5799 1002 5837
rect 956 5765 962 5799
rect 996 5765 1002 5799
rect 956 5727 1002 5765
rect 956 5693 962 5727
rect 996 5693 1002 5727
rect 956 5655 1002 5693
rect 956 5621 962 5655
rect 996 5621 1002 5655
rect 956 5606 1002 5621
rect 1052 6591 1098 6606
rect 1052 6557 1058 6591
rect 1092 6557 1098 6591
rect 1052 6519 1098 6557
rect 1052 6485 1058 6519
rect 1092 6485 1098 6519
rect 1052 6447 1098 6485
rect 1052 6413 1058 6447
rect 1092 6413 1098 6447
rect 1052 6375 1098 6413
rect 1052 6341 1058 6375
rect 1092 6341 1098 6375
rect 1052 6303 1098 6341
rect 1052 6269 1058 6303
rect 1092 6269 1098 6303
rect 1052 6231 1098 6269
rect 1052 6197 1058 6231
rect 1092 6197 1098 6231
rect 1052 6159 1098 6197
rect 1052 6125 1058 6159
rect 1092 6125 1098 6159
rect 1052 6087 1098 6125
rect 1052 6053 1058 6087
rect 1092 6053 1098 6087
rect 1052 6015 1098 6053
rect 1052 5981 1058 6015
rect 1092 5981 1098 6015
rect 1052 5943 1098 5981
rect 1052 5909 1058 5943
rect 1092 5909 1098 5943
rect 1052 5871 1098 5909
rect 1052 5837 1058 5871
rect 1092 5837 1098 5871
rect 1052 5799 1098 5837
rect 1052 5765 1058 5799
rect 1092 5765 1098 5799
rect 1052 5727 1098 5765
rect 1052 5693 1058 5727
rect 1092 5693 1098 5727
rect 1052 5655 1098 5693
rect 1052 5621 1058 5655
rect 1092 5621 1098 5655
rect 1052 5606 1098 5621
rect 1148 6591 1194 6606
rect 1148 6557 1154 6591
rect 1188 6557 1194 6591
rect 1148 6519 1194 6557
rect 1148 6485 1154 6519
rect 1188 6485 1194 6519
rect 1148 6447 1194 6485
rect 1148 6413 1154 6447
rect 1188 6413 1194 6447
rect 1148 6375 1194 6413
rect 1148 6341 1154 6375
rect 1188 6341 1194 6375
rect 1148 6303 1194 6341
rect 1148 6269 1154 6303
rect 1188 6269 1194 6303
rect 1148 6231 1194 6269
rect 1148 6197 1154 6231
rect 1188 6197 1194 6231
rect 1148 6159 1194 6197
rect 1148 6125 1154 6159
rect 1188 6125 1194 6159
rect 1148 6087 1194 6125
rect 1148 6053 1154 6087
rect 1188 6053 1194 6087
rect 1148 6015 1194 6053
rect 1148 5981 1154 6015
rect 1188 5981 1194 6015
rect 1148 5943 1194 5981
rect 1148 5909 1154 5943
rect 1188 5909 1194 5943
rect 1148 5871 1194 5909
rect 1148 5837 1154 5871
rect 1188 5837 1194 5871
rect 1148 5799 1194 5837
rect 1148 5765 1154 5799
rect 1188 5765 1194 5799
rect 1148 5727 1194 5765
rect 1148 5693 1154 5727
rect 1188 5693 1194 5727
rect 1148 5655 1194 5693
rect 1148 5621 1154 5655
rect 1188 5621 1194 5655
rect 1148 5606 1194 5621
rect 1244 6591 1290 6606
rect 1244 6557 1250 6591
rect 1284 6557 1290 6591
rect 1244 6519 1290 6557
rect 1244 6485 1250 6519
rect 1284 6485 1290 6519
rect 1244 6447 1290 6485
rect 1244 6413 1250 6447
rect 1284 6413 1290 6447
rect 1244 6375 1290 6413
rect 1244 6341 1250 6375
rect 1284 6341 1290 6375
rect 1244 6303 1290 6341
rect 1244 6269 1250 6303
rect 1284 6269 1290 6303
rect 1244 6231 1290 6269
rect 1244 6197 1250 6231
rect 1284 6197 1290 6231
rect 1244 6159 1290 6197
rect 1244 6125 1250 6159
rect 1284 6125 1290 6159
rect 1244 6087 1290 6125
rect 1244 6053 1250 6087
rect 1284 6053 1290 6087
rect 1244 6015 1290 6053
rect 1244 5981 1250 6015
rect 1284 5981 1290 6015
rect 1244 5943 1290 5981
rect 1244 5909 1250 5943
rect 1284 5909 1290 5943
rect 1244 5871 1290 5909
rect 1244 5837 1250 5871
rect 1284 5837 1290 5871
rect 1244 5799 1290 5837
rect 1244 5765 1250 5799
rect 1284 5765 1290 5799
rect 1244 5727 1290 5765
rect 1244 5693 1250 5727
rect 1284 5693 1290 5727
rect 1244 5655 1290 5693
rect 1244 5621 1250 5655
rect 1284 5621 1290 5655
rect 1244 5606 1290 5621
rect 1340 6591 1386 6606
rect 1340 6557 1346 6591
rect 1380 6557 1386 6591
rect 1340 6519 1386 6557
rect 1340 6485 1346 6519
rect 1380 6485 1386 6519
rect 1340 6447 1386 6485
rect 1340 6413 1346 6447
rect 1380 6413 1386 6447
rect 1340 6375 1386 6413
rect 1340 6341 1346 6375
rect 1380 6341 1386 6375
rect 1340 6303 1386 6341
rect 1340 6269 1346 6303
rect 1380 6269 1386 6303
rect 1340 6231 1386 6269
rect 1340 6197 1346 6231
rect 1380 6197 1386 6231
rect 1340 6159 1386 6197
rect 1340 6125 1346 6159
rect 1380 6125 1386 6159
rect 1340 6087 1386 6125
rect 1340 6053 1346 6087
rect 1380 6053 1386 6087
rect 1340 6015 1386 6053
rect 1340 5981 1346 6015
rect 1380 5981 1386 6015
rect 1340 5943 1386 5981
rect 1340 5909 1346 5943
rect 1380 5909 1386 5943
rect 1340 5871 1386 5909
rect 1340 5837 1346 5871
rect 1380 5837 1386 5871
rect 1340 5799 1386 5837
rect 1340 5765 1346 5799
rect 1380 5765 1386 5799
rect 1340 5727 1386 5765
rect 1340 5693 1346 5727
rect 1380 5693 1386 5727
rect 1340 5655 1386 5693
rect 1340 5621 1346 5655
rect 1380 5621 1386 5655
rect 1340 5606 1386 5621
rect 1954 6587 2000 6602
rect 1954 6553 1960 6587
rect 1994 6553 2000 6587
rect 1954 6515 2000 6553
rect 1954 6481 1960 6515
rect 1994 6481 2000 6515
rect 1954 6443 2000 6481
rect 1954 6409 1960 6443
rect 1994 6409 2000 6443
rect 1954 6371 2000 6409
rect 1954 6337 1960 6371
rect 1994 6337 2000 6371
rect 1954 6299 2000 6337
rect 1954 6265 1960 6299
rect 1994 6265 2000 6299
rect 1954 6227 2000 6265
rect 1954 6193 1960 6227
rect 1994 6193 2000 6227
rect 1954 6155 2000 6193
rect 1954 6121 1960 6155
rect 1994 6121 2000 6155
rect 1954 6083 2000 6121
rect 1954 6049 1960 6083
rect 1994 6049 2000 6083
rect 1954 6011 2000 6049
rect 1954 5977 1960 6011
rect 1994 5977 2000 6011
rect 1954 5939 2000 5977
rect 1954 5905 1960 5939
rect 1994 5905 2000 5939
rect 1954 5867 2000 5905
rect 1954 5833 1960 5867
rect 1994 5833 2000 5867
rect 1954 5795 2000 5833
rect 1954 5761 1960 5795
rect 1994 5761 2000 5795
rect 1954 5723 2000 5761
rect 1954 5689 1960 5723
rect 1994 5689 2000 5723
rect 1954 5651 2000 5689
rect 1954 5617 1960 5651
rect 1994 5617 2000 5651
rect 1954 5602 2000 5617
rect 2050 6587 2096 6602
rect 2050 6553 2056 6587
rect 2090 6553 2096 6587
rect 2050 6515 2096 6553
rect 2050 6481 2056 6515
rect 2090 6481 2096 6515
rect 2050 6443 2096 6481
rect 2050 6409 2056 6443
rect 2090 6409 2096 6443
rect 2050 6371 2096 6409
rect 2050 6337 2056 6371
rect 2090 6337 2096 6371
rect 2050 6299 2096 6337
rect 2050 6265 2056 6299
rect 2090 6265 2096 6299
rect 2050 6227 2096 6265
rect 2050 6193 2056 6227
rect 2090 6193 2096 6227
rect 2050 6155 2096 6193
rect 2050 6121 2056 6155
rect 2090 6121 2096 6155
rect 2050 6083 2096 6121
rect 2050 6049 2056 6083
rect 2090 6049 2096 6083
rect 2050 6011 2096 6049
rect 2050 5977 2056 6011
rect 2090 5977 2096 6011
rect 2050 5939 2096 5977
rect 2050 5905 2056 5939
rect 2090 5905 2096 5939
rect 2050 5867 2096 5905
rect 2050 5833 2056 5867
rect 2090 5833 2096 5867
rect 2050 5795 2096 5833
rect 2050 5761 2056 5795
rect 2090 5761 2096 5795
rect 2050 5723 2096 5761
rect 2050 5689 2056 5723
rect 2090 5689 2096 5723
rect 2050 5651 2096 5689
rect 2050 5617 2056 5651
rect 2090 5617 2096 5651
rect 2050 5602 2096 5617
rect 2146 6587 2192 6602
rect 2146 6553 2152 6587
rect 2186 6553 2192 6587
rect 2146 6515 2192 6553
rect 2146 6481 2152 6515
rect 2186 6481 2192 6515
rect 2146 6443 2192 6481
rect 2146 6409 2152 6443
rect 2186 6409 2192 6443
rect 2146 6371 2192 6409
rect 2146 6337 2152 6371
rect 2186 6337 2192 6371
rect 2146 6299 2192 6337
rect 2146 6265 2152 6299
rect 2186 6265 2192 6299
rect 2146 6227 2192 6265
rect 2146 6193 2152 6227
rect 2186 6193 2192 6227
rect 2146 6155 2192 6193
rect 2146 6121 2152 6155
rect 2186 6121 2192 6155
rect 2146 6083 2192 6121
rect 2146 6049 2152 6083
rect 2186 6049 2192 6083
rect 2146 6011 2192 6049
rect 2146 5977 2152 6011
rect 2186 5977 2192 6011
rect 2146 5939 2192 5977
rect 2146 5905 2152 5939
rect 2186 5905 2192 5939
rect 2146 5867 2192 5905
rect 2146 5833 2152 5867
rect 2186 5833 2192 5867
rect 2146 5795 2192 5833
rect 2146 5761 2152 5795
rect 2186 5761 2192 5795
rect 2146 5723 2192 5761
rect 2146 5689 2152 5723
rect 2186 5689 2192 5723
rect 2146 5651 2192 5689
rect 2146 5617 2152 5651
rect 2186 5617 2192 5651
rect 2146 5602 2192 5617
rect 2242 6587 2288 6602
rect 2242 6553 2248 6587
rect 2282 6553 2288 6587
rect 2242 6515 2288 6553
rect 2242 6481 2248 6515
rect 2282 6481 2288 6515
rect 2242 6443 2288 6481
rect 2242 6409 2248 6443
rect 2282 6409 2288 6443
rect 2242 6371 2288 6409
rect 2242 6337 2248 6371
rect 2282 6337 2288 6371
rect 2242 6299 2288 6337
rect 2242 6265 2248 6299
rect 2282 6265 2288 6299
rect 2242 6227 2288 6265
rect 2242 6193 2248 6227
rect 2282 6193 2288 6227
rect 2242 6155 2288 6193
rect 2242 6121 2248 6155
rect 2282 6121 2288 6155
rect 2242 6083 2288 6121
rect 2242 6049 2248 6083
rect 2282 6049 2288 6083
rect 2242 6011 2288 6049
rect 2242 5977 2248 6011
rect 2282 5977 2288 6011
rect 2242 5939 2288 5977
rect 2242 5905 2248 5939
rect 2282 5905 2288 5939
rect 2242 5867 2288 5905
rect 2242 5833 2248 5867
rect 2282 5833 2288 5867
rect 2242 5795 2288 5833
rect 2242 5761 2248 5795
rect 2282 5761 2288 5795
rect 2242 5723 2288 5761
rect 2242 5689 2248 5723
rect 2282 5689 2288 5723
rect 2242 5651 2288 5689
rect 2242 5617 2248 5651
rect 2282 5617 2288 5651
rect 2242 5602 2288 5617
rect 2338 6587 2384 6602
rect 2338 6553 2344 6587
rect 2378 6553 2384 6587
rect 2338 6515 2384 6553
rect 2338 6481 2344 6515
rect 2378 6481 2384 6515
rect 2338 6443 2384 6481
rect 2338 6409 2344 6443
rect 2378 6409 2384 6443
rect 2338 6371 2384 6409
rect 2338 6337 2344 6371
rect 2378 6337 2384 6371
rect 2338 6299 2384 6337
rect 2338 6265 2344 6299
rect 2378 6265 2384 6299
rect 2338 6227 2384 6265
rect 2338 6193 2344 6227
rect 2378 6193 2384 6227
rect 2338 6155 2384 6193
rect 2338 6121 2344 6155
rect 2378 6121 2384 6155
rect 2338 6083 2384 6121
rect 2338 6049 2344 6083
rect 2378 6049 2384 6083
rect 2338 6011 2384 6049
rect 2338 5977 2344 6011
rect 2378 5977 2384 6011
rect 2338 5939 2384 5977
rect 2338 5905 2344 5939
rect 2378 5905 2384 5939
rect 2338 5867 2384 5905
rect 2338 5833 2344 5867
rect 2378 5833 2384 5867
rect 2338 5795 2384 5833
rect 2338 5761 2344 5795
rect 2378 5761 2384 5795
rect 2338 5723 2384 5761
rect 2338 5689 2344 5723
rect 2378 5689 2384 5723
rect 2338 5651 2384 5689
rect 2338 5617 2344 5651
rect 2378 5617 2384 5651
rect 2338 5602 2384 5617
rect 2434 6587 2480 6602
rect 2434 6553 2440 6587
rect 2474 6553 2480 6587
rect 2434 6515 2480 6553
rect 2434 6481 2440 6515
rect 2474 6481 2480 6515
rect 2434 6443 2480 6481
rect 2434 6409 2440 6443
rect 2474 6409 2480 6443
rect 2434 6371 2480 6409
rect 2434 6337 2440 6371
rect 2474 6337 2480 6371
rect 2434 6299 2480 6337
rect 2434 6265 2440 6299
rect 2474 6265 2480 6299
rect 2434 6227 2480 6265
rect 2434 6193 2440 6227
rect 2474 6193 2480 6227
rect 2434 6155 2480 6193
rect 2434 6121 2440 6155
rect 2474 6121 2480 6155
rect 2434 6083 2480 6121
rect 2434 6049 2440 6083
rect 2474 6049 2480 6083
rect 2434 6011 2480 6049
rect 2434 5977 2440 6011
rect 2474 5977 2480 6011
rect 2434 5939 2480 5977
rect 2434 5905 2440 5939
rect 2474 5905 2480 5939
rect 2434 5867 2480 5905
rect 2434 5833 2440 5867
rect 2474 5833 2480 5867
rect 2434 5795 2480 5833
rect 2434 5761 2440 5795
rect 2474 5761 2480 5795
rect 2434 5723 2480 5761
rect 2434 5689 2440 5723
rect 2474 5689 2480 5723
rect 2434 5651 2480 5689
rect 2434 5617 2440 5651
rect 2474 5617 2480 5651
rect 2434 5602 2480 5617
rect 2530 6587 2576 6602
rect 2530 6553 2536 6587
rect 2570 6553 2576 6587
rect 2530 6515 2576 6553
rect 2530 6481 2536 6515
rect 2570 6481 2576 6515
rect 2530 6443 2576 6481
rect 2530 6409 2536 6443
rect 2570 6409 2576 6443
rect 2530 6371 2576 6409
rect 2530 6337 2536 6371
rect 2570 6337 2576 6371
rect 2530 6299 2576 6337
rect 2530 6265 2536 6299
rect 2570 6265 2576 6299
rect 2530 6227 2576 6265
rect 2530 6193 2536 6227
rect 2570 6193 2576 6227
rect 2530 6155 2576 6193
rect 2530 6121 2536 6155
rect 2570 6121 2576 6155
rect 2530 6083 2576 6121
rect 2530 6049 2536 6083
rect 2570 6049 2576 6083
rect 2530 6011 2576 6049
rect 2530 5977 2536 6011
rect 2570 5977 2576 6011
rect 2530 5939 2576 5977
rect 2530 5905 2536 5939
rect 2570 5905 2576 5939
rect 2530 5867 2576 5905
rect 2530 5833 2536 5867
rect 2570 5833 2576 5867
rect 2530 5795 2576 5833
rect 2530 5761 2536 5795
rect 2570 5761 2576 5795
rect 2530 5723 2576 5761
rect 2530 5689 2536 5723
rect 2570 5689 2576 5723
rect 2530 5651 2576 5689
rect 2530 5617 2536 5651
rect 2570 5617 2576 5651
rect 2530 5602 2576 5617
rect 2626 6587 2672 6602
rect 2626 6553 2632 6587
rect 2666 6553 2672 6587
rect 2626 6515 2672 6553
rect 2626 6481 2632 6515
rect 2666 6481 2672 6515
rect 2626 6443 2672 6481
rect 2626 6409 2632 6443
rect 2666 6409 2672 6443
rect 2626 6371 2672 6409
rect 2626 6337 2632 6371
rect 2666 6337 2672 6371
rect 2626 6299 2672 6337
rect 2626 6265 2632 6299
rect 2666 6265 2672 6299
rect 2626 6227 2672 6265
rect 2626 6193 2632 6227
rect 2666 6193 2672 6227
rect 2626 6155 2672 6193
rect 2626 6121 2632 6155
rect 2666 6121 2672 6155
rect 2626 6083 2672 6121
rect 2626 6049 2632 6083
rect 2666 6049 2672 6083
rect 2626 6011 2672 6049
rect 2626 5977 2632 6011
rect 2666 5977 2672 6011
rect 2626 5939 2672 5977
rect 2626 5905 2632 5939
rect 2666 5905 2672 5939
rect 2626 5867 2672 5905
rect 2626 5833 2632 5867
rect 2666 5833 2672 5867
rect 2626 5795 2672 5833
rect 2626 5761 2632 5795
rect 2666 5761 2672 5795
rect 2626 5723 2672 5761
rect 2626 5689 2632 5723
rect 2666 5689 2672 5723
rect 2626 5651 2672 5689
rect 2626 5617 2632 5651
rect 2666 5617 2672 5651
rect 2626 5602 2672 5617
rect 2722 6587 2768 6602
rect 2722 6553 2728 6587
rect 2762 6553 2768 6587
rect 2722 6515 2768 6553
rect 2722 6481 2728 6515
rect 2762 6481 2768 6515
rect 2722 6443 2768 6481
rect 2722 6409 2728 6443
rect 2762 6409 2768 6443
rect 2722 6371 2768 6409
rect 2722 6337 2728 6371
rect 2762 6337 2768 6371
rect 2722 6299 2768 6337
rect 2722 6265 2728 6299
rect 2762 6265 2768 6299
rect 2722 6227 2768 6265
rect 2722 6193 2728 6227
rect 2762 6193 2768 6227
rect 2722 6155 2768 6193
rect 2722 6121 2728 6155
rect 2762 6121 2768 6155
rect 2722 6083 2768 6121
rect 2722 6049 2728 6083
rect 2762 6049 2768 6083
rect 2722 6011 2768 6049
rect 2722 5977 2728 6011
rect 2762 5977 2768 6011
rect 2722 5939 2768 5977
rect 2722 5905 2728 5939
rect 2762 5905 2768 5939
rect 2722 5867 2768 5905
rect 2722 5833 2728 5867
rect 2762 5833 2768 5867
rect 2722 5795 2768 5833
rect 2722 5761 2728 5795
rect 2762 5761 2768 5795
rect 2722 5723 2768 5761
rect 2722 5689 2728 5723
rect 2762 5689 2768 5723
rect 2722 5651 2768 5689
rect 2722 5617 2728 5651
rect 2762 5617 2768 5651
rect 2722 5602 2768 5617
rect 3144 6575 3190 6590
rect 3144 6541 3150 6575
rect 3184 6541 3190 6575
rect 3144 6503 3190 6541
rect 3144 6469 3150 6503
rect 3184 6469 3190 6503
rect 3144 6431 3190 6469
rect 3144 6397 3150 6431
rect 3184 6397 3190 6431
rect 3144 6359 3190 6397
rect 3144 6325 3150 6359
rect 3184 6325 3190 6359
rect 3144 6287 3190 6325
rect 3144 6253 3150 6287
rect 3184 6253 3190 6287
rect 3144 6215 3190 6253
rect 3144 6181 3150 6215
rect 3184 6181 3190 6215
rect 3144 6143 3190 6181
rect 3144 6109 3150 6143
rect 3184 6109 3190 6143
rect 3144 6071 3190 6109
rect 3144 6037 3150 6071
rect 3184 6037 3190 6071
rect 3144 5999 3190 6037
rect 3144 5965 3150 5999
rect 3184 5965 3190 5999
rect 3144 5927 3190 5965
rect 3144 5893 3150 5927
rect 3184 5893 3190 5927
rect 3144 5855 3190 5893
rect 3144 5821 3150 5855
rect 3184 5821 3190 5855
rect 3144 5783 3190 5821
rect 3144 5749 3150 5783
rect 3184 5749 3190 5783
rect 3144 5711 3190 5749
rect 3144 5677 3150 5711
rect 3184 5677 3190 5711
rect 3144 5639 3190 5677
rect 3144 5605 3150 5639
rect 3184 5605 3190 5639
rect 3144 5590 3190 5605
rect 3240 6575 3286 6590
rect 3240 6541 3246 6575
rect 3280 6541 3286 6575
rect 3240 6503 3286 6541
rect 3240 6469 3246 6503
rect 3280 6469 3286 6503
rect 3240 6431 3286 6469
rect 3240 6397 3246 6431
rect 3280 6397 3286 6431
rect 3240 6359 3286 6397
rect 3240 6325 3246 6359
rect 3280 6325 3286 6359
rect 3240 6287 3286 6325
rect 3240 6253 3246 6287
rect 3280 6253 3286 6287
rect 3240 6215 3286 6253
rect 3240 6181 3246 6215
rect 3280 6181 3286 6215
rect 3240 6143 3286 6181
rect 3240 6109 3246 6143
rect 3280 6109 3286 6143
rect 3240 6071 3286 6109
rect 3240 6037 3246 6071
rect 3280 6037 3286 6071
rect 3240 5999 3286 6037
rect 3240 5965 3246 5999
rect 3280 5965 3286 5999
rect 3240 5927 3286 5965
rect 3240 5893 3246 5927
rect 3280 5893 3286 5927
rect 3240 5855 3286 5893
rect 3240 5821 3246 5855
rect 3280 5821 3286 5855
rect 3240 5783 3286 5821
rect 3240 5749 3246 5783
rect 3280 5749 3286 5783
rect 3240 5711 3286 5749
rect 3240 5677 3246 5711
rect 3280 5677 3286 5711
rect 3240 5639 3286 5677
rect 3240 5605 3246 5639
rect 3280 5605 3286 5639
rect 3240 5590 3286 5605
rect 3336 6575 3382 6590
rect 3336 6541 3342 6575
rect 3376 6541 3382 6575
rect 3336 6503 3382 6541
rect 3336 6469 3342 6503
rect 3376 6469 3382 6503
rect 3336 6431 3382 6469
rect 3336 6397 3342 6431
rect 3376 6397 3382 6431
rect 3336 6359 3382 6397
rect 3336 6325 3342 6359
rect 3376 6325 3382 6359
rect 3336 6287 3382 6325
rect 3336 6253 3342 6287
rect 3376 6253 3382 6287
rect 3336 6215 3382 6253
rect 3336 6181 3342 6215
rect 3376 6181 3382 6215
rect 3336 6143 3382 6181
rect 3336 6109 3342 6143
rect 3376 6109 3382 6143
rect 3336 6071 3382 6109
rect 3336 6037 3342 6071
rect 3376 6037 3382 6071
rect 3336 5999 3382 6037
rect 3336 5965 3342 5999
rect 3376 5965 3382 5999
rect 3336 5927 3382 5965
rect 3336 5893 3342 5927
rect 3376 5893 3382 5927
rect 3336 5855 3382 5893
rect 3336 5821 3342 5855
rect 3376 5821 3382 5855
rect 3336 5783 3382 5821
rect 3336 5749 3342 5783
rect 3376 5749 3382 5783
rect 3336 5711 3382 5749
rect 3336 5677 3342 5711
rect 3376 5677 3382 5711
rect 3336 5639 3382 5677
rect 3336 5605 3342 5639
rect 3376 5605 3382 5639
rect 3336 5590 3382 5605
rect 3432 6575 3478 6590
rect 3432 6541 3438 6575
rect 3472 6541 3478 6575
rect 3432 6503 3478 6541
rect 3432 6469 3438 6503
rect 3472 6469 3478 6503
rect 3432 6431 3478 6469
rect 3432 6397 3438 6431
rect 3472 6397 3478 6431
rect 3432 6359 3478 6397
rect 3432 6325 3438 6359
rect 3472 6325 3478 6359
rect 3432 6287 3478 6325
rect 3432 6253 3438 6287
rect 3472 6253 3478 6287
rect 3432 6215 3478 6253
rect 3432 6181 3438 6215
rect 3472 6181 3478 6215
rect 3432 6143 3478 6181
rect 3432 6109 3438 6143
rect 3472 6109 3478 6143
rect 3432 6071 3478 6109
rect 3432 6037 3438 6071
rect 3472 6037 3478 6071
rect 3432 5999 3478 6037
rect 3432 5965 3438 5999
rect 3472 5965 3478 5999
rect 3432 5927 3478 5965
rect 3432 5893 3438 5927
rect 3472 5893 3478 5927
rect 3432 5855 3478 5893
rect 3432 5821 3438 5855
rect 3472 5821 3478 5855
rect 3432 5783 3478 5821
rect 3432 5749 3438 5783
rect 3472 5749 3478 5783
rect 3432 5711 3478 5749
rect 3432 5677 3438 5711
rect 3472 5677 3478 5711
rect 3432 5639 3478 5677
rect 3432 5605 3438 5639
rect 3472 5605 3478 5639
rect 3432 5590 3478 5605
rect 3528 6575 3574 6590
rect 3528 6541 3534 6575
rect 3568 6541 3574 6575
rect 3528 6503 3574 6541
rect 3528 6469 3534 6503
rect 3568 6469 3574 6503
rect 3528 6431 3574 6469
rect 3528 6397 3534 6431
rect 3568 6397 3574 6431
rect 3528 6359 3574 6397
rect 3528 6325 3534 6359
rect 3568 6325 3574 6359
rect 3528 6287 3574 6325
rect 3528 6253 3534 6287
rect 3568 6253 3574 6287
rect 3528 6215 3574 6253
rect 3528 6181 3534 6215
rect 3568 6181 3574 6215
rect 3528 6143 3574 6181
rect 3528 6109 3534 6143
rect 3568 6109 3574 6143
rect 3528 6071 3574 6109
rect 3528 6037 3534 6071
rect 3568 6037 3574 6071
rect 3528 5999 3574 6037
rect 3528 5965 3534 5999
rect 3568 5965 3574 5999
rect 3528 5927 3574 5965
rect 3528 5893 3534 5927
rect 3568 5893 3574 5927
rect 3528 5855 3574 5893
rect 3528 5821 3534 5855
rect 3568 5821 3574 5855
rect 3528 5783 3574 5821
rect 3528 5749 3534 5783
rect 3568 5749 3574 5783
rect 3528 5711 3574 5749
rect 3528 5677 3534 5711
rect 3568 5677 3574 5711
rect 3528 5639 3574 5677
rect 3528 5605 3534 5639
rect 3568 5605 3574 5639
rect 3528 5590 3574 5605
rect 3624 6575 3670 6590
rect 3624 6541 3630 6575
rect 3664 6541 3670 6575
rect 3624 6503 3670 6541
rect 3624 6469 3630 6503
rect 3664 6469 3670 6503
rect 3624 6431 3670 6469
rect 3624 6397 3630 6431
rect 3664 6397 3670 6431
rect 3624 6359 3670 6397
rect 3624 6325 3630 6359
rect 3664 6325 3670 6359
rect 3624 6287 3670 6325
rect 3624 6253 3630 6287
rect 3664 6253 3670 6287
rect 3624 6215 3670 6253
rect 3624 6181 3630 6215
rect 3664 6181 3670 6215
rect 3624 6143 3670 6181
rect 3624 6109 3630 6143
rect 3664 6109 3670 6143
rect 3624 6071 3670 6109
rect 3624 6037 3630 6071
rect 3664 6037 3670 6071
rect 3624 5999 3670 6037
rect 3624 5965 3630 5999
rect 3664 5965 3670 5999
rect 3624 5927 3670 5965
rect 3624 5893 3630 5927
rect 3664 5893 3670 5927
rect 3624 5855 3670 5893
rect 3624 5821 3630 5855
rect 3664 5821 3670 5855
rect 3624 5783 3670 5821
rect 3624 5749 3630 5783
rect 3664 5749 3670 5783
rect 3624 5711 3670 5749
rect 3624 5677 3630 5711
rect 3664 5677 3670 5711
rect 3624 5639 3670 5677
rect 3624 5605 3630 5639
rect 3664 5605 3670 5639
rect 3624 5590 3670 5605
rect 3720 6575 3766 6590
rect 3720 6541 3726 6575
rect 3760 6541 3766 6575
rect 3720 6503 3766 6541
rect 3720 6469 3726 6503
rect 3760 6469 3766 6503
rect 3720 6431 3766 6469
rect 3720 6397 3726 6431
rect 3760 6397 3766 6431
rect 3720 6359 3766 6397
rect 3720 6325 3726 6359
rect 3760 6325 3766 6359
rect 3720 6287 3766 6325
rect 3720 6253 3726 6287
rect 3760 6253 3766 6287
rect 3720 6215 3766 6253
rect 3720 6181 3726 6215
rect 3760 6181 3766 6215
rect 3720 6143 3766 6181
rect 3720 6109 3726 6143
rect 3760 6109 3766 6143
rect 3720 6071 3766 6109
rect 3720 6037 3726 6071
rect 3760 6037 3766 6071
rect 3720 5999 3766 6037
rect 3720 5965 3726 5999
rect 3760 5965 3766 5999
rect 3720 5927 3766 5965
rect 3720 5893 3726 5927
rect 3760 5893 3766 5927
rect 3720 5855 3766 5893
rect 3720 5821 3726 5855
rect 3760 5821 3766 5855
rect 3720 5783 3766 5821
rect 3720 5749 3726 5783
rect 3760 5749 3766 5783
rect 3720 5711 3766 5749
rect 3720 5677 3726 5711
rect 3760 5677 3766 5711
rect 3720 5639 3766 5677
rect 3720 5605 3726 5639
rect 3760 5605 3766 5639
rect 3720 5590 3766 5605
rect 3816 6575 3862 6590
rect 3816 6541 3822 6575
rect 3856 6541 3862 6575
rect 3816 6503 3862 6541
rect 3816 6469 3822 6503
rect 3856 6469 3862 6503
rect 3816 6431 3862 6469
rect 3816 6397 3822 6431
rect 3856 6397 3862 6431
rect 3816 6359 3862 6397
rect 3816 6325 3822 6359
rect 3856 6325 3862 6359
rect 3816 6287 3862 6325
rect 3816 6253 3822 6287
rect 3856 6253 3862 6287
rect 3816 6215 3862 6253
rect 3816 6181 3822 6215
rect 3856 6181 3862 6215
rect 3816 6143 3862 6181
rect 3816 6109 3822 6143
rect 3856 6109 3862 6143
rect 3816 6071 3862 6109
rect 3816 6037 3822 6071
rect 3856 6037 3862 6071
rect 3816 5999 3862 6037
rect 3816 5965 3822 5999
rect 3856 5965 3862 5999
rect 3816 5927 3862 5965
rect 3816 5893 3822 5927
rect 3856 5893 3862 5927
rect 3816 5855 3862 5893
rect 3816 5821 3822 5855
rect 3856 5821 3862 5855
rect 3816 5783 3862 5821
rect 3816 5749 3822 5783
rect 3856 5749 3862 5783
rect 3816 5711 3862 5749
rect 3816 5677 3822 5711
rect 3856 5677 3862 5711
rect 3816 5639 3862 5677
rect 3816 5605 3822 5639
rect 3856 5605 3862 5639
rect 3816 5590 3862 5605
rect 3912 6575 3958 6590
rect 3912 6541 3918 6575
rect 3952 6541 3958 6575
rect 3912 6503 3958 6541
rect 3912 6469 3918 6503
rect 3952 6469 3958 6503
rect 3912 6431 3958 6469
rect 3912 6397 3918 6431
rect 3952 6397 3958 6431
rect 3912 6359 3958 6397
rect 3912 6325 3918 6359
rect 3952 6325 3958 6359
rect 3912 6287 3958 6325
rect 3912 6253 3918 6287
rect 3952 6253 3958 6287
rect 3912 6215 3958 6253
rect 3912 6181 3918 6215
rect 3952 6181 3958 6215
rect 3912 6143 3958 6181
rect 3912 6109 3918 6143
rect 3952 6109 3958 6143
rect 3912 6071 3958 6109
rect 3912 6037 3918 6071
rect 3952 6037 3958 6071
rect 3912 5999 3958 6037
rect 3912 5965 3918 5999
rect 3952 5965 3958 5999
rect 3912 5927 3958 5965
rect 3912 5893 3918 5927
rect 3952 5893 3958 5927
rect 3912 5855 3958 5893
rect 3912 5821 3918 5855
rect 3952 5821 3958 5855
rect 3912 5783 3958 5821
rect 3912 5749 3918 5783
rect 3952 5749 3958 5783
rect 3912 5711 3958 5749
rect 3912 5677 3918 5711
rect 3952 5677 3958 5711
rect 3912 5639 3958 5677
rect 3912 5605 3918 5639
rect 3952 5605 3958 5639
rect 3912 5590 3958 5605
rect 4008 6575 4054 6590
rect 4008 6541 4014 6575
rect 4048 6541 4054 6575
rect 4008 6503 4054 6541
rect 4008 6469 4014 6503
rect 4048 6469 4054 6503
rect 4008 6431 4054 6469
rect 4008 6397 4014 6431
rect 4048 6397 4054 6431
rect 4008 6359 4054 6397
rect 4008 6325 4014 6359
rect 4048 6325 4054 6359
rect 4008 6287 4054 6325
rect 4008 6253 4014 6287
rect 4048 6253 4054 6287
rect 4008 6215 4054 6253
rect 4008 6181 4014 6215
rect 4048 6181 4054 6215
rect 4008 6143 4054 6181
rect 4008 6109 4014 6143
rect 4048 6109 4054 6143
rect 4008 6071 4054 6109
rect 4008 6037 4014 6071
rect 4048 6037 4054 6071
rect 4008 5999 4054 6037
rect 4008 5965 4014 5999
rect 4048 5965 4054 5999
rect 4008 5927 4054 5965
rect 4008 5893 4014 5927
rect 4048 5893 4054 5927
rect 4008 5855 4054 5893
rect 4008 5821 4014 5855
rect 4048 5821 4054 5855
rect 4008 5783 4054 5821
rect 4008 5749 4014 5783
rect 4048 5749 4054 5783
rect 4008 5711 4054 5749
rect 4008 5677 4014 5711
rect 4048 5677 4054 5711
rect 4008 5639 4054 5677
rect 4008 5605 4014 5639
rect 4048 5605 4054 5639
rect 4008 5590 4054 5605
rect 4104 6575 4150 6590
rect 4104 6541 4110 6575
rect 4144 6541 4150 6575
rect 4104 6503 4150 6541
rect 4104 6469 4110 6503
rect 4144 6469 4150 6503
rect 4104 6431 4150 6469
rect 4104 6397 4110 6431
rect 4144 6397 4150 6431
rect 4104 6359 4150 6397
rect 4104 6325 4110 6359
rect 4144 6325 4150 6359
rect 4104 6287 4150 6325
rect 4104 6253 4110 6287
rect 4144 6253 4150 6287
rect 4104 6215 4150 6253
rect 4104 6181 4110 6215
rect 4144 6181 4150 6215
rect 4104 6143 4150 6181
rect 4104 6109 4110 6143
rect 4144 6109 4150 6143
rect 4104 6071 4150 6109
rect 4104 6037 4110 6071
rect 4144 6037 4150 6071
rect 4104 5999 4150 6037
rect 4104 5965 4110 5999
rect 4144 5965 4150 5999
rect 4104 5927 4150 5965
rect 4104 5893 4110 5927
rect 4144 5893 4150 5927
rect 4104 5855 4150 5893
rect 4104 5821 4110 5855
rect 4144 5821 4150 5855
rect 4104 5783 4150 5821
rect 4104 5749 4110 5783
rect 4144 5749 4150 5783
rect 4104 5711 4150 5749
rect 4104 5677 4110 5711
rect 4144 5677 4150 5711
rect 4104 5639 4150 5677
rect 4104 5605 4110 5639
rect 4144 5605 4150 5639
rect 4104 5590 4150 5605
rect 4200 6575 4246 6590
rect 4200 6541 4206 6575
rect 4240 6541 4246 6575
rect 4200 6503 4246 6541
rect 4200 6469 4206 6503
rect 4240 6469 4246 6503
rect 4200 6431 4246 6469
rect 4200 6397 4206 6431
rect 4240 6397 4246 6431
rect 4200 6359 4246 6397
rect 4200 6325 4206 6359
rect 4240 6325 4246 6359
rect 4200 6287 4246 6325
rect 4200 6253 4206 6287
rect 4240 6253 4246 6287
rect 4200 6215 4246 6253
rect 4200 6181 4206 6215
rect 4240 6181 4246 6215
rect 4200 6143 4246 6181
rect 4200 6109 4206 6143
rect 4240 6109 4246 6143
rect 4200 6071 4246 6109
rect 4200 6037 4206 6071
rect 4240 6037 4246 6071
rect 4200 5999 4246 6037
rect 4200 5965 4206 5999
rect 4240 5965 4246 5999
rect 4200 5927 4246 5965
rect 4200 5893 4206 5927
rect 4240 5893 4246 5927
rect 4200 5855 4246 5893
rect 4200 5821 4206 5855
rect 4240 5821 4246 5855
rect 4200 5783 4246 5821
rect 4200 5749 4206 5783
rect 4240 5749 4246 5783
rect 4200 5711 4246 5749
rect 4200 5677 4206 5711
rect 4240 5677 4246 5711
rect 4200 5639 4246 5677
rect 4200 5605 4206 5639
rect 4240 5605 4246 5639
rect 4200 5590 4246 5605
rect 4296 6575 4342 6590
rect 4296 6541 4302 6575
rect 4336 6541 4342 6575
rect 4296 6503 4342 6541
rect 4296 6469 4302 6503
rect 4336 6469 4342 6503
rect 4296 6431 4342 6469
rect 4296 6397 4302 6431
rect 4336 6397 4342 6431
rect 4296 6359 4342 6397
rect 4296 6325 4302 6359
rect 4336 6325 4342 6359
rect 4296 6287 4342 6325
rect 4296 6253 4302 6287
rect 4336 6253 4342 6287
rect 4296 6215 4342 6253
rect 4296 6181 4302 6215
rect 4336 6181 4342 6215
rect 4296 6143 4342 6181
rect 4296 6109 4302 6143
rect 4336 6109 4342 6143
rect 4296 6071 4342 6109
rect 4296 6037 4302 6071
rect 4336 6037 4342 6071
rect 4296 5999 4342 6037
rect 4296 5965 4302 5999
rect 4336 5965 4342 5999
rect 4296 5927 4342 5965
rect 4296 5893 4302 5927
rect 4336 5893 4342 5927
rect 4296 5855 4342 5893
rect 4296 5821 4302 5855
rect 4336 5821 4342 5855
rect 4296 5783 4342 5821
rect 4296 5749 4302 5783
rect 4336 5749 4342 5783
rect 4296 5711 4342 5749
rect 4296 5677 4302 5711
rect 4336 5677 4342 5711
rect 4296 5639 4342 5677
rect 4296 5605 4302 5639
rect 4336 5605 4342 5639
rect 4296 5590 4342 5605
rect 4910 6571 4956 6586
rect 4910 6537 4916 6571
rect 4950 6537 4956 6571
rect 4910 6499 4956 6537
rect 4910 6465 4916 6499
rect 4950 6465 4956 6499
rect 4910 6427 4956 6465
rect 4910 6393 4916 6427
rect 4950 6393 4956 6427
rect 4910 6355 4956 6393
rect 4910 6321 4916 6355
rect 4950 6321 4956 6355
rect 4910 6283 4956 6321
rect 4910 6249 4916 6283
rect 4950 6249 4956 6283
rect 4910 6211 4956 6249
rect 4910 6177 4916 6211
rect 4950 6177 4956 6211
rect 4910 6139 4956 6177
rect 4910 6105 4916 6139
rect 4950 6105 4956 6139
rect 4910 6067 4956 6105
rect 4910 6033 4916 6067
rect 4950 6033 4956 6067
rect 4910 5995 4956 6033
rect 4910 5961 4916 5995
rect 4950 5961 4956 5995
rect 4910 5923 4956 5961
rect 4910 5889 4916 5923
rect 4950 5889 4956 5923
rect 4910 5851 4956 5889
rect 4910 5817 4916 5851
rect 4950 5817 4956 5851
rect 4910 5779 4956 5817
rect 4910 5745 4916 5779
rect 4950 5745 4956 5779
rect 4910 5707 4956 5745
rect 4910 5673 4916 5707
rect 4950 5673 4956 5707
rect 4910 5635 4956 5673
rect 4910 5601 4916 5635
rect 4950 5601 4956 5635
rect 4910 5586 4956 5601
rect 5006 6571 5052 6586
rect 5006 6537 5012 6571
rect 5046 6537 5052 6571
rect 5006 6499 5052 6537
rect 5006 6465 5012 6499
rect 5046 6465 5052 6499
rect 5006 6427 5052 6465
rect 5006 6393 5012 6427
rect 5046 6393 5052 6427
rect 5006 6355 5052 6393
rect 5006 6321 5012 6355
rect 5046 6321 5052 6355
rect 5006 6283 5052 6321
rect 5006 6249 5012 6283
rect 5046 6249 5052 6283
rect 5006 6211 5052 6249
rect 5006 6177 5012 6211
rect 5046 6177 5052 6211
rect 5006 6139 5052 6177
rect 5006 6105 5012 6139
rect 5046 6105 5052 6139
rect 5006 6067 5052 6105
rect 5006 6033 5012 6067
rect 5046 6033 5052 6067
rect 5006 5995 5052 6033
rect 5006 5961 5012 5995
rect 5046 5961 5052 5995
rect 5006 5923 5052 5961
rect 5006 5889 5012 5923
rect 5046 5889 5052 5923
rect 5006 5851 5052 5889
rect 5006 5817 5012 5851
rect 5046 5817 5052 5851
rect 5006 5779 5052 5817
rect 5006 5745 5012 5779
rect 5046 5745 5052 5779
rect 5006 5707 5052 5745
rect 5006 5673 5012 5707
rect 5046 5673 5052 5707
rect 5006 5635 5052 5673
rect 5006 5601 5012 5635
rect 5046 5601 5052 5635
rect 5006 5586 5052 5601
rect 5102 6571 5148 6586
rect 5102 6537 5108 6571
rect 5142 6537 5148 6571
rect 5102 6499 5148 6537
rect 5102 6465 5108 6499
rect 5142 6465 5148 6499
rect 5102 6427 5148 6465
rect 5102 6393 5108 6427
rect 5142 6393 5148 6427
rect 5102 6355 5148 6393
rect 5102 6321 5108 6355
rect 5142 6321 5148 6355
rect 5102 6283 5148 6321
rect 5102 6249 5108 6283
rect 5142 6249 5148 6283
rect 5102 6211 5148 6249
rect 5102 6177 5108 6211
rect 5142 6177 5148 6211
rect 5102 6139 5148 6177
rect 5102 6105 5108 6139
rect 5142 6105 5148 6139
rect 5102 6067 5148 6105
rect 5102 6033 5108 6067
rect 5142 6033 5148 6067
rect 5102 5995 5148 6033
rect 5102 5961 5108 5995
rect 5142 5961 5148 5995
rect 5102 5923 5148 5961
rect 5102 5889 5108 5923
rect 5142 5889 5148 5923
rect 5102 5851 5148 5889
rect 5102 5817 5108 5851
rect 5142 5817 5148 5851
rect 5102 5779 5148 5817
rect 5102 5745 5108 5779
rect 5142 5745 5148 5779
rect 5102 5707 5148 5745
rect 5102 5673 5108 5707
rect 5142 5673 5148 5707
rect 5102 5635 5148 5673
rect 5102 5601 5108 5635
rect 5142 5601 5148 5635
rect 5102 5586 5148 5601
rect 5198 6571 5244 6586
rect 5198 6537 5204 6571
rect 5238 6537 5244 6571
rect 5198 6499 5244 6537
rect 5198 6465 5204 6499
rect 5238 6465 5244 6499
rect 5198 6427 5244 6465
rect 5198 6393 5204 6427
rect 5238 6393 5244 6427
rect 5198 6355 5244 6393
rect 5198 6321 5204 6355
rect 5238 6321 5244 6355
rect 5198 6283 5244 6321
rect 5198 6249 5204 6283
rect 5238 6249 5244 6283
rect 5198 6211 5244 6249
rect 5198 6177 5204 6211
rect 5238 6177 5244 6211
rect 5198 6139 5244 6177
rect 5198 6105 5204 6139
rect 5238 6105 5244 6139
rect 5198 6067 5244 6105
rect 5198 6033 5204 6067
rect 5238 6033 5244 6067
rect 5198 5995 5244 6033
rect 5198 5961 5204 5995
rect 5238 5961 5244 5995
rect 5198 5923 5244 5961
rect 5198 5889 5204 5923
rect 5238 5889 5244 5923
rect 5198 5851 5244 5889
rect 5198 5817 5204 5851
rect 5238 5817 5244 5851
rect 5198 5779 5244 5817
rect 5198 5745 5204 5779
rect 5238 5745 5244 5779
rect 5198 5707 5244 5745
rect 5198 5673 5204 5707
rect 5238 5673 5244 5707
rect 5198 5635 5244 5673
rect 5198 5601 5204 5635
rect 5238 5601 5244 5635
rect 5198 5586 5244 5601
rect 5294 6571 5340 6586
rect 5294 6537 5300 6571
rect 5334 6537 5340 6571
rect 5294 6499 5340 6537
rect 5294 6465 5300 6499
rect 5334 6465 5340 6499
rect 5294 6427 5340 6465
rect 5294 6393 5300 6427
rect 5334 6393 5340 6427
rect 5294 6355 5340 6393
rect 5294 6321 5300 6355
rect 5334 6321 5340 6355
rect 5294 6283 5340 6321
rect 5294 6249 5300 6283
rect 5334 6249 5340 6283
rect 5294 6211 5340 6249
rect 5294 6177 5300 6211
rect 5334 6177 5340 6211
rect 5294 6139 5340 6177
rect 5294 6105 5300 6139
rect 5334 6105 5340 6139
rect 5294 6067 5340 6105
rect 5294 6033 5300 6067
rect 5334 6033 5340 6067
rect 5294 5995 5340 6033
rect 5294 5961 5300 5995
rect 5334 5961 5340 5995
rect 5294 5923 5340 5961
rect 5294 5889 5300 5923
rect 5334 5889 5340 5923
rect 5294 5851 5340 5889
rect 5294 5817 5300 5851
rect 5334 5817 5340 5851
rect 5294 5779 5340 5817
rect 5294 5745 5300 5779
rect 5334 5745 5340 5779
rect 5294 5707 5340 5745
rect 5294 5673 5300 5707
rect 5334 5673 5340 5707
rect 5294 5635 5340 5673
rect 5294 5601 5300 5635
rect 5334 5601 5340 5635
rect 5294 5586 5340 5601
rect 5390 6571 5436 6586
rect 5390 6537 5396 6571
rect 5430 6537 5436 6571
rect 5390 6499 5436 6537
rect 5390 6465 5396 6499
rect 5430 6465 5436 6499
rect 5390 6427 5436 6465
rect 5390 6393 5396 6427
rect 5430 6393 5436 6427
rect 5390 6355 5436 6393
rect 5390 6321 5396 6355
rect 5430 6321 5436 6355
rect 5390 6283 5436 6321
rect 5390 6249 5396 6283
rect 5430 6249 5436 6283
rect 5390 6211 5436 6249
rect 5390 6177 5396 6211
rect 5430 6177 5436 6211
rect 5390 6139 5436 6177
rect 5390 6105 5396 6139
rect 5430 6105 5436 6139
rect 5390 6067 5436 6105
rect 5390 6033 5396 6067
rect 5430 6033 5436 6067
rect 5390 5995 5436 6033
rect 5390 5961 5396 5995
rect 5430 5961 5436 5995
rect 5390 5923 5436 5961
rect 5390 5889 5396 5923
rect 5430 5889 5436 5923
rect 5390 5851 5436 5889
rect 5390 5817 5396 5851
rect 5430 5817 5436 5851
rect 5390 5779 5436 5817
rect 5390 5745 5396 5779
rect 5430 5745 5436 5779
rect 5390 5707 5436 5745
rect 5390 5673 5396 5707
rect 5430 5673 5436 5707
rect 5390 5635 5436 5673
rect 5390 5601 5396 5635
rect 5430 5601 5436 5635
rect 5390 5586 5436 5601
rect 5486 6571 5532 6586
rect 5486 6537 5492 6571
rect 5526 6537 5532 6571
rect 5486 6499 5532 6537
rect 5486 6465 5492 6499
rect 5526 6465 5532 6499
rect 5486 6427 5532 6465
rect 5486 6393 5492 6427
rect 5526 6393 5532 6427
rect 5486 6355 5532 6393
rect 5486 6321 5492 6355
rect 5526 6321 5532 6355
rect 5486 6283 5532 6321
rect 5486 6249 5492 6283
rect 5526 6249 5532 6283
rect 5486 6211 5532 6249
rect 5486 6177 5492 6211
rect 5526 6177 5532 6211
rect 5486 6139 5532 6177
rect 5486 6105 5492 6139
rect 5526 6105 5532 6139
rect 5486 6067 5532 6105
rect 5486 6033 5492 6067
rect 5526 6033 5532 6067
rect 5486 5995 5532 6033
rect 5486 5961 5492 5995
rect 5526 5961 5532 5995
rect 5486 5923 5532 5961
rect 5486 5889 5492 5923
rect 5526 5889 5532 5923
rect 5486 5851 5532 5889
rect 5486 5817 5492 5851
rect 5526 5817 5532 5851
rect 5486 5779 5532 5817
rect 5486 5745 5492 5779
rect 5526 5745 5532 5779
rect 5486 5707 5532 5745
rect 5486 5673 5492 5707
rect 5526 5673 5532 5707
rect 5486 5635 5532 5673
rect 5486 5601 5492 5635
rect 5526 5601 5532 5635
rect 5486 5586 5532 5601
rect 5582 6571 5628 6586
rect 5582 6537 5588 6571
rect 5622 6537 5628 6571
rect 5582 6499 5628 6537
rect 5582 6465 5588 6499
rect 5622 6465 5628 6499
rect 5582 6427 5628 6465
rect 5582 6393 5588 6427
rect 5622 6393 5628 6427
rect 5582 6355 5628 6393
rect 5582 6321 5588 6355
rect 5622 6321 5628 6355
rect 5582 6283 5628 6321
rect 5582 6249 5588 6283
rect 5622 6249 5628 6283
rect 5582 6211 5628 6249
rect 5582 6177 5588 6211
rect 5622 6177 5628 6211
rect 5582 6139 5628 6177
rect 5582 6105 5588 6139
rect 5622 6105 5628 6139
rect 5582 6067 5628 6105
rect 5582 6033 5588 6067
rect 5622 6033 5628 6067
rect 5582 5995 5628 6033
rect 5582 5961 5588 5995
rect 5622 5961 5628 5995
rect 5582 5923 5628 5961
rect 5582 5889 5588 5923
rect 5622 5889 5628 5923
rect 5582 5851 5628 5889
rect 5582 5817 5588 5851
rect 5622 5817 5628 5851
rect 5582 5779 5628 5817
rect 5582 5745 5588 5779
rect 5622 5745 5628 5779
rect 5582 5707 5628 5745
rect 5582 5673 5588 5707
rect 5622 5673 5628 5707
rect 5582 5635 5628 5673
rect 5582 5601 5588 5635
rect 5622 5601 5628 5635
rect 5582 5586 5628 5601
rect 5678 6571 5724 6586
rect 5678 6537 5684 6571
rect 5718 6537 5724 6571
rect 5678 6499 5724 6537
rect 5678 6465 5684 6499
rect 5718 6465 5724 6499
rect 5678 6427 5724 6465
rect 5678 6393 5684 6427
rect 5718 6393 5724 6427
rect 5678 6355 5724 6393
rect 5678 6321 5684 6355
rect 5718 6321 5724 6355
rect 5678 6283 5724 6321
rect 5678 6249 5684 6283
rect 5718 6249 5724 6283
rect 5678 6211 5724 6249
rect 5678 6177 5684 6211
rect 5718 6177 5724 6211
rect 5678 6139 5724 6177
rect 5678 6105 5684 6139
rect 5718 6105 5724 6139
rect 5678 6067 5724 6105
rect 5678 6033 5684 6067
rect 5718 6033 5724 6067
rect 5678 5995 5724 6033
rect 5678 5961 5684 5995
rect 5718 5961 5724 5995
rect 5678 5923 5724 5961
rect 5678 5889 5684 5923
rect 5718 5889 5724 5923
rect 5678 5851 5724 5889
rect 5678 5817 5684 5851
rect 5718 5817 5724 5851
rect 5678 5779 5724 5817
rect 5678 5745 5684 5779
rect 5718 5745 5724 5779
rect 5678 5707 5724 5745
rect 5678 5673 5684 5707
rect 5718 5673 5724 5707
rect 5678 5635 5724 5673
rect 5678 5601 5684 5635
rect 5718 5601 5724 5635
rect 5678 5586 5724 5601
rect 6174 6575 6220 6590
rect 6174 6541 6180 6575
rect 6214 6541 6220 6575
rect 6174 6503 6220 6541
rect 6174 6469 6180 6503
rect 6214 6469 6220 6503
rect 6174 6431 6220 6469
rect 6174 6397 6180 6431
rect 6214 6397 6220 6431
rect 6174 6359 6220 6397
rect 6174 6325 6180 6359
rect 6214 6325 6220 6359
rect 6174 6287 6220 6325
rect 6174 6253 6180 6287
rect 6214 6253 6220 6287
rect 6174 6215 6220 6253
rect 6174 6181 6180 6215
rect 6214 6181 6220 6215
rect 6174 6143 6220 6181
rect 6174 6109 6180 6143
rect 6214 6109 6220 6143
rect 6174 6071 6220 6109
rect 6174 6037 6180 6071
rect 6214 6037 6220 6071
rect 6174 5999 6220 6037
rect 6174 5965 6180 5999
rect 6214 5965 6220 5999
rect 6174 5927 6220 5965
rect 6174 5893 6180 5927
rect 6214 5893 6220 5927
rect 6174 5855 6220 5893
rect 6174 5821 6180 5855
rect 6214 5821 6220 5855
rect 6174 5783 6220 5821
rect 6174 5749 6180 5783
rect 6214 5749 6220 5783
rect 6174 5711 6220 5749
rect 6174 5677 6180 5711
rect 6214 5677 6220 5711
rect 6174 5639 6220 5677
rect 6174 5605 6180 5639
rect 6214 5605 6220 5639
rect 6174 5590 6220 5605
rect 6270 6575 6316 6590
rect 6270 6541 6276 6575
rect 6310 6541 6316 6575
rect 6270 6503 6316 6541
rect 6270 6469 6276 6503
rect 6310 6469 6316 6503
rect 6270 6431 6316 6469
rect 6270 6397 6276 6431
rect 6310 6397 6316 6431
rect 6270 6359 6316 6397
rect 6270 6325 6276 6359
rect 6310 6325 6316 6359
rect 6270 6287 6316 6325
rect 6270 6253 6276 6287
rect 6310 6253 6316 6287
rect 6270 6215 6316 6253
rect 6270 6181 6276 6215
rect 6310 6181 6316 6215
rect 6270 6143 6316 6181
rect 6270 6109 6276 6143
rect 6310 6109 6316 6143
rect 6270 6071 6316 6109
rect 6270 6037 6276 6071
rect 6310 6037 6316 6071
rect 6270 5999 6316 6037
rect 6270 5965 6276 5999
rect 6310 5965 6316 5999
rect 6270 5927 6316 5965
rect 6270 5893 6276 5927
rect 6310 5893 6316 5927
rect 6270 5855 6316 5893
rect 6270 5821 6276 5855
rect 6310 5821 6316 5855
rect 6270 5783 6316 5821
rect 6270 5749 6276 5783
rect 6310 5749 6316 5783
rect 6270 5711 6316 5749
rect 6270 5677 6276 5711
rect 6310 5677 6316 5711
rect 6270 5639 6316 5677
rect 6270 5605 6276 5639
rect 6310 5605 6316 5639
rect 6270 5590 6316 5605
rect 6366 6575 6412 6590
rect 6366 6541 6372 6575
rect 6406 6541 6412 6575
rect 6366 6503 6412 6541
rect 6366 6469 6372 6503
rect 6406 6469 6412 6503
rect 6366 6431 6412 6469
rect 6366 6397 6372 6431
rect 6406 6397 6412 6431
rect 6366 6359 6412 6397
rect 6366 6325 6372 6359
rect 6406 6325 6412 6359
rect 6366 6287 6412 6325
rect 6366 6253 6372 6287
rect 6406 6253 6412 6287
rect 6366 6215 6412 6253
rect 6366 6181 6372 6215
rect 6406 6181 6412 6215
rect 6366 6143 6412 6181
rect 6366 6109 6372 6143
rect 6406 6109 6412 6143
rect 6366 6071 6412 6109
rect 6366 6037 6372 6071
rect 6406 6037 6412 6071
rect 6366 5999 6412 6037
rect 6366 5965 6372 5999
rect 6406 5965 6412 5999
rect 6366 5927 6412 5965
rect 6366 5893 6372 5927
rect 6406 5893 6412 5927
rect 6366 5855 6412 5893
rect 6366 5821 6372 5855
rect 6406 5821 6412 5855
rect 6366 5783 6412 5821
rect 6366 5749 6372 5783
rect 6406 5749 6412 5783
rect 6366 5711 6412 5749
rect 6366 5677 6372 5711
rect 6406 5677 6412 5711
rect 6366 5639 6412 5677
rect 6366 5605 6372 5639
rect 6406 5605 6412 5639
rect 6366 5590 6412 5605
rect 6462 6575 6508 6590
rect 6462 6541 6468 6575
rect 6502 6541 6508 6575
rect 6462 6503 6508 6541
rect 6462 6469 6468 6503
rect 6502 6469 6508 6503
rect 6462 6431 6508 6469
rect 6462 6397 6468 6431
rect 6502 6397 6508 6431
rect 6462 6359 6508 6397
rect 6462 6325 6468 6359
rect 6502 6325 6508 6359
rect 6462 6287 6508 6325
rect 6462 6253 6468 6287
rect 6502 6253 6508 6287
rect 6462 6215 6508 6253
rect 6462 6181 6468 6215
rect 6502 6181 6508 6215
rect 6462 6143 6508 6181
rect 6462 6109 6468 6143
rect 6502 6109 6508 6143
rect 6462 6071 6508 6109
rect 6462 6037 6468 6071
rect 6502 6037 6508 6071
rect 6462 5999 6508 6037
rect 6462 5965 6468 5999
rect 6502 5965 6508 5999
rect 6462 5927 6508 5965
rect 6462 5893 6468 5927
rect 6502 5893 6508 5927
rect 6462 5855 6508 5893
rect 6462 5821 6468 5855
rect 6502 5821 6508 5855
rect 6462 5783 6508 5821
rect 6462 5749 6468 5783
rect 6502 5749 6508 5783
rect 6462 5711 6508 5749
rect 6462 5677 6468 5711
rect 6502 5677 6508 5711
rect 6462 5639 6508 5677
rect 6462 5605 6468 5639
rect 6502 5605 6508 5639
rect 6462 5590 6508 5605
rect 6558 6575 6604 6590
rect 6558 6541 6564 6575
rect 6598 6541 6604 6575
rect 6558 6503 6604 6541
rect 6558 6469 6564 6503
rect 6598 6469 6604 6503
rect 6558 6431 6604 6469
rect 6558 6397 6564 6431
rect 6598 6397 6604 6431
rect 6558 6359 6604 6397
rect 6558 6325 6564 6359
rect 6598 6325 6604 6359
rect 6558 6287 6604 6325
rect 6558 6253 6564 6287
rect 6598 6253 6604 6287
rect 6558 6215 6604 6253
rect 6558 6181 6564 6215
rect 6598 6181 6604 6215
rect 6558 6143 6604 6181
rect 6558 6109 6564 6143
rect 6598 6109 6604 6143
rect 6558 6071 6604 6109
rect 6558 6037 6564 6071
rect 6598 6037 6604 6071
rect 6558 5999 6604 6037
rect 6558 5965 6564 5999
rect 6598 5965 6604 5999
rect 6558 5927 6604 5965
rect 6558 5893 6564 5927
rect 6598 5893 6604 5927
rect 6558 5855 6604 5893
rect 6558 5821 6564 5855
rect 6598 5821 6604 5855
rect 6558 5783 6604 5821
rect 6558 5749 6564 5783
rect 6598 5749 6604 5783
rect 6558 5711 6604 5749
rect 6558 5677 6564 5711
rect 6598 5677 6604 5711
rect 6558 5639 6604 5677
rect 6558 5605 6564 5639
rect 6598 5605 6604 5639
rect 6558 5590 6604 5605
rect 6654 6575 6700 6590
rect 6654 6541 6660 6575
rect 6694 6541 6700 6575
rect 6654 6503 6700 6541
rect 6654 6469 6660 6503
rect 6694 6469 6700 6503
rect 6654 6431 6700 6469
rect 6654 6397 6660 6431
rect 6694 6397 6700 6431
rect 6654 6359 6700 6397
rect 6654 6325 6660 6359
rect 6694 6325 6700 6359
rect 6654 6287 6700 6325
rect 6654 6253 6660 6287
rect 6694 6253 6700 6287
rect 6654 6215 6700 6253
rect 6654 6181 6660 6215
rect 6694 6181 6700 6215
rect 6654 6143 6700 6181
rect 6654 6109 6660 6143
rect 6694 6109 6700 6143
rect 6654 6071 6700 6109
rect 6654 6037 6660 6071
rect 6694 6037 6700 6071
rect 6654 5999 6700 6037
rect 6654 5965 6660 5999
rect 6694 5965 6700 5999
rect 6654 5927 6700 5965
rect 6654 5893 6660 5927
rect 6694 5893 6700 5927
rect 6654 5855 6700 5893
rect 6654 5821 6660 5855
rect 6694 5821 6700 5855
rect 6654 5783 6700 5821
rect 6654 5749 6660 5783
rect 6694 5749 6700 5783
rect 6654 5711 6700 5749
rect 6654 5677 6660 5711
rect 6694 5677 6700 5711
rect 6654 5639 6700 5677
rect 6654 5605 6660 5639
rect 6694 5605 6700 5639
rect 6654 5590 6700 5605
rect 6750 6575 6796 6590
rect 6750 6541 6756 6575
rect 6790 6541 6796 6575
rect 6750 6503 6796 6541
rect 6750 6469 6756 6503
rect 6790 6469 6796 6503
rect 6750 6431 6796 6469
rect 6750 6397 6756 6431
rect 6790 6397 6796 6431
rect 6750 6359 6796 6397
rect 6750 6325 6756 6359
rect 6790 6325 6796 6359
rect 6750 6287 6796 6325
rect 6750 6253 6756 6287
rect 6790 6253 6796 6287
rect 6750 6215 6796 6253
rect 6750 6181 6756 6215
rect 6790 6181 6796 6215
rect 6750 6143 6796 6181
rect 6750 6109 6756 6143
rect 6790 6109 6796 6143
rect 6750 6071 6796 6109
rect 6750 6037 6756 6071
rect 6790 6037 6796 6071
rect 6750 5999 6796 6037
rect 6750 5965 6756 5999
rect 6790 5965 6796 5999
rect 6750 5927 6796 5965
rect 6750 5893 6756 5927
rect 6790 5893 6796 5927
rect 6750 5855 6796 5893
rect 6750 5821 6756 5855
rect 6790 5821 6796 5855
rect 6750 5783 6796 5821
rect 6750 5749 6756 5783
rect 6790 5749 6796 5783
rect 6750 5711 6796 5749
rect 6750 5677 6756 5711
rect 6790 5677 6796 5711
rect 6750 5639 6796 5677
rect 6750 5605 6756 5639
rect 6790 5605 6796 5639
rect 6750 5590 6796 5605
rect 6846 6575 6892 6590
rect 6846 6541 6852 6575
rect 6886 6541 6892 6575
rect 6846 6503 6892 6541
rect 6846 6469 6852 6503
rect 6886 6469 6892 6503
rect 6846 6431 6892 6469
rect 6846 6397 6852 6431
rect 6886 6397 6892 6431
rect 6846 6359 6892 6397
rect 6846 6325 6852 6359
rect 6886 6325 6892 6359
rect 6846 6287 6892 6325
rect 6846 6253 6852 6287
rect 6886 6253 6892 6287
rect 6846 6215 6892 6253
rect 6846 6181 6852 6215
rect 6886 6181 6892 6215
rect 6846 6143 6892 6181
rect 6846 6109 6852 6143
rect 6886 6109 6892 6143
rect 6846 6071 6892 6109
rect 6846 6037 6852 6071
rect 6886 6037 6892 6071
rect 6846 5999 6892 6037
rect 6846 5965 6852 5999
rect 6886 5965 6892 5999
rect 6846 5927 6892 5965
rect 6846 5893 6852 5927
rect 6886 5893 6892 5927
rect 6846 5855 6892 5893
rect 6846 5821 6852 5855
rect 6886 5821 6892 5855
rect 6846 5783 6892 5821
rect 6846 5749 6852 5783
rect 6886 5749 6892 5783
rect 6846 5711 6892 5749
rect 6846 5677 6852 5711
rect 6886 5677 6892 5711
rect 6846 5639 6892 5677
rect 6846 5605 6852 5639
rect 6886 5605 6892 5639
rect 6846 5590 6892 5605
rect 6942 6575 6988 6590
rect 6942 6541 6948 6575
rect 6982 6541 6988 6575
rect 6942 6503 6988 6541
rect 6942 6469 6948 6503
rect 6982 6469 6988 6503
rect 6942 6431 6988 6469
rect 6942 6397 6948 6431
rect 6982 6397 6988 6431
rect 6942 6359 6988 6397
rect 6942 6325 6948 6359
rect 6982 6325 6988 6359
rect 6942 6287 6988 6325
rect 6942 6253 6948 6287
rect 6982 6253 6988 6287
rect 6942 6215 6988 6253
rect 6942 6181 6948 6215
rect 6982 6181 6988 6215
rect 6942 6143 6988 6181
rect 6942 6109 6948 6143
rect 6982 6109 6988 6143
rect 6942 6071 6988 6109
rect 6942 6037 6948 6071
rect 6982 6037 6988 6071
rect 6942 5999 6988 6037
rect 6942 5965 6948 5999
rect 6982 5965 6988 5999
rect 6942 5927 6988 5965
rect 6942 5893 6948 5927
rect 6982 5893 6988 5927
rect 6942 5855 6988 5893
rect 6942 5821 6948 5855
rect 6982 5821 6988 5855
rect 6942 5783 6988 5821
rect 6942 5749 6948 5783
rect 6982 5749 6988 5783
rect 6942 5711 6988 5749
rect 6942 5677 6948 5711
rect 6982 5677 6988 5711
rect 6942 5639 6988 5677
rect 6942 5605 6948 5639
rect 6982 5605 6988 5639
rect 6942 5590 6988 5605
rect 7038 6575 7084 6590
rect 7038 6541 7044 6575
rect 7078 6541 7084 6575
rect 7038 6503 7084 6541
rect 7038 6469 7044 6503
rect 7078 6469 7084 6503
rect 7038 6431 7084 6469
rect 7038 6397 7044 6431
rect 7078 6397 7084 6431
rect 7038 6359 7084 6397
rect 7038 6325 7044 6359
rect 7078 6325 7084 6359
rect 7038 6287 7084 6325
rect 7038 6253 7044 6287
rect 7078 6253 7084 6287
rect 7038 6215 7084 6253
rect 7038 6181 7044 6215
rect 7078 6181 7084 6215
rect 7038 6143 7084 6181
rect 7038 6109 7044 6143
rect 7078 6109 7084 6143
rect 7038 6071 7084 6109
rect 7038 6037 7044 6071
rect 7078 6037 7084 6071
rect 7038 5999 7084 6037
rect 7038 5965 7044 5999
rect 7078 5965 7084 5999
rect 7038 5927 7084 5965
rect 7038 5893 7044 5927
rect 7078 5893 7084 5927
rect 7038 5855 7084 5893
rect 7038 5821 7044 5855
rect 7078 5821 7084 5855
rect 7038 5783 7084 5821
rect 7038 5749 7044 5783
rect 7078 5749 7084 5783
rect 7038 5711 7084 5749
rect 7038 5677 7044 5711
rect 7078 5677 7084 5711
rect 7038 5639 7084 5677
rect 7038 5605 7044 5639
rect 7078 5605 7084 5639
rect 7038 5590 7084 5605
rect 7134 6575 7180 6590
rect 7134 6541 7140 6575
rect 7174 6541 7180 6575
rect 7134 6503 7180 6541
rect 7134 6469 7140 6503
rect 7174 6469 7180 6503
rect 7134 6431 7180 6469
rect 7134 6397 7140 6431
rect 7174 6397 7180 6431
rect 7134 6359 7180 6397
rect 7134 6325 7140 6359
rect 7174 6325 7180 6359
rect 7134 6287 7180 6325
rect 7134 6253 7140 6287
rect 7174 6253 7180 6287
rect 7134 6215 7180 6253
rect 7134 6181 7140 6215
rect 7174 6181 7180 6215
rect 7134 6143 7180 6181
rect 7134 6109 7140 6143
rect 7174 6109 7180 6143
rect 7134 6071 7180 6109
rect 7134 6037 7140 6071
rect 7174 6037 7180 6071
rect 7134 5999 7180 6037
rect 7134 5965 7140 5999
rect 7174 5965 7180 5999
rect 7134 5927 7180 5965
rect 7134 5893 7140 5927
rect 7174 5893 7180 5927
rect 7134 5855 7180 5893
rect 7134 5821 7140 5855
rect 7174 5821 7180 5855
rect 7134 5783 7180 5821
rect 7134 5749 7140 5783
rect 7174 5749 7180 5783
rect 7134 5711 7180 5749
rect 7134 5677 7140 5711
rect 7174 5677 7180 5711
rect 7134 5639 7180 5677
rect 7134 5605 7140 5639
rect 7174 5605 7180 5639
rect 7134 5590 7180 5605
rect 7230 6575 7276 6590
rect 7230 6541 7236 6575
rect 7270 6541 7276 6575
rect 7230 6503 7276 6541
rect 7230 6469 7236 6503
rect 7270 6469 7276 6503
rect 7230 6431 7276 6469
rect 7230 6397 7236 6431
rect 7270 6397 7276 6431
rect 7230 6359 7276 6397
rect 7230 6325 7236 6359
rect 7270 6325 7276 6359
rect 7230 6287 7276 6325
rect 7230 6253 7236 6287
rect 7270 6253 7276 6287
rect 7230 6215 7276 6253
rect 7230 6181 7236 6215
rect 7270 6181 7276 6215
rect 7230 6143 7276 6181
rect 7230 6109 7236 6143
rect 7270 6109 7276 6143
rect 7230 6071 7276 6109
rect 7230 6037 7236 6071
rect 7270 6037 7276 6071
rect 7230 5999 7276 6037
rect 7230 5965 7236 5999
rect 7270 5965 7276 5999
rect 7230 5927 7276 5965
rect 7230 5893 7236 5927
rect 7270 5893 7276 5927
rect 7230 5855 7276 5893
rect 7230 5821 7236 5855
rect 7270 5821 7276 5855
rect 7230 5783 7276 5821
rect 7230 5749 7236 5783
rect 7270 5749 7276 5783
rect 7230 5711 7276 5749
rect 7230 5677 7236 5711
rect 7270 5677 7276 5711
rect 7230 5639 7276 5677
rect 7230 5605 7236 5639
rect 7270 5605 7276 5639
rect 7230 5590 7276 5605
rect 7326 6575 7372 6590
rect 7326 6541 7332 6575
rect 7366 6541 7372 6575
rect 7326 6503 7372 6541
rect 7326 6469 7332 6503
rect 7366 6469 7372 6503
rect 7326 6431 7372 6469
rect 7326 6397 7332 6431
rect 7366 6397 7372 6431
rect 7326 6359 7372 6397
rect 7326 6325 7332 6359
rect 7366 6325 7372 6359
rect 7326 6287 7372 6325
rect 7326 6253 7332 6287
rect 7366 6253 7372 6287
rect 7326 6215 7372 6253
rect 7326 6181 7332 6215
rect 7366 6181 7372 6215
rect 7326 6143 7372 6181
rect 7326 6109 7332 6143
rect 7366 6109 7372 6143
rect 7326 6071 7372 6109
rect 7326 6037 7332 6071
rect 7366 6037 7372 6071
rect 7326 5999 7372 6037
rect 7326 5965 7332 5999
rect 7366 5965 7372 5999
rect 7326 5927 7372 5965
rect 7326 5893 7332 5927
rect 7366 5893 7372 5927
rect 7326 5855 7372 5893
rect 7326 5821 7332 5855
rect 7366 5821 7372 5855
rect 7326 5783 7372 5821
rect 7326 5749 7332 5783
rect 7366 5749 7372 5783
rect 7326 5711 7372 5749
rect 7326 5677 7332 5711
rect 7366 5677 7372 5711
rect 7326 5639 7372 5677
rect 7326 5605 7332 5639
rect 7366 5605 7372 5639
rect 7326 5590 7372 5605
rect 7940 6571 7986 6586
rect 7940 6537 7946 6571
rect 7980 6537 7986 6571
rect 7940 6499 7986 6537
rect 7940 6465 7946 6499
rect 7980 6465 7986 6499
rect 7940 6427 7986 6465
rect 7940 6393 7946 6427
rect 7980 6393 7986 6427
rect 7940 6355 7986 6393
rect 7940 6321 7946 6355
rect 7980 6321 7986 6355
rect 7940 6283 7986 6321
rect 7940 6249 7946 6283
rect 7980 6249 7986 6283
rect 7940 6211 7986 6249
rect 7940 6177 7946 6211
rect 7980 6177 7986 6211
rect 7940 6139 7986 6177
rect 7940 6105 7946 6139
rect 7980 6105 7986 6139
rect 7940 6067 7986 6105
rect 7940 6033 7946 6067
rect 7980 6033 7986 6067
rect 7940 5995 7986 6033
rect 7940 5961 7946 5995
rect 7980 5961 7986 5995
rect 7940 5923 7986 5961
rect 7940 5889 7946 5923
rect 7980 5889 7986 5923
rect 7940 5851 7986 5889
rect 7940 5817 7946 5851
rect 7980 5817 7986 5851
rect 7940 5779 7986 5817
rect 7940 5745 7946 5779
rect 7980 5745 7986 5779
rect 7940 5707 7986 5745
rect 7940 5673 7946 5707
rect 7980 5673 7986 5707
rect 7940 5635 7986 5673
rect 7940 5601 7946 5635
rect 7980 5601 7986 5635
rect 7940 5586 7986 5601
rect 8036 6571 8082 6586
rect 8036 6537 8042 6571
rect 8076 6537 8082 6571
rect 8036 6499 8082 6537
rect 8036 6465 8042 6499
rect 8076 6465 8082 6499
rect 8036 6427 8082 6465
rect 8036 6393 8042 6427
rect 8076 6393 8082 6427
rect 8036 6355 8082 6393
rect 8036 6321 8042 6355
rect 8076 6321 8082 6355
rect 8036 6283 8082 6321
rect 8036 6249 8042 6283
rect 8076 6249 8082 6283
rect 8036 6211 8082 6249
rect 8036 6177 8042 6211
rect 8076 6177 8082 6211
rect 8036 6139 8082 6177
rect 8036 6105 8042 6139
rect 8076 6105 8082 6139
rect 8036 6067 8082 6105
rect 8036 6033 8042 6067
rect 8076 6033 8082 6067
rect 8036 5995 8082 6033
rect 8036 5961 8042 5995
rect 8076 5961 8082 5995
rect 8036 5923 8082 5961
rect 8036 5889 8042 5923
rect 8076 5889 8082 5923
rect 8036 5851 8082 5889
rect 8036 5817 8042 5851
rect 8076 5817 8082 5851
rect 8036 5779 8082 5817
rect 8036 5745 8042 5779
rect 8076 5745 8082 5779
rect 8036 5707 8082 5745
rect 8036 5673 8042 5707
rect 8076 5673 8082 5707
rect 8036 5635 8082 5673
rect 8036 5601 8042 5635
rect 8076 5601 8082 5635
rect 8036 5586 8082 5601
rect 8132 6571 8178 6586
rect 8132 6537 8138 6571
rect 8172 6537 8178 6571
rect 8132 6499 8178 6537
rect 8132 6465 8138 6499
rect 8172 6465 8178 6499
rect 8132 6427 8178 6465
rect 8132 6393 8138 6427
rect 8172 6393 8178 6427
rect 8132 6355 8178 6393
rect 8132 6321 8138 6355
rect 8172 6321 8178 6355
rect 8132 6283 8178 6321
rect 8132 6249 8138 6283
rect 8172 6249 8178 6283
rect 8132 6211 8178 6249
rect 8132 6177 8138 6211
rect 8172 6177 8178 6211
rect 8132 6139 8178 6177
rect 8132 6105 8138 6139
rect 8172 6105 8178 6139
rect 8132 6067 8178 6105
rect 8132 6033 8138 6067
rect 8172 6033 8178 6067
rect 8132 5995 8178 6033
rect 8132 5961 8138 5995
rect 8172 5961 8178 5995
rect 8132 5923 8178 5961
rect 8132 5889 8138 5923
rect 8172 5889 8178 5923
rect 8132 5851 8178 5889
rect 8132 5817 8138 5851
rect 8172 5817 8178 5851
rect 8132 5779 8178 5817
rect 8132 5745 8138 5779
rect 8172 5745 8178 5779
rect 8132 5707 8178 5745
rect 8132 5673 8138 5707
rect 8172 5673 8178 5707
rect 8132 5635 8178 5673
rect 8132 5601 8138 5635
rect 8172 5601 8178 5635
rect 8132 5586 8178 5601
rect 8228 6571 8274 6586
rect 8228 6537 8234 6571
rect 8268 6537 8274 6571
rect 8228 6499 8274 6537
rect 8228 6465 8234 6499
rect 8268 6465 8274 6499
rect 8228 6427 8274 6465
rect 8228 6393 8234 6427
rect 8268 6393 8274 6427
rect 8228 6355 8274 6393
rect 8228 6321 8234 6355
rect 8268 6321 8274 6355
rect 8228 6283 8274 6321
rect 8228 6249 8234 6283
rect 8268 6249 8274 6283
rect 8228 6211 8274 6249
rect 8228 6177 8234 6211
rect 8268 6177 8274 6211
rect 8228 6139 8274 6177
rect 8228 6105 8234 6139
rect 8268 6105 8274 6139
rect 8228 6067 8274 6105
rect 8228 6033 8234 6067
rect 8268 6033 8274 6067
rect 8228 5995 8274 6033
rect 8228 5961 8234 5995
rect 8268 5961 8274 5995
rect 8228 5923 8274 5961
rect 8228 5889 8234 5923
rect 8268 5889 8274 5923
rect 8228 5851 8274 5889
rect 8228 5817 8234 5851
rect 8268 5817 8274 5851
rect 8228 5779 8274 5817
rect 8228 5745 8234 5779
rect 8268 5745 8274 5779
rect 8228 5707 8274 5745
rect 8228 5673 8234 5707
rect 8268 5673 8274 5707
rect 8228 5635 8274 5673
rect 8228 5601 8234 5635
rect 8268 5601 8274 5635
rect 8228 5586 8274 5601
rect 8324 6571 8370 6586
rect 8324 6537 8330 6571
rect 8364 6537 8370 6571
rect 8324 6499 8370 6537
rect 8324 6465 8330 6499
rect 8364 6465 8370 6499
rect 8324 6427 8370 6465
rect 8324 6393 8330 6427
rect 8364 6393 8370 6427
rect 8324 6355 8370 6393
rect 8324 6321 8330 6355
rect 8364 6321 8370 6355
rect 8324 6283 8370 6321
rect 8324 6249 8330 6283
rect 8364 6249 8370 6283
rect 8324 6211 8370 6249
rect 8324 6177 8330 6211
rect 8364 6177 8370 6211
rect 8324 6139 8370 6177
rect 8324 6105 8330 6139
rect 8364 6105 8370 6139
rect 8324 6067 8370 6105
rect 8324 6033 8330 6067
rect 8364 6033 8370 6067
rect 8324 5995 8370 6033
rect 8324 5961 8330 5995
rect 8364 5961 8370 5995
rect 8324 5923 8370 5961
rect 8324 5889 8330 5923
rect 8364 5889 8370 5923
rect 8324 5851 8370 5889
rect 8324 5817 8330 5851
rect 8364 5817 8370 5851
rect 8324 5779 8370 5817
rect 8324 5745 8330 5779
rect 8364 5745 8370 5779
rect 8324 5707 8370 5745
rect 8324 5673 8330 5707
rect 8364 5673 8370 5707
rect 8324 5635 8370 5673
rect 8324 5601 8330 5635
rect 8364 5601 8370 5635
rect 8324 5586 8370 5601
rect 8420 6571 8466 6586
rect 8420 6537 8426 6571
rect 8460 6537 8466 6571
rect 8420 6499 8466 6537
rect 8420 6465 8426 6499
rect 8460 6465 8466 6499
rect 8420 6427 8466 6465
rect 8420 6393 8426 6427
rect 8460 6393 8466 6427
rect 8420 6355 8466 6393
rect 8420 6321 8426 6355
rect 8460 6321 8466 6355
rect 8420 6283 8466 6321
rect 8420 6249 8426 6283
rect 8460 6249 8466 6283
rect 8420 6211 8466 6249
rect 8420 6177 8426 6211
rect 8460 6177 8466 6211
rect 8420 6139 8466 6177
rect 8420 6105 8426 6139
rect 8460 6105 8466 6139
rect 8420 6067 8466 6105
rect 8420 6033 8426 6067
rect 8460 6033 8466 6067
rect 8420 5995 8466 6033
rect 8420 5961 8426 5995
rect 8460 5961 8466 5995
rect 8420 5923 8466 5961
rect 8420 5889 8426 5923
rect 8460 5889 8466 5923
rect 8420 5851 8466 5889
rect 8420 5817 8426 5851
rect 8460 5817 8466 5851
rect 8420 5779 8466 5817
rect 8420 5745 8426 5779
rect 8460 5745 8466 5779
rect 8420 5707 8466 5745
rect 8420 5673 8426 5707
rect 8460 5673 8466 5707
rect 8420 5635 8466 5673
rect 8420 5601 8426 5635
rect 8460 5601 8466 5635
rect 8420 5586 8466 5601
rect 8516 6571 8562 6586
rect 8516 6537 8522 6571
rect 8556 6537 8562 6571
rect 8516 6499 8562 6537
rect 8516 6465 8522 6499
rect 8556 6465 8562 6499
rect 8516 6427 8562 6465
rect 8516 6393 8522 6427
rect 8556 6393 8562 6427
rect 8516 6355 8562 6393
rect 8516 6321 8522 6355
rect 8556 6321 8562 6355
rect 8516 6283 8562 6321
rect 8516 6249 8522 6283
rect 8556 6249 8562 6283
rect 8516 6211 8562 6249
rect 8516 6177 8522 6211
rect 8556 6177 8562 6211
rect 8516 6139 8562 6177
rect 8516 6105 8522 6139
rect 8556 6105 8562 6139
rect 8516 6067 8562 6105
rect 8516 6033 8522 6067
rect 8556 6033 8562 6067
rect 8516 5995 8562 6033
rect 8516 5961 8522 5995
rect 8556 5961 8562 5995
rect 8516 5923 8562 5961
rect 8516 5889 8522 5923
rect 8556 5889 8562 5923
rect 8516 5851 8562 5889
rect 8516 5817 8522 5851
rect 8556 5817 8562 5851
rect 8516 5779 8562 5817
rect 8516 5745 8522 5779
rect 8556 5745 8562 5779
rect 8516 5707 8562 5745
rect 8516 5673 8522 5707
rect 8556 5673 8562 5707
rect 8516 5635 8562 5673
rect 8516 5601 8522 5635
rect 8556 5601 8562 5635
rect 8516 5586 8562 5601
rect 8612 6571 8658 6586
rect 8612 6537 8618 6571
rect 8652 6537 8658 6571
rect 8612 6499 8658 6537
rect 8612 6465 8618 6499
rect 8652 6465 8658 6499
rect 8612 6427 8658 6465
rect 8612 6393 8618 6427
rect 8652 6393 8658 6427
rect 8612 6355 8658 6393
rect 8612 6321 8618 6355
rect 8652 6321 8658 6355
rect 8612 6283 8658 6321
rect 8612 6249 8618 6283
rect 8652 6249 8658 6283
rect 8612 6211 8658 6249
rect 8612 6177 8618 6211
rect 8652 6177 8658 6211
rect 8612 6139 8658 6177
rect 8612 6105 8618 6139
rect 8652 6105 8658 6139
rect 8612 6067 8658 6105
rect 8612 6033 8618 6067
rect 8652 6033 8658 6067
rect 8612 5995 8658 6033
rect 8612 5961 8618 5995
rect 8652 5961 8658 5995
rect 8612 5923 8658 5961
rect 8612 5889 8618 5923
rect 8652 5889 8658 5923
rect 8612 5851 8658 5889
rect 8612 5817 8618 5851
rect 8652 5817 8658 5851
rect 8612 5779 8658 5817
rect 8612 5745 8618 5779
rect 8652 5745 8658 5779
rect 8612 5707 8658 5745
rect 8612 5673 8618 5707
rect 8652 5673 8658 5707
rect 8612 5635 8658 5673
rect 8612 5601 8618 5635
rect 8652 5601 8658 5635
rect 8612 5586 8658 5601
rect 8708 6571 8754 6586
rect 8708 6537 8714 6571
rect 8748 6537 8754 6571
rect 8708 6499 8754 6537
rect 8708 6465 8714 6499
rect 8748 6465 8754 6499
rect 8708 6427 8754 6465
rect 8708 6393 8714 6427
rect 8748 6393 8754 6427
rect 8708 6355 8754 6393
rect 8708 6321 8714 6355
rect 8748 6321 8754 6355
rect 8708 6283 8754 6321
rect 8708 6249 8714 6283
rect 8748 6249 8754 6283
rect 8708 6211 8754 6249
rect 8708 6177 8714 6211
rect 8748 6177 8754 6211
rect 8708 6139 8754 6177
rect 8708 6105 8714 6139
rect 8748 6105 8754 6139
rect 8708 6067 8754 6105
rect 8708 6033 8714 6067
rect 8748 6033 8754 6067
rect 8708 5995 8754 6033
rect 8708 5961 8714 5995
rect 8748 5961 8754 5995
rect 8708 5923 8754 5961
rect 8708 5889 8714 5923
rect 8748 5889 8754 5923
rect 8708 5851 8754 5889
rect 8708 5817 8714 5851
rect 8748 5817 8754 5851
rect 8708 5779 8754 5817
rect 8708 5745 8714 5779
rect 8748 5745 8754 5779
rect 8708 5707 8754 5745
rect 8708 5673 8714 5707
rect 8748 5673 8754 5707
rect 8708 5635 8754 5673
rect 8708 5601 8714 5635
rect 8748 5601 8754 5635
rect 8708 5586 8754 5601
rect 9262 6573 9308 6588
rect 9262 6539 9268 6573
rect 9302 6539 9308 6573
rect 9262 6501 9308 6539
rect 9262 6467 9268 6501
rect 9302 6467 9308 6501
rect 9262 6429 9308 6467
rect 9262 6395 9268 6429
rect 9302 6395 9308 6429
rect 9262 6357 9308 6395
rect 9262 6323 9268 6357
rect 9302 6323 9308 6357
rect 9262 6285 9308 6323
rect 9262 6251 9268 6285
rect 9302 6251 9308 6285
rect 9262 6213 9308 6251
rect 9262 6179 9268 6213
rect 9302 6179 9308 6213
rect 9262 6141 9308 6179
rect 9262 6107 9268 6141
rect 9302 6107 9308 6141
rect 9262 6069 9308 6107
rect 9262 6035 9268 6069
rect 9302 6035 9308 6069
rect 9262 5997 9308 6035
rect 9262 5963 9268 5997
rect 9302 5963 9308 5997
rect 9262 5925 9308 5963
rect 9262 5891 9268 5925
rect 9302 5891 9308 5925
rect 9262 5853 9308 5891
rect 9262 5819 9268 5853
rect 9302 5819 9308 5853
rect 9262 5781 9308 5819
rect 9262 5747 9268 5781
rect 9302 5747 9308 5781
rect 9262 5709 9308 5747
rect 9262 5675 9268 5709
rect 9302 5675 9308 5709
rect 9262 5637 9308 5675
rect 9262 5603 9268 5637
rect 9302 5603 9308 5637
rect 9262 5588 9308 5603
rect 9358 6573 9404 6588
rect 9358 6539 9364 6573
rect 9398 6539 9404 6573
rect 9358 6501 9404 6539
rect 9358 6467 9364 6501
rect 9398 6467 9404 6501
rect 9358 6429 9404 6467
rect 9358 6395 9364 6429
rect 9398 6395 9404 6429
rect 9358 6357 9404 6395
rect 9358 6323 9364 6357
rect 9398 6323 9404 6357
rect 9358 6285 9404 6323
rect 9358 6251 9364 6285
rect 9398 6251 9404 6285
rect 9358 6213 9404 6251
rect 9358 6179 9364 6213
rect 9398 6179 9404 6213
rect 9358 6141 9404 6179
rect 9358 6107 9364 6141
rect 9398 6107 9404 6141
rect 9358 6069 9404 6107
rect 9358 6035 9364 6069
rect 9398 6035 9404 6069
rect 9358 5997 9404 6035
rect 9358 5963 9364 5997
rect 9398 5963 9404 5997
rect 9358 5925 9404 5963
rect 9358 5891 9364 5925
rect 9398 5891 9404 5925
rect 9358 5853 9404 5891
rect 9358 5819 9364 5853
rect 9398 5819 9404 5853
rect 9358 5781 9404 5819
rect 9358 5747 9364 5781
rect 9398 5747 9404 5781
rect 9358 5709 9404 5747
rect 9358 5675 9364 5709
rect 9398 5675 9404 5709
rect 9358 5637 9404 5675
rect 9358 5603 9364 5637
rect 9398 5603 9404 5637
rect 9358 5588 9404 5603
rect 9454 6573 9500 6588
rect 9454 6539 9460 6573
rect 9494 6539 9500 6573
rect 9454 6501 9500 6539
rect 9454 6467 9460 6501
rect 9494 6467 9500 6501
rect 9454 6429 9500 6467
rect 9454 6395 9460 6429
rect 9494 6395 9500 6429
rect 9454 6357 9500 6395
rect 9454 6323 9460 6357
rect 9494 6323 9500 6357
rect 9454 6285 9500 6323
rect 9454 6251 9460 6285
rect 9494 6251 9500 6285
rect 9454 6213 9500 6251
rect 9454 6179 9460 6213
rect 9494 6179 9500 6213
rect 9454 6141 9500 6179
rect 9454 6107 9460 6141
rect 9494 6107 9500 6141
rect 9454 6069 9500 6107
rect 9454 6035 9460 6069
rect 9494 6035 9500 6069
rect 9454 5997 9500 6035
rect 9454 5963 9460 5997
rect 9494 5963 9500 5997
rect 9454 5925 9500 5963
rect 9454 5891 9460 5925
rect 9494 5891 9500 5925
rect 9454 5853 9500 5891
rect 9454 5819 9460 5853
rect 9494 5819 9500 5853
rect 9454 5781 9500 5819
rect 9454 5747 9460 5781
rect 9494 5747 9500 5781
rect 9454 5709 9500 5747
rect 9454 5675 9460 5709
rect 9494 5675 9500 5709
rect 9454 5637 9500 5675
rect 9454 5603 9460 5637
rect 9494 5603 9500 5637
rect 9454 5588 9500 5603
rect 9550 6573 9596 6588
rect 9550 6539 9556 6573
rect 9590 6539 9596 6573
rect 9550 6501 9596 6539
rect 9550 6467 9556 6501
rect 9590 6467 9596 6501
rect 9550 6429 9596 6467
rect 9550 6395 9556 6429
rect 9590 6395 9596 6429
rect 9550 6357 9596 6395
rect 9550 6323 9556 6357
rect 9590 6323 9596 6357
rect 9550 6285 9596 6323
rect 9550 6251 9556 6285
rect 9590 6251 9596 6285
rect 9550 6213 9596 6251
rect 9550 6179 9556 6213
rect 9590 6179 9596 6213
rect 9550 6141 9596 6179
rect 9550 6107 9556 6141
rect 9590 6107 9596 6141
rect 9550 6069 9596 6107
rect 9550 6035 9556 6069
rect 9590 6035 9596 6069
rect 9550 5997 9596 6035
rect 9550 5963 9556 5997
rect 9590 5963 9596 5997
rect 9550 5925 9596 5963
rect 9550 5891 9556 5925
rect 9590 5891 9596 5925
rect 9550 5853 9596 5891
rect 9550 5819 9556 5853
rect 9590 5819 9596 5853
rect 9550 5781 9596 5819
rect 9550 5747 9556 5781
rect 9590 5747 9596 5781
rect 9550 5709 9596 5747
rect 9550 5675 9556 5709
rect 9590 5675 9596 5709
rect 9550 5637 9596 5675
rect 9550 5603 9556 5637
rect 9590 5603 9596 5637
rect 9550 5588 9596 5603
rect 9646 6573 9692 6588
rect 9646 6539 9652 6573
rect 9686 6539 9692 6573
rect 9646 6501 9692 6539
rect 9646 6467 9652 6501
rect 9686 6467 9692 6501
rect 9646 6429 9692 6467
rect 9646 6395 9652 6429
rect 9686 6395 9692 6429
rect 9646 6357 9692 6395
rect 9646 6323 9652 6357
rect 9686 6323 9692 6357
rect 9646 6285 9692 6323
rect 9646 6251 9652 6285
rect 9686 6251 9692 6285
rect 9646 6213 9692 6251
rect 9646 6179 9652 6213
rect 9686 6179 9692 6213
rect 9646 6141 9692 6179
rect 9646 6107 9652 6141
rect 9686 6107 9692 6141
rect 9646 6069 9692 6107
rect 9646 6035 9652 6069
rect 9686 6035 9692 6069
rect 9646 5997 9692 6035
rect 9646 5963 9652 5997
rect 9686 5963 9692 5997
rect 9646 5925 9692 5963
rect 9646 5891 9652 5925
rect 9686 5891 9692 5925
rect 9646 5853 9692 5891
rect 9646 5819 9652 5853
rect 9686 5819 9692 5853
rect 9646 5781 9692 5819
rect 9646 5747 9652 5781
rect 9686 5747 9692 5781
rect 9646 5709 9692 5747
rect 9646 5675 9652 5709
rect 9686 5675 9692 5709
rect 9646 5637 9692 5675
rect 9646 5603 9652 5637
rect 9686 5603 9692 5637
rect 9646 5588 9692 5603
rect 9742 6573 9788 6588
rect 9742 6539 9748 6573
rect 9782 6539 9788 6573
rect 9742 6501 9788 6539
rect 9742 6467 9748 6501
rect 9782 6467 9788 6501
rect 9742 6429 9788 6467
rect 9742 6395 9748 6429
rect 9782 6395 9788 6429
rect 9742 6357 9788 6395
rect 9742 6323 9748 6357
rect 9782 6323 9788 6357
rect 9742 6285 9788 6323
rect 9742 6251 9748 6285
rect 9782 6251 9788 6285
rect 9742 6213 9788 6251
rect 9742 6179 9748 6213
rect 9782 6179 9788 6213
rect 9742 6141 9788 6179
rect 9742 6107 9748 6141
rect 9782 6107 9788 6141
rect 9742 6069 9788 6107
rect 9742 6035 9748 6069
rect 9782 6035 9788 6069
rect 9742 5997 9788 6035
rect 9742 5963 9748 5997
rect 9782 5963 9788 5997
rect 9742 5925 9788 5963
rect 9742 5891 9748 5925
rect 9782 5891 9788 5925
rect 9742 5853 9788 5891
rect 9742 5819 9748 5853
rect 9782 5819 9788 5853
rect 9742 5781 9788 5819
rect 9742 5747 9748 5781
rect 9782 5747 9788 5781
rect 9742 5709 9788 5747
rect 9742 5675 9748 5709
rect 9782 5675 9788 5709
rect 9742 5637 9788 5675
rect 9742 5603 9748 5637
rect 9782 5603 9788 5637
rect 9742 5588 9788 5603
rect 9838 6573 9884 6588
rect 9838 6539 9844 6573
rect 9878 6539 9884 6573
rect 9838 6501 9884 6539
rect 9838 6467 9844 6501
rect 9878 6467 9884 6501
rect 9838 6429 9884 6467
rect 9838 6395 9844 6429
rect 9878 6395 9884 6429
rect 9838 6357 9884 6395
rect 9838 6323 9844 6357
rect 9878 6323 9884 6357
rect 9838 6285 9884 6323
rect 9838 6251 9844 6285
rect 9878 6251 9884 6285
rect 9838 6213 9884 6251
rect 9838 6179 9844 6213
rect 9878 6179 9884 6213
rect 9838 6141 9884 6179
rect 9838 6107 9844 6141
rect 9878 6107 9884 6141
rect 9838 6069 9884 6107
rect 9838 6035 9844 6069
rect 9878 6035 9884 6069
rect 9838 5997 9884 6035
rect 9838 5963 9844 5997
rect 9878 5963 9884 5997
rect 9838 5925 9884 5963
rect 9838 5891 9844 5925
rect 9878 5891 9884 5925
rect 9838 5853 9884 5891
rect 9838 5819 9844 5853
rect 9878 5819 9884 5853
rect 9838 5781 9884 5819
rect 9838 5747 9844 5781
rect 9878 5747 9884 5781
rect 9838 5709 9884 5747
rect 9838 5675 9844 5709
rect 9878 5675 9884 5709
rect 9838 5637 9884 5675
rect 9838 5603 9844 5637
rect 9878 5603 9884 5637
rect 9838 5588 9884 5603
rect 9934 6573 9980 6588
rect 9934 6539 9940 6573
rect 9974 6539 9980 6573
rect 9934 6501 9980 6539
rect 9934 6467 9940 6501
rect 9974 6467 9980 6501
rect 9934 6429 9980 6467
rect 9934 6395 9940 6429
rect 9974 6395 9980 6429
rect 9934 6357 9980 6395
rect 9934 6323 9940 6357
rect 9974 6323 9980 6357
rect 9934 6285 9980 6323
rect 9934 6251 9940 6285
rect 9974 6251 9980 6285
rect 9934 6213 9980 6251
rect 9934 6179 9940 6213
rect 9974 6179 9980 6213
rect 9934 6141 9980 6179
rect 9934 6107 9940 6141
rect 9974 6107 9980 6141
rect 9934 6069 9980 6107
rect 9934 6035 9940 6069
rect 9974 6035 9980 6069
rect 9934 5997 9980 6035
rect 9934 5963 9940 5997
rect 9974 5963 9980 5997
rect 9934 5925 9980 5963
rect 9934 5891 9940 5925
rect 9974 5891 9980 5925
rect 9934 5853 9980 5891
rect 9934 5819 9940 5853
rect 9974 5819 9980 5853
rect 9934 5781 9980 5819
rect 9934 5747 9940 5781
rect 9974 5747 9980 5781
rect 9934 5709 9980 5747
rect 9934 5675 9940 5709
rect 9974 5675 9980 5709
rect 9934 5637 9980 5675
rect 9934 5603 9940 5637
rect 9974 5603 9980 5637
rect 9934 5588 9980 5603
rect 10030 6573 10076 6588
rect 10030 6539 10036 6573
rect 10070 6539 10076 6573
rect 10030 6501 10076 6539
rect 10030 6467 10036 6501
rect 10070 6467 10076 6501
rect 10030 6429 10076 6467
rect 10030 6395 10036 6429
rect 10070 6395 10076 6429
rect 10030 6357 10076 6395
rect 10030 6323 10036 6357
rect 10070 6323 10076 6357
rect 10030 6285 10076 6323
rect 10030 6251 10036 6285
rect 10070 6251 10076 6285
rect 10030 6213 10076 6251
rect 10030 6179 10036 6213
rect 10070 6179 10076 6213
rect 10030 6141 10076 6179
rect 10030 6107 10036 6141
rect 10070 6107 10076 6141
rect 10030 6069 10076 6107
rect 10030 6035 10036 6069
rect 10070 6035 10076 6069
rect 10030 5997 10076 6035
rect 10030 5963 10036 5997
rect 10070 5963 10076 5997
rect 10030 5925 10076 5963
rect 10030 5891 10036 5925
rect 10070 5891 10076 5925
rect 10030 5853 10076 5891
rect 10030 5819 10036 5853
rect 10070 5819 10076 5853
rect 10030 5781 10076 5819
rect 10030 5747 10036 5781
rect 10070 5747 10076 5781
rect 10030 5709 10076 5747
rect 10030 5675 10036 5709
rect 10070 5675 10076 5709
rect 10030 5637 10076 5675
rect 10030 5603 10036 5637
rect 10070 5603 10076 5637
rect 10030 5588 10076 5603
rect 10126 6573 10172 6588
rect 10126 6539 10132 6573
rect 10166 6539 10172 6573
rect 10126 6501 10172 6539
rect 10126 6467 10132 6501
rect 10166 6467 10172 6501
rect 10126 6429 10172 6467
rect 10126 6395 10132 6429
rect 10166 6395 10172 6429
rect 10126 6357 10172 6395
rect 10126 6323 10132 6357
rect 10166 6323 10172 6357
rect 10126 6285 10172 6323
rect 10126 6251 10132 6285
rect 10166 6251 10172 6285
rect 10126 6213 10172 6251
rect 10126 6179 10132 6213
rect 10166 6179 10172 6213
rect 10126 6141 10172 6179
rect 10126 6107 10132 6141
rect 10166 6107 10172 6141
rect 10126 6069 10172 6107
rect 10126 6035 10132 6069
rect 10166 6035 10172 6069
rect 10126 5997 10172 6035
rect 10126 5963 10132 5997
rect 10166 5963 10172 5997
rect 10126 5925 10172 5963
rect 10126 5891 10132 5925
rect 10166 5891 10172 5925
rect 10126 5853 10172 5891
rect 10126 5819 10132 5853
rect 10166 5819 10172 5853
rect 10126 5781 10172 5819
rect 10126 5747 10132 5781
rect 10166 5747 10172 5781
rect 10126 5709 10172 5747
rect 10126 5675 10132 5709
rect 10166 5675 10172 5709
rect 10126 5637 10172 5675
rect 10126 5603 10132 5637
rect 10166 5603 10172 5637
rect 10126 5588 10172 5603
rect 10222 6573 10268 6588
rect 10222 6539 10228 6573
rect 10262 6539 10268 6573
rect 10222 6501 10268 6539
rect 10222 6467 10228 6501
rect 10262 6467 10268 6501
rect 10222 6429 10268 6467
rect 10222 6395 10228 6429
rect 10262 6395 10268 6429
rect 10222 6357 10268 6395
rect 10222 6323 10228 6357
rect 10262 6323 10268 6357
rect 10222 6285 10268 6323
rect 10222 6251 10228 6285
rect 10262 6251 10268 6285
rect 10222 6213 10268 6251
rect 10222 6179 10228 6213
rect 10262 6179 10268 6213
rect 10222 6141 10268 6179
rect 10222 6107 10228 6141
rect 10262 6107 10268 6141
rect 10222 6069 10268 6107
rect 10222 6035 10228 6069
rect 10262 6035 10268 6069
rect 10222 5997 10268 6035
rect 10222 5963 10228 5997
rect 10262 5963 10268 5997
rect 10222 5925 10268 5963
rect 10222 5891 10228 5925
rect 10262 5891 10268 5925
rect 10222 5853 10268 5891
rect 10222 5819 10228 5853
rect 10262 5819 10268 5853
rect 10222 5781 10268 5819
rect 10222 5747 10228 5781
rect 10262 5747 10268 5781
rect 10222 5709 10268 5747
rect 10222 5675 10228 5709
rect 10262 5675 10268 5709
rect 10222 5637 10268 5675
rect 10222 5603 10228 5637
rect 10262 5603 10268 5637
rect 10222 5588 10268 5603
rect 10318 6573 10364 6588
rect 10318 6539 10324 6573
rect 10358 6539 10364 6573
rect 10318 6501 10364 6539
rect 10318 6467 10324 6501
rect 10358 6467 10364 6501
rect 10318 6429 10364 6467
rect 10318 6395 10324 6429
rect 10358 6395 10364 6429
rect 10318 6357 10364 6395
rect 10318 6323 10324 6357
rect 10358 6323 10364 6357
rect 10318 6285 10364 6323
rect 10318 6251 10324 6285
rect 10358 6251 10364 6285
rect 10318 6213 10364 6251
rect 10318 6179 10324 6213
rect 10358 6179 10364 6213
rect 10318 6141 10364 6179
rect 10318 6107 10324 6141
rect 10358 6107 10364 6141
rect 10318 6069 10364 6107
rect 10318 6035 10324 6069
rect 10358 6035 10364 6069
rect 10318 5997 10364 6035
rect 10318 5963 10324 5997
rect 10358 5963 10364 5997
rect 10318 5925 10364 5963
rect 10318 5891 10324 5925
rect 10358 5891 10364 5925
rect 10318 5853 10364 5891
rect 10318 5819 10324 5853
rect 10358 5819 10364 5853
rect 10318 5781 10364 5819
rect 10318 5747 10324 5781
rect 10358 5747 10364 5781
rect 10318 5709 10364 5747
rect 10318 5675 10324 5709
rect 10358 5675 10364 5709
rect 10318 5637 10364 5675
rect 10318 5603 10324 5637
rect 10358 5603 10364 5637
rect 10318 5588 10364 5603
rect 10414 6573 10460 6588
rect 10414 6539 10420 6573
rect 10454 6539 10460 6573
rect 10414 6501 10460 6539
rect 10414 6467 10420 6501
rect 10454 6467 10460 6501
rect 10414 6429 10460 6467
rect 10414 6395 10420 6429
rect 10454 6395 10460 6429
rect 10414 6357 10460 6395
rect 10414 6323 10420 6357
rect 10454 6323 10460 6357
rect 10414 6285 10460 6323
rect 10414 6251 10420 6285
rect 10454 6251 10460 6285
rect 10414 6213 10460 6251
rect 10414 6179 10420 6213
rect 10454 6179 10460 6213
rect 10414 6141 10460 6179
rect 10414 6107 10420 6141
rect 10454 6107 10460 6141
rect 10414 6069 10460 6107
rect 10414 6035 10420 6069
rect 10454 6035 10460 6069
rect 10414 5997 10460 6035
rect 10414 5963 10420 5997
rect 10454 5963 10460 5997
rect 10414 5925 10460 5963
rect 10414 5891 10420 5925
rect 10454 5891 10460 5925
rect 10414 5853 10460 5891
rect 10414 5819 10420 5853
rect 10454 5819 10460 5853
rect 10414 5781 10460 5819
rect 10414 5747 10420 5781
rect 10454 5747 10460 5781
rect 10414 5709 10460 5747
rect 10414 5675 10420 5709
rect 10454 5675 10460 5709
rect 10414 5637 10460 5675
rect 10414 5603 10420 5637
rect 10454 5603 10460 5637
rect 10414 5588 10460 5603
rect 11028 6569 11074 6584
rect 11028 6535 11034 6569
rect 11068 6535 11074 6569
rect 11028 6497 11074 6535
rect 11028 6463 11034 6497
rect 11068 6463 11074 6497
rect 11028 6425 11074 6463
rect 11028 6391 11034 6425
rect 11068 6391 11074 6425
rect 11028 6353 11074 6391
rect 11028 6319 11034 6353
rect 11068 6319 11074 6353
rect 11028 6281 11074 6319
rect 11028 6247 11034 6281
rect 11068 6247 11074 6281
rect 11028 6209 11074 6247
rect 11028 6175 11034 6209
rect 11068 6175 11074 6209
rect 11028 6137 11074 6175
rect 11028 6103 11034 6137
rect 11068 6103 11074 6137
rect 11028 6065 11074 6103
rect 11028 6031 11034 6065
rect 11068 6031 11074 6065
rect 11028 5993 11074 6031
rect 11028 5959 11034 5993
rect 11068 5959 11074 5993
rect 11028 5921 11074 5959
rect 11028 5887 11034 5921
rect 11068 5887 11074 5921
rect 11028 5849 11074 5887
rect 11028 5815 11034 5849
rect 11068 5815 11074 5849
rect 11028 5777 11074 5815
rect 11028 5743 11034 5777
rect 11068 5743 11074 5777
rect 11028 5705 11074 5743
rect 11028 5671 11034 5705
rect 11068 5671 11074 5705
rect 11028 5633 11074 5671
rect 11028 5599 11034 5633
rect 11068 5599 11074 5633
rect 11028 5584 11074 5599
rect 11124 6569 11170 6584
rect 11124 6535 11130 6569
rect 11164 6535 11170 6569
rect 11124 6497 11170 6535
rect 11124 6463 11130 6497
rect 11164 6463 11170 6497
rect 11124 6425 11170 6463
rect 11124 6391 11130 6425
rect 11164 6391 11170 6425
rect 11124 6353 11170 6391
rect 11124 6319 11130 6353
rect 11164 6319 11170 6353
rect 11124 6281 11170 6319
rect 11124 6247 11130 6281
rect 11164 6247 11170 6281
rect 11124 6209 11170 6247
rect 11124 6175 11130 6209
rect 11164 6175 11170 6209
rect 11124 6137 11170 6175
rect 11124 6103 11130 6137
rect 11164 6103 11170 6137
rect 11124 6065 11170 6103
rect 11124 6031 11130 6065
rect 11164 6031 11170 6065
rect 11124 5993 11170 6031
rect 11124 5959 11130 5993
rect 11164 5959 11170 5993
rect 11124 5921 11170 5959
rect 11124 5887 11130 5921
rect 11164 5887 11170 5921
rect 11124 5849 11170 5887
rect 11124 5815 11130 5849
rect 11164 5815 11170 5849
rect 11124 5777 11170 5815
rect 11124 5743 11130 5777
rect 11164 5743 11170 5777
rect 11124 5705 11170 5743
rect 11124 5671 11130 5705
rect 11164 5671 11170 5705
rect 11124 5633 11170 5671
rect 11124 5599 11130 5633
rect 11164 5599 11170 5633
rect 11124 5584 11170 5599
rect 11220 6569 11266 6584
rect 11220 6535 11226 6569
rect 11260 6535 11266 6569
rect 11220 6497 11266 6535
rect 11220 6463 11226 6497
rect 11260 6463 11266 6497
rect 11220 6425 11266 6463
rect 11220 6391 11226 6425
rect 11260 6391 11266 6425
rect 11220 6353 11266 6391
rect 11220 6319 11226 6353
rect 11260 6319 11266 6353
rect 11220 6281 11266 6319
rect 11220 6247 11226 6281
rect 11260 6247 11266 6281
rect 11220 6209 11266 6247
rect 11220 6175 11226 6209
rect 11260 6175 11266 6209
rect 11220 6137 11266 6175
rect 11220 6103 11226 6137
rect 11260 6103 11266 6137
rect 11220 6065 11266 6103
rect 11220 6031 11226 6065
rect 11260 6031 11266 6065
rect 11220 5993 11266 6031
rect 11220 5959 11226 5993
rect 11260 5959 11266 5993
rect 11220 5921 11266 5959
rect 11220 5887 11226 5921
rect 11260 5887 11266 5921
rect 11220 5849 11266 5887
rect 11220 5815 11226 5849
rect 11260 5815 11266 5849
rect 11220 5777 11266 5815
rect 11220 5743 11226 5777
rect 11260 5743 11266 5777
rect 11220 5705 11266 5743
rect 11220 5671 11226 5705
rect 11260 5671 11266 5705
rect 11220 5633 11266 5671
rect 11220 5599 11226 5633
rect 11260 5599 11266 5633
rect 11220 5584 11266 5599
rect 11316 6569 11362 6584
rect 11316 6535 11322 6569
rect 11356 6535 11362 6569
rect 11316 6497 11362 6535
rect 11316 6463 11322 6497
rect 11356 6463 11362 6497
rect 11316 6425 11362 6463
rect 11316 6391 11322 6425
rect 11356 6391 11362 6425
rect 11316 6353 11362 6391
rect 11316 6319 11322 6353
rect 11356 6319 11362 6353
rect 11316 6281 11362 6319
rect 11316 6247 11322 6281
rect 11356 6247 11362 6281
rect 11316 6209 11362 6247
rect 11316 6175 11322 6209
rect 11356 6175 11362 6209
rect 11316 6137 11362 6175
rect 11316 6103 11322 6137
rect 11356 6103 11362 6137
rect 11316 6065 11362 6103
rect 11316 6031 11322 6065
rect 11356 6031 11362 6065
rect 11316 5993 11362 6031
rect 11316 5959 11322 5993
rect 11356 5959 11362 5993
rect 11316 5921 11362 5959
rect 11316 5887 11322 5921
rect 11356 5887 11362 5921
rect 11316 5849 11362 5887
rect 11316 5815 11322 5849
rect 11356 5815 11362 5849
rect 11316 5777 11362 5815
rect 11316 5743 11322 5777
rect 11356 5743 11362 5777
rect 11316 5705 11362 5743
rect 11316 5671 11322 5705
rect 11356 5671 11362 5705
rect 11316 5633 11362 5671
rect 11316 5599 11322 5633
rect 11356 5599 11362 5633
rect 11316 5584 11362 5599
rect 11412 6569 11458 6584
rect 11412 6535 11418 6569
rect 11452 6535 11458 6569
rect 11412 6497 11458 6535
rect 11412 6463 11418 6497
rect 11452 6463 11458 6497
rect 11412 6425 11458 6463
rect 11412 6391 11418 6425
rect 11452 6391 11458 6425
rect 11412 6353 11458 6391
rect 11412 6319 11418 6353
rect 11452 6319 11458 6353
rect 11412 6281 11458 6319
rect 11412 6247 11418 6281
rect 11452 6247 11458 6281
rect 11412 6209 11458 6247
rect 11412 6175 11418 6209
rect 11452 6175 11458 6209
rect 11412 6137 11458 6175
rect 11412 6103 11418 6137
rect 11452 6103 11458 6137
rect 11412 6065 11458 6103
rect 11412 6031 11418 6065
rect 11452 6031 11458 6065
rect 11412 5993 11458 6031
rect 11412 5959 11418 5993
rect 11452 5959 11458 5993
rect 11412 5921 11458 5959
rect 11412 5887 11418 5921
rect 11452 5887 11458 5921
rect 11412 5849 11458 5887
rect 11412 5815 11418 5849
rect 11452 5815 11458 5849
rect 11412 5777 11458 5815
rect 11412 5743 11418 5777
rect 11452 5743 11458 5777
rect 11412 5705 11458 5743
rect 11412 5671 11418 5705
rect 11452 5671 11458 5705
rect 11412 5633 11458 5671
rect 11412 5599 11418 5633
rect 11452 5599 11458 5633
rect 11412 5584 11458 5599
rect 11508 6569 11554 6584
rect 11508 6535 11514 6569
rect 11548 6535 11554 6569
rect 11508 6497 11554 6535
rect 11508 6463 11514 6497
rect 11548 6463 11554 6497
rect 11508 6425 11554 6463
rect 11508 6391 11514 6425
rect 11548 6391 11554 6425
rect 11508 6353 11554 6391
rect 11508 6319 11514 6353
rect 11548 6319 11554 6353
rect 11508 6281 11554 6319
rect 11508 6247 11514 6281
rect 11548 6247 11554 6281
rect 11508 6209 11554 6247
rect 11508 6175 11514 6209
rect 11548 6175 11554 6209
rect 11508 6137 11554 6175
rect 11508 6103 11514 6137
rect 11548 6103 11554 6137
rect 11508 6065 11554 6103
rect 11508 6031 11514 6065
rect 11548 6031 11554 6065
rect 11508 5993 11554 6031
rect 11508 5959 11514 5993
rect 11548 5959 11554 5993
rect 11508 5921 11554 5959
rect 11508 5887 11514 5921
rect 11548 5887 11554 5921
rect 11508 5849 11554 5887
rect 11508 5815 11514 5849
rect 11548 5815 11554 5849
rect 11508 5777 11554 5815
rect 11508 5743 11514 5777
rect 11548 5743 11554 5777
rect 11508 5705 11554 5743
rect 11508 5671 11514 5705
rect 11548 5671 11554 5705
rect 11508 5633 11554 5671
rect 11508 5599 11514 5633
rect 11548 5599 11554 5633
rect 11508 5584 11554 5599
rect 11604 6569 11650 6584
rect 11604 6535 11610 6569
rect 11644 6535 11650 6569
rect 11604 6497 11650 6535
rect 11604 6463 11610 6497
rect 11644 6463 11650 6497
rect 11604 6425 11650 6463
rect 11604 6391 11610 6425
rect 11644 6391 11650 6425
rect 11604 6353 11650 6391
rect 11604 6319 11610 6353
rect 11644 6319 11650 6353
rect 11604 6281 11650 6319
rect 11604 6247 11610 6281
rect 11644 6247 11650 6281
rect 11604 6209 11650 6247
rect 11604 6175 11610 6209
rect 11644 6175 11650 6209
rect 11604 6137 11650 6175
rect 11604 6103 11610 6137
rect 11644 6103 11650 6137
rect 11604 6065 11650 6103
rect 11604 6031 11610 6065
rect 11644 6031 11650 6065
rect 11604 5993 11650 6031
rect 11604 5959 11610 5993
rect 11644 5959 11650 5993
rect 11604 5921 11650 5959
rect 11604 5887 11610 5921
rect 11644 5887 11650 5921
rect 11604 5849 11650 5887
rect 11604 5815 11610 5849
rect 11644 5815 11650 5849
rect 11604 5777 11650 5815
rect 11604 5743 11610 5777
rect 11644 5743 11650 5777
rect 11604 5705 11650 5743
rect 11604 5671 11610 5705
rect 11644 5671 11650 5705
rect 11604 5633 11650 5671
rect 11604 5599 11610 5633
rect 11644 5599 11650 5633
rect 11604 5584 11650 5599
rect 11700 6569 11746 6584
rect 11700 6535 11706 6569
rect 11740 6535 11746 6569
rect 11700 6497 11746 6535
rect 11700 6463 11706 6497
rect 11740 6463 11746 6497
rect 11700 6425 11746 6463
rect 11700 6391 11706 6425
rect 11740 6391 11746 6425
rect 11700 6353 11746 6391
rect 11700 6319 11706 6353
rect 11740 6319 11746 6353
rect 11700 6281 11746 6319
rect 11700 6247 11706 6281
rect 11740 6247 11746 6281
rect 11700 6209 11746 6247
rect 11700 6175 11706 6209
rect 11740 6175 11746 6209
rect 11700 6137 11746 6175
rect 11700 6103 11706 6137
rect 11740 6103 11746 6137
rect 11700 6065 11746 6103
rect 11700 6031 11706 6065
rect 11740 6031 11746 6065
rect 11700 5993 11746 6031
rect 11700 5959 11706 5993
rect 11740 5959 11746 5993
rect 11700 5921 11746 5959
rect 11700 5887 11706 5921
rect 11740 5887 11746 5921
rect 11700 5849 11746 5887
rect 11700 5815 11706 5849
rect 11740 5815 11746 5849
rect 11700 5777 11746 5815
rect 11700 5743 11706 5777
rect 11740 5743 11746 5777
rect 11700 5705 11746 5743
rect 11700 5671 11706 5705
rect 11740 5671 11746 5705
rect 11700 5633 11746 5671
rect 11700 5599 11706 5633
rect 11740 5599 11746 5633
rect 11700 5584 11746 5599
rect 11796 6569 11842 6584
rect 11796 6535 11802 6569
rect 11836 6535 11842 6569
rect 11796 6497 11842 6535
rect 11796 6463 11802 6497
rect 11836 6463 11842 6497
rect 11796 6425 11842 6463
rect 11796 6391 11802 6425
rect 11836 6391 11842 6425
rect 11796 6353 11842 6391
rect 11796 6319 11802 6353
rect 11836 6319 11842 6353
rect 11796 6281 11842 6319
rect 11796 6247 11802 6281
rect 11836 6247 11842 6281
rect 11796 6209 11842 6247
rect 11796 6175 11802 6209
rect 11836 6175 11842 6209
rect 11796 6137 11842 6175
rect 11796 6103 11802 6137
rect 11836 6103 11842 6137
rect 11796 6065 11842 6103
rect 11796 6031 11802 6065
rect 11836 6031 11842 6065
rect 11796 5993 11842 6031
rect 11796 5959 11802 5993
rect 11836 5959 11842 5993
rect 11796 5921 11842 5959
rect 11796 5887 11802 5921
rect 11836 5887 11842 5921
rect 11796 5849 11842 5887
rect 11796 5815 11802 5849
rect 11836 5815 11842 5849
rect 11796 5777 11842 5815
rect 11796 5743 11802 5777
rect 11836 5743 11842 5777
rect 11796 5705 11842 5743
rect 11796 5671 11802 5705
rect 11836 5671 11842 5705
rect 11796 5633 11842 5671
rect 11796 5599 11802 5633
rect 11836 5599 11842 5633
rect 11796 5584 11842 5599
rect 12418 6547 12464 6562
rect 12418 6513 12424 6547
rect 12458 6513 12464 6547
rect 12418 6475 12464 6513
rect 12418 6441 12424 6475
rect 12458 6441 12464 6475
rect 12418 6403 12464 6441
rect 12418 6369 12424 6403
rect 12458 6369 12464 6403
rect 12418 6331 12464 6369
rect 12418 6297 12424 6331
rect 12458 6297 12464 6331
rect 12418 6259 12464 6297
rect 12418 6225 12424 6259
rect 12458 6225 12464 6259
rect 12418 6187 12464 6225
rect 12418 6153 12424 6187
rect 12458 6153 12464 6187
rect 12418 6115 12464 6153
rect 12418 6081 12424 6115
rect 12458 6081 12464 6115
rect 12418 6043 12464 6081
rect 12418 6009 12424 6043
rect 12458 6009 12464 6043
rect 12418 5971 12464 6009
rect 12418 5937 12424 5971
rect 12458 5937 12464 5971
rect 12418 5899 12464 5937
rect 12418 5865 12424 5899
rect 12458 5865 12464 5899
rect 12418 5827 12464 5865
rect 12418 5793 12424 5827
rect 12458 5793 12464 5827
rect 12418 5755 12464 5793
rect 12418 5721 12424 5755
rect 12458 5721 12464 5755
rect 12418 5683 12464 5721
rect 12418 5649 12424 5683
rect 12458 5649 12464 5683
rect 12418 5611 12464 5649
rect 12418 5577 12424 5611
rect 12458 5577 12464 5611
rect 12418 5562 12464 5577
rect 12514 6547 12560 6562
rect 12514 6513 12520 6547
rect 12554 6513 12560 6547
rect 12514 6475 12560 6513
rect 12514 6441 12520 6475
rect 12554 6441 12560 6475
rect 12514 6403 12560 6441
rect 12514 6369 12520 6403
rect 12554 6369 12560 6403
rect 12514 6331 12560 6369
rect 12514 6297 12520 6331
rect 12554 6297 12560 6331
rect 12514 6259 12560 6297
rect 12514 6225 12520 6259
rect 12554 6225 12560 6259
rect 12514 6187 12560 6225
rect 12514 6153 12520 6187
rect 12554 6153 12560 6187
rect 12514 6115 12560 6153
rect 12514 6081 12520 6115
rect 12554 6081 12560 6115
rect 12514 6043 12560 6081
rect 12514 6009 12520 6043
rect 12554 6009 12560 6043
rect 12514 5971 12560 6009
rect 12514 5937 12520 5971
rect 12554 5937 12560 5971
rect 12514 5899 12560 5937
rect 12514 5865 12520 5899
rect 12554 5865 12560 5899
rect 12514 5827 12560 5865
rect 12514 5793 12520 5827
rect 12554 5793 12560 5827
rect 12514 5755 12560 5793
rect 12514 5721 12520 5755
rect 12554 5721 12560 5755
rect 12514 5683 12560 5721
rect 12514 5649 12520 5683
rect 12554 5649 12560 5683
rect 12514 5611 12560 5649
rect 12514 5577 12520 5611
rect 12554 5577 12560 5611
rect 12514 5562 12560 5577
rect 12610 6547 12656 6562
rect 12610 6513 12616 6547
rect 12650 6513 12656 6547
rect 12610 6475 12656 6513
rect 12610 6441 12616 6475
rect 12650 6441 12656 6475
rect 12610 6403 12656 6441
rect 12610 6369 12616 6403
rect 12650 6369 12656 6403
rect 12610 6331 12656 6369
rect 12610 6297 12616 6331
rect 12650 6297 12656 6331
rect 12610 6259 12656 6297
rect 12610 6225 12616 6259
rect 12650 6225 12656 6259
rect 12610 6187 12656 6225
rect 12610 6153 12616 6187
rect 12650 6153 12656 6187
rect 12610 6115 12656 6153
rect 12610 6081 12616 6115
rect 12650 6081 12656 6115
rect 12610 6043 12656 6081
rect 12610 6009 12616 6043
rect 12650 6009 12656 6043
rect 12610 5971 12656 6009
rect 12610 5937 12616 5971
rect 12650 5937 12656 5971
rect 12610 5899 12656 5937
rect 12610 5865 12616 5899
rect 12650 5865 12656 5899
rect 12610 5827 12656 5865
rect 12610 5793 12616 5827
rect 12650 5793 12656 5827
rect 12610 5755 12656 5793
rect 12610 5721 12616 5755
rect 12650 5721 12656 5755
rect 12610 5683 12656 5721
rect 12610 5649 12616 5683
rect 12650 5649 12656 5683
rect 12610 5611 12656 5649
rect 12610 5577 12616 5611
rect 12650 5577 12656 5611
rect 12610 5562 12656 5577
rect 12706 6547 12752 6562
rect 12706 6513 12712 6547
rect 12746 6513 12752 6547
rect 12706 6475 12752 6513
rect 12706 6441 12712 6475
rect 12746 6441 12752 6475
rect 12706 6403 12752 6441
rect 12706 6369 12712 6403
rect 12746 6369 12752 6403
rect 12706 6331 12752 6369
rect 12706 6297 12712 6331
rect 12746 6297 12752 6331
rect 12706 6259 12752 6297
rect 12706 6225 12712 6259
rect 12746 6225 12752 6259
rect 12706 6187 12752 6225
rect 12706 6153 12712 6187
rect 12746 6153 12752 6187
rect 12706 6115 12752 6153
rect 12706 6081 12712 6115
rect 12746 6081 12752 6115
rect 12706 6043 12752 6081
rect 12706 6009 12712 6043
rect 12746 6009 12752 6043
rect 12706 5971 12752 6009
rect 12706 5937 12712 5971
rect 12746 5937 12752 5971
rect 12706 5899 12752 5937
rect 12706 5865 12712 5899
rect 12746 5865 12752 5899
rect 12706 5827 12752 5865
rect 12706 5793 12712 5827
rect 12746 5793 12752 5827
rect 12706 5755 12752 5793
rect 12706 5721 12712 5755
rect 12746 5721 12752 5755
rect 12706 5683 12752 5721
rect 12706 5649 12712 5683
rect 12746 5649 12752 5683
rect 12706 5611 12752 5649
rect 12706 5577 12712 5611
rect 12746 5577 12752 5611
rect 12706 5562 12752 5577
rect 12802 6547 12848 6562
rect 12802 6513 12808 6547
rect 12842 6513 12848 6547
rect 12802 6475 12848 6513
rect 12802 6441 12808 6475
rect 12842 6441 12848 6475
rect 12802 6403 12848 6441
rect 12802 6369 12808 6403
rect 12842 6369 12848 6403
rect 12802 6331 12848 6369
rect 12802 6297 12808 6331
rect 12842 6297 12848 6331
rect 12802 6259 12848 6297
rect 12802 6225 12808 6259
rect 12842 6225 12848 6259
rect 12802 6187 12848 6225
rect 12802 6153 12808 6187
rect 12842 6153 12848 6187
rect 12802 6115 12848 6153
rect 12802 6081 12808 6115
rect 12842 6081 12848 6115
rect 12802 6043 12848 6081
rect 12802 6009 12808 6043
rect 12842 6009 12848 6043
rect 12802 5971 12848 6009
rect 12802 5937 12808 5971
rect 12842 5937 12848 5971
rect 12802 5899 12848 5937
rect 12802 5865 12808 5899
rect 12842 5865 12848 5899
rect 12802 5827 12848 5865
rect 12802 5793 12808 5827
rect 12842 5793 12848 5827
rect 12802 5755 12848 5793
rect 12802 5721 12808 5755
rect 12842 5721 12848 5755
rect 12802 5683 12848 5721
rect 12802 5649 12808 5683
rect 12842 5649 12848 5683
rect 12802 5611 12848 5649
rect 12802 5577 12808 5611
rect 12842 5577 12848 5611
rect 12802 5562 12848 5577
rect 12898 6547 12944 6562
rect 12898 6513 12904 6547
rect 12938 6513 12944 6547
rect 12898 6475 12944 6513
rect 12898 6441 12904 6475
rect 12938 6441 12944 6475
rect 12898 6403 12944 6441
rect 12898 6369 12904 6403
rect 12938 6369 12944 6403
rect 12898 6331 12944 6369
rect 12898 6297 12904 6331
rect 12938 6297 12944 6331
rect 12898 6259 12944 6297
rect 12898 6225 12904 6259
rect 12938 6225 12944 6259
rect 12898 6187 12944 6225
rect 12898 6153 12904 6187
rect 12938 6153 12944 6187
rect 12898 6115 12944 6153
rect 12898 6081 12904 6115
rect 12938 6081 12944 6115
rect 12898 6043 12944 6081
rect 12898 6009 12904 6043
rect 12938 6009 12944 6043
rect 12898 5971 12944 6009
rect 12898 5937 12904 5971
rect 12938 5937 12944 5971
rect 12898 5899 12944 5937
rect 12898 5865 12904 5899
rect 12938 5865 12944 5899
rect 12898 5827 12944 5865
rect 12898 5793 12904 5827
rect 12938 5793 12944 5827
rect 12898 5755 12944 5793
rect 12898 5721 12904 5755
rect 12938 5721 12944 5755
rect 12898 5683 12944 5721
rect 12898 5649 12904 5683
rect 12938 5649 12944 5683
rect 12898 5611 12944 5649
rect 12898 5577 12904 5611
rect 12938 5577 12944 5611
rect 12898 5562 12944 5577
rect 12994 6547 13040 6562
rect 12994 6513 13000 6547
rect 13034 6513 13040 6547
rect 12994 6475 13040 6513
rect 12994 6441 13000 6475
rect 13034 6441 13040 6475
rect 12994 6403 13040 6441
rect 12994 6369 13000 6403
rect 13034 6369 13040 6403
rect 12994 6331 13040 6369
rect 12994 6297 13000 6331
rect 13034 6297 13040 6331
rect 12994 6259 13040 6297
rect 12994 6225 13000 6259
rect 13034 6225 13040 6259
rect 12994 6187 13040 6225
rect 12994 6153 13000 6187
rect 13034 6153 13040 6187
rect 12994 6115 13040 6153
rect 12994 6081 13000 6115
rect 13034 6081 13040 6115
rect 12994 6043 13040 6081
rect 12994 6009 13000 6043
rect 13034 6009 13040 6043
rect 12994 5971 13040 6009
rect 12994 5937 13000 5971
rect 13034 5937 13040 5971
rect 12994 5899 13040 5937
rect 12994 5865 13000 5899
rect 13034 5865 13040 5899
rect 12994 5827 13040 5865
rect 12994 5793 13000 5827
rect 13034 5793 13040 5827
rect 12994 5755 13040 5793
rect 12994 5721 13000 5755
rect 13034 5721 13040 5755
rect 12994 5683 13040 5721
rect 12994 5649 13000 5683
rect 13034 5649 13040 5683
rect 12994 5611 13040 5649
rect 12994 5577 13000 5611
rect 13034 5577 13040 5611
rect 12994 5562 13040 5577
rect 13090 6547 13136 6562
rect 13090 6513 13096 6547
rect 13130 6513 13136 6547
rect 13090 6475 13136 6513
rect 13090 6441 13096 6475
rect 13130 6441 13136 6475
rect 13090 6403 13136 6441
rect 13090 6369 13096 6403
rect 13130 6369 13136 6403
rect 13090 6331 13136 6369
rect 13090 6297 13096 6331
rect 13130 6297 13136 6331
rect 13090 6259 13136 6297
rect 13090 6225 13096 6259
rect 13130 6225 13136 6259
rect 13090 6187 13136 6225
rect 13090 6153 13096 6187
rect 13130 6153 13136 6187
rect 13090 6115 13136 6153
rect 13090 6081 13096 6115
rect 13130 6081 13136 6115
rect 13090 6043 13136 6081
rect 13090 6009 13096 6043
rect 13130 6009 13136 6043
rect 13090 5971 13136 6009
rect 13090 5937 13096 5971
rect 13130 5937 13136 5971
rect 13090 5899 13136 5937
rect 13090 5865 13096 5899
rect 13130 5865 13136 5899
rect 13090 5827 13136 5865
rect 13090 5793 13096 5827
rect 13130 5793 13136 5827
rect 13090 5755 13136 5793
rect 13090 5721 13096 5755
rect 13130 5721 13136 5755
rect 13090 5683 13136 5721
rect 13090 5649 13096 5683
rect 13130 5649 13136 5683
rect 13090 5611 13136 5649
rect 13090 5577 13096 5611
rect 13130 5577 13136 5611
rect 13090 5562 13136 5577
rect 13186 6547 13232 6562
rect 13186 6513 13192 6547
rect 13226 6513 13232 6547
rect 13186 6475 13232 6513
rect 13186 6441 13192 6475
rect 13226 6441 13232 6475
rect 13186 6403 13232 6441
rect 13186 6369 13192 6403
rect 13226 6369 13232 6403
rect 13186 6331 13232 6369
rect 13186 6297 13192 6331
rect 13226 6297 13232 6331
rect 13186 6259 13232 6297
rect 13186 6225 13192 6259
rect 13226 6225 13232 6259
rect 13186 6187 13232 6225
rect 13186 6153 13192 6187
rect 13226 6153 13232 6187
rect 13186 6115 13232 6153
rect 13186 6081 13192 6115
rect 13226 6081 13232 6115
rect 13186 6043 13232 6081
rect 13186 6009 13192 6043
rect 13226 6009 13232 6043
rect 13186 5971 13232 6009
rect 13186 5937 13192 5971
rect 13226 5937 13232 5971
rect 13186 5899 13232 5937
rect 13186 5865 13192 5899
rect 13226 5865 13232 5899
rect 13186 5827 13232 5865
rect 13186 5793 13192 5827
rect 13226 5793 13232 5827
rect 13186 5755 13232 5793
rect 13186 5721 13192 5755
rect 13226 5721 13232 5755
rect 13186 5683 13232 5721
rect 13186 5649 13192 5683
rect 13226 5649 13232 5683
rect 13186 5611 13232 5649
rect 13186 5577 13192 5611
rect 13226 5577 13232 5611
rect 13186 5562 13232 5577
rect 13282 6547 13328 6562
rect 13282 6513 13288 6547
rect 13322 6513 13328 6547
rect 13282 6475 13328 6513
rect 13282 6441 13288 6475
rect 13322 6441 13328 6475
rect 13282 6403 13328 6441
rect 13282 6369 13288 6403
rect 13322 6369 13328 6403
rect 13282 6331 13328 6369
rect 13282 6297 13288 6331
rect 13322 6297 13328 6331
rect 13282 6259 13328 6297
rect 13282 6225 13288 6259
rect 13322 6225 13328 6259
rect 13282 6187 13328 6225
rect 13282 6153 13288 6187
rect 13322 6153 13328 6187
rect 13282 6115 13328 6153
rect 13282 6081 13288 6115
rect 13322 6081 13328 6115
rect 13282 6043 13328 6081
rect 13282 6009 13288 6043
rect 13322 6009 13328 6043
rect 13282 5971 13328 6009
rect 13282 5937 13288 5971
rect 13322 5937 13328 5971
rect 13282 5899 13328 5937
rect 13282 5865 13288 5899
rect 13322 5865 13328 5899
rect 13282 5827 13328 5865
rect 13282 5793 13288 5827
rect 13322 5793 13328 5827
rect 13282 5755 13328 5793
rect 13282 5721 13288 5755
rect 13322 5721 13328 5755
rect 13282 5683 13328 5721
rect 13282 5649 13288 5683
rect 13322 5649 13328 5683
rect 13282 5611 13328 5649
rect 13282 5577 13288 5611
rect 13322 5577 13328 5611
rect 13282 5562 13328 5577
rect 13378 6547 13424 6562
rect 13378 6513 13384 6547
rect 13418 6513 13424 6547
rect 13378 6475 13424 6513
rect 13378 6441 13384 6475
rect 13418 6441 13424 6475
rect 13378 6403 13424 6441
rect 13378 6369 13384 6403
rect 13418 6369 13424 6403
rect 13378 6331 13424 6369
rect 13378 6297 13384 6331
rect 13418 6297 13424 6331
rect 13378 6259 13424 6297
rect 13378 6225 13384 6259
rect 13418 6225 13424 6259
rect 13378 6187 13424 6225
rect 13378 6153 13384 6187
rect 13418 6153 13424 6187
rect 13378 6115 13424 6153
rect 13378 6081 13384 6115
rect 13418 6081 13424 6115
rect 13378 6043 13424 6081
rect 13378 6009 13384 6043
rect 13418 6009 13424 6043
rect 13378 5971 13424 6009
rect 13378 5937 13384 5971
rect 13418 5937 13424 5971
rect 13378 5899 13424 5937
rect 13378 5865 13384 5899
rect 13418 5865 13424 5899
rect 13378 5827 13424 5865
rect 13378 5793 13384 5827
rect 13418 5793 13424 5827
rect 13378 5755 13424 5793
rect 13378 5721 13384 5755
rect 13418 5721 13424 5755
rect 13378 5683 13424 5721
rect 13378 5649 13384 5683
rect 13418 5649 13424 5683
rect 13378 5611 13424 5649
rect 13378 5577 13384 5611
rect 13418 5577 13424 5611
rect 13378 5562 13424 5577
rect 13474 6547 13520 6562
rect 13474 6513 13480 6547
rect 13514 6513 13520 6547
rect 13474 6475 13520 6513
rect 13474 6441 13480 6475
rect 13514 6441 13520 6475
rect 13474 6403 13520 6441
rect 13474 6369 13480 6403
rect 13514 6369 13520 6403
rect 13474 6331 13520 6369
rect 13474 6297 13480 6331
rect 13514 6297 13520 6331
rect 13474 6259 13520 6297
rect 13474 6225 13480 6259
rect 13514 6225 13520 6259
rect 13474 6187 13520 6225
rect 13474 6153 13480 6187
rect 13514 6153 13520 6187
rect 13474 6115 13520 6153
rect 13474 6081 13480 6115
rect 13514 6081 13520 6115
rect 13474 6043 13520 6081
rect 13474 6009 13480 6043
rect 13514 6009 13520 6043
rect 13474 5971 13520 6009
rect 13474 5937 13480 5971
rect 13514 5937 13520 5971
rect 13474 5899 13520 5937
rect 13474 5865 13480 5899
rect 13514 5865 13520 5899
rect 13474 5827 13520 5865
rect 13474 5793 13480 5827
rect 13514 5793 13520 5827
rect 13474 5755 13520 5793
rect 13474 5721 13480 5755
rect 13514 5721 13520 5755
rect 13474 5683 13520 5721
rect 13474 5649 13480 5683
rect 13514 5649 13520 5683
rect 13474 5611 13520 5649
rect 13474 5577 13480 5611
rect 13514 5577 13520 5611
rect 13474 5562 13520 5577
rect 13570 6547 13616 6562
rect 13570 6513 13576 6547
rect 13610 6513 13616 6547
rect 13570 6475 13616 6513
rect 13570 6441 13576 6475
rect 13610 6441 13616 6475
rect 13570 6403 13616 6441
rect 13570 6369 13576 6403
rect 13610 6369 13616 6403
rect 13570 6331 13616 6369
rect 13570 6297 13576 6331
rect 13610 6297 13616 6331
rect 13570 6259 13616 6297
rect 13570 6225 13576 6259
rect 13610 6225 13616 6259
rect 13570 6187 13616 6225
rect 13570 6153 13576 6187
rect 13610 6153 13616 6187
rect 13570 6115 13616 6153
rect 13570 6081 13576 6115
rect 13610 6081 13616 6115
rect 13570 6043 13616 6081
rect 13570 6009 13576 6043
rect 13610 6009 13616 6043
rect 13570 5971 13616 6009
rect 13570 5937 13576 5971
rect 13610 5937 13616 5971
rect 13570 5899 13616 5937
rect 13570 5865 13576 5899
rect 13610 5865 13616 5899
rect 13570 5827 13616 5865
rect 13570 5793 13576 5827
rect 13610 5793 13616 5827
rect 13570 5755 13616 5793
rect 13570 5721 13576 5755
rect 13610 5721 13616 5755
rect 13570 5683 13616 5721
rect 13570 5649 13576 5683
rect 13610 5649 13616 5683
rect 13570 5611 13616 5649
rect 13570 5577 13576 5611
rect 13610 5577 13616 5611
rect 13570 5562 13616 5577
rect 14184 6543 14230 6558
rect 14184 6509 14190 6543
rect 14224 6509 14230 6543
rect 14184 6471 14230 6509
rect 14184 6437 14190 6471
rect 14224 6437 14230 6471
rect 14184 6399 14230 6437
rect 14184 6365 14190 6399
rect 14224 6365 14230 6399
rect 14184 6327 14230 6365
rect 14184 6293 14190 6327
rect 14224 6293 14230 6327
rect 14184 6255 14230 6293
rect 14184 6221 14190 6255
rect 14224 6221 14230 6255
rect 14184 6183 14230 6221
rect 14184 6149 14190 6183
rect 14224 6149 14230 6183
rect 14184 6111 14230 6149
rect 14184 6077 14190 6111
rect 14224 6077 14230 6111
rect 14184 6039 14230 6077
rect 14184 6005 14190 6039
rect 14224 6005 14230 6039
rect 14184 5967 14230 6005
rect 14184 5933 14190 5967
rect 14224 5933 14230 5967
rect 14184 5895 14230 5933
rect 14184 5861 14190 5895
rect 14224 5861 14230 5895
rect 14184 5823 14230 5861
rect 14184 5789 14190 5823
rect 14224 5789 14230 5823
rect 14184 5751 14230 5789
rect 14184 5717 14190 5751
rect 14224 5717 14230 5751
rect 14184 5679 14230 5717
rect 14184 5645 14190 5679
rect 14224 5645 14230 5679
rect 14184 5607 14230 5645
rect 14184 5573 14190 5607
rect 14224 5573 14230 5607
rect 14184 5558 14230 5573
rect 14280 6543 14326 6558
rect 14280 6509 14286 6543
rect 14320 6509 14326 6543
rect 14280 6471 14326 6509
rect 14280 6437 14286 6471
rect 14320 6437 14326 6471
rect 14280 6399 14326 6437
rect 14280 6365 14286 6399
rect 14320 6365 14326 6399
rect 14280 6327 14326 6365
rect 14280 6293 14286 6327
rect 14320 6293 14326 6327
rect 14280 6255 14326 6293
rect 14280 6221 14286 6255
rect 14320 6221 14326 6255
rect 14280 6183 14326 6221
rect 14280 6149 14286 6183
rect 14320 6149 14326 6183
rect 14280 6111 14326 6149
rect 14280 6077 14286 6111
rect 14320 6077 14326 6111
rect 14280 6039 14326 6077
rect 14280 6005 14286 6039
rect 14320 6005 14326 6039
rect 14280 5967 14326 6005
rect 14280 5933 14286 5967
rect 14320 5933 14326 5967
rect 14280 5895 14326 5933
rect 14280 5861 14286 5895
rect 14320 5861 14326 5895
rect 14280 5823 14326 5861
rect 14280 5789 14286 5823
rect 14320 5789 14326 5823
rect 14280 5751 14326 5789
rect 14280 5717 14286 5751
rect 14320 5717 14326 5751
rect 14280 5679 14326 5717
rect 14280 5645 14286 5679
rect 14320 5645 14326 5679
rect 14280 5607 14326 5645
rect 14280 5573 14286 5607
rect 14320 5573 14326 5607
rect 14280 5558 14326 5573
rect 14376 6543 14422 6558
rect 14376 6509 14382 6543
rect 14416 6509 14422 6543
rect 14376 6471 14422 6509
rect 14376 6437 14382 6471
rect 14416 6437 14422 6471
rect 14376 6399 14422 6437
rect 14376 6365 14382 6399
rect 14416 6365 14422 6399
rect 14376 6327 14422 6365
rect 14376 6293 14382 6327
rect 14416 6293 14422 6327
rect 14376 6255 14422 6293
rect 14376 6221 14382 6255
rect 14416 6221 14422 6255
rect 14376 6183 14422 6221
rect 14376 6149 14382 6183
rect 14416 6149 14422 6183
rect 14376 6111 14422 6149
rect 14376 6077 14382 6111
rect 14416 6077 14422 6111
rect 14376 6039 14422 6077
rect 14376 6005 14382 6039
rect 14416 6005 14422 6039
rect 14376 5967 14422 6005
rect 14376 5933 14382 5967
rect 14416 5933 14422 5967
rect 14376 5895 14422 5933
rect 14376 5861 14382 5895
rect 14416 5861 14422 5895
rect 14376 5823 14422 5861
rect 14376 5789 14382 5823
rect 14416 5789 14422 5823
rect 14376 5751 14422 5789
rect 14376 5717 14382 5751
rect 14416 5717 14422 5751
rect 14376 5679 14422 5717
rect 14376 5645 14382 5679
rect 14416 5645 14422 5679
rect 14376 5607 14422 5645
rect 14376 5573 14382 5607
rect 14416 5573 14422 5607
rect 14376 5558 14422 5573
rect 14472 6543 14518 6558
rect 14472 6509 14478 6543
rect 14512 6509 14518 6543
rect 14472 6471 14518 6509
rect 14472 6437 14478 6471
rect 14512 6437 14518 6471
rect 14472 6399 14518 6437
rect 14472 6365 14478 6399
rect 14512 6365 14518 6399
rect 14472 6327 14518 6365
rect 14472 6293 14478 6327
rect 14512 6293 14518 6327
rect 14472 6255 14518 6293
rect 14472 6221 14478 6255
rect 14512 6221 14518 6255
rect 14472 6183 14518 6221
rect 14472 6149 14478 6183
rect 14512 6149 14518 6183
rect 14472 6111 14518 6149
rect 14472 6077 14478 6111
rect 14512 6077 14518 6111
rect 14472 6039 14518 6077
rect 14472 6005 14478 6039
rect 14512 6005 14518 6039
rect 14472 5967 14518 6005
rect 14472 5933 14478 5967
rect 14512 5933 14518 5967
rect 14472 5895 14518 5933
rect 14472 5861 14478 5895
rect 14512 5861 14518 5895
rect 14472 5823 14518 5861
rect 14472 5789 14478 5823
rect 14512 5789 14518 5823
rect 14472 5751 14518 5789
rect 14472 5717 14478 5751
rect 14512 5717 14518 5751
rect 14472 5679 14518 5717
rect 14472 5645 14478 5679
rect 14512 5645 14518 5679
rect 14472 5607 14518 5645
rect 14472 5573 14478 5607
rect 14512 5573 14518 5607
rect 14472 5558 14518 5573
rect 14568 6543 14614 6558
rect 14568 6509 14574 6543
rect 14608 6509 14614 6543
rect 14568 6471 14614 6509
rect 14568 6437 14574 6471
rect 14608 6437 14614 6471
rect 14568 6399 14614 6437
rect 14568 6365 14574 6399
rect 14608 6365 14614 6399
rect 14568 6327 14614 6365
rect 14568 6293 14574 6327
rect 14608 6293 14614 6327
rect 14568 6255 14614 6293
rect 14568 6221 14574 6255
rect 14608 6221 14614 6255
rect 14568 6183 14614 6221
rect 14568 6149 14574 6183
rect 14608 6149 14614 6183
rect 14568 6111 14614 6149
rect 14568 6077 14574 6111
rect 14608 6077 14614 6111
rect 14568 6039 14614 6077
rect 14568 6005 14574 6039
rect 14608 6005 14614 6039
rect 14568 5967 14614 6005
rect 14568 5933 14574 5967
rect 14608 5933 14614 5967
rect 14568 5895 14614 5933
rect 14568 5861 14574 5895
rect 14608 5861 14614 5895
rect 14568 5823 14614 5861
rect 14568 5789 14574 5823
rect 14608 5789 14614 5823
rect 14568 5751 14614 5789
rect 14568 5717 14574 5751
rect 14608 5717 14614 5751
rect 14568 5679 14614 5717
rect 14568 5645 14574 5679
rect 14608 5645 14614 5679
rect 14568 5607 14614 5645
rect 14568 5573 14574 5607
rect 14608 5573 14614 5607
rect 14568 5558 14614 5573
rect 14664 6543 14710 6558
rect 14664 6509 14670 6543
rect 14704 6509 14710 6543
rect 14664 6471 14710 6509
rect 14664 6437 14670 6471
rect 14704 6437 14710 6471
rect 14664 6399 14710 6437
rect 14664 6365 14670 6399
rect 14704 6365 14710 6399
rect 14664 6327 14710 6365
rect 14664 6293 14670 6327
rect 14704 6293 14710 6327
rect 14664 6255 14710 6293
rect 14664 6221 14670 6255
rect 14704 6221 14710 6255
rect 14664 6183 14710 6221
rect 14664 6149 14670 6183
rect 14704 6149 14710 6183
rect 14664 6111 14710 6149
rect 14664 6077 14670 6111
rect 14704 6077 14710 6111
rect 14664 6039 14710 6077
rect 14664 6005 14670 6039
rect 14704 6005 14710 6039
rect 14664 5967 14710 6005
rect 14664 5933 14670 5967
rect 14704 5933 14710 5967
rect 14664 5895 14710 5933
rect 14664 5861 14670 5895
rect 14704 5861 14710 5895
rect 14664 5823 14710 5861
rect 14664 5789 14670 5823
rect 14704 5789 14710 5823
rect 14664 5751 14710 5789
rect 14664 5717 14670 5751
rect 14704 5717 14710 5751
rect 14664 5679 14710 5717
rect 14664 5645 14670 5679
rect 14704 5645 14710 5679
rect 14664 5607 14710 5645
rect 14664 5573 14670 5607
rect 14704 5573 14710 5607
rect 14664 5558 14710 5573
rect 14760 6543 14806 6558
rect 14760 6509 14766 6543
rect 14800 6509 14806 6543
rect 14760 6471 14806 6509
rect 14760 6437 14766 6471
rect 14800 6437 14806 6471
rect 14760 6399 14806 6437
rect 14760 6365 14766 6399
rect 14800 6365 14806 6399
rect 14760 6327 14806 6365
rect 14760 6293 14766 6327
rect 14800 6293 14806 6327
rect 14760 6255 14806 6293
rect 14760 6221 14766 6255
rect 14800 6221 14806 6255
rect 14760 6183 14806 6221
rect 14760 6149 14766 6183
rect 14800 6149 14806 6183
rect 14760 6111 14806 6149
rect 14760 6077 14766 6111
rect 14800 6077 14806 6111
rect 14760 6039 14806 6077
rect 14760 6005 14766 6039
rect 14800 6005 14806 6039
rect 14760 5967 14806 6005
rect 14760 5933 14766 5967
rect 14800 5933 14806 5967
rect 14760 5895 14806 5933
rect 14760 5861 14766 5895
rect 14800 5861 14806 5895
rect 14760 5823 14806 5861
rect 14760 5789 14766 5823
rect 14800 5789 14806 5823
rect 14760 5751 14806 5789
rect 14760 5717 14766 5751
rect 14800 5717 14806 5751
rect 14760 5679 14806 5717
rect 14760 5645 14766 5679
rect 14800 5645 14806 5679
rect 14760 5607 14806 5645
rect 14760 5573 14766 5607
rect 14800 5573 14806 5607
rect 14760 5558 14806 5573
rect 14856 6543 14902 6558
rect 14856 6509 14862 6543
rect 14896 6509 14902 6543
rect 14856 6471 14902 6509
rect 14856 6437 14862 6471
rect 14896 6437 14902 6471
rect 14856 6399 14902 6437
rect 14856 6365 14862 6399
rect 14896 6365 14902 6399
rect 14856 6327 14902 6365
rect 14856 6293 14862 6327
rect 14896 6293 14902 6327
rect 14856 6255 14902 6293
rect 14856 6221 14862 6255
rect 14896 6221 14902 6255
rect 14856 6183 14902 6221
rect 14856 6149 14862 6183
rect 14896 6149 14902 6183
rect 14856 6111 14902 6149
rect 14856 6077 14862 6111
rect 14896 6077 14902 6111
rect 14856 6039 14902 6077
rect 14856 6005 14862 6039
rect 14896 6005 14902 6039
rect 14856 5967 14902 6005
rect 14856 5933 14862 5967
rect 14896 5933 14902 5967
rect 14856 5895 14902 5933
rect 14856 5861 14862 5895
rect 14896 5861 14902 5895
rect 14856 5823 14902 5861
rect 14856 5789 14862 5823
rect 14896 5789 14902 5823
rect 14856 5751 14902 5789
rect 14856 5717 14862 5751
rect 14896 5717 14902 5751
rect 14856 5679 14902 5717
rect 14856 5645 14862 5679
rect 14896 5645 14902 5679
rect 14856 5607 14902 5645
rect 14856 5573 14862 5607
rect 14896 5573 14902 5607
rect 14856 5558 14902 5573
rect 14952 6543 14998 6558
rect 14952 6509 14958 6543
rect 14992 6509 14998 6543
rect 14952 6471 14998 6509
rect 14952 6437 14958 6471
rect 14992 6437 14998 6471
rect 14952 6399 14998 6437
rect 14952 6365 14958 6399
rect 14992 6365 14998 6399
rect 14952 6327 14998 6365
rect 14952 6293 14958 6327
rect 14992 6293 14998 6327
rect 14952 6255 14998 6293
rect 15582 6345 15676 6356
rect 15582 6293 15603 6345
rect 15655 6293 15676 6345
rect 15582 6282 15676 6293
rect 14952 6221 14958 6255
rect 14992 6221 14998 6255
rect 14952 6183 14998 6221
rect 14952 6149 14958 6183
rect 14992 6149 14998 6183
rect 14952 6111 14998 6149
rect 15592 6182 15666 6282
rect 15592 6148 15614 6182
rect 15648 6148 15666 6182
rect 15592 6126 15666 6148
rect 14952 6077 14958 6111
rect 14992 6077 14998 6111
rect 14952 6039 14998 6077
rect 14952 6005 14958 6039
rect 14992 6005 14998 6039
rect 14952 5967 14998 6005
rect 14952 5933 14958 5967
rect 14992 5933 14998 5967
rect 14952 5895 14998 5933
rect 14952 5861 14958 5895
rect 14992 5861 14998 5895
rect 14952 5823 14998 5861
rect 14952 5789 14958 5823
rect 14992 5789 14998 5823
rect 14952 5751 14998 5789
rect 14952 5717 14958 5751
rect 14992 5717 14998 5751
rect 14952 5679 14998 5717
rect 14952 5645 14958 5679
rect 14992 5645 14998 5679
rect 14952 5607 14998 5645
rect 14952 5573 14958 5607
rect 14992 5573 14998 5607
rect 14952 5558 14998 5573
rect 15512 5879 15558 5926
rect 15512 5845 15518 5879
rect 15552 5845 15558 5879
rect 15512 5807 15558 5845
rect 15512 5773 15518 5807
rect 15552 5773 15558 5807
rect 15512 5735 15558 5773
rect 15512 5701 15518 5735
rect 15552 5701 15558 5735
rect 15512 5663 15558 5701
rect 15512 5629 15518 5663
rect 15552 5629 15558 5663
rect 15512 5591 15558 5629
rect 15512 5557 15518 5591
rect 15552 5557 15558 5591
rect 15512 5519 15558 5557
rect 15512 5485 15518 5519
rect 15552 5485 15558 5519
rect 15512 5447 15558 5485
rect 858 5406 942 5420
rect 858 5372 880 5406
rect 914 5372 942 5406
rect 858 5264 942 5372
rect 2312 5410 2408 5430
rect 2312 5376 2344 5410
rect 2378 5376 2408 5410
rect 2312 5264 2408 5376
rect 858 5190 2408 5264
rect 3802 5390 3898 5408
rect 3802 5356 3836 5390
rect 3870 5356 3898 5390
rect 3802 5248 3898 5356
rect 5262 5394 5364 5414
rect 5262 5360 5300 5394
rect 5334 5360 5364 5394
rect 5262 5248 5364 5360
rect 1570 5124 1624 5190
rect 3800 5164 5364 5248
rect 6828 5390 6930 5420
rect 6828 5356 6866 5390
rect 6900 5356 6930 5390
rect 6828 5268 6930 5356
rect 8290 5394 8396 5414
rect 8290 5360 8330 5394
rect 8364 5360 8396 5394
rect 8290 5268 8396 5360
rect 6828 5170 8396 5268
rect 9920 5388 10026 5400
rect 9920 5354 9954 5388
rect 9988 5354 10026 5388
rect 9920 5270 10026 5354
rect 11370 5392 11494 5414
rect 11370 5358 11418 5392
rect 11452 5358 11494 5392
rect 15512 5413 15518 5447
rect 15552 5413 15558 5447
rect 11370 5270 11494 5358
rect 1570 5090 1580 5124
rect 1614 5090 1624 5124
rect 1570 5074 1624 5090
rect 4526 5108 4580 5164
rect 4526 5074 4536 5108
rect 4570 5074 4580 5108
rect 4526 5058 4580 5074
rect 7556 5108 7610 5170
rect 9920 5156 11494 5270
rect 13070 5362 13194 5380
rect 13070 5328 13110 5362
rect 13144 5328 13194 5362
rect 13070 5236 13194 5328
rect 14528 5366 14650 5386
rect 14528 5332 14574 5366
rect 14608 5332 14650 5366
rect 14528 5236 14650 5332
rect 7556 5074 7566 5108
rect 7600 5074 7610 5108
rect 7556 5058 7610 5074
rect 10644 5106 10698 5156
rect 13070 5122 14650 5236
rect 15512 5375 15558 5413
rect 15512 5341 15518 5375
rect 15552 5341 15558 5375
rect 15512 5303 15558 5341
rect 15512 5269 15518 5303
rect 15552 5269 15558 5303
rect 15512 5231 15558 5269
rect 15512 5197 15518 5231
rect 15552 5197 15558 5231
rect 15512 5159 15558 5197
rect 15512 5125 15518 5159
rect 15552 5125 15558 5159
rect 10644 5072 10654 5106
rect 10688 5072 10698 5106
rect 10644 5056 10698 5072
rect 13800 5080 13854 5122
rect 13800 5046 13810 5080
rect 13844 5046 13854 5080
rect 13800 5030 13854 5046
rect 15512 5087 15558 5125
rect 15512 5053 15518 5087
rect 15552 5053 15558 5087
rect 15512 5015 15558 5053
rect 15512 4981 15518 5015
rect 15552 4981 15558 5015
rect -1126 4769 -402 4792
rect -1126 4735 -1067 4769
rect -1033 4735 -402 4769
rect -1126 4630 -402 4735
rect 1478 4929 1524 4944
rect 1478 4895 1484 4929
rect 1518 4895 1524 4929
rect 1478 4857 1524 4895
rect 1478 4823 1484 4857
rect 1518 4823 1524 4857
rect 1478 4785 1524 4823
rect 1478 4751 1484 4785
rect 1518 4751 1524 4785
rect 1478 4713 1524 4751
rect 1478 4679 1484 4713
rect 1518 4679 1524 4713
rect 1478 4641 1524 4679
rect -1906 3354 -1896 3462
rect -1782 3442 -1772 3462
rect -1782 3434 -1546 3442
rect -1782 3428 -1544 3434
rect -1782 3394 -1590 3428
rect -1556 3394 -1544 3428
rect -1782 3388 -1544 3394
rect -1782 3380 -1546 3388
rect -1782 3372 -1590 3380
rect -1782 3354 -1772 3372
rect -1126 3324 -1020 4630
rect 1478 4607 1484 4641
rect 1518 4607 1524 4641
rect 1478 4569 1524 4607
rect 1478 4535 1484 4569
rect 1518 4535 1524 4569
rect 1478 4497 1524 4535
rect 1478 4463 1484 4497
rect 1518 4463 1524 4497
rect 1478 4425 1524 4463
rect 1478 4391 1484 4425
rect 1518 4391 1524 4425
rect 1478 4353 1524 4391
rect 1478 4319 1484 4353
rect 1518 4319 1524 4353
rect 1478 4281 1524 4319
rect 1478 4247 1484 4281
rect 1518 4247 1524 4281
rect 1478 4209 1524 4247
rect 1478 4175 1484 4209
rect 1518 4175 1524 4209
rect 1478 4137 1524 4175
rect 1478 4103 1484 4137
rect 1518 4103 1524 4137
rect 1478 4065 1524 4103
rect 1478 4031 1484 4065
rect 1518 4031 1524 4065
rect 1478 3993 1524 4031
rect 1478 3959 1484 3993
rect 1518 3959 1524 3993
rect 1478 3944 1524 3959
rect 1574 4929 1620 4944
rect 1574 4895 1580 4929
rect 1614 4895 1620 4929
rect 1574 4857 1620 4895
rect 1574 4823 1580 4857
rect 1614 4823 1620 4857
rect 1574 4785 1620 4823
rect 1574 4751 1580 4785
rect 1614 4751 1620 4785
rect 1574 4713 1620 4751
rect 1574 4679 1580 4713
rect 1614 4679 1620 4713
rect 1574 4641 1620 4679
rect 1574 4607 1580 4641
rect 1614 4607 1620 4641
rect 1574 4569 1620 4607
rect 1574 4535 1580 4569
rect 1614 4535 1620 4569
rect 1574 4497 1620 4535
rect 1574 4463 1580 4497
rect 1614 4463 1620 4497
rect 1574 4425 1620 4463
rect 1574 4391 1580 4425
rect 1614 4391 1620 4425
rect 1574 4353 1620 4391
rect 1574 4319 1580 4353
rect 1614 4319 1620 4353
rect 1574 4281 1620 4319
rect 1574 4247 1580 4281
rect 1614 4247 1620 4281
rect 1574 4209 1620 4247
rect 1574 4175 1580 4209
rect 1614 4175 1620 4209
rect 1574 4137 1620 4175
rect 1574 4103 1580 4137
rect 1614 4103 1620 4137
rect 1574 4065 1620 4103
rect 1574 4031 1580 4065
rect 1614 4031 1620 4065
rect 1574 3993 1620 4031
rect 1574 3959 1580 3993
rect 1614 3959 1620 3993
rect 1574 3944 1620 3959
rect 1670 4929 1716 4944
rect 1670 4895 1676 4929
rect 1710 4895 1716 4929
rect 1670 4857 1716 4895
rect 1670 4823 1676 4857
rect 1710 4823 1716 4857
rect 1670 4785 1716 4823
rect 1670 4751 1676 4785
rect 1710 4751 1716 4785
rect 1670 4713 1716 4751
rect 1670 4679 1676 4713
rect 1710 4679 1716 4713
rect 1670 4641 1716 4679
rect 1670 4607 1676 4641
rect 1710 4607 1716 4641
rect 1670 4569 1716 4607
rect 1670 4535 1676 4569
rect 1710 4535 1716 4569
rect 1670 4497 1716 4535
rect 1670 4463 1676 4497
rect 1710 4463 1716 4497
rect 1670 4425 1716 4463
rect 1670 4391 1676 4425
rect 1710 4391 1716 4425
rect 1670 4353 1716 4391
rect 1670 4319 1676 4353
rect 1710 4319 1716 4353
rect 1670 4281 1716 4319
rect 1670 4247 1676 4281
rect 1710 4247 1716 4281
rect 1670 4209 1716 4247
rect 1670 4175 1676 4209
rect 1710 4175 1716 4209
rect 1670 4137 1716 4175
rect 1670 4103 1676 4137
rect 1710 4103 1716 4137
rect 1670 4065 1716 4103
rect 1670 4031 1676 4065
rect 1710 4031 1716 4065
rect 1670 3993 1716 4031
rect 1670 3959 1676 3993
rect 1710 3959 1716 3993
rect 1670 3944 1716 3959
rect 1766 4929 1812 4944
rect 1766 4895 1772 4929
rect 1806 4895 1812 4929
rect 1766 4857 1812 4895
rect 1766 4823 1772 4857
rect 1806 4823 1812 4857
rect 1766 4785 1812 4823
rect 1766 4751 1772 4785
rect 1806 4751 1812 4785
rect 1766 4713 1812 4751
rect 1766 4679 1772 4713
rect 1806 4679 1812 4713
rect 1766 4641 1812 4679
rect 1766 4607 1772 4641
rect 1806 4607 1812 4641
rect 1766 4569 1812 4607
rect 1766 4535 1772 4569
rect 1806 4535 1812 4569
rect 1766 4497 1812 4535
rect 1766 4463 1772 4497
rect 1806 4463 1812 4497
rect 1766 4425 1812 4463
rect 1766 4391 1772 4425
rect 1806 4391 1812 4425
rect 1766 4353 1812 4391
rect 1766 4319 1772 4353
rect 1806 4319 1812 4353
rect 1766 4281 1812 4319
rect 1766 4247 1772 4281
rect 1806 4247 1812 4281
rect 1766 4209 1812 4247
rect 1766 4175 1772 4209
rect 1806 4175 1812 4209
rect 1766 4137 1812 4175
rect 1766 4103 1772 4137
rect 1806 4103 1812 4137
rect 1766 4065 1812 4103
rect 1766 4031 1772 4065
rect 1806 4031 1812 4065
rect 1766 3993 1812 4031
rect 1766 3959 1772 3993
rect 1806 3959 1812 3993
rect 1766 3944 1812 3959
rect 1862 4929 1908 4944
rect 1862 4895 1868 4929
rect 1902 4895 1908 4929
rect 15512 4943 15558 4981
rect 1862 4857 1908 4895
rect 1862 4823 1868 4857
rect 1902 4823 1908 4857
rect 1862 4785 1908 4823
rect 1862 4751 1868 4785
rect 1902 4751 1908 4785
rect 1862 4713 1908 4751
rect 1862 4679 1868 4713
rect 1902 4679 1908 4713
rect 1862 4641 1908 4679
rect 1862 4607 1868 4641
rect 1902 4607 1908 4641
rect 1862 4569 1908 4607
rect 1862 4535 1868 4569
rect 1902 4535 1908 4569
rect 1862 4497 1908 4535
rect 1862 4463 1868 4497
rect 1902 4463 1908 4497
rect 1862 4425 1908 4463
rect 1862 4391 1868 4425
rect 1902 4391 1908 4425
rect 1862 4353 1908 4391
rect 1862 4319 1868 4353
rect 1902 4319 1908 4353
rect 1862 4281 1908 4319
rect 1862 4247 1868 4281
rect 1902 4247 1908 4281
rect 1862 4209 1908 4247
rect 1862 4175 1868 4209
rect 1902 4175 1908 4209
rect 1862 4137 1908 4175
rect 1862 4103 1868 4137
rect 1902 4103 1908 4137
rect 1862 4065 1908 4103
rect 1862 4031 1868 4065
rect 1902 4031 1908 4065
rect 1862 3993 1908 4031
rect 1862 3959 1868 3993
rect 1902 3959 1908 3993
rect 1862 3944 1908 3959
rect 4434 4913 4480 4928
rect 4434 4879 4440 4913
rect 4474 4879 4480 4913
rect 4434 4841 4480 4879
rect 4434 4807 4440 4841
rect 4474 4807 4480 4841
rect 4434 4769 4480 4807
rect 4434 4735 4440 4769
rect 4474 4735 4480 4769
rect 4434 4697 4480 4735
rect 4434 4663 4440 4697
rect 4474 4663 4480 4697
rect 4434 4625 4480 4663
rect 4434 4591 4440 4625
rect 4474 4591 4480 4625
rect 4434 4553 4480 4591
rect 4434 4519 4440 4553
rect 4474 4519 4480 4553
rect 4434 4481 4480 4519
rect 4434 4447 4440 4481
rect 4474 4447 4480 4481
rect 4434 4409 4480 4447
rect 4434 4375 4440 4409
rect 4474 4375 4480 4409
rect 4434 4337 4480 4375
rect 4434 4303 4440 4337
rect 4474 4303 4480 4337
rect 4434 4265 4480 4303
rect 4434 4231 4440 4265
rect 4474 4231 4480 4265
rect 4434 4193 4480 4231
rect 4434 4159 4440 4193
rect 4474 4159 4480 4193
rect 4434 4121 4480 4159
rect 4434 4087 4440 4121
rect 4474 4087 4480 4121
rect 4434 4049 4480 4087
rect 4434 4015 4440 4049
rect 4474 4015 4480 4049
rect 4434 3977 4480 4015
rect 4434 3943 4440 3977
rect 4474 3943 4480 3977
rect 4434 3928 4480 3943
rect 4530 4913 4576 4928
rect 4530 4879 4536 4913
rect 4570 4879 4576 4913
rect 4530 4841 4576 4879
rect 4530 4807 4536 4841
rect 4570 4807 4576 4841
rect 4530 4769 4576 4807
rect 4530 4735 4536 4769
rect 4570 4735 4576 4769
rect 4530 4697 4576 4735
rect 4530 4663 4536 4697
rect 4570 4663 4576 4697
rect 4530 4625 4576 4663
rect 4530 4591 4536 4625
rect 4570 4591 4576 4625
rect 4530 4553 4576 4591
rect 4530 4519 4536 4553
rect 4570 4519 4576 4553
rect 4530 4481 4576 4519
rect 4530 4447 4536 4481
rect 4570 4447 4576 4481
rect 4530 4409 4576 4447
rect 4530 4375 4536 4409
rect 4570 4375 4576 4409
rect 4530 4337 4576 4375
rect 4530 4303 4536 4337
rect 4570 4303 4576 4337
rect 4530 4265 4576 4303
rect 4530 4231 4536 4265
rect 4570 4231 4576 4265
rect 4530 4193 4576 4231
rect 4530 4159 4536 4193
rect 4570 4159 4576 4193
rect 4530 4121 4576 4159
rect 4530 4087 4536 4121
rect 4570 4087 4576 4121
rect 4530 4049 4576 4087
rect 4530 4015 4536 4049
rect 4570 4015 4576 4049
rect 4530 3977 4576 4015
rect 4530 3943 4536 3977
rect 4570 3943 4576 3977
rect 4530 3928 4576 3943
rect 4626 4913 4672 4928
rect 4626 4879 4632 4913
rect 4666 4879 4672 4913
rect 4626 4841 4672 4879
rect 4626 4807 4632 4841
rect 4666 4807 4672 4841
rect 4626 4769 4672 4807
rect 4626 4735 4632 4769
rect 4666 4735 4672 4769
rect 4626 4697 4672 4735
rect 4626 4663 4632 4697
rect 4666 4663 4672 4697
rect 4626 4625 4672 4663
rect 4626 4591 4632 4625
rect 4666 4591 4672 4625
rect 4626 4553 4672 4591
rect 4626 4519 4632 4553
rect 4666 4519 4672 4553
rect 4626 4481 4672 4519
rect 4626 4447 4632 4481
rect 4666 4447 4672 4481
rect 4626 4409 4672 4447
rect 4626 4375 4632 4409
rect 4666 4375 4672 4409
rect 4626 4337 4672 4375
rect 4626 4303 4632 4337
rect 4666 4303 4672 4337
rect 4626 4265 4672 4303
rect 4626 4231 4632 4265
rect 4666 4231 4672 4265
rect 4626 4193 4672 4231
rect 4626 4159 4632 4193
rect 4666 4159 4672 4193
rect 4626 4121 4672 4159
rect 4626 4087 4632 4121
rect 4666 4087 4672 4121
rect 4626 4049 4672 4087
rect 4626 4015 4632 4049
rect 4666 4015 4672 4049
rect 4626 3977 4672 4015
rect 4626 3943 4632 3977
rect 4666 3943 4672 3977
rect 4626 3928 4672 3943
rect 4722 4913 4768 4928
rect 4722 4879 4728 4913
rect 4762 4879 4768 4913
rect 4722 4841 4768 4879
rect 4722 4807 4728 4841
rect 4762 4807 4768 4841
rect 4722 4769 4768 4807
rect 4722 4735 4728 4769
rect 4762 4735 4768 4769
rect 4722 4697 4768 4735
rect 4722 4663 4728 4697
rect 4762 4663 4768 4697
rect 4722 4625 4768 4663
rect 4722 4591 4728 4625
rect 4762 4591 4768 4625
rect 4722 4553 4768 4591
rect 4722 4519 4728 4553
rect 4762 4519 4768 4553
rect 4722 4481 4768 4519
rect 4722 4447 4728 4481
rect 4762 4447 4768 4481
rect 4722 4409 4768 4447
rect 4722 4375 4728 4409
rect 4762 4375 4768 4409
rect 4722 4337 4768 4375
rect 4722 4303 4728 4337
rect 4762 4303 4768 4337
rect 4722 4265 4768 4303
rect 4722 4231 4728 4265
rect 4762 4231 4768 4265
rect 4722 4193 4768 4231
rect 4722 4159 4728 4193
rect 4762 4159 4768 4193
rect 4722 4121 4768 4159
rect 4722 4087 4728 4121
rect 4762 4087 4768 4121
rect 4722 4049 4768 4087
rect 4722 4015 4728 4049
rect 4762 4015 4768 4049
rect 4722 3977 4768 4015
rect 4722 3943 4728 3977
rect 4762 3943 4768 3977
rect 4722 3928 4768 3943
rect 4818 4913 4864 4928
rect 4818 4879 4824 4913
rect 4858 4879 4864 4913
rect 4818 4841 4864 4879
rect 4818 4807 4824 4841
rect 4858 4807 4864 4841
rect 4818 4769 4864 4807
rect 4818 4735 4824 4769
rect 4858 4735 4864 4769
rect 4818 4697 4864 4735
rect 4818 4663 4824 4697
rect 4858 4663 4864 4697
rect 4818 4625 4864 4663
rect 4818 4591 4824 4625
rect 4858 4591 4864 4625
rect 4818 4553 4864 4591
rect 4818 4519 4824 4553
rect 4858 4519 4864 4553
rect 4818 4481 4864 4519
rect 4818 4447 4824 4481
rect 4858 4447 4864 4481
rect 4818 4409 4864 4447
rect 4818 4375 4824 4409
rect 4858 4375 4864 4409
rect 4818 4337 4864 4375
rect 4818 4303 4824 4337
rect 4858 4303 4864 4337
rect 4818 4265 4864 4303
rect 4818 4231 4824 4265
rect 4858 4231 4864 4265
rect 4818 4193 4864 4231
rect 4818 4159 4824 4193
rect 4858 4159 4864 4193
rect 4818 4121 4864 4159
rect 4818 4087 4824 4121
rect 4858 4087 4864 4121
rect 4818 4049 4864 4087
rect 4818 4015 4824 4049
rect 4858 4015 4864 4049
rect 4818 3977 4864 4015
rect 4818 3943 4824 3977
rect 4858 3943 4864 3977
rect 4818 3928 4864 3943
rect 7464 4913 7510 4928
rect 7464 4879 7470 4913
rect 7504 4879 7510 4913
rect 7464 4841 7510 4879
rect 7464 4807 7470 4841
rect 7504 4807 7510 4841
rect 7464 4769 7510 4807
rect 7464 4735 7470 4769
rect 7504 4735 7510 4769
rect 7464 4697 7510 4735
rect 7464 4663 7470 4697
rect 7504 4663 7510 4697
rect 7464 4625 7510 4663
rect 7464 4591 7470 4625
rect 7504 4591 7510 4625
rect 7464 4553 7510 4591
rect 7464 4519 7470 4553
rect 7504 4519 7510 4553
rect 7464 4481 7510 4519
rect 7464 4447 7470 4481
rect 7504 4447 7510 4481
rect 7464 4409 7510 4447
rect 7464 4375 7470 4409
rect 7504 4375 7510 4409
rect 7464 4337 7510 4375
rect 7464 4303 7470 4337
rect 7504 4303 7510 4337
rect 7464 4265 7510 4303
rect 7464 4231 7470 4265
rect 7504 4231 7510 4265
rect 7464 4193 7510 4231
rect 7464 4159 7470 4193
rect 7504 4159 7510 4193
rect 7464 4121 7510 4159
rect 7464 4087 7470 4121
rect 7504 4087 7510 4121
rect 7464 4049 7510 4087
rect 7464 4015 7470 4049
rect 7504 4015 7510 4049
rect 7464 3977 7510 4015
rect 7464 3943 7470 3977
rect 7504 3943 7510 3977
rect 7464 3928 7510 3943
rect 7560 4913 7606 4928
rect 7560 4879 7566 4913
rect 7600 4879 7606 4913
rect 7560 4841 7606 4879
rect 7560 4807 7566 4841
rect 7600 4807 7606 4841
rect 7560 4769 7606 4807
rect 7560 4735 7566 4769
rect 7600 4735 7606 4769
rect 7560 4697 7606 4735
rect 7560 4663 7566 4697
rect 7600 4663 7606 4697
rect 7560 4625 7606 4663
rect 7560 4591 7566 4625
rect 7600 4591 7606 4625
rect 7560 4553 7606 4591
rect 7560 4519 7566 4553
rect 7600 4519 7606 4553
rect 7560 4481 7606 4519
rect 7560 4447 7566 4481
rect 7600 4447 7606 4481
rect 7560 4409 7606 4447
rect 7560 4375 7566 4409
rect 7600 4375 7606 4409
rect 7560 4337 7606 4375
rect 7560 4303 7566 4337
rect 7600 4303 7606 4337
rect 7560 4265 7606 4303
rect 7560 4231 7566 4265
rect 7600 4231 7606 4265
rect 7560 4193 7606 4231
rect 7560 4159 7566 4193
rect 7600 4159 7606 4193
rect 7560 4121 7606 4159
rect 7560 4087 7566 4121
rect 7600 4087 7606 4121
rect 7560 4049 7606 4087
rect 7560 4015 7566 4049
rect 7600 4015 7606 4049
rect 7560 3977 7606 4015
rect 7560 3943 7566 3977
rect 7600 3943 7606 3977
rect 7560 3928 7606 3943
rect 7656 4913 7702 4928
rect 7656 4879 7662 4913
rect 7696 4879 7702 4913
rect 7656 4841 7702 4879
rect 7656 4807 7662 4841
rect 7696 4807 7702 4841
rect 7656 4769 7702 4807
rect 7656 4735 7662 4769
rect 7696 4735 7702 4769
rect 7656 4697 7702 4735
rect 7656 4663 7662 4697
rect 7696 4663 7702 4697
rect 7656 4625 7702 4663
rect 7656 4591 7662 4625
rect 7696 4591 7702 4625
rect 7656 4553 7702 4591
rect 7656 4519 7662 4553
rect 7696 4519 7702 4553
rect 7656 4481 7702 4519
rect 7656 4447 7662 4481
rect 7696 4447 7702 4481
rect 7656 4409 7702 4447
rect 7656 4375 7662 4409
rect 7696 4375 7702 4409
rect 7656 4337 7702 4375
rect 7656 4303 7662 4337
rect 7696 4303 7702 4337
rect 7656 4265 7702 4303
rect 7656 4231 7662 4265
rect 7696 4231 7702 4265
rect 7656 4193 7702 4231
rect 7656 4159 7662 4193
rect 7696 4159 7702 4193
rect 7656 4121 7702 4159
rect 7656 4087 7662 4121
rect 7696 4087 7702 4121
rect 7656 4049 7702 4087
rect 7656 4015 7662 4049
rect 7696 4015 7702 4049
rect 7656 3977 7702 4015
rect 7656 3943 7662 3977
rect 7696 3943 7702 3977
rect 7656 3928 7702 3943
rect 7752 4913 7798 4928
rect 7752 4879 7758 4913
rect 7792 4879 7798 4913
rect 7752 4841 7798 4879
rect 7752 4807 7758 4841
rect 7792 4807 7798 4841
rect 7752 4769 7798 4807
rect 7752 4735 7758 4769
rect 7792 4735 7798 4769
rect 7752 4697 7798 4735
rect 7752 4663 7758 4697
rect 7792 4663 7798 4697
rect 7752 4625 7798 4663
rect 7752 4591 7758 4625
rect 7792 4591 7798 4625
rect 7752 4553 7798 4591
rect 7752 4519 7758 4553
rect 7792 4519 7798 4553
rect 7752 4481 7798 4519
rect 7752 4447 7758 4481
rect 7792 4447 7798 4481
rect 7752 4409 7798 4447
rect 7752 4375 7758 4409
rect 7792 4375 7798 4409
rect 7752 4337 7798 4375
rect 7752 4303 7758 4337
rect 7792 4303 7798 4337
rect 7752 4265 7798 4303
rect 7752 4231 7758 4265
rect 7792 4231 7798 4265
rect 7752 4193 7798 4231
rect 7752 4159 7758 4193
rect 7792 4159 7798 4193
rect 7752 4121 7798 4159
rect 7752 4087 7758 4121
rect 7792 4087 7798 4121
rect 7752 4049 7798 4087
rect 7752 4015 7758 4049
rect 7792 4015 7798 4049
rect 7752 3977 7798 4015
rect 7752 3943 7758 3977
rect 7792 3943 7798 3977
rect 7752 3928 7798 3943
rect 7848 4913 7894 4928
rect 7848 4879 7854 4913
rect 7888 4879 7894 4913
rect 7848 4841 7894 4879
rect 7848 4807 7854 4841
rect 7888 4807 7894 4841
rect 7848 4769 7894 4807
rect 7848 4735 7854 4769
rect 7888 4735 7894 4769
rect 7848 4697 7894 4735
rect 7848 4663 7854 4697
rect 7888 4663 7894 4697
rect 7848 4625 7894 4663
rect 7848 4591 7854 4625
rect 7888 4591 7894 4625
rect 7848 4553 7894 4591
rect 7848 4519 7854 4553
rect 7888 4519 7894 4553
rect 7848 4481 7894 4519
rect 7848 4447 7854 4481
rect 7888 4447 7894 4481
rect 7848 4409 7894 4447
rect 7848 4375 7854 4409
rect 7888 4375 7894 4409
rect 7848 4337 7894 4375
rect 7848 4303 7854 4337
rect 7888 4303 7894 4337
rect 7848 4265 7894 4303
rect 7848 4231 7854 4265
rect 7888 4231 7894 4265
rect 7848 4193 7894 4231
rect 7848 4159 7854 4193
rect 7888 4159 7894 4193
rect 7848 4121 7894 4159
rect 7848 4087 7854 4121
rect 7888 4087 7894 4121
rect 7848 4049 7894 4087
rect 7848 4015 7854 4049
rect 7888 4015 7894 4049
rect 7848 3977 7894 4015
rect 7848 3943 7854 3977
rect 7888 3943 7894 3977
rect 7848 3928 7894 3943
rect 10552 4911 10598 4926
rect 10552 4877 10558 4911
rect 10592 4877 10598 4911
rect 10552 4839 10598 4877
rect 10552 4805 10558 4839
rect 10592 4805 10598 4839
rect 10552 4767 10598 4805
rect 10552 4733 10558 4767
rect 10592 4733 10598 4767
rect 10552 4695 10598 4733
rect 10552 4661 10558 4695
rect 10592 4661 10598 4695
rect 10552 4623 10598 4661
rect 10552 4589 10558 4623
rect 10592 4589 10598 4623
rect 10552 4551 10598 4589
rect 10552 4517 10558 4551
rect 10592 4517 10598 4551
rect 10552 4479 10598 4517
rect 10552 4445 10558 4479
rect 10592 4445 10598 4479
rect 10552 4407 10598 4445
rect 10552 4373 10558 4407
rect 10592 4373 10598 4407
rect 10552 4335 10598 4373
rect 10552 4301 10558 4335
rect 10592 4301 10598 4335
rect 10552 4263 10598 4301
rect 10552 4229 10558 4263
rect 10592 4229 10598 4263
rect 10552 4191 10598 4229
rect 10552 4157 10558 4191
rect 10592 4157 10598 4191
rect 10552 4119 10598 4157
rect 10552 4085 10558 4119
rect 10592 4085 10598 4119
rect 10552 4047 10598 4085
rect 10552 4013 10558 4047
rect 10592 4013 10598 4047
rect 10552 3975 10598 4013
rect 10552 3941 10558 3975
rect 10592 3941 10598 3975
rect 10552 3926 10598 3941
rect 10648 4911 10694 4926
rect 10648 4877 10654 4911
rect 10688 4877 10694 4911
rect 10648 4839 10694 4877
rect 10648 4805 10654 4839
rect 10688 4805 10694 4839
rect 10648 4767 10694 4805
rect 10648 4733 10654 4767
rect 10688 4733 10694 4767
rect 10648 4695 10694 4733
rect 10648 4661 10654 4695
rect 10688 4661 10694 4695
rect 10648 4623 10694 4661
rect 10648 4589 10654 4623
rect 10688 4589 10694 4623
rect 10648 4551 10694 4589
rect 10648 4517 10654 4551
rect 10688 4517 10694 4551
rect 10648 4479 10694 4517
rect 10648 4445 10654 4479
rect 10688 4445 10694 4479
rect 10648 4407 10694 4445
rect 10648 4373 10654 4407
rect 10688 4373 10694 4407
rect 10648 4335 10694 4373
rect 10648 4301 10654 4335
rect 10688 4301 10694 4335
rect 10648 4263 10694 4301
rect 10648 4229 10654 4263
rect 10688 4229 10694 4263
rect 10648 4191 10694 4229
rect 10648 4157 10654 4191
rect 10688 4157 10694 4191
rect 10648 4119 10694 4157
rect 10648 4085 10654 4119
rect 10688 4085 10694 4119
rect 10648 4047 10694 4085
rect 10648 4013 10654 4047
rect 10688 4013 10694 4047
rect 10648 3975 10694 4013
rect 10648 3941 10654 3975
rect 10688 3941 10694 3975
rect 10648 3926 10694 3941
rect 10744 4911 10790 4926
rect 10744 4877 10750 4911
rect 10784 4877 10790 4911
rect 10744 4839 10790 4877
rect 10744 4805 10750 4839
rect 10784 4805 10790 4839
rect 10744 4767 10790 4805
rect 10744 4733 10750 4767
rect 10784 4733 10790 4767
rect 10744 4695 10790 4733
rect 10744 4661 10750 4695
rect 10784 4661 10790 4695
rect 10744 4623 10790 4661
rect 10744 4589 10750 4623
rect 10784 4589 10790 4623
rect 10744 4551 10790 4589
rect 10744 4517 10750 4551
rect 10784 4517 10790 4551
rect 10744 4479 10790 4517
rect 10744 4445 10750 4479
rect 10784 4445 10790 4479
rect 10744 4407 10790 4445
rect 10744 4373 10750 4407
rect 10784 4373 10790 4407
rect 10744 4335 10790 4373
rect 10744 4301 10750 4335
rect 10784 4301 10790 4335
rect 10744 4263 10790 4301
rect 10744 4229 10750 4263
rect 10784 4229 10790 4263
rect 10744 4191 10790 4229
rect 10744 4157 10750 4191
rect 10784 4157 10790 4191
rect 10744 4119 10790 4157
rect 10744 4085 10750 4119
rect 10784 4085 10790 4119
rect 10744 4047 10790 4085
rect 10744 4013 10750 4047
rect 10784 4013 10790 4047
rect 10744 3975 10790 4013
rect 10744 3941 10750 3975
rect 10784 3941 10790 3975
rect 10744 3926 10790 3941
rect 10840 4911 10886 4926
rect 10840 4877 10846 4911
rect 10880 4877 10886 4911
rect 10840 4839 10886 4877
rect 10840 4805 10846 4839
rect 10880 4805 10886 4839
rect 10840 4767 10886 4805
rect 10840 4733 10846 4767
rect 10880 4733 10886 4767
rect 10840 4695 10886 4733
rect 10840 4661 10846 4695
rect 10880 4661 10886 4695
rect 10840 4623 10886 4661
rect 10840 4589 10846 4623
rect 10880 4589 10886 4623
rect 10840 4551 10886 4589
rect 10840 4517 10846 4551
rect 10880 4517 10886 4551
rect 10840 4479 10886 4517
rect 10840 4445 10846 4479
rect 10880 4445 10886 4479
rect 10840 4407 10886 4445
rect 10840 4373 10846 4407
rect 10880 4373 10886 4407
rect 10840 4335 10886 4373
rect 10840 4301 10846 4335
rect 10880 4301 10886 4335
rect 10840 4263 10886 4301
rect 10840 4229 10846 4263
rect 10880 4229 10886 4263
rect 10840 4191 10886 4229
rect 10840 4157 10846 4191
rect 10880 4157 10886 4191
rect 10840 4119 10886 4157
rect 10840 4085 10846 4119
rect 10880 4085 10886 4119
rect 10840 4047 10886 4085
rect 10840 4013 10846 4047
rect 10880 4013 10886 4047
rect 10840 3975 10886 4013
rect 10840 3941 10846 3975
rect 10880 3941 10886 3975
rect 10840 3926 10886 3941
rect 10936 4911 10982 4926
rect 10936 4877 10942 4911
rect 10976 4877 10982 4911
rect 15512 4909 15518 4943
rect 15552 4909 15558 4943
rect 10936 4839 10982 4877
rect 10936 4805 10942 4839
rect 10976 4805 10982 4839
rect 10936 4767 10982 4805
rect 10936 4733 10942 4767
rect 10976 4733 10982 4767
rect 10936 4695 10982 4733
rect 10936 4661 10942 4695
rect 10976 4661 10982 4695
rect 10936 4623 10982 4661
rect 10936 4589 10942 4623
rect 10976 4589 10982 4623
rect 10936 4551 10982 4589
rect 10936 4517 10942 4551
rect 10976 4517 10982 4551
rect 10936 4479 10982 4517
rect 10936 4445 10942 4479
rect 10976 4445 10982 4479
rect 10936 4407 10982 4445
rect 10936 4373 10942 4407
rect 10976 4373 10982 4407
rect 10936 4335 10982 4373
rect 10936 4301 10942 4335
rect 10976 4301 10982 4335
rect 10936 4263 10982 4301
rect 10936 4229 10942 4263
rect 10976 4229 10982 4263
rect 10936 4191 10982 4229
rect 10936 4157 10942 4191
rect 10976 4157 10982 4191
rect 10936 4119 10982 4157
rect 10936 4085 10942 4119
rect 10976 4085 10982 4119
rect 10936 4047 10982 4085
rect 10936 4013 10942 4047
rect 10976 4013 10982 4047
rect 10936 3975 10982 4013
rect 10936 3941 10942 3975
rect 10976 3941 10982 3975
rect 10936 3926 10982 3941
rect 13708 4885 13754 4900
rect 13708 4851 13714 4885
rect 13748 4851 13754 4885
rect 13708 4813 13754 4851
rect 13708 4779 13714 4813
rect 13748 4779 13754 4813
rect 13708 4741 13754 4779
rect 13708 4707 13714 4741
rect 13748 4707 13754 4741
rect 13708 4669 13754 4707
rect 13708 4635 13714 4669
rect 13748 4635 13754 4669
rect 13708 4597 13754 4635
rect 13708 4563 13714 4597
rect 13748 4563 13754 4597
rect 13708 4525 13754 4563
rect 13708 4491 13714 4525
rect 13748 4491 13754 4525
rect 13708 4453 13754 4491
rect 13708 4419 13714 4453
rect 13748 4419 13754 4453
rect 13708 4381 13754 4419
rect 13708 4347 13714 4381
rect 13748 4347 13754 4381
rect 13708 4309 13754 4347
rect 13708 4275 13714 4309
rect 13748 4275 13754 4309
rect 13708 4237 13754 4275
rect 13708 4203 13714 4237
rect 13748 4203 13754 4237
rect 13708 4165 13754 4203
rect 13708 4131 13714 4165
rect 13748 4131 13754 4165
rect 13708 4093 13754 4131
rect 13708 4059 13714 4093
rect 13748 4059 13754 4093
rect 13708 4021 13754 4059
rect 13708 3987 13714 4021
rect 13748 3987 13754 4021
rect 13708 3949 13754 3987
rect 13708 3915 13714 3949
rect 13748 3915 13754 3949
rect 13708 3900 13754 3915
rect 13804 4885 13850 4900
rect 13804 4851 13810 4885
rect 13844 4851 13850 4885
rect 13804 4813 13850 4851
rect 13804 4779 13810 4813
rect 13844 4779 13850 4813
rect 13804 4741 13850 4779
rect 13804 4707 13810 4741
rect 13844 4707 13850 4741
rect 13804 4669 13850 4707
rect 13804 4635 13810 4669
rect 13844 4635 13850 4669
rect 13804 4597 13850 4635
rect 13804 4563 13810 4597
rect 13844 4563 13850 4597
rect 13804 4525 13850 4563
rect 13804 4491 13810 4525
rect 13844 4491 13850 4525
rect 13804 4453 13850 4491
rect 13804 4419 13810 4453
rect 13844 4419 13850 4453
rect 13804 4381 13850 4419
rect 13804 4347 13810 4381
rect 13844 4347 13850 4381
rect 13804 4309 13850 4347
rect 13804 4275 13810 4309
rect 13844 4275 13850 4309
rect 13804 4237 13850 4275
rect 13804 4203 13810 4237
rect 13844 4203 13850 4237
rect 13804 4165 13850 4203
rect 13804 4131 13810 4165
rect 13844 4131 13850 4165
rect 13804 4093 13850 4131
rect 13804 4059 13810 4093
rect 13844 4059 13850 4093
rect 13804 4021 13850 4059
rect 13804 3987 13810 4021
rect 13844 3987 13850 4021
rect 13804 3949 13850 3987
rect 13804 3915 13810 3949
rect 13844 3915 13850 3949
rect 13804 3900 13850 3915
rect 13900 4885 13946 4900
rect 13900 4851 13906 4885
rect 13940 4851 13946 4885
rect 13900 4813 13946 4851
rect 13900 4779 13906 4813
rect 13940 4779 13946 4813
rect 13900 4741 13946 4779
rect 13900 4707 13906 4741
rect 13940 4707 13946 4741
rect 13900 4669 13946 4707
rect 13900 4635 13906 4669
rect 13940 4635 13946 4669
rect 13900 4597 13946 4635
rect 13900 4563 13906 4597
rect 13940 4563 13946 4597
rect 13900 4525 13946 4563
rect 13900 4491 13906 4525
rect 13940 4491 13946 4525
rect 13900 4453 13946 4491
rect 13900 4419 13906 4453
rect 13940 4419 13946 4453
rect 13900 4381 13946 4419
rect 13900 4347 13906 4381
rect 13940 4347 13946 4381
rect 13900 4309 13946 4347
rect 13900 4275 13906 4309
rect 13940 4275 13946 4309
rect 13900 4237 13946 4275
rect 13900 4203 13906 4237
rect 13940 4203 13946 4237
rect 13900 4165 13946 4203
rect 13900 4131 13906 4165
rect 13940 4131 13946 4165
rect 13900 4093 13946 4131
rect 13900 4059 13906 4093
rect 13940 4059 13946 4093
rect 13900 4021 13946 4059
rect 13900 3987 13906 4021
rect 13940 3987 13946 4021
rect 13900 3949 13946 3987
rect 13900 3915 13906 3949
rect 13940 3915 13946 3949
rect 13900 3900 13946 3915
rect 13996 4885 14042 4900
rect 13996 4851 14002 4885
rect 14036 4851 14042 4885
rect 13996 4813 14042 4851
rect 13996 4779 14002 4813
rect 14036 4779 14042 4813
rect 13996 4741 14042 4779
rect 13996 4707 14002 4741
rect 14036 4707 14042 4741
rect 13996 4669 14042 4707
rect 13996 4635 14002 4669
rect 14036 4635 14042 4669
rect 13996 4597 14042 4635
rect 13996 4563 14002 4597
rect 14036 4563 14042 4597
rect 13996 4525 14042 4563
rect 13996 4491 14002 4525
rect 14036 4491 14042 4525
rect 13996 4453 14042 4491
rect 13996 4419 14002 4453
rect 14036 4419 14042 4453
rect 13996 4381 14042 4419
rect 13996 4347 14002 4381
rect 14036 4347 14042 4381
rect 13996 4309 14042 4347
rect 13996 4275 14002 4309
rect 14036 4275 14042 4309
rect 13996 4237 14042 4275
rect 13996 4203 14002 4237
rect 14036 4203 14042 4237
rect 13996 4165 14042 4203
rect 13996 4131 14002 4165
rect 14036 4131 14042 4165
rect 13996 4093 14042 4131
rect 13996 4059 14002 4093
rect 14036 4059 14042 4093
rect 13996 4021 14042 4059
rect 13996 3987 14002 4021
rect 14036 3987 14042 4021
rect 13996 3949 14042 3987
rect 13996 3915 14002 3949
rect 14036 3915 14042 3949
rect 13996 3900 14042 3915
rect 14092 4885 14138 4900
rect 14092 4851 14098 4885
rect 14132 4851 14138 4885
rect 14092 4813 14138 4851
rect 14092 4779 14098 4813
rect 14132 4779 14138 4813
rect 14092 4741 14138 4779
rect 14092 4707 14098 4741
rect 14132 4707 14138 4741
rect 14092 4669 14138 4707
rect 14092 4635 14098 4669
rect 14132 4635 14138 4669
rect 14092 4597 14138 4635
rect 14092 4563 14098 4597
rect 14132 4563 14138 4597
rect 14092 4525 14138 4563
rect 14092 4491 14098 4525
rect 14132 4491 14138 4525
rect 14092 4453 14138 4491
rect 14092 4419 14098 4453
rect 14132 4419 14138 4453
rect 14092 4381 14138 4419
rect 14092 4347 14098 4381
rect 14132 4347 14138 4381
rect 14092 4309 14138 4347
rect 14092 4275 14098 4309
rect 14132 4275 14138 4309
rect 14092 4237 14138 4275
rect 14092 4203 14098 4237
rect 14132 4203 14138 4237
rect 14092 4165 14138 4203
rect 14092 4131 14098 4165
rect 14132 4131 14138 4165
rect 14092 4093 14138 4131
rect 14092 4059 14098 4093
rect 14132 4059 14138 4093
rect 14092 4021 14138 4059
rect 14092 3987 14098 4021
rect 14132 3987 14138 4021
rect 14092 3949 14138 3987
rect 14092 3915 14098 3949
rect 14132 3915 14138 3949
rect 15512 4871 15558 4909
rect 15512 4837 15518 4871
rect 15552 4837 15558 4871
rect 15512 4799 15558 4837
rect 15512 4765 15518 4799
rect 15552 4765 15558 4799
rect 15512 4727 15558 4765
rect 15512 4693 15518 4727
rect 15552 4693 15558 4727
rect 15512 4655 15558 4693
rect 15512 4621 15518 4655
rect 15552 4621 15558 4655
rect 15512 4583 15558 4621
rect 15512 4549 15518 4583
rect 15552 4549 15558 4583
rect 15512 4511 15558 4549
rect 15512 4477 15518 4511
rect 15552 4477 15558 4511
rect 15512 4439 15558 4477
rect 15512 4405 15518 4439
rect 15552 4405 15558 4439
rect 15512 4367 15558 4405
rect 15512 4333 15518 4367
rect 15552 4333 15558 4367
rect 15512 4295 15558 4333
rect 15512 4261 15518 4295
rect 15552 4261 15558 4295
rect 15512 4223 15558 4261
rect 15512 4189 15518 4223
rect 15552 4189 15558 4223
rect 15512 4151 15558 4189
rect 15512 4117 15518 4151
rect 15552 4117 15558 4151
rect 15512 4079 15558 4117
rect 15512 4045 15518 4079
rect 15552 4045 15558 4079
rect 15512 4007 15558 4045
rect 15512 3973 15518 4007
rect 15552 3973 15558 4007
rect 15512 3926 15558 3973
rect 15608 5879 15654 5926
rect 15608 5845 15614 5879
rect 15648 5845 15654 5879
rect 15608 5807 15654 5845
rect 15608 5773 15614 5807
rect 15648 5773 15654 5807
rect 15608 5735 15654 5773
rect 15608 5701 15614 5735
rect 15648 5701 15654 5735
rect 15608 5663 15654 5701
rect 15608 5629 15614 5663
rect 15648 5629 15654 5663
rect 15608 5591 15654 5629
rect 15608 5557 15614 5591
rect 15648 5557 15654 5591
rect 15608 5519 15654 5557
rect 15608 5485 15614 5519
rect 15648 5485 15654 5519
rect 15608 5447 15654 5485
rect 15608 5413 15614 5447
rect 15648 5413 15654 5447
rect 15608 5375 15654 5413
rect 15608 5341 15614 5375
rect 15648 5341 15654 5375
rect 15608 5303 15654 5341
rect 15608 5269 15614 5303
rect 15648 5269 15654 5303
rect 15608 5231 15654 5269
rect 15608 5197 15614 5231
rect 15648 5197 15654 5231
rect 15608 5159 15654 5197
rect 15608 5125 15614 5159
rect 15648 5125 15654 5159
rect 15608 5087 15654 5125
rect 15608 5053 15614 5087
rect 15648 5053 15654 5087
rect 15608 5015 15654 5053
rect 15608 4981 15614 5015
rect 15648 4981 15654 5015
rect 15608 4943 15654 4981
rect 15608 4909 15614 4943
rect 15648 4909 15654 4943
rect 15608 4871 15654 4909
rect 15608 4837 15614 4871
rect 15648 4837 15654 4871
rect 15608 4799 15654 4837
rect 15608 4765 15614 4799
rect 15648 4765 15654 4799
rect 15608 4727 15654 4765
rect 15608 4693 15614 4727
rect 15648 4693 15654 4727
rect 15608 4655 15654 4693
rect 15608 4621 15614 4655
rect 15648 4621 15654 4655
rect 15608 4583 15654 4621
rect 15608 4549 15614 4583
rect 15648 4549 15654 4583
rect 15608 4511 15654 4549
rect 15608 4477 15614 4511
rect 15648 4477 15654 4511
rect 15608 4439 15654 4477
rect 15608 4405 15614 4439
rect 15648 4405 15654 4439
rect 15608 4367 15654 4405
rect 15608 4333 15614 4367
rect 15648 4333 15654 4367
rect 15608 4295 15654 4333
rect 15608 4261 15614 4295
rect 15648 4261 15654 4295
rect 15608 4223 15654 4261
rect 15608 4189 15614 4223
rect 15648 4189 15654 4223
rect 15608 4151 15654 4189
rect 15608 4117 15614 4151
rect 15648 4117 15654 4151
rect 15608 4079 15654 4117
rect 15608 4045 15614 4079
rect 15648 4045 15654 4079
rect 15608 4007 15654 4045
rect 15608 3973 15614 4007
rect 15648 3973 15654 4007
rect 15608 3926 15654 3973
rect 15704 5879 15750 5926
rect 15704 5845 15710 5879
rect 15744 5845 15750 5879
rect 15704 5807 15750 5845
rect 15704 5773 15710 5807
rect 15744 5773 15750 5807
rect 15704 5735 15750 5773
rect 15704 5701 15710 5735
rect 15744 5701 15750 5735
rect 15704 5663 15750 5701
rect 15704 5629 15710 5663
rect 15744 5629 15750 5663
rect 15704 5591 15750 5629
rect 15704 5557 15710 5591
rect 15744 5557 15750 5591
rect 15704 5519 15750 5557
rect 15704 5485 15710 5519
rect 15744 5485 15750 5519
rect 15704 5447 15750 5485
rect 15704 5413 15710 5447
rect 15744 5413 15750 5447
rect 15704 5375 15750 5413
rect 15704 5341 15710 5375
rect 15744 5341 15750 5375
rect 15704 5303 15750 5341
rect 15704 5269 15710 5303
rect 15744 5269 15750 5303
rect 15704 5231 15750 5269
rect 15704 5197 15710 5231
rect 15744 5197 15750 5231
rect 15704 5159 15750 5197
rect 15704 5125 15710 5159
rect 15744 5125 15750 5159
rect 15704 5087 15750 5125
rect 15704 5053 15710 5087
rect 15744 5053 15750 5087
rect 15704 5015 15750 5053
rect 15704 4981 15710 5015
rect 15744 4981 15750 5015
rect 15704 4943 15750 4981
rect 15704 4909 15710 4943
rect 15744 4909 15750 4943
rect 15704 4871 15750 4909
rect 15704 4837 15710 4871
rect 15744 4837 15750 4871
rect 15704 4799 15750 4837
rect 15704 4765 15710 4799
rect 15744 4765 15750 4799
rect 15704 4727 15750 4765
rect 15704 4693 15710 4727
rect 15744 4693 15750 4727
rect 15704 4655 15750 4693
rect 15704 4621 15710 4655
rect 15744 4621 15750 4655
rect 15704 4583 15750 4621
rect 15704 4549 15710 4583
rect 15744 4549 15750 4583
rect 15704 4511 15750 4549
rect 15704 4477 15710 4511
rect 15744 4477 15750 4511
rect 15704 4439 15750 4477
rect 15704 4405 15710 4439
rect 15744 4405 15750 4439
rect 15704 4367 15750 4405
rect 15704 4333 15710 4367
rect 15744 4333 15750 4367
rect 15704 4295 15750 4333
rect 15704 4261 15710 4295
rect 15744 4261 15750 4295
rect 15704 4223 15750 4261
rect 15704 4189 15710 4223
rect 15744 4189 15750 4223
rect 15704 4151 15750 4189
rect 15704 4117 15710 4151
rect 15744 4117 15750 4151
rect 15704 4079 15750 4117
rect 15704 4045 15710 4079
rect 15744 4045 15750 4079
rect 15704 4007 15750 4045
rect 15704 3973 15710 4007
rect 15744 3973 15750 4007
rect 15704 3926 15750 3973
rect 14092 3900 14138 3915
rect 15332 3794 15394 3798
rect 1842 3790 2168 3792
rect 1566 3783 1624 3788
rect 1760 3787 2168 3790
rect 1566 3777 1626 3783
rect 1566 3743 1580 3777
rect 1614 3743 1626 3777
rect 1760 3777 2101 3787
rect 1566 3737 1626 3743
rect 1662 3754 1724 3770
rect 1566 3730 1624 3737
rect -1126 3290 -1110 3324
rect -1076 3290 -1020 3324
rect -1126 3276 -1020 3290
rect 1662 3720 1676 3754
rect 1710 3720 1724 3754
rect 1760 3743 1772 3777
rect 1806 3743 2101 3777
rect 1760 3735 2101 3743
rect 2153 3735 2168 3787
rect 11054 3774 11064 3780
rect 1760 3732 2168 3735
rect 1842 3730 2168 3732
rect 4522 3767 4580 3772
rect 4714 3769 5000 3774
rect 4522 3761 4582 3767
rect -1692 3221 -1646 3236
rect -1692 3187 -1686 3221
rect -1652 3187 -1646 3221
rect -1692 3149 -1646 3187
rect -1692 3115 -1686 3149
rect -1652 3115 -1646 3149
rect -1692 3077 -1646 3115
rect -1692 3043 -1686 3077
rect -1652 3043 -1646 3077
rect -1692 3005 -1646 3043
rect -1692 2971 -1686 3005
rect -1652 2971 -1646 3005
rect -1692 2933 -1646 2971
rect -1692 2899 -1686 2933
rect -1652 2899 -1646 2933
rect -1692 2861 -1646 2899
rect -1692 2827 -1686 2861
rect -1652 2827 -1646 2861
rect -1692 2789 -1646 2827
rect -1692 2755 -1686 2789
rect -1652 2755 -1646 2789
rect -1692 2717 -1646 2755
rect -1692 2683 -1686 2717
rect -1652 2683 -1646 2717
rect -1692 2645 -1646 2683
rect -1692 2611 -1686 2645
rect -1652 2611 -1646 2645
rect -1692 2573 -1646 2611
rect -1692 2539 -1686 2573
rect -1652 2539 -1646 2573
rect -1692 2501 -1646 2539
rect -1692 2467 -1686 2501
rect -1652 2467 -1646 2501
rect -1692 2429 -1646 2467
rect -1692 2395 -1686 2429
rect -1652 2395 -1646 2429
rect -1692 2357 -1646 2395
rect -1692 2323 -1686 2357
rect -1652 2323 -1646 2357
rect -1692 2285 -1646 2323
rect -1692 2251 -1686 2285
rect -1652 2251 -1646 2285
rect -1692 2236 -1646 2251
rect -1596 3221 -1550 3236
rect -1596 3187 -1590 3221
rect -1556 3187 -1550 3221
rect -1596 3149 -1550 3187
rect -1596 3115 -1590 3149
rect -1556 3115 -1550 3149
rect -1596 3077 -1550 3115
rect -1596 3043 -1590 3077
rect -1556 3043 -1550 3077
rect -1596 3005 -1550 3043
rect -1596 2971 -1590 3005
rect -1556 2971 -1550 3005
rect -1596 2933 -1550 2971
rect -1596 2899 -1590 2933
rect -1556 2899 -1550 2933
rect -1596 2861 -1550 2899
rect -1596 2827 -1590 2861
rect -1556 2827 -1550 2861
rect -1596 2789 -1550 2827
rect -1596 2755 -1590 2789
rect -1556 2755 -1550 2789
rect -1596 2717 -1550 2755
rect -1596 2683 -1590 2717
rect -1556 2683 -1550 2717
rect -1596 2645 -1550 2683
rect -1596 2611 -1590 2645
rect -1556 2611 -1550 2645
rect -1596 2573 -1550 2611
rect -1596 2539 -1590 2573
rect -1556 2539 -1550 2573
rect -1596 2501 -1550 2539
rect -1596 2467 -1590 2501
rect -1556 2467 -1550 2501
rect -1596 2429 -1550 2467
rect -1596 2395 -1590 2429
rect -1556 2395 -1550 2429
rect -1596 2357 -1550 2395
rect -1596 2323 -1590 2357
rect -1556 2323 -1550 2357
rect -1596 2285 -1550 2323
rect -1596 2251 -1590 2285
rect -1556 2251 -1550 2285
rect -1596 2236 -1550 2251
rect -1500 3221 -1454 3236
rect -1500 3187 -1494 3221
rect -1460 3187 -1454 3221
rect -1500 3149 -1454 3187
rect -1500 3115 -1494 3149
rect -1460 3115 -1454 3149
rect -1500 3077 -1454 3115
rect -1500 3043 -1494 3077
rect -1460 3043 -1454 3077
rect -1500 3005 -1454 3043
rect -1500 2971 -1494 3005
rect -1460 2971 -1454 3005
rect -1500 2933 -1454 2971
rect -1500 2899 -1494 2933
rect -1460 2899 -1454 2933
rect -1500 2861 -1454 2899
rect -1500 2827 -1494 2861
rect -1460 2827 -1454 2861
rect -1500 2789 -1454 2827
rect -1500 2755 -1494 2789
rect -1460 2755 -1454 2789
rect -1500 2717 -1454 2755
rect -1500 2683 -1494 2717
rect -1460 2683 -1454 2717
rect -1500 2645 -1454 2683
rect -1500 2611 -1494 2645
rect -1460 2611 -1454 2645
rect -1500 2573 -1454 2611
rect -1500 2539 -1494 2573
rect -1460 2539 -1454 2573
rect -1500 2501 -1454 2539
rect -1500 2467 -1494 2501
rect -1460 2467 -1454 2501
rect -1500 2429 -1454 2467
rect -1500 2395 -1494 2429
rect -1460 2395 -1454 2429
rect -1500 2357 -1454 2395
rect -1500 2323 -1494 2357
rect -1460 2323 -1454 2357
rect -1500 2285 -1454 2323
rect -1500 2251 -1494 2285
rect -1460 2251 -1454 2285
rect -1500 2236 -1454 2251
rect -1404 3221 -1358 3236
rect -1404 3187 -1398 3221
rect -1364 3187 -1358 3221
rect -1404 3149 -1358 3187
rect -1404 3115 -1398 3149
rect -1364 3115 -1358 3149
rect -1404 3077 -1358 3115
rect -1404 3043 -1398 3077
rect -1364 3043 -1358 3077
rect -1404 3005 -1358 3043
rect -1404 2971 -1398 3005
rect -1364 2971 -1358 3005
rect -1404 2933 -1358 2971
rect -1404 2899 -1398 2933
rect -1364 2899 -1358 2933
rect -1404 2861 -1358 2899
rect -1404 2827 -1398 2861
rect -1364 2827 -1358 2861
rect -1404 2789 -1358 2827
rect -1404 2755 -1398 2789
rect -1364 2755 -1358 2789
rect -1404 2717 -1358 2755
rect -1404 2683 -1398 2717
rect -1364 2683 -1358 2717
rect -1404 2645 -1358 2683
rect -1404 2611 -1398 2645
rect -1364 2611 -1358 2645
rect -1404 2573 -1358 2611
rect -1404 2539 -1398 2573
rect -1364 2539 -1358 2573
rect -1404 2501 -1358 2539
rect -1404 2467 -1398 2501
rect -1364 2467 -1358 2501
rect -1404 2429 -1358 2467
rect -1404 2395 -1398 2429
rect -1364 2395 -1358 2429
rect -1404 2357 -1358 2395
rect -1404 2323 -1398 2357
rect -1364 2323 -1358 2357
rect -1404 2285 -1358 2323
rect -1404 2251 -1398 2285
rect -1364 2251 -1358 2285
rect -1404 2236 -1358 2251
rect -1308 3221 -1262 3236
rect -1308 3187 -1302 3221
rect -1268 3187 -1262 3221
rect -1308 3149 -1262 3187
rect -1308 3115 -1302 3149
rect -1268 3115 -1262 3149
rect -1308 3077 -1262 3115
rect -1308 3043 -1302 3077
rect -1268 3043 -1262 3077
rect -1308 3005 -1262 3043
rect -1308 2971 -1302 3005
rect -1268 2971 -1262 3005
rect -1308 2933 -1262 2971
rect -1308 2899 -1302 2933
rect -1268 2899 -1262 2933
rect -1308 2861 -1262 2899
rect -1308 2827 -1302 2861
rect -1268 2827 -1262 2861
rect -1308 2789 -1262 2827
rect -1308 2755 -1302 2789
rect -1268 2755 -1262 2789
rect -1308 2717 -1262 2755
rect -1308 2683 -1302 2717
rect -1268 2683 -1262 2717
rect -1308 2645 -1262 2683
rect -1308 2611 -1302 2645
rect -1268 2611 -1262 2645
rect -1308 2573 -1262 2611
rect -1308 2539 -1302 2573
rect -1268 2539 -1262 2573
rect -1308 2501 -1262 2539
rect -1308 2467 -1302 2501
rect -1268 2467 -1262 2501
rect -1308 2429 -1262 2467
rect -1308 2395 -1302 2429
rect -1268 2395 -1262 2429
rect -1308 2357 -1262 2395
rect -1308 2323 -1302 2357
rect -1268 2323 -1262 2357
rect -1308 2285 -1262 2323
rect -1308 2251 -1302 2285
rect -1268 2251 -1262 2285
rect -1308 2236 -1262 2251
rect -1212 3221 -1166 3236
rect -1212 3187 -1206 3221
rect -1172 3187 -1166 3221
rect -1212 3149 -1166 3187
rect -1212 3115 -1206 3149
rect -1172 3115 -1166 3149
rect -1212 3077 -1166 3115
rect -1212 3043 -1206 3077
rect -1172 3043 -1166 3077
rect -1212 3005 -1166 3043
rect -1212 2971 -1206 3005
rect -1172 2971 -1166 3005
rect -1212 2933 -1166 2971
rect -1212 2899 -1206 2933
rect -1172 2899 -1166 2933
rect -1212 2861 -1166 2899
rect -1212 2827 -1206 2861
rect -1172 2827 -1166 2861
rect -1212 2789 -1166 2827
rect -1212 2755 -1206 2789
rect -1172 2755 -1166 2789
rect -1212 2717 -1166 2755
rect -1212 2683 -1206 2717
rect -1172 2683 -1166 2717
rect -1212 2645 -1166 2683
rect -1212 2611 -1206 2645
rect -1172 2611 -1166 2645
rect -1212 2573 -1166 2611
rect -1212 2539 -1206 2573
rect -1172 2539 -1166 2573
rect -1212 2501 -1166 2539
rect -1212 2467 -1206 2501
rect -1172 2467 -1166 2501
rect -1212 2429 -1166 2467
rect -1212 2395 -1206 2429
rect -1172 2395 -1166 2429
rect -1212 2357 -1166 2395
rect -1212 2323 -1206 2357
rect -1172 2323 -1166 2357
rect -1212 2285 -1166 2323
rect -1212 2251 -1206 2285
rect -1172 2251 -1166 2285
rect -1212 2236 -1166 2251
rect -1116 3221 -1070 3236
rect -1116 3187 -1110 3221
rect -1076 3187 -1070 3221
rect -1116 3149 -1070 3187
rect -1116 3115 -1110 3149
rect -1076 3115 -1070 3149
rect -1116 3077 -1070 3115
rect -1116 3043 -1110 3077
rect -1076 3043 -1070 3077
rect -1116 3005 -1070 3043
rect -1116 2971 -1110 3005
rect -1076 2971 -1070 3005
rect -1116 2933 -1070 2971
rect -1116 2899 -1110 2933
rect -1076 2899 -1070 2933
rect -1116 2861 -1070 2899
rect -1116 2827 -1110 2861
rect -1076 2827 -1070 2861
rect -1116 2789 -1070 2827
rect -1116 2755 -1110 2789
rect -1076 2755 -1070 2789
rect -1116 2717 -1070 2755
rect -1116 2683 -1110 2717
rect -1076 2683 -1070 2717
rect -1116 2645 -1070 2683
rect -1116 2611 -1110 2645
rect -1076 2611 -1070 2645
rect -1116 2573 -1070 2611
rect -1116 2539 -1110 2573
rect -1076 2539 -1070 2573
rect -1116 2501 -1070 2539
rect -1116 2467 -1110 2501
rect -1076 2467 -1070 2501
rect -1116 2429 -1070 2467
rect -1116 2395 -1110 2429
rect -1076 2395 -1070 2429
rect -1116 2357 -1070 2395
rect -1116 2323 -1110 2357
rect -1076 2323 -1070 2357
rect -1116 2285 -1070 2323
rect -1116 2251 -1110 2285
rect -1076 2251 -1070 2285
rect -1116 2236 -1070 2251
rect -1020 3221 -974 3236
rect -1020 3187 -1014 3221
rect -980 3187 -974 3221
rect -1020 3149 -974 3187
rect -1020 3115 -1014 3149
rect -980 3115 -974 3149
rect -1020 3077 -974 3115
rect -1020 3043 -1014 3077
rect -980 3043 -974 3077
rect -1020 3005 -974 3043
rect -1020 2971 -1014 3005
rect -980 2971 -974 3005
rect -1020 2933 -974 2971
rect -1020 2899 -1014 2933
rect -980 2899 -974 2933
rect -1020 2861 -974 2899
rect -1020 2827 -1014 2861
rect -980 2827 -974 2861
rect -1020 2789 -974 2827
rect -1020 2755 -1014 2789
rect -980 2755 -974 2789
rect -1020 2717 -974 2755
rect -1020 2683 -1014 2717
rect -980 2683 -974 2717
rect -1020 2645 -974 2683
rect -1020 2611 -1014 2645
rect -980 2611 -974 2645
rect -1020 2573 -974 2611
rect -1020 2539 -1014 2573
rect -980 2539 -974 2573
rect -1020 2501 -974 2539
rect -1020 2467 -1014 2501
rect -980 2467 -974 2501
rect -1020 2429 -974 2467
rect -1020 2395 -1014 2429
rect -980 2395 -974 2429
rect -1020 2357 -974 2395
rect -1020 2323 -1014 2357
rect -980 2323 -974 2357
rect -1020 2285 -974 2323
rect -1020 2251 -1014 2285
rect -980 2251 -974 2285
rect -1020 2236 -974 2251
rect -924 3221 -878 3236
rect -924 3187 -918 3221
rect -884 3187 -878 3221
rect -924 3149 -878 3187
rect -924 3115 -918 3149
rect -884 3115 -878 3149
rect -924 3077 -878 3115
rect -924 3043 -918 3077
rect -884 3043 -878 3077
rect -924 3005 -878 3043
rect 1662 3086 1724 3720
rect 4522 3727 4536 3761
rect 4570 3727 4582 3761
rect 4714 3761 4933 3769
rect 4522 3721 4582 3727
rect 4618 3738 4680 3754
rect 4522 3714 4580 3721
rect 4618 3704 4632 3738
rect 4666 3704 4680 3738
rect 4714 3727 4728 3761
rect 4762 3727 4933 3761
rect 4714 3717 4933 3727
rect 4985 3717 5000 3769
rect 4714 3712 5000 3717
rect 5598 3761 7614 3774
rect 5598 3727 7566 3761
rect 7600 3727 7614 3761
rect 7744 3761 8364 3774
rect 5598 3712 7614 3727
rect 7648 3738 7710 3754
rect 3658 3305 3720 3320
rect 3658 3253 3663 3305
rect 3715 3253 3720 3305
rect 3658 3086 3720 3253
rect 1662 3024 4244 3086
rect -924 2971 -918 3005
rect -884 2971 -878 3005
rect -924 2933 -878 2971
rect 1394 3013 1626 3018
rect 1394 2961 1409 3013
rect 1461 3002 1626 3013
rect 1461 2968 1578 3002
rect 1612 2968 1626 3002
rect 1461 2961 1626 2968
rect 1394 2956 1626 2961
rect 1662 2994 1724 3024
rect 1662 2960 1674 2994
rect 1708 2960 1724 2994
rect 1662 2948 1724 2960
rect -924 2899 -918 2933
rect -884 2899 -878 2933
rect -924 2861 -878 2899
rect -924 2827 -918 2861
rect -884 2827 -878 2861
rect -924 2789 -878 2827
rect -924 2755 -918 2789
rect -884 2755 -878 2789
rect -924 2717 -878 2755
rect -924 2683 -918 2717
rect -884 2683 -878 2717
rect -924 2645 -878 2683
rect -924 2611 -918 2645
rect -884 2611 -878 2645
rect -924 2573 -878 2611
rect -924 2539 -918 2573
rect -884 2539 -878 2573
rect -924 2501 -878 2539
rect -924 2467 -918 2501
rect -884 2467 -878 2501
rect -924 2429 -878 2467
rect -924 2395 -918 2429
rect -884 2395 -878 2429
rect -924 2357 -878 2395
rect -924 2323 -918 2357
rect -884 2323 -878 2357
rect -924 2285 -878 2323
rect -924 2251 -918 2285
rect -884 2251 -878 2285
rect -924 2236 -878 2251
rect 1476 2815 1522 2830
rect 1476 2781 1482 2815
rect 1516 2781 1522 2815
rect 1476 2743 1522 2781
rect 1476 2709 1482 2743
rect 1516 2709 1522 2743
rect 1476 2671 1522 2709
rect 1476 2637 1482 2671
rect 1516 2637 1522 2671
rect 1476 2599 1522 2637
rect 1476 2565 1482 2599
rect 1516 2565 1522 2599
rect 1476 2527 1522 2565
rect 1476 2493 1482 2527
rect 1516 2493 1522 2527
rect 1476 2455 1522 2493
rect 1476 2421 1482 2455
rect 1516 2421 1522 2455
rect 1476 2383 1522 2421
rect 1476 2349 1482 2383
rect 1516 2349 1522 2383
rect 1476 2311 1522 2349
rect 1476 2277 1482 2311
rect 1516 2277 1522 2311
rect 1476 2239 1522 2277
rect 1476 2205 1482 2239
rect 1516 2205 1522 2239
rect -1110 2172 -1048 2190
rect -1110 2138 -1097 2172
rect -1063 2138 -1048 2172
rect -1110 1298 -1048 2138
rect 1476 2167 1522 2205
rect 1476 2133 1482 2167
rect 1516 2133 1522 2167
rect 1476 2095 1522 2133
rect 1476 2061 1482 2095
rect 1516 2061 1522 2095
rect 1476 2023 1522 2061
rect 1476 1989 1482 2023
rect 1516 1989 1522 2023
rect 1476 1951 1522 1989
rect 1476 1917 1482 1951
rect 1516 1917 1522 1951
rect 1476 1879 1522 1917
rect 1476 1845 1482 1879
rect 1516 1845 1522 1879
rect 1476 1830 1522 1845
rect 1572 2815 1618 2830
rect 1572 2781 1578 2815
rect 1612 2781 1618 2815
rect 1572 2743 1618 2781
rect 1572 2709 1578 2743
rect 1612 2709 1618 2743
rect 1572 2671 1618 2709
rect 1572 2637 1578 2671
rect 1612 2637 1618 2671
rect 1572 2599 1618 2637
rect 1572 2565 1578 2599
rect 1612 2565 1618 2599
rect 1572 2527 1618 2565
rect 1572 2493 1578 2527
rect 1612 2493 1618 2527
rect 1572 2455 1618 2493
rect 1572 2421 1578 2455
rect 1612 2421 1618 2455
rect 1572 2383 1618 2421
rect 1572 2349 1578 2383
rect 1612 2349 1618 2383
rect 1572 2311 1618 2349
rect 1572 2277 1578 2311
rect 1612 2277 1618 2311
rect 1572 2239 1618 2277
rect 1572 2205 1578 2239
rect 1612 2205 1618 2239
rect 1572 2167 1618 2205
rect 1572 2133 1578 2167
rect 1612 2133 1618 2167
rect 1572 2095 1618 2133
rect 1572 2061 1578 2095
rect 1612 2061 1618 2095
rect 1572 2023 1618 2061
rect 1572 1989 1578 2023
rect 1612 1989 1618 2023
rect 1572 1951 1618 1989
rect 1572 1917 1578 1951
rect 1612 1917 1618 1951
rect 1572 1879 1618 1917
rect 1572 1845 1578 1879
rect 1612 1845 1618 1879
rect 1572 1830 1618 1845
rect 1668 2815 1714 2830
rect 1668 2781 1674 2815
rect 1708 2781 1714 2815
rect 1668 2743 1714 2781
rect 1668 2709 1674 2743
rect 1708 2709 1714 2743
rect 1668 2671 1714 2709
rect 1668 2637 1674 2671
rect 1708 2637 1714 2671
rect 1668 2599 1714 2637
rect 1668 2565 1674 2599
rect 1708 2565 1714 2599
rect 1668 2527 1714 2565
rect 1668 2493 1674 2527
rect 1708 2493 1714 2527
rect 1668 2455 1714 2493
rect 1668 2421 1674 2455
rect 1708 2421 1714 2455
rect 1668 2383 1714 2421
rect 1668 2349 1674 2383
rect 1708 2349 1714 2383
rect 1668 2311 1714 2349
rect 1668 2277 1674 2311
rect 1708 2277 1714 2311
rect 1668 2239 1714 2277
rect 1668 2205 1674 2239
rect 1708 2205 1714 2239
rect 1668 2167 1714 2205
rect 1668 2133 1674 2167
rect 1708 2133 1714 2167
rect 1668 2095 1714 2133
rect 1668 2061 1674 2095
rect 1708 2061 1714 2095
rect 1668 2023 1714 2061
rect 1668 1989 1674 2023
rect 1708 1989 1714 2023
rect 1668 1951 1714 1989
rect 1668 1917 1674 1951
rect 1708 1917 1714 1951
rect 1668 1879 1714 1917
rect 1668 1845 1674 1879
rect 1708 1845 1714 1879
rect 1668 1830 1714 1845
rect 1764 2815 1810 2830
rect 1764 2781 1770 2815
rect 1804 2781 1810 2815
rect 1764 2743 1810 2781
rect 1764 2709 1770 2743
rect 1804 2709 1810 2743
rect 1764 2671 1810 2709
rect 1764 2637 1770 2671
rect 1804 2637 1810 2671
rect 1764 2599 1810 2637
rect 1764 2565 1770 2599
rect 1804 2565 1810 2599
rect 1764 2527 1810 2565
rect 1764 2493 1770 2527
rect 1804 2493 1810 2527
rect 1764 2455 1810 2493
rect 1764 2421 1770 2455
rect 1804 2421 1810 2455
rect 1764 2383 1810 2421
rect 1764 2349 1770 2383
rect 1804 2349 1810 2383
rect 1764 2311 1810 2349
rect 1764 2277 1770 2311
rect 1804 2277 1810 2311
rect 1764 2239 1810 2277
rect 1764 2205 1770 2239
rect 1804 2205 1810 2239
rect 1764 2167 1810 2205
rect 1764 2133 1770 2167
rect 1804 2133 1810 2167
rect 1764 2095 1810 2133
rect 1764 2061 1770 2095
rect 1804 2061 1810 2095
rect 1764 2023 1810 2061
rect 1764 1989 1770 2023
rect 1804 1989 1810 2023
rect 1764 1951 1810 1989
rect 1764 1917 1770 1951
rect 1804 1917 1810 1951
rect 1764 1879 1810 1917
rect 1764 1845 1770 1879
rect 1804 1845 1810 1879
rect 1764 1830 1810 1845
rect 1860 2815 1906 2830
rect 1860 2781 1866 2815
rect 1900 2781 1906 2815
rect 1860 2743 1906 2781
rect 1860 2709 1866 2743
rect 1900 2709 1906 2743
rect 1860 2671 1906 2709
rect 1860 2637 1866 2671
rect 1900 2637 1906 2671
rect 1860 2599 1906 2637
rect 1860 2565 1866 2599
rect 1900 2565 1906 2599
rect 1860 2527 1906 2565
rect 1860 2493 1866 2527
rect 1900 2493 1906 2527
rect 1860 2455 1906 2493
rect 1860 2421 1866 2455
rect 1900 2421 1906 2455
rect 1860 2383 1906 2421
rect 1860 2349 1866 2383
rect 1900 2349 1906 2383
rect 1860 2311 1906 2349
rect 1860 2277 1866 2311
rect 1900 2277 1906 2311
rect 2232 2360 2294 3024
rect 4182 3000 4244 3024
rect 4618 3068 4680 3704
rect 5600 3215 5662 3712
rect 7648 3704 7662 3738
rect 7696 3704 7710 3738
rect 7744 3727 7758 3761
rect 7792 3727 8364 3761
rect 7744 3712 8364 3727
rect 10008 3767 10698 3772
rect 10008 3715 10023 3767
rect 10075 3765 10698 3767
rect 10075 3759 10700 3765
rect 10075 3725 10654 3759
rect 10688 3725 10700 3759
rect 10830 3759 11064 3774
rect 10075 3719 10700 3725
rect 10736 3736 10798 3752
rect 10075 3715 10698 3719
rect 7648 3532 7710 3704
rect 7122 3479 7710 3532
rect 7122 3427 7127 3479
rect 7179 3470 7710 3479
rect 7179 3427 7184 3470
rect 7122 3412 7184 3427
rect 5600 3163 5605 3215
rect 5657 3163 5662 3215
rect 5600 3148 5662 3163
rect 7284 3158 7346 3170
rect 7276 3092 7286 3158
rect 7374 3092 7384 3158
rect 4618 3006 7200 3068
rect 4182 2992 4560 3000
rect 4182 2986 4580 2992
rect 4182 2952 4534 2986
rect 4568 2952 4580 2986
rect 4182 2946 4580 2952
rect 4618 2978 4680 3006
rect 4182 2938 4560 2946
rect 4618 2944 4630 2978
rect 4664 2944 4680 2978
rect 4618 2932 4680 2944
rect 4432 2799 4478 2814
rect 4432 2765 4438 2799
rect 4472 2765 4478 2799
rect 4432 2727 4478 2765
rect 4432 2693 4438 2727
rect 4472 2693 4478 2727
rect 4432 2655 4478 2693
rect 2550 2592 2642 2622
rect 2550 2540 2570 2592
rect 2622 2540 2642 2592
rect 2550 2428 2642 2540
rect 2550 2394 2579 2428
rect 2613 2394 2642 2428
rect 2550 2388 2642 2394
rect 4432 2621 4438 2655
rect 4472 2621 4478 2655
rect 4432 2583 4478 2621
rect 4432 2549 4438 2583
rect 4472 2549 4478 2583
rect 4432 2511 4478 2549
rect 4432 2477 4438 2511
rect 4472 2477 4478 2511
rect 4432 2439 4478 2477
rect 4432 2405 4438 2439
rect 4472 2405 4478 2439
rect 4432 2367 4478 2405
rect 2232 2350 2438 2360
rect 2232 2316 2392 2350
rect 2426 2316 2438 2350
rect 2232 2298 2438 2316
rect 4432 2333 4438 2367
rect 4472 2333 4478 2367
rect 1860 2239 1906 2277
rect 4432 2295 4478 2333
rect 1860 2205 1866 2239
rect 1900 2205 1906 2239
rect 1860 2167 1906 2205
rect 1860 2133 1866 2167
rect 1900 2133 1906 2167
rect 1860 2095 1906 2133
rect 1860 2061 1866 2095
rect 1900 2061 1906 2095
rect 2494 2229 2540 2276
rect 2494 2195 2500 2229
rect 2534 2195 2540 2229
rect 2494 2157 2540 2195
rect 2494 2123 2500 2157
rect 2534 2123 2540 2157
rect 2494 2076 2540 2123
rect 2652 2229 2698 2276
rect 2652 2195 2658 2229
rect 2692 2195 2698 2229
rect 2652 2157 2698 2195
rect 2652 2123 2658 2157
rect 2692 2123 2698 2157
rect 2652 2076 2698 2123
rect 4432 2261 4438 2295
rect 4472 2261 4478 2295
rect 4432 2223 4478 2261
rect 4432 2189 4438 2223
rect 4472 2189 4478 2223
rect 4432 2151 4478 2189
rect 4432 2117 4438 2151
rect 4472 2117 4478 2151
rect 4432 2079 4478 2117
rect 1860 2023 1906 2061
rect 1860 1989 1866 2023
rect 1900 1989 1906 2023
rect 1860 1951 1906 1989
rect 1860 1917 1866 1951
rect 1900 1917 1906 1951
rect 1860 1879 1906 1917
rect 1860 1845 1866 1879
rect 1900 1845 1906 1879
rect 1860 1830 1906 1845
rect 4432 2045 4438 2079
rect 4472 2045 4478 2079
rect 4432 2007 4478 2045
rect 4432 1973 4438 2007
rect 4472 1973 4478 2007
rect 4432 1935 4478 1973
rect 4432 1901 4438 1935
rect 4472 1901 4478 1935
rect 4432 1863 4478 1901
rect 4432 1829 4438 1863
rect 4472 1829 4478 1863
rect 4432 1814 4478 1829
rect 4528 2799 4574 2814
rect 4528 2765 4534 2799
rect 4568 2765 4574 2799
rect 4528 2727 4574 2765
rect 4528 2693 4534 2727
rect 4568 2693 4574 2727
rect 4528 2655 4574 2693
rect 4528 2621 4534 2655
rect 4568 2621 4574 2655
rect 4528 2583 4574 2621
rect 4528 2549 4534 2583
rect 4568 2549 4574 2583
rect 4528 2511 4574 2549
rect 4528 2477 4534 2511
rect 4568 2477 4574 2511
rect 4528 2439 4574 2477
rect 4528 2405 4534 2439
rect 4568 2405 4574 2439
rect 4528 2367 4574 2405
rect 4528 2333 4534 2367
rect 4568 2333 4574 2367
rect 4528 2295 4574 2333
rect 4528 2261 4534 2295
rect 4568 2261 4574 2295
rect 4528 2223 4574 2261
rect 4528 2189 4534 2223
rect 4568 2189 4574 2223
rect 4528 2151 4574 2189
rect 4528 2117 4534 2151
rect 4568 2117 4574 2151
rect 4528 2079 4574 2117
rect 4528 2045 4534 2079
rect 4568 2045 4574 2079
rect 4528 2007 4574 2045
rect 4528 1973 4534 2007
rect 4568 1973 4574 2007
rect 4528 1935 4574 1973
rect 4528 1901 4534 1935
rect 4568 1901 4574 1935
rect 4528 1863 4574 1901
rect 4528 1829 4534 1863
rect 4568 1829 4574 1863
rect 4528 1814 4574 1829
rect 4624 2799 4670 2814
rect 4624 2765 4630 2799
rect 4664 2765 4670 2799
rect 4624 2727 4670 2765
rect 4624 2693 4630 2727
rect 4664 2693 4670 2727
rect 4624 2655 4670 2693
rect 4624 2621 4630 2655
rect 4664 2621 4670 2655
rect 4624 2583 4670 2621
rect 4624 2549 4630 2583
rect 4664 2549 4670 2583
rect 4624 2511 4670 2549
rect 4624 2477 4630 2511
rect 4664 2477 4670 2511
rect 4624 2439 4670 2477
rect 4624 2405 4630 2439
rect 4664 2405 4670 2439
rect 4624 2367 4670 2405
rect 4624 2333 4630 2367
rect 4664 2333 4670 2367
rect 4624 2295 4670 2333
rect 4624 2261 4630 2295
rect 4664 2261 4670 2295
rect 4624 2223 4670 2261
rect 4624 2189 4630 2223
rect 4664 2189 4670 2223
rect 4624 2151 4670 2189
rect 4624 2117 4630 2151
rect 4664 2117 4670 2151
rect 4624 2079 4670 2117
rect 4624 2045 4630 2079
rect 4664 2045 4670 2079
rect 4624 2007 4670 2045
rect 4624 1973 4630 2007
rect 4664 1973 4670 2007
rect 4624 1935 4670 1973
rect 4624 1901 4630 1935
rect 4664 1901 4670 1935
rect 4624 1863 4670 1901
rect 4624 1829 4630 1863
rect 4664 1829 4670 1863
rect 4624 1814 4670 1829
rect 4720 2799 4766 2814
rect 4720 2765 4726 2799
rect 4760 2765 4766 2799
rect 4720 2727 4766 2765
rect 4720 2693 4726 2727
rect 4760 2693 4766 2727
rect 4720 2655 4766 2693
rect 4720 2621 4726 2655
rect 4760 2621 4766 2655
rect 4720 2583 4766 2621
rect 4720 2549 4726 2583
rect 4760 2549 4766 2583
rect 4720 2511 4766 2549
rect 4720 2477 4726 2511
rect 4760 2477 4766 2511
rect 4720 2439 4766 2477
rect 4720 2405 4726 2439
rect 4760 2405 4766 2439
rect 4720 2367 4766 2405
rect 4720 2333 4726 2367
rect 4760 2333 4766 2367
rect 4720 2295 4766 2333
rect 4720 2261 4726 2295
rect 4760 2261 4766 2295
rect 4720 2223 4766 2261
rect 4720 2189 4726 2223
rect 4760 2189 4766 2223
rect 4720 2151 4766 2189
rect 4720 2117 4726 2151
rect 4760 2117 4766 2151
rect 4720 2079 4766 2117
rect 4720 2045 4726 2079
rect 4760 2045 4766 2079
rect 4720 2007 4766 2045
rect 4720 1973 4726 2007
rect 4760 1973 4766 2007
rect 4720 1935 4766 1973
rect 4720 1901 4726 1935
rect 4760 1901 4766 1935
rect 4720 1863 4766 1901
rect 4720 1829 4726 1863
rect 4760 1829 4766 1863
rect 4720 1814 4766 1829
rect 4816 2799 4862 2814
rect 4816 2765 4822 2799
rect 4856 2765 4862 2799
rect 4816 2727 4862 2765
rect 4816 2693 4822 2727
rect 4856 2693 4862 2727
rect 4816 2655 4862 2693
rect 4816 2621 4822 2655
rect 4856 2621 4862 2655
rect 4816 2583 4862 2621
rect 4816 2549 4822 2583
rect 4856 2549 4862 2583
rect 4816 2511 4862 2549
rect 4816 2477 4822 2511
rect 4856 2477 4862 2511
rect 4816 2439 4862 2477
rect 4816 2405 4822 2439
rect 4856 2405 4862 2439
rect 4816 2367 4862 2405
rect 4816 2333 4822 2367
rect 4856 2333 4862 2367
rect 4816 2295 4862 2333
rect 5132 2360 5194 3006
rect 7138 3000 7200 3006
rect 7284 3000 7346 3092
rect 7648 3048 7710 3470
rect 8298 3408 8360 3712
rect 10008 3710 10698 3715
rect 10736 3702 10750 3736
rect 10784 3702 10798 3736
rect 10830 3725 10846 3759
rect 10880 3725 11064 3759
rect 10830 3710 11064 3725
rect 11054 3706 11064 3710
rect 11150 3706 11160 3780
rect 13560 3739 13854 3748
rect 13560 3733 13856 3739
rect 8672 3592 8682 3676
rect 8752 3652 8762 3676
rect 10736 3652 10798 3702
rect 8752 3596 10798 3652
rect 8752 3592 8762 3596
rect 10404 3471 10466 3486
rect 10404 3419 10409 3471
rect 10461 3419 10466 3471
rect 10404 3408 10466 3419
rect 8298 3352 8746 3408
rect 8850 3352 10466 3408
rect 8298 3350 10466 3352
rect 8298 3346 10464 3350
rect 7138 2992 7608 3000
rect 7648 2998 10260 3048
rect 10736 3046 10798 3596
rect 13560 3699 13810 3733
rect 13844 3699 13856 3733
rect 13988 3733 14642 3750
rect 13560 3693 13856 3699
rect 13892 3710 13954 3726
rect 13560 3684 13854 3693
rect 13076 3471 13138 3486
rect 13560 3474 13628 3684
rect 13076 3419 13081 3471
rect 13133 3419 13138 3471
rect 13076 3300 13138 3419
rect 13426 3464 13628 3474
rect 13426 3412 13436 3464
rect 13498 3412 13628 3464
rect 13426 3410 13628 3412
rect 13892 3676 13906 3710
rect 13940 3676 13954 3710
rect 13988 3699 14002 3733
rect 14036 3699 14642 3733
rect 15326 3732 15336 3794
rect 15398 3779 15614 3794
rect 15398 3745 15566 3779
rect 15600 3745 15614 3779
rect 15398 3732 15614 3745
rect 15698 3760 15760 3772
rect 13988 3684 14642 3699
rect 13892 3300 13954 3676
rect 13076 3238 13954 3300
rect 13892 3174 13954 3238
rect 13892 3112 14296 3174
rect 7138 2986 7610 2992
rect 7138 2952 7564 2986
rect 7598 2952 7610 2986
rect 7138 2946 7610 2952
rect 7648 2986 10698 2998
rect 7648 2978 7710 2986
rect 7138 2938 7608 2946
rect 7648 2944 7660 2978
rect 7694 2944 7710 2978
rect 7648 2932 7710 2944
rect 7462 2799 7508 2814
rect 7462 2765 7468 2799
rect 7502 2765 7508 2799
rect 7462 2727 7508 2765
rect 7462 2693 7468 2727
rect 7502 2693 7508 2727
rect 7462 2655 7508 2693
rect 5550 2592 5642 2622
rect 5550 2540 5570 2592
rect 5622 2540 5642 2592
rect 5550 2428 5642 2540
rect 5550 2394 5579 2428
rect 5613 2394 5642 2428
rect 5550 2388 5642 2394
rect 7462 2621 7468 2655
rect 7502 2621 7508 2655
rect 7462 2583 7508 2621
rect 7462 2549 7468 2583
rect 7502 2549 7508 2583
rect 7462 2511 7508 2549
rect 7462 2477 7468 2511
rect 7502 2477 7508 2511
rect 7462 2439 7508 2477
rect 7462 2405 7468 2439
rect 7502 2405 7508 2439
rect 7462 2367 7508 2405
rect 5132 2350 5438 2360
rect 5132 2316 5392 2350
rect 5426 2316 5438 2350
rect 5132 2298 5438 2316
rect 7462 2333 7468 2367
rect 7502 2333 7508 2367
rect 4816 2261 4822 2295
rect 4856 2261 4862 2295
rect 7462 2295 7508 2333
rect 4816 2223 4862 2261
rect 4816 2189 4822 2223
rect 4856 2189 4862 2223
rect 4816 2151 4862 2189
rect 4816 2117 4822 2151
rect 4856 2117 4862 2151
rect 4816 2079 4862 2117
rect 4816 2045 4822 2079
rect 4856 2045 4862 2079
rect 5494 2229 5540 2276
rect 5494 2195 5500 2229
rect 5534 2195 5540 2229
rect 5494 2157 5540 2195
rect 5494 2123 5500 2157
rect 5534 2123 5540 2157
rect 5494 2076 5540 2123
rect 5652 2229 5698 2276
rect 5652 2195 5658 2229
rect 5692 2195 5698 2229
rect 5652 2157 5698 2195
rect 5652 2123 5658 2157
rect 5692 2123 5698 2157
rect 5652 2076 5698 2123
rect 7462 2261 7468 2295
rect 7502 2261 7508 2295
rect 7462 2223 7508 2261
rect 7462 2189 7468 2223
rect 7502 2189 7508 2223
rect 7462 2151 7508 2189
rect 7462 2117 7468 2151
rect 7502 2117 7508 2151
rect 7462 2079 7508 2117
rect 4816 2007 4862 2045
rect 4816 1973 4822 2007
rect 4856 1973 4862 2007
rect 4816 1935 4862 1973
rect 4816 1901 4822 1935
rect 4856 1901 4862 1935
rect 4816 1863 4862 1901
rect 4816 1829 4822 1863
rect 4856 1829 4862 1863
rect 4816 1814 4862 1829
rect 7462 2045 7468 2079
rect 7502 2045 7508 2079
rect 7462 2007 7508 2045
rect 7462 1973 7468 2007
rect 7502 1973 7508 2007
rect 7462 1935 7508 1973
rect 7462 1901 7468 1935
rect 7502 1901 7508 1935
rect 7462 1863 7508 1901
rect 7462 1829 7468 1863
rect 7502 1829 7508 1863
rect 7462 1814 7508 1829
rect 7558 2799 7604 2814
rect 7558 2765 7564 2799
rect 7598 2765 7604 2799
rect 7558 2727 7604 2765
rect 7558 2693 7564 2727
rect 7598 2693 7604 2727
rect 7558 2655 7604 2693
rect 7558 2621 7564 2655
rect 7598 2621 7604 2655
rect 7558 2583 7604 2621
rect 7558 2549 7564 2583
rect 7598 2549 7604 2583
rect 7558 2511 7604 2549
rect 7558 2477 7564 2511
rect 7598 2477 7604 2511
rect 7558 2439 7604 2477
rect 7558 2405 7564 2439
rect 7598 2405 7604 2439
rect 7558 2367 7604 2405
rect 7558 2333 7564 2367
rect 7598 2333 7604 2367
rect 7558 2295 7604 2333
rect 7558 2261 7564 2295
rect 7598 2261 7604 2295
rect 7558 2223 7604 2261
rect 7558 2189 7564 2223
rect 7598 2189 7604 2223
rect 7558 2151 7604 2189
rect 7558 2117 7564 2151
rect 7598 2117 7604 2151
rect 7558 2079 7604 2117
rect 7558 2045 7564 2079
rect 7598 2045 7604 2079
rect 7558 2007 7604 2045
rect 7558 1973 7564 2007
rect 7598 1973 7604 2007
rect 7558 1935 7604 1973
rect 7558 1901 7564 1935
rect 7598 1901 7604 1935
rect 7558 1863 7604 1901
rect 7558 1829 7564 1863
rect 7598 1829 7604 1863
rect 7558 1814 7604 1829
rect 7654 2799 7700 2814
rect 7654 2765 7660 2799
rect 7694 2765 7700 2799
rect 7654 2727 7700 2765
rect 7654 2693 7660 2727
rect 7694 2693 7700 2727
rect 7654 2655 7700 2693
rect 7654 2621 7660 2655
rect 7694 2621 7700 2655
rect 7654 2583 7700 2621
rect 7654 2549 7660 2583
rect 7694 2549 7700 2583
rect 7654 2511 7700 2549
rect 7654 2477 7660 2511
rect 7694 2477 7700 2511
rect 7654 2439 7700 2477
rect 7654 2405 7660 2439
rect 7694 2405 7700 2439
rect 7654 2367 7700 2405
rect 7654 2333 7660 2367
rect 7694 2333 7700 2367
rect 7654 2295 7700 2333
rect 7654 2261 7660 2295
rect 7694 2261 7700 2295
rect 7654 2223 7700 2261
rect 7654 2189 7660 2223
rect 7694 2189 7700 2223
rect 7654 2151 7700 2189
rect 7654 2117 7660 2151
rect 7694 2117 7700 2151
rect 7654 2079 7700 2117
rect 7654 2045 7660 2079
rect 7694 2045 7700 2079
rect 7654 2007 7700 2045
rect 7654 1973 7660 2007
rect 7694 1973 7700 2007
rect 7654 1935 7700 1973
rect 7654 1901 7660 1935
rect 7694 1901 7700 1935
rect 7654 1863 7700 1901
rect 7654 1829 7660 1863
rect 7694 1829 7700 1863
rect 7654 1814 7700 1829
rect 7750 2799 7796 2814
rect 7750 2765 7756 2799
rect 7790 2765 7796 2799
rect 7750 2727 7796 2765
rect 7750 2693 7756 2727
rect 7790 2693 7796 2727
rect 7750 2655 7796 2693
rect 7750 2621 7756 2655
rect 7790 2621 7796 2655
rect 7750 2583 7796 2621
rect 7750 2549 7756 2583
rect 7790 2549 7796 2583
rect 7750 2511 7796 2549
rect 7750 2477 7756 2511
rect 7790 2477 7796 2511
rect 7750 2439 7796 2477
rect 7750 2405 7756 2439
rect 7790 2405 7796 2439
rect 7750 2367 7796 2405
rect 7750 2333 7756 2367
rect 7790 2333 7796 2367
rect 7750 2295 7796 2333
rect 7750 2261 7756 2295
rect 7790 2261 7796 2295
rect 7750 2223 7796 2261
rect 7750 2189 7756 2223
rect 7790 2189 7796 2223
rect 7750 2151 7796 2189
rect 7750 2117 7756 2151
rect 7790 2117 7796 2151
rect 7750 2079 7796 2117
rect 7750 2045 7756 2079
rect 7790 2045 7796 2079
rect 7750 2007 7796 2045
rect 7750 1973 7756 2007
rect 7790 1973 7796 2007
rect 7750 1935 7796 1973
rect 7750 1901 7756 1935
rect 7790 1901 7796 1935
rect 7750 1863 7796 1901
rect 7750 1829 7756 1863
rect 7790 1829 7796 1863
rect 7750 1814 7796 1829
rect 7846 2799 7892 2814
rect 7846 2765 7852 2799
rect 7886 2765 7892 2799
rect 7846 2727 7892 2765
rect 7846 2693 7852 2727
rect 7886 2693 7892 2727
rect 7846 2655 7892 2693
rect 7846 2621 7852 2655
rect 7886 2621 7892 2655
rect 7846 2583 7892 2621
rect 7846 2549 7852 2583
rect 7886 2549 7892 2583
rect 7846 2511 7892 2549
rect 7846 2477 7852 2511
rect 7886 2477 7892 2511
rect 7846 2439 7892 2477
rect 7846 2405 7852 2439
rect 7886 2405 7892 2439
rect 7846 2367 7892 2405
rect 7846 2333 7852 2367
rect 7886 2333 7892 2367
rect 7846 2295 7892 2333
rect 8232 2360 8294 2986
rect 10196 2984 10698 2986
rect 10196 2950 10652 2984
rect 10686 2950 10698 2984
rect 10196 2936 10698 2950
rect 10736 2984 13522 3046
rect 10736 2976 10798 2984
rect 10736 2942 10748 2976
rect 10782 2942 10798 2976
rect 10736 2930 10798 2942
rect 10550 2797 10596 2812
rect 10550 2763 10556 2797
rect 10590 2763 10596 2797
rect 10550 2725 10596 2763
rect 10550 2691 10556 2725
rect 10590 2691 10596 2725
rect 10550 2653 10596 2691
rect 8550 2597 8644 2628
rect 8550 2545 8571 2597
rect 8623 2545 8644 2597
rect 8550 2514 8644 2545
rect 10550 2619 10556 2653
rect 10590 2619 10596 2653
rect 10550 2581 10596 2619
rect 10550 2547 10556 2581
rect 10590 2547 10596 2581
rect 8550 2428 8642 2514
rect 8550 2394 8579 2428
rect 8613 2394 8642 2428
rect 8550 2388 8642 2394
rect 10550 2509 10596 2547
rect 10550 2475 10556 2509
rect 10590 2475 10596 2509
rect 10550 2437 10596 2475
rect 10550 2403 10556 2437
rect 10590 2403 10596 2437
rect 10550 2365 10596 2403
rect 8232 2350 8440 2360
rect 8232 2316 8392 2350
rect 8426 2316 8440 2350
rect 8232 2298 8440 2316
rect 10550 2331 10556 2365
rect 10590 2331 10596 2365
rect 7846 2261 7852 2295
rect 7886 2261 7892 2295
rect 10550 2293 10596 2331
rect 7846 2223 7892 2261
rect 7846 2189 7852 2223
rect 7886 2189 7892 2223
rect 7846 2151 7892 2189
rect 7846 2117 7852 2151
rect 7886 2117 7892 2151
rect 7846 2079 7892 2117
rect 7846 2045 7852 2079
rect 7886 2045 7892 2079
rect 8494 2229 8540 2276
rect 8494 2195 8500 2229
rect 8534 2195 8540 2229
rect 8494 2157 8540 2195
rect 8494 2123 8500 2157
rect 8534 2123 8540 2157
rect 8494 2076 8540 2123
rect 8652 2229 8698 2276
rect 8652 2195 8658 2229
rect 8692 2195 8698 2229
rect 8652 2157 8698 2195
rect 8652 2123 8658 2157
rect 8692 2123 8698 2157
rect 8652 2076 8698 2123
rect 10550 2259 10556 2293
rect 10590 2259 10596 2293
rect 10550 2221 10596 2259
rect 10550 2187 10556 2221
rect 10590 2187 10596 2221
rect 10550 2149 10596 2187
rect 10550 2115 10556 2149
rect 10590 2115 10596 2149
rect 10550 2077 10596 2115
rect 7846 2007 7892 2045
rect 7846 1973 7852 2007
rect 7886 1973 7892 2007
rect 7846 1935 7892 1973
rect 7846 1901 7852 1935
rect 7886 1901 7892 1935
rect 7846 1863 7892 1901
rect 7846 1829 7852 1863
rect 7886 1829 7892 1863
rect 7846 1814 7892 1829
rect 10550 2043 10556 2077
rect 10590 2043 10596 2077
rect 10550 2005 10596 2043
rect 10550 1971 10556 2005
rect 10590 1971 10596 2005
rect 10550 1933 10596 1971
rect 10550 1899 10556 1933
rect 10590 1899 10596 1933
rect 10550 1861 10596 1899
rect 10550 1827 10556 1861
rect 10590 1827 10596 1861
rect 10550 1812 10596 1827
rect 10646 2797 10692 2812
rect 10646 2763 10652 2797
rect 10686 2763 10692 2797
rect 10646 2725 10692 2763
rect 10646 2691 10652 2725
rect 10686 2691 10692 2725
rect 10646 2653 10692 2691
rect 10646 2619 10652 2653
rect 10686 2619 10692 2653
rect 10646 2581 10692 2619
rect 10646 2547 10652 2581
rect 10686 2547 10692 2581
rect 10646 2509 10692 2547
rect 10646 2475 10652 2509
rect 10686 2475 10692 2509
rect 10646 2437 10692 2475
rect 10646 2403 10652 2437
rect 10686 2403 10692 2437
rect 10646 2365 10692 2403
rect 10646 2331 10652 2365
rect 10686 2331 10692 2365
rect 10646 2293 10692 2331
rect 10646 2259 10652 2293
rect 10686 2259 10692 2293
rect 10646 2221 10692 2259
rect 10646 2187 10652 2221
rect 10686 2187 10692 2221
rect 10646 2149 10692 2187
rect 10646 2115 10652 2149
rect 10686 2115 10692 2149
rect 10646 2077 10692 2115
rect 10646 2043 10652 2077
rect 10686 2043 10692 2077
rect 10646 2005 10692 2043
rect 10646 1971 10652 2005
rect 10686 1971 10692 2005
rect 10646 1933 10692 1971
rect 10646 1899 10652 1933
rect 10686 1899 10692 1933
rect 10646 1861 10692 1899
rect 10646 1827 10652 1861
rect 10686 1827 10692 1861
rect 10646 1812 10692 1827
rect 10742 2797 10788 2812
rect 10742 2763 10748 2797
rect 10782 2763 10788 2797
rect 10742 2725 10788 2763
rect 10742 2691 10748 2725
rect 10782 2691 10788 2725
rect 10742 2653 10788 2691
rect 10742 2619 10748 2653
rect 10782 2619 10788 2653
rect 10742 2581 10788 2619
rect 10742 2547 10748 2581
rect 10782 2547 10788 2581
rect 10742 2509 10788 2547
rect 10742 2475 10748 2509
rect 10782 2475 10788 2509
rect 10742 2437 10788 2475
rect 10742 2403 10748 2437
rect 10782 2403 10788 2437
rect 10742 2365 10788 2403
rect 10742 2331 10748 2365
rect 10782 2331 10788 2365
rect 10742 2293 10788 2331
rect 10742 2259 10748 2293
rect 10782 2259 10788 2293
rect 10742 2221 10788 2259
rect 10742 2187 10748 2221
rect 10782 2187 10788 2221
rect 10742 2149 10788 2187
rect 10742 2115 10748 2149
rect 10782 2115 10788 2149
rect 10742 2077 10788 2115
rect 10742 2043 10748 2077
rect 10782 2043 10788 2077
rect 10742 2005 10788 2043
rect 10742 1971 10748 2005
rect 10782 1971 10788 2005
rect 10742 1933 10788 1971
rect 10742 1899 10748 1933
rect 10782 1899 10788 1933
rect 10742 1861 10788 1899
rect 10742 1827 10748 1861
rect 10782 1827 10788 1861
rect 10742 1812 10788 1827
rect 10838 2797 10884 2812
rect 10838 2763 10844 2797
rect 10878 2763 10884 2797
rect 10838 2725 10884 2763
rect 10838 2691 10844 2725
rect 10878 2691 10884 2725
rect 10838 2653 10884 2691
rect 10838 2619 10844 2653
rect 10878 2619 10884 2653
rect 10838 2581 10884 2619
rect 10838 2547 10844 2581
rect 10878 2547 10884 2581
rect 10838 2509 10884 2547
rect 10838 2475 10844 2509
rect 10878 2475 10884 2509
rect 10838 2437 10884 2475
rect 10838 2403 10844 2437
rect 10878 2403 10884 2437
rect 10838 2365 10884 2403
rect 10838 2331 10844 2365
rect 10878 2331 10884 2365
rect 10838 2293 10884 2331
rect 10838 2259 10844 2293
rect 10878 2259 10884 2293
rect 10838 2221 10884 2259
rect 10838 2187 10844 2221
rect 10878 2187 10884 2221
rect 10838 2149 10884 2187
rect 10838 2115 10844 2149
rect 10878 2115 10884 2149
rect 10838 2077 10884 2115
rect 10838 2043 10844 2077
rect 10878 2043 10884 2077
rect 10838 2005 10884 2043
rect 10838 1971 10844 2005
rect 10878 1971 10884 2005
rect 10838 1933 10884 1971
rect 10838 1899 10844 1933
rect 10878 1899 10884 1933
rect 10838 1861 10884 1899
rect 10838 1827 10844 1861
rect 10878 1827 10884 1861
rect 10838 1812 10884 1827
rect 10934 2797 10980 2812
rect 10934 2763 10940 2797
rect 10974 2763 10980 2797
rect 10934 2725 10980 2763
rect 10934 2691 10940 2725
rect 10974 2691 10980 2725
rect 10934 2653 10980 2691
rect 10934 2619 10940 2653
rect 10974 2619 10980 2653
rect 10934 2581 10980 2619
rect 10934 2547 10940 2581
rect 10974 2547 10980 2581
rect 10934 2509 10980 2547
rect 10934 2475 10940 2509
rect 10974 2475 10980 2509
rect 10934 2437 10980 2475
rect 10934 2403 10940 2437
rect 10974 2403 10980 2437
rect 10934 2365 10980 2403
rect 10934 2331 10940 2365
rect 10974 2331 10980 2365
rect 10934 2293 10980 2331
rect 11232 2360 11294 2984
rect 13460 2972 13522 2984
rect 13460 2958 13856 2972
rect 13460 2924 13808 2958
rect 13842 2924 13856 2958
rect 13460 2910 13856 2924
rect 13892 2950 13954 3112
rect 13892 2916 13904 2950
rect 13938 2916 13954 2950
rect 13892 2904 13954 2916
rect 13706 2771 13752 2786
rect 13706 2737 13712 2771
rect 13746 2737 13752 2771
rect 13706 2699 13752 2737
rect 13706 2665 13712 2699
rect 13746 2665 13752 2699
rect 13706 2627 13752 2665
rect 11550 2568 11642 2598
rect 11550 2516 11570 2568
rect 11622 2516 11642 2568
rect 11550 2428 11642 2516
rect 11550 2394 11579 2428
rect 11613 2394 11642 2428
rect 11550 2388 11642 2394
rect 13706 2593 13712 2627
rect 13746 2593 13752 2627
rect 13706 2555 13752 2593
rect 13706 2521 13712 2555
rect 13746 2521 13752 2555
rect 13706 2483 13752 2521
rect 13706 2449 13712 2483
rect 13746 2449 13752 2483
rect 13706 2411 13752 2449
rect 13706 2377 13712 2411
rect 13746 2377 13752 2411
rect 11232 2350 11440 2360
rect 11232 2316 11392 2350
rect 11426 2316 11440 2350
rect 11232 2298 11440 2316
rect 13706 2339 13752 2377
rect 13706 2305 13712 2339
rect 13746 2305 13752 2339
rect 10934 2259 10940 2293
rect 10974 2259 10980 2293
rect 10934 2221 10980 2259
rect 10934 2187 10940 2221
rect 10974 2187 10980 2221
rect 10934 2149 10980 2187
rect 10934 2115 10940 2149
rect 10974 2115 10980 2149
rect 10934 2077 10980 2115
rect 10934 2043 10940 2077
rect 10974 2043 10980 2077
rect 11494 2229 11540 2276
rect 11494 2195 11500 2229
rect 11534 2195 11540 2229
rect 11494 2157 11540 2195
rect 11494 2123 11500 2157
rect 11534 2123 11540 2157
rect 11494 2076 11540 2123
rect 11652 2229 11698 2276
rect 11652 2195 11658 2229
rect 11692 2195 11698 2229
rect 11652 2157 11698 2195
rect 11652 2123 11658 2157
rect 11692 2123 11698 2157
rect 11652 2076 11698 2123
rect 13706 2267 13752 2305
rect 13706 2233 13712 2267
rect 13746 2233 13752 2267
rect 13706 2195 13752 2233
rect 13706 2161 13712 2195
rect 13746 2161 13752 2195
rect 13706 2123 13752 2161
rect 13706 2089 13712 2123
rect 13746 2089 13752 2123
rect 10934 2005 10980 2043
rect 10934 1971 10940 2005
rect 10974 1971 10980 2005
rect 10934 1933 10980 1971
rect 10934 1899 10940 1933
rect 10974 1899 10980 1933
rect 10934 1861 10980 1899
rect 10934 1827 10940 1861
rect 10974 1827 10980 1861
rect 10934 1812 10980 1827
rect 13706 2051 13752 2089
rect 13706 2017 13712 2051
rect 13746 2017 13752 2051
rect 13706 1979 13752 2017
rect 13706 1945 13712 1979
rect 13746 1945 13752 1979
rect 13706 1907 13752 1945
rect 13706 1873 13712 1907
rect 13746 1873 13752 1907
rect 13706 1835 13752 1873
rect 13706 1801 13712 1835
rect 13746 1801 13752 1835
rect 13706 1786 13752 1801
rect 13802 2771 13848 2786
rect 13802 2737 13808 2771
rect 13842 2737 13848 2771
rect 13802 2699 13848 2737
rect 13802 2665 13808 2699
rect 13842 2665 13848 2699
rect 13802 2627 13848 2665
rect 13802 2593 13808 2627
rect 13842 2593 13848 2627
rect 13802 2555 13848 2593
rect 13802 2521 13808 2555
rect 13842 2521 13848 2555
rect 13802 2483 13848 2521
rect 13802 2449 13808 2483
rect 13842 2449 13848 2483
rect 13802 2411 13848 2449
rect 13802 2377 13808 2411
rect 13842 2377 13848 2411
rect 13802 2339 13848 2377
rect 13802 2305 13808 2339
rect 13842 2305 13848 2339
rect 13802 2267 13848 2305
rect 13802 2233 13808 2267
rect 13842 2233 13848 2267
rect 13802 2195 13848 2233
rect 13802 2161 13808 2195
rect 13842 2161 13848 2195
rect 13802 2123 13848 2161
rect 13802 2089 13808 2123
rect 13842 2089 13848 2123
rect 13802 2051 13848 2089
rect 13802 2017 13808 2051
rect 13842 2017 13848 2051
rect 13802 1979 13848 2017
rect 13802 1945 13808 1979
rect 13842 1945 13848 1979
rect 13802 1907 13848 1945
rect 13802 1873 13808 1907
rect 13842 1873 13848 1907
rect 13802 1835 13848 1873
rect 13802 1801 13808 1835
rect 13842 1801 13848 1835
rect 13802 1786 13848 1801
rect 13898 2771 13944 2786
rect 13898 2737 13904 2771
rect 13938 2737 13944 2771
rect 13898 2699 13944 2737
rect 13898 2665 13904 2699
rect 13938 2665 13944 2699
rect 13898 2627 13944 2665
rect 13898 2593 13904 2627
rect 13938 2593 13944 2627
rect 13898 2555 13944 2593
rect 13898 2521 13904 2555
rect 13938 2521 13944 2555
rect 13898 2483 13944 2521
rect 13898 2449 13904 2483
rect 13938 2449 13944 2483
rect 13898 2411 13944 2449
rect 13898 2377 13904 2411
rect 13938 2377 13944 2411
rect 13898 2339 13944 2377
rect 13898 2305 13904 2339
rect 13938 2305 13944 2339
rect 13898 2267 13944 2305
rect 13898 2233 13904 2267
rect 13938 2233 13944 2267
rect 13898 2195 13944 2233
rect 13898 2161 13904 2195
rect 13938 2161 13944 2195
rect 13898 2123 13944 2161
rect 13898 2089 13904 2123
rect 13938 2089 13944 2123
rect 13898 2051 13944 2089
rect 13898 2017 13904 2051
rect 13938 2017 13944 2051
rect 13898 1979 13944 2017
rect 13898 1945 13904 1979
rect 13938 1945 13944 1979
rect 13898 1907 13944 1945
rect 13898 1873 13904 1907
rect 13938 1873 13944 1907
rect 13898 1835 13944 1873
rect 13898 1801 13904 1835
rect 13938 1801 13944 1835
rect 13898 1786 13944 1801
rect 13994 2771 14040 2786
rect 13994 2737 14000 2771
rect 14034 2737 14040 2771
rect 13994 2699 14040 2737
rect 13994 2665 14000 2699
rect 14034 2665 14040 2699
rect 13994 2627 14040 2665
rect 13994 2593 14000 2627
rect 14034 2593 14040 2627
rect 13994 2555 14040 2593
rect 13994 2521 14000 2555
rect 14034 2521 14040 2555
rect 13994 2483 14040 2521
rect 13994 2449 14000 2483
rect 14034 2449 14040 2483
rect 13994 2411 14040 2449
rect 13994 2377 14000 2411
rect 14034 2377 14040 2411
rect 13994 2339 14040 2377
rect 13994 2305 14000 2339
rect 14034 2305 14040 2339
rect 13994 2267 14040 2305
rect 13994 2233 14000 2267
rect 14034 2233 14040 2267
rect 13994 2195 14040 2233
rect 13994 2161 14000 2195
rect 14034 2161 14040 2195
rect 13994 2123 14040 2161
rect 13994 2089 14000 2123
rect 14034 2089 14040 2123
rect 13994 2051 14040 2089
rect 13994 2017 14000 2051
rect 14034 2017 14040 2051
rect 13994 1979 14040 2017
rect 13994 1945 14000 1979
rect 14034 1945 14040 1979
rect 13994 1907 14040 1945
rect 13994 1873 14000 1907
rect 14034 1873 14040 1907
rect 13994 1835 14040 1873
rect 13994 1801 14000 1835
rect 14034 1801 14040 1835
rect 13994 1786 14040 1801
rect 14090 2771 14136 2786
rect 14090 2737 14096 2771
rect 14130 2737 14136 2771
rect 14090 2699 14136 2737
rect 14090 2665 14096 2699
rect 14130 2665 14136 2699
rect 14090 2627 14136 2665
rect 14090 2593 14096 2627
rect 14130 2593 14136 2627
rect 14090 2555 14136 2593
rect 14090 2521 14096 2555
rect 14130 2521 14136 2555
rect 14090 2483 14136 2521
rect 14090 2449 14096 2483
rect 14130 2449 14136 2483
rect 14090 2411 14136 2449
rect 14090 2377 14096 2411
rect 14130 2377 14136 2411
rect 14090 2339 14136 2377
rect 14090 2305 14096 2339
rect 14130 2305 14136 2339
rect 14090 2267 14136 2305
rect 14232 2360 14294 3112
rect 14550 2428 14642 3684
rect 14550 2394 14579 2428
rect 14613 2394 14642 2428
rect 14550 2388 14642 2394
rect 14232 2350 14442 2360
rect 14232 2316 14392 2350
rect 14426 2316 14442 2350
rect 14232 2298 14442 2316
rect 14090 2233 14096 2267
rect 14130 2233 14136 2267
rect 14090 2195 14136 2233
rect 14090 2161 14096 2195
rect 14130 2161 14136 2195
rect 14090 2123 14136 2161
rect 14090 2089 14096 2123
rect 14130 2089 14136 2123
rect 14090 2051 14136 2089
rect 14494 2229 14540 2276
rect 14494 2195 14500 2229
rect 14534 2195 14540 2229
rect 14494 2157 14540 2195
rect 14494 2123 14500 2157
rect 14534 2123 14540 2157
rect 14494 2076 14540 2123
rect 14652 2229 14698 2276
rect 14652 2195 14658 2229
rect 14692 2195 14698 2229
rect 14652 2157 14698 2195
rect 14652 2123 14658 2157
rect 14692 2123 14698 2157
rect 14652 2076 14698 2123
rect 14090 2017 14096 2051
rect 14130 2017 14136 2051
rect 14090 1979 14136 2017
rect 14090 1945 14096 1979
rect 14130 1945 14136 1979
rect 14090 1907 14136 1945
rect 14090 1873 14096 1907
rect 14130 1873 14136 1907
rect 14090 1835 14136 1873
rect 14090 1801 14096 1835
rect 14130 1801 14136 1835
rect 14090 1786 14136 1801
rect 1566 1696 1624 1708
rect 1566 1662 1578 1696
rect 1612 1662 1624 1696
rect 1566 1626 1624 1662
rect 4522 1680 4580 1692
rect 4522 1646 4534 1680
rect 4568 1646 4580 1680
rect 706 1546 2456 1626
rect 4522 1614 4580 1646
rect 7552 1680 7610 1692
rect 7552 1646 7564 1680
rect 7598 1646 7610 1680
rect 3674 1612 5408 1614
rect 706 1458 798 1546
rect 706 1424 734 1458
rect 768 1424 798 1458
rect 706 1404 798 1424
rect 2382 1452 2456 1546
rect 2382 1418 2400 1452
rect 2434 1418 2456 1452
rect 2382 1404 2456 1418
rect 3672 1530 5408 1612
rect 7552 1610 7610 1646
rect 10640 1678 10698 1690
rect 10640 1644 10652 1678
rect 10686 1644 10698 1678
rect 10640 1612 10698 1644
rect 13796 1652 13854 1664
rect 13796 1618 13808 1652
rect 13842 1618 13854 1652
rect 3672 1442 3746 1530
rect 3672 1408 3690 1442
rect 3724 1408 3746 1442
rect 3672 1390 3746 1408
rect 5332 1436 5408 1530
rect 5332 1402 5356 1436
rect 5390 1402 5408 1436
rect 5332 1388 5408 1402
rect 6700 1524 8436 1610
rect 6700 1442 6776 1524
rect 6700 1408 6720 1442
rect 6754 1408 6776 1442
rect 6700 1384 6776 1408
rect 8360 1436 8436 1524
rect 8360 1402 8386 1436
rect 8420 1402 8436 1436
rect 8360 1378 8436 1402
rect 9788 1526 11530 1612
rect 13796 1592 13854 1618
rect 9788 1440 9864 1526
rect 9788 1406 9808 1440
rect 9842 1406 9864 1440
rect 9788 1380 9864 1406
rect 11452 1434 11530 1526
rect 11452 1400 11474 1434
rect 11508 1400 11530 1434
rect 11452 1388 11530 1400
rect 12940 1510 14684 1592
rect 12940 1414 13018 1510
rect 12940 1380 12964 1414
rect 12998 1380 13018 1414
rect 12940 1354 13018 1380
rect 14608 1408 14684 1510
rect 14608 1374 14630 1408
rect 14664 1374 14684 1408
rect 14608 1358 14684 1374
rect 15332 1380 15394 3732
rect 15698 3726 15710 3760
rect 15744 3726 15760 3760
rect 15452 1692 15514 1736
rect 15446 1596 15456 1692
rect 15538 1596 15548 1692
rect 15452 1492 15514 1596
rect 15452 1458 15466 1492
rect 15500 1458 15514 1492
rect 15452 1444 15514 1458
rect 15332 1370 15468 1380
rect -1110 1264 -1095 1298
rect -1061 1264 -1048 1298
rect -1110 1256 -1048 1264
rect -916 1298 -420 1354
rect 15332 1336 15422 1370
rect 15456 1336 15468 1370
rect 15332 1328 15468 1336
rect 15332 1326 15394 1328
rect -916 1264 -899 1298
rect -865 1264 -420 1298
rect -916 1238 -420 1264
rect -1692 1051 -1646 1066
rect -1692 1017 -1686 1051
rect -1652 1017 -1646 1051
rect -1692 979 -1646 1017
rect -1692 945 -1686 979
rect -1652 945 -1646 979
rect -1692 907 -1646 945
rect -1692 873 -1686 907
rect -1652 873 -1646 907
rect -1692 835 -1646 873
rect -1692 801 -1686 835
rect -1652 801 -1646 835
rect -1692 763 -1646 801
rect -1692 729 -1686 763
rect -1652 729 -1646 763
rect -1692 691 -1646 729
rect -1692 657 -1686 691
rect -1652 657 -1646 691
rect -1692 619 -1646 657
rect -1692 585 -1686 619
rect -1652 585 -1646 619
rect -1692 547 -1646 585
rect -1692 513 -1686 547
rect -1652 513 -1646 547
rect -1692 475 -1646 513
rect -1692 441 -1686 475
rect -1652 441 -1646 475
rect -1692 403 -1646 441
rect -1692 369 -1686 403
rect -1652 369 -1646 403
rect -1692 331 -1646 369
rect -1692 297 -1686 331
rect -1652 297 -1646 331
rect -1692 259 -1646 297
rect -1692 225 -1686 259
rect -1652 225 -1646 259
rect -1692 187 -1646 225
rect -1692 153 -1686 187
rect -1652 153 -1646 187
rect -1692 115 -1646 153
rect -1692 81 -1686 115
rect -1652 81 -1646 115
rect -1692 66 -1646 81
rect -1594 1051 -1548 1066
rect -1594 1017 -1588 1051
rect -1554 1017 -1548 1051
rect -1594 979 -1548 1017
rect -1594 945 -1588 979
rect -1554 945 -1548 979
rect -1594 907 -1548 945
rect -1594 873 -1588 907
rect -1554 873 -1548 907
rect -1594 835 -1548 873
rect -1594 801 -1588 835
rect -1554 801 -1548 835
rect -1594 763 -1548 801
rect -1594 729 -1588 763
rect -1554 729 -1548 763
rect -1594 691 -1548 729
rect -1594 657 -1588 691
rect -1554 657 -1548 691
rect -1594 619 -1548 657
rect -1594 585 -1588 619
rect -1554 585 -1548 619
rect -1594 547 -1548 585
rect -1594 513 -1588 547
rect -1554 513 -1548 547
rect -1594 475 -1548 513
rect -1594 441 -1588 475
rect -1554 441 -1548 475
rect -1594 403 -1548 441
rect -1594 369 -1588 403
rect -1554 369 -1548 403
rect -1594 331 -1548 369
rect -1594 297 -1588 331
rect -1554 297 -1548 331
rect -1594 259 -1548 297
rect -1594 225 -1588 259
rect -1554 225 -1548 259
rect -1594 187 -1548 225
rect -1594 153 -1588 187
rect -1554 153 -1548 187
rect -1594 115 -1548 153
rect -1594 81 -1588 115
rect -1554 81 -1548 115
rect -1594 66 -1548 81
rect -1496 1051 -1450 1066
rect -1496 1017 -1490 1051
rect -1456 1017 -1450 1051
rect -1496 979 -1450 1017
rect -1496 945 -1490 979
rect -1456 945 -1450 979
rect -1496 907 -1450 945
rect -1496 873 -1490 907
rect -1456 873 -1450 907
rect -1496 835 -1450 873
rect -1496 801 -1490 835
rect -1456 801 -1450 835
rect -1496 763 -1450 801
rect -1496 729 -1490 763
rect -1456 729 -1450 763
rect -1496 691 -1450 729
rect -1496 657 -1490 691
rect -1456 657 -1450 691
rect -1496 619 -1450 657
rect -1496 585 -1490 619
rect -1456 585 -1450 619
rect -1496 547 -1450 585
rect -1496 513 -1490 547
rect -1456 513 -1450 547
rect -1496 475 -1450 513
rect -1496 441 -1490 475
rect -1456 441 -1450 475
rect -1496 403 -1450 441
rect -1496 369 -1490 403
rect -1456 369 -1450 403
rect -1496 331 -1450 369
rect -1496 297 -1490 331
rect -1456 297 -1450 331
rect -1496 259 -1450 297
rect -1496 225 -1490 259
rect -1456 225 -1450 259
rect -1496 187 -1450 225
rect -1496 153 -1490 187
rect -1456 153 -1450 187
rect -1496 115 -1450 153
rect -1496 81 -1490 115
rect -1456 81 -1450 115
rect -1496 66 -1450 81
rect -1398 1051 -1352 1066
rect -1398 1017 -1392 1051
rect -1358 1017 -1352 1051
rect -1398 979 -1352 1017
rect -1398 945 -1392 979
rect -1358 945 -1352 979
rect -1398 907 -1352 945
rect -1398 873 -1392 907
rect -1358 873 -1352 907
rect -1398 835 -1352 873
rect -1398 801 -1392 835
rect -1358 801 -1352 835
rect -1398 763 -1352 801
rect -1398 729 -1392 763
rect -1358 729 -1352 763
rect -1398 691 -1352 729
rect -1398 657 -1392 691
rect -1358 657 -1352 691
rect -1398 619 -1352 657
rect -1398 585 -1392 619
rect -1358 585 -1352 619
rect -1398 547 -1352 585
rect -1398 513 -1392 547
rect -1358 513 -1352 547
rect -1398 475 -1352 513
rect -1398 441 -1392 475
rect -1358 441 -1352 475
rect -1398 403 -1352 441
rect -1398 369 -1392 403
rect -1358 369 -1352 403
rect -1398 331 -1352 369
rect -1398 297 -1392 331
rect -1358 297 -1352 331
rect -1398 259 -1352 297
rect -1398 225 -1392 259
rect -1358 225 -1352 259
rect -1398 187 -1352 225
rect -1398 153 -1392 187
rect -1358 153 -1352 187
rect -1398 115 -1352 153
rect -1398 81 -1392 115
rect -1358 81 -1352 115
rect -1398 66 -1352 81
rect -1300 1051 -1254 1066
rect -1300 1017 -1294 1051
rect -1260 1017 -1254 1051
rect -1300 979 -1254 1017
rect -1300 945 -1294 979
rect -1260 945 -1254 979
rect -1300 907 -1254 945
rect -1300 873 -1294 907
rect -1260 873 -1254 907
rect -1300 835 -1254 873
rect -1300 801 -1294 835
rect -1260 801 -1254 835
rect -1300 763 -1254 801
rect -1300 729 -1294 763
rect -1260 729 -1254 763
rect -1300 691 -1254 729
rect -1300 657 -1294 691
rect -1260 657 -1254 691
rect -1300 619 -1254 657
rect -1300 585 -1294 619
rect -1260 585 -1254 619
rect -1300 547 -1254 585
rect -1300 513 -1294 547
rect -1260 513 -1254 547
rect -1300 475 -1254 513
rect -1300 441 -1294 475
rect -1260 441 -1254 475
rect -1300 403 -1254 441
rect -1300 369 -1294 403
rect -1260 369 -1254 403
rect -1300 331 -1254 369
rect -1300 297 -1294 331
rect -1260 297 -1254 331
rect -1300 259 -1254 297
rect -1300 225 -1294 259
rect -1260 225 -1254 259
rect -1300 187 -1254 225
rect -1300 153 -1294 187
rect -1260 153 -1254 187
rect -1300 115 -1254 153
rect -1300 81 -1294 115
rect -1260 81 -1254 115
rect -1300 66 -1254 81
rect -1202 1051 -1156 1066
rect -1202 1017 -1196 1051
rect -1162 1017 -1156 1051
rect -1202 979 -1156 1017
rect -1202 945 -1196 979
rect -1162 945 -1156 979
rect -1202 907 -1156 945
rect -1202 873 -1196 907
rect -1162 873 -1156 907
rect -1202 835 -1156 873
rect -1202 801 -1196 835
rect -1162 801 -1156 835
rect -1202 763 -1156 801
rect -1202 729 -1196 763
rect -1162 729 -1156 763
rect -1202 691 -1156 729
rect -1202 657 -1196 691
rect -1162 657 -1156 691
rect -1202 619 -1156 657
rect -1202 585 -1196 619
rect -1162 585 -1156 619
rect -1202 547 -1156 585
rect -1202 513 -1196 547
rect -1162 513 -1156 547
rect -1202 475 -1156 513
rect -1202 441 -1196 475
rect -1162 441 -1156 475
rect -1202 403 -1156 441
rect -1202 369 -1196 403
rect -1162 369 -1156 403
rect -1202 331 -1156 369
rect -1202 297 -1196 331
rect -1162 297 -1156 331
rect -1202 259 -1156 297
rect -1202 225 -1196 259
rect -1162 225 -1156 259
rect -1202 187 -1156 225
rect -1202 153 -1196 187
rect -1162 153 -1156 187
rect -1202 115 -1156 153
rect -1202 81 -1196 115
rect -1162 81 -1156 115
rect -1202 66 -1156 81
rect -1104 1051 -1058 1066
rect -1104 1017 -1098 1051
rect -1064 1017 -1058 1051
rect -1104 979 -1058 1017
rect -1104 945 -1098 979
rect -1064 945 -1058 979
rect -1104 907 -1058 945
rect -1104 873 -1098 907
rect -1064 873 -1058 907
rect -1104 835 -1058 873
rect -1104 801 -1098 835
rect -1064 801 -1058 835
rect -1104 763 -1058 801
rect -1104 729 -1098 763
rect -1064 729 -1058 763
rect -1104 691 -1058 729
rect -1104 657 -1098 691
rect -1064 657 -1058 691
rect -1104 619 -1058 657
rect -1104 585 -1098 619
rect -1064 585 -1058 619
rect -1104 547 -1058 585
rect -1104 513 -1098 547
rect -1064 513 -1058 547
rect -1104 475 -1058 513
rect -1104 441 -1098 475
rect -1064 441 -1058 475
rect -1104 403 -1058 441
rect -1104 369 -1098 403
rect -1064 369 -1058 403
rect -1104 331 -1058 369
rect -1104 297 -1098 331
rect -1064 297 -1058 331
rect -1104 259 -1058 297
rect -1104 225 -1098 259
rect -1064 225 -1058 259
rect -1104 187 -1058 225
rect -1104 153 -1098 187
rect -1064 153 -1058 187
rect -1104 115 -1058 153
rect -1104 81 -1098 115
rect -1064 81 -1058 115
rect -1104 66 -1058 81
rect -1006 1051 -960 1066
rect -1006 1017 -1000 1051
rect -966 1017 -960 1051
rect -1006 979 -960 1017
rect -1006 945 -1000 979
rect -966 945 -960 979
rect -1006 907 -960 945
rect -1006 873 -1000 907
rect -966 873 -960 907
rect -1006 835 -960 873
rect -1006 801 -1000 835
rect -966 801 -960 835
rect -1006 763 -960 801
rect -1006 729 -1000 763
rect -966 729 -960 763
rect -1006 691 -960 729
rect -1006 657 -1000 691
rect -966 657 -960 691
rect -1006 619 -960 657
rect -1006 585 -1000 619
rect -966 585 -960 619
rect -1006 547 -960 585
rect -1006 513 -1000 547
rect -966 513 -960 547
rect -1006 475 -960 513
rect -1006 441 -1000 475
rect -966 441 -960 475
rect -1006 403 -960 441
rect -1006 369 -1000 403
rect -966 369 -960 403
rect -1006 331 -960 369
rect -1006 297 -1000 331
rect -966 297 -960 331
rect -1006 259 -960 297
rect -1006 225 -1000 259
rect -966 225 -960 259
rect -1006 187 -960 225
rect -1006 153 -1000 187
rect -966 153 -960 187
rect -1006 115 -960 153
rect -1006 81 -1000 115
rect -966 81 -960 115
rect -1006 66 -960 81
rect -908 1051 -862 1066
rect -908 1017 -902 1051
rect -868 1017 -862 1051
rect -908 979 -862 1017
rect -908 945 -902 979
rect -868 945 -862 979
rect -908 907 -862 945
rect -908 873 -902 907
rect -868 873 -862 907
rect -908 835 -862 873
rect -908 801 -902 835
rect -868 801 -862 835
rect -908 763 -862 801
rect -908 729 -902 763
rect -868 729 -862 763
rect -908 691 -862 729
rect -908 657 -902 691
rect -868 657 -862 691
rect -908 619 -862 657
rect -908 585 -902 619
rect -868 585 -862 619
rect -908 547 -862 585
rect -908 513 -902 547
rect -868 513 -862 547
rect -908 475 -862 513
rect -908 441 -902 475
rect -868 441 -862 475
rect -908 403 -862 441
rect -908 369 -902 403
rect -868 369 -862 403
rect -908 331 -862 369
rect -908 297 -902 331
rect -868 297 -862 331
rect -908 259 -862 297
rect -908 225 -902 259
rect -868 225 -862 259
rect -908 187 -862 225
rect -908 153 -902 187
rect -868 153 -862 187
rect -908 115 -862 153
rect -908 81 -902 115
rect -868 81 -862 115
rect -908 66 -862 81
rect -560 -126 -420 1238
rect 152 1253 198 1268
rect 152 1219 158 1253
rect 192 1219 198 1253
rect 152 1181 198 1219
rect 152 1147 158 1181
rect 192 1147 198 1181
rect 152 1109 198 1147
rect 152 1075 158 1109
rect 192 1075 198 1109
rect 152 1037 198 1075
rect 152 1003 158 1037
rect 192 1003 198 1037
rect 152 965 198 1003
rect 152 931 158 965
rect 192 931 198 965
rect 152 893 198 931
rect 152 859 158 893
rect 192 859 198 893
rect 152 821 198 859
rect 152 787 158 821
rect 192 787 198 821
rect 152 749 198 787
rect 152 715 158 749
rect 192 715 198 749
rect 152 677 198 715
rect 152 643 158 677
rect 192 643 198 677
rect 152 605 198 643
rect 152 571 158 605
rect 192 571 198 605
rect 152 533 198 571
rect 152 499 158 533
rect 192 499 198 533
rect 152 461 198 499
rect 152 427 158 461
rect 192 427 198 461
rect 152 389 198 427
rect 152 355 158 389
rect 192 355 198 389
rect 152 317 198 355
rect 152 283 158 317
rect 192 283 198 317
rect 152 268 198 283
rect 248 1253 294 1268
rect 248 1219 254 1253
rect 288 1219 294 1253
rect 248 1181 294 1219
rect 248 1147 254 1181
rect 288 1147 294 1181
rect 248 1109 294 1147
rect 248 1075 254 1109
rect 288 1075 294 1109
rect 248 1037 294 1075
rect 248 1003 254 1037
rect 288 1003 294 1037
rect 248 965 294 1003
rect 248 931 254 965
rect 288 931 294 965
rect 248 893 294 931
rect 248 859 254 893
rect 288 859 294 893
rect 248 821 294 859
rect 248 787 254 821
rect 288 787 294 821
rect 248 749 294 787
rect 248 715 254 749
rect 288 715 294 749
rect 248 677 294 715
rect 248 643 254 677
rect 288 643 294 677
rect 248 605 294 643
rect 248 571 254 605
rect 288 571 294 605
rect 248 533 294 571
rect 248 499 254 533
rect 288 499 294 533
rect 248 461 294 499
rect 248 427 254 461
rect 288 427 294 461
rect 248 389 294 427
rect 248 355 254 389
rect 288 355 294 389
rect 248 317 294 355
rect 248 283 254 317
rect 288 283 294 317
rect 248 268 294 283
rect 344 1253 390 1268
rect 344 1219 350 1253
rect 384 1219 390 1253
rect 344 1181 390 1219
rect 344 1147 350 1181
rect 384 1147 390 1181
rect 344 1109 390 1147
rect 344 1075 350 1109
rect 384 1075 390 1109
rect 344 1037 390 1075
rect 344 1003 350 1037
rect 384 1003 390 1037
rect 344 965 390 1003
rect 344 931 350 965
rect 384 931 390 965
rect 344 893 390 931
rect 344 859 350 893
rect 384 859 390 893
rect 344 821 390 859
rect 344 787 350 821
rect 384 787 390 821
rect 344 749 390 787
rect 344 715 350 749
rect 384 715 390 749
rect 344 677 390 715
rect 344 643 350 677
rect 384 643 390 677
rect 344 605 390 643
rect 344 571 350 605
rect 384 571 390 605
rect 344 533 390 571
rect 344 499 350 533
rect 384 499 390 533
rect 344 461 390 499
rect 344 427 350 461
rect 384 427 390 461
rect 344 389 390 427
rect 344 355 350 389
rect 384 355 390 389
rect 344 317 390 355
rect 344 283 350 317
rect 384 283 390 317
rect 344 268 390 283
rect 440 1253 486 1268
rect 440 1219 446 1253
rect 480 1219 486 1253
rect 440 1181 486 1219
rect 440 1147 446 1181
rect 480 1147 486 1181
rect 440 1109 486 1147
rect 440 1075 446 1109
rect 480 1075 486 1109
rect 440 1037 486 1075
rect 440 1003 446 1037
rect 480 1003 486 1037
rect 440 965 486 1003
rect 440 931 446 965
rect 480 931 486 965
rect 440 893 486 931
rect 440 859 446 893
rect 480 859 486 893
rect 440 821 486 859
rect 440 787 446 821
rect 480 787 486 821
rect 440 749 486 787
rect 440 715 446 749
rect 480 715 486 749
rect 440 677 486 715
rect 440 643 446 677
rect 480 643 486 677
rect 440 605 486 643
rect 440 571 446 605
rect 480 571 486 605
rect 440 533 486 571
rect 440 499 446 533
rect 480 499 486 533
rect 440 461 486 499
rect 440 427 446 461
rect 480 427 486 461
rect 440 389 486 427
rect 440 355 446 389
rect 480 355 486 389
rect 440 317 486 355
rect 440 283 446 317
rect 480 283 486 317
rect 440 268 486 283
rect 536 1253 582 1268
rect 536 1219 542 1253
rect 576 1219 582 1253
rect 536 1181 582 1219
rect 536 1147 542 1181
rect 576 1147 582 1181
rect 536 1109 582 1147
rect 536 1075 542 1109
rect 576 1075 582 1109
rect 536 1037 582 1075
rect 536 1003 542 1037
rect 576 1003 582 1037
rect 536 965 582 1003
rect 536 931 542 965
rect 576 931 582 965
rect 536 893 582 931
rect 536 859 542 893
rect 576 859 582 893
rect 536 821 582 859
rect 536 787 542 821
rect 576 787 582 821
rect 536 749 582 787
rect 536 715 542 749
rect 576 715 582 749
rect 536 677 582 715
rect 536 643 542 677
rect 576 643 582 677
rect 536 605 582 643
rect 536 571 542 605
rect 576 571 582 605
rect 536 533 582 571
rect 536 499 542 533
rect 576 499 582 533
rect 536 461 582 499
rect 536 427 542 461
rect 576 427 582 461
rect 536 389 582 427
rect 536 355 542 389
rect 576 355 582 389
rect 536 317 582 355
rect 536 283 542 317
rect 576 283 582 317
rect 536 268 582 283
rect 632 1253 678 1268
rect 632 1219 638 1253
rect 672 1219 678 1253
rect 632 1181 678 1219
rect 632 1147 638 1181
rect 672 1147 678 1181
rect 632 1109 678 1147
rect 632 1075 638 1109
rect 672 1075 678 1109
rect 632 1037 678 1075
rect 632 1003 638 1037
rect 672 1003 678 1037
rect 632 965 678 1003
rect 632 931 638 965
rect 672 931 678 965
rect 632 893 678 931
rect 632 859 638 893
rect 672 859 678 893
rect 632 821 678 859
rect 632 787 638 821
rect 672 787 678 821
rect 632 749 678 787
rect 632 715 638 749
rect 672 715 678 749
rect 632 677 678 715
rect 632 643 638 677
rect 672 643 678 677
rect 632 605 678 643
rect 632 571 638 605
rect 672 571 678 605
rect 632 533 678 571
rect 632 499 638 533
rect 672 499 678 533
rect 632 461 678 499
rect 632 427 638 461
rect 672 427 678 461
rect 632 389 678 427
rect 632 355 638 389
rect 672 355 678 389
rect 632 317 678 355
rect 632 283 638 317
rect 672 283 678 317
rect 632 268 678 283
rect 728 1253 774 1268
rect 728 1219 734 1253
rect 768 1219 774 1253
rect 728 1181 774 1219
rect 728 1147 734 1181
rect 768 1147 774 1181
rect 728 1109 774 1147
rect 728 1075 734 1109
rect 768 1075 774 1109
rect 728 1037 774 1075
rect 728 1003 734 1037
rect 768 1003 774 1037
rect 728 965 774 1003
rect 728 931 734 965
rect 768 931 774 965
rect 728 893 774 931
rect 728 859 734 893
rect 768 859 774 893
rect 728 821 774 859
rect 728 787 734 821
rect 768 787 774 821
rect 728 749 774 787
rect 728 715 734 749
rect 768 715 774 749
rect 728 677 774 715
rect 728 643 734 677
rect 768 643 774 677
rect 728 605 774 643
rect 728 571 734 605
rect 768 571 774 605
rect 728 533 774 571
rect 728 499 734 533
rect 768 499 774 533
rect 728 461 774 499
rect 728 427 734 461
rect 768 427 774 461
rect 728 389 774 427
rect 728 355 734 389
rect 768 355 774 389
rect 728 317 774 355
rect 728 283 734 317
rect 768 283 774 317
rect 728 268 774 283
rect 824 1253 870 1268
rect 824 1219 830 1253
rect 864 1219 870 1253
rect 824 1181 870 1219
rect 824 1147 830 1181
rect 864 1147 870 1181
rect 824 1109 870 1147
rect 824 1075 830 1109
rect 864 1075 870 1109
rect 824 1037 870 1075
rect 824 1003 830 1037
rect 864 1003 870 1037
rect 824 965 870 1003
rect 824 931 830 965
rect 864 931 870 965
rect 824 893 870 931
rect 824 859 830 893
rect 864 859 870 893
rect 824 821 870 859
rect 824 787 830 821
rect 864 787 870 821
rect 824 749 870 787
rect 824 715 830 749
rect 864 715 870 749
rect 824 677 870 715
rect 824 643 830 677
rect 864 643 870 677
rect 824 605 870 643
rect 824 571 830 605
rect 864 571 870 605
rect 824 533 870 571
rect 824 499 830 533
rect 864 499 870 533
rect 824 461 870 499
rect 824 427 830 461
rect 864 427 870 461
rect 824 389 870 427
rect 824 355 830 389
rect 864 355 870 389
rect 824 317 870 355
rect 824 283 830 317
rect 864 283 870 317
rect 824 268 870 283
rect 920 1253 966 1268
rect 920 1219 926 1253
rect 960 1219 966 1253
rect 920 1181 966 1219
rect 920 1147 926 1181
rect 960 1147 966 1181
rect 920 1109 966 1147
rect 920 1075 926 1109
rect 960 1075 966 1109
rect 920 1037 966 1075
rect 920 1003 926 1037
rect 960 1003 966 1037
rect 920 965 966 1003
rect 920 931 926 965
rect 960 931 966 965
rect 920 893 966 931
rect 920 859 926 893
rect 960 859 966 893
rect 920 821 966 859
rect 920 787 926 821
rect 960 787 966 821
rect 920 749 966 787
rect 920 715 926 749
rect 960 715 966 749
rect 920 677 966 715
rect 920 643 926 677
rect 960 643 966 677
rect 920 605 966 643
rect 920 571 926 605
rect 960 571 966 605
rect 920 533 966 571
rect 920 499 926 533
rect 960 499 966 533
rect 920 461 966 499
rect 920 427 926 461
rect 960 427 966 461
rect 920 389 966 427
rect 920 355 926 389
rect 960 355 966 389
rect 920 317 966 355
rect 920 283 926 317
rect 960 283 966 317
rect 920 268 966 283
rect 1016 1253 1062 1268
rect 1016 1219 1022 1253
rect 1056 1219 1062 1253
rect 1016 1181 1062 1219
rect 1016 1147 1022 1181
rect 1056 1147 1062 1181
rect 1016 1109 1062 1147
rect 1016 1075 1022 1109
rect 1056 1075 1062 1109
rect 1016 1037 1062 1075
rect 1016 1003 1022 1037
rect 1056 1003 1062 1037
rect 1016 965 1062 1003
rect 1016 931 1022 965
rect 1056 931 1062 965
rect 1016 893 1062 931
rect 1016 859 1022 893
rect 1056 859 1062 893
rect 1016 821 1062 859
rect 1016 787 1022 821
rect 1056 787 1062 821
rect 1016 749 1062 787
rect 1016 715 1022 749
rect 1056 715 1062 749
rect 1016 677 1062 715
rect 1016 643 1022 677
rect 1056 643 1062 677
rect 1016 605 1062 643
rect 1016 571 1022 605
rect 1056 571 1062 605
rect 1016 533 1062 571
rect 1016 499 1022 533
rect 1056 499 1062 533
rect 1016 461 1062 499
rect 1016 427 1022 461
rect 1056 427 1062 461
rect 1016 389 1062 427
rect 1016 355 1022 389
rect 1056 355 1062 389
rect 1016 317 1062 355
rect 1016 283 1022 317
rect 1056 283 1062 317
rect 1016 268 1062 283
rect 1112 1253 1158 1268
rect 1112 1219 1118 1253
rect 1152 1219 1158 1253
rect 1112 1181 1158 1219
rect 1112 1147 1118 1181
rect 1152 1147 1158 1181
rect 1112 1109 1158 1147
rect 1112 1075 1118 1109
rect 1152 1075 1158 1109
rect 1112 1037 1158 1075
rect 1112 1003 1118 1037
rect 1152 1003 1158 1037
rect 1112 965 1158 1003
rect 1112 931 1118 965
rect 1152 931 1158 965
rect 1112 893 1158 931
rect 1112 859 1118 893
rect 1152 859 1158 893
rect 1112 821 1158 859
rect 1112 787 1118 821
rect 1152 787 1158 821
rect 1112 749 1158 787
rect 1112 715 1118 749
rect 1152 715 1158 749
rect 1112 677 1158 715
rect 1112 643 1118 677
rect 1152 643 1158 677
rect 1112 605 1158 643
rect 1112 571 1118 605
rect 1152 571 1158 605
rect 1112 533 1158 571
rect 1112 499 1118 533
rect 1152 499 1158 533
rect 1112 461 1158 499
rect 1112 427 1118 461
rect 1152 427 1158 461
rect 1112 389 1158 427
rect 1112 355 1118 389
rect 1152 355 1158 389
rect 1112 317 1158 355
rect 1112 283 1118 317
rect 1152 283 1158 317
rect 1112 268 1158 283
rect 1208 1253 1254 1268
rect 1208 1219 1214 1253
rect 1248 1219 1254 1253
rect 1208 1181 1254 1219
rect 1208 1147 1214 1181
rect 1248 1147 1254 1181
rect 1208 1109 1254 1147
rect 1208 1075 1214 1109
rect 1248 1075 1254 1109
rect 1208 1037 1254 1075
rect 1208 1003 1214 1037
rect 1248 1003 1254 1037
rect 1208 965 1254 1003
rect 1208 931 1214 965
rect 1248 931 1254 965
rect 1208 893 1254 931
rect 1208 859 1214 893
rect 1248 859 1254 893
rect 1208 821 1254 859
rect 1208 787 1214 821
rect 1248 787 1254 821
rect 1208 749 1254 787
rect 1208 715 1214 749
rect 1248 715 1254 749
rect 1208 677 1254 715
rect 1208 643 1214 677
rect 1248 643 1254 677
rect 1208 605 1254 643
rect 1208 571 1214 605
rect 1248 571 1254 605
rect 1208 533 1254 571
rect 1208 499 1214 533
rect 1248 499 1254 533
rect 1208 461 1254 499
rect 1208 427 1214 461
rect 1248 427 1254 461
rect 1208 389 1254 427
rect 1208 355 1214 389
rect 1248 355 1254 389
rect 1208 317 1254 355
rect 1208 283 1214 317
rect 1248 283 1254 317
rect 1208 268 1254 283
rect 1304 1253 1350 1268
rect 1304 1219 1310 1253
rect 1344 1219 1350 1253
rect 1304 1181 1350 1219
rect 1304 1147 1310 1181
rect 1344 1147 1350 1181
rect 1304 1109 1350 1147
rect 1304 1075 1310 1109
rect 1344 1075 1350 1109
rect 1304 1037 1350 1075
rect 1304 1003 1310 1037
rect 1344 1003 1350 1037
rect 1304 965 1350 1003
rect 1304 931 1310 965
rect 1344 931 1350 965
rect 1304 893 1350 931
rect 1304 859 1310 893
rect 1344 859 1350 893
rect 1304 821 1350 859
rect 1304 787 1310 821
rect 1344 787 1350 821
rect 1304 749 1350 787
rect 1304 715 1310 749
rect 1344 715 1350 749
rect 1304 677 1350 715
rect 1304 643 1310 677
rect 1344 643 1350 677
rect 1304 605 1350 643
rect 1304 571 1310 605
rect 1344 571 1350 605
rect 1304 533 1350 571
rect 1304 499 1310 533
rect 1344 499 1350 533
rect 1304 461 1350 499
rect 1304 427 1310 461
rect 1344 427 1350 461
rect 1304 389 1350 427
rect 1304 355 1310 389
rect 1344 355 1350 389
rect 1304 317 1350 355
rect 1304 283 1310 317
rect 1344 283 1350 317
rect 1304 268 1350 283
rect 1920 1253 1966 1268
rect 1920 1219 1926 1253
rect 1960 1219 1966 1253
rect 1920 1181 1966 1219
rect 1920 1147 1926 1181
rect 1960 1147 1966 1181
rect 1920 1109 1966 1147
rect 1920 1075 1926 1109
rect 1960 1075 1966 1109
rect 1920 1037 1966 1075
rect 1920 1003 1926 1037
rect 1960 1003 1966 1037
rect 1920 965 1966 1003
rect 1920 931 1926 965
rect 1960 931 1966 965
rect 1920 893 1966 931
rect 1920 859 1926 893
rect 1960 859 1966 893
rect 1920 821 1966 859
rect 1920 787 1926 821
rect 1960 787 1966 821
rect 1920 749 1966 787
rect 1920 715 1926 749
rect 1960 715 1966 749
rect 1920 677 1966 715
rect 1920 643 1926 677
rect 1960 643 1966 677
rect 1920 605 1966 643
rect 1920 571 1926 605
rect 1960 571 1966 605
rect 1920 533 1966 571
rect 1920 499 1926 533
rect 1960 499 1966 533
rect 1920 461 1966 499
rect 1920 427 1926 461
rect 1960 427 1966 461
rect 1920 389 1966 427
rect 1920 355 1926 389
rect 1960 355 1966 389
rect 1920 317 1966 355
rect 1920 283 1926 317
rect 1960 283 1966 317
rect 1920 268 1966 283
rect 2016 1253 2062 1268
rect 2016 1219 2022 1253
rect 2056 1219 2062 1253
rect 2016 1181 2062 1219
rect 2016 1147 2022 1181
rect 2056 1147 2062 1181
rect 2016 1109 2062 1147
rect 2016 1075 2022 1109
rect 2056 1075 2062 1109
rect 2016 1037 2062 1075
rect 2016 1003 2022 1037
rect 2056 1003 2062 1037
rect 2016 965 2062 1003
rect 2016 931 2022 965
rect 2056 931 2062 965
rect 2016 893 2062 931
rect 2016 859 2022 893
rect 2056 859 2062 893
rect 2016 821 2062 859
rect 2016 787 2022 821
rect 2056 787 2062 821
rect 2016 749 2062 787
rect 2016 715 2022 749
rect 2056 715 2062 749
rect 2016 677 2062 715
rect 2016 643 2022 677
rect 2056 643 2062 677
rect 2016 605 2062 643
rect 2016 571 2022 605
rect 2056 571 2062 605
rect 2016 533 2062 571
rect 2016 499 2022 533
rect 2056 499 2062 533
rect 2016 461 2062 499
rect 2016 427 2022 461
rect 2056 427 2062 461
rect 2016 389 2062 427
rect 2016 355 2022 389
rect 2056 355 2062 389
rect 2016 317 2062 355
rect 2016 283 2022 317
rect 2056 283 2062 317
rect 2016 268 2062 283
rect 2112 1253 2158 1268
rect 2112 1219 2118 1253
rect 2152 1219 2158 1253
rect 2112 1181 2158 1219
rect 2112 1147 2118 1181
rect 2152 1147 2158 1181
rect 2112 1109 2158 1147
rect 2112 1075 2118 1109
rect 2152 1075 2158 1109
rect 2112 1037 2158 1075
rect 2112 1003 2118 1037
rect 2152 1003 2158 1037
rect 2112 965 2158 1003
rect 2112 931 2118 965
rect 2152 931 2158 965
rect 2112 893 2158 931
rect 2112 859 2118 893
rect 2152 859 2158 893
rect 2112 821 2158 859
rect 2112 787 2118 821
rect 2152 787 2158 821
rect 2112 749 2158 787
rect 2112 715 2118 749
rect 2152 715 2158 749
rect 2112 677 2158 715
rect 2112 643 2118 677
rect 2152 643 2158 677
rect 2112 605 2158 643
rect 2112 571 2118 605
rect 2152 571 2158 605
rect 2112 533 2158 571
rect 2112 499 2118 533
rect 2152 499 2158 533
rect 2112 461 2158 499
rect 2112 427 2118 461
rect 2152 427 2158 461
rect 2112 389 2158 427
rect 2112 355 2118 389
rect 2152 355 2158 389
rect 2112 317 2158 355
rect 2112 283 2118 317
rect 2152 283 2158 317
rect 2112 268 2158 283
rect 2208 1253 2254 1268
rect 2208 1219 2214 1253
rect 2248 1219 2254 1253
rect 2208 1181 2254 1219
rect 2208 1147 2214 1181
rect 2248 1147 2254 1181
rect 2208 1109 2254 1147
rect 2208 1075 2214 1109
rect 2248 1075 2254 1109
rect 2208 1037 2254 1075
rect 2208 1003 2214 1037
rect 2248 1003 2254 1037
rect 2208 965 2254 1003
rect 2208 931 2214 965
rect 2248 931 2254 965
rect 2208 893 2254 931
rect 2208 859 2214 893
rect 2248 859 2254 893
rect 2208 821 2254 859
rect 2208 787 2214 821
rect 2248 787 2254 821
rect 2208 749 2254 787
rect 2208 715 2214 749
rect 2248 715 2254 749
rect 2208 677 2254 715
rect 2208 643 2214 677
rect 2248 643 2254 677
rect 2208 605 2254 643
rect 2208 571 2214 605
rect 2248 571 2254 605
rect 2208 533 2254 571
rect 2208 499 2214 533
rect 2248 499 2254 533
rect 2208 461 2254 499
rect 2208 427 2214 461
rect 2248 427 2254 461
rect 2208 389 2254 427
rect 2208 355 2214 389
rect 2248 355 2254 389
rect 2208 317 2254 355
rect 2208 283 2214 317
rect 2248 283 2254 317
rect 2208 268 2254 283
rect 2304 1253 2350 1268
rect 2304 1219 2310 1253
rect 2344 1219 2350 1253
rect 2304 1181 2350 1219
rect 2304 1147 2310 1181
rect 2344 1147 2350 1181
rect 2304 1109 2350 1147
rect 2304 1075 2310 1109
rect 2344 1075 2350 1109
rect 2304 1037 2350 1075
rect 2304 1003 2310 1037
rect 2344 1003 2350 1037
rect 2304 965 2350 1003
rect 2304 931 2310 965
rect 2344 931 2350 965
rect 2304 893 2350 931
rect 2304 859 2310 893
rect 2344 859 2350 893
rect 2304 821 2350 859
rect 2304 787 2310 821
rect 2344 787 2350 821
rect 2304 749 2350 787
rect 2304 715 2310 749
rect 2344 715 2350 749
rect 2304 677 2350 715
rect 2304 643 2310 677
rect 2344 643 2350 677
rect 2304 605 2350 643
rect 2304 571 2310 605
rect 2344 571 2350 605
rect 2304 533 2350 571
rect 2304 499 2310 533
rect 2344 499 2350 533
rect 2304 461 2350 499
rect 2304 427 2310 461
rect 2344 427 2350 461
rect 2304 389 2350 427
rect 2304 355 2310 389
rect 2344 355 2350 389
rect 2304 317 2350 355
rect 2304 283 2310 317
rect 2344 283 2350 317
rect 2304 268 2350 283
rect 2400 1253 2446 1268
rect 2400 1219 2406 1253
rect 2440 1219 2446 1253
rect 2400 1181 2446 1219
rect 2400 1147 2406 1181
rect 2440 1147 2446 1181
rect 2400 1109 2446 1147
rect 2400 1075 2406 1109
rect 2440 1075 2446 1109
rect 2400 1037 2446 1075
rect 2400 1003 2406 1037
rect 2440 1003 2446 1037
rect 2400 965 2446 1003
rect 2400 931 2406 965
rect 2440 931 2446 965
rect 2400 893 2446 931
rect 2400 859 2406 893
rect 2440 859 2446 893
rect 2400 821 2446 859
rect 2400 787 2406 821
rect 2440 787 2446 821
rect 2400 749 2446 787
rect 2400 715 2406 749
rect 2440 715 2446 749
rect 2400 677 2446 715
rect 2400 643 2406 677
rect 2440 643 2446 677
rect 2400 605 2446 643
rect 2400 571 2406 605
rect 2440 571 2446 605
rect 2400 533 2446 571
rect 2400 499 2406 533
rect 2440 499 2446 533
rect 2400 461 2446 499
rect 2400 427 2406 461
rect 2440 427 2446 461
rect 2400 389 2446 427
rect 2400 355 2406 389
rect 2440 355 2446 389
rect 2400 317 2446 355
rect 2400 283 2406 317
rect 2440 283 2446 317
rect 2400 268 2446 283
rect 2496 1253 2542 1268
rect 2496 1219 2502 1253
rect 2536 1219 2542 1253
rect 2496 1181 2542 1219
rect 2496 1147 2502 1181
rect 2536 1147 2542 1181
rect 2496 1109 2542 1147
rect 2496 1075 2502 1109
rect 2536 1075 2542 1109
rect 2496 1037 2542 1075
rect 2496 1003 2502 1037
rect 2536 1003 2542 1037
rect 2496 965 2542 1003
rect 2496 931 2502 965
rect 2536 931 2542 965
rect 2496 893 2542 931
rect 2496 859 2502 893
rect 2536 859 2542 893
rect 2496 821 2542 859
rect 2496 787 2502 821
rect 2536 787 2542 821
rect 2496 749 2542 787
rect 2496 715 2502 749
rect 2536 715 2542 749
rect 2496 677 2542 715
rect 2496 643 2502 677
rect 2536 643 2542 677
rect 2496 605 2542 643
rect 2496 571 2502 605
rect 2536 571 2542 605
rect 2496 533 2542 571
rect 2496 499 2502 533
rect 2536 499 2542 533
rect 2496 461 2542 499
rect 2496 427 2502 461
rect 2536 427 2542 461
rect 2496 389 2542 427
rect 2496 355 2502 389
rect 2536 355 2542 389
rect 2496 317 2542 355
rect 2496 283 2502 317
rect 2536 283 2542 317
rect 2496 268 2542 283
rect 2592 1253 2638 1268
rect 2592 1219 2598 1253
rect 2632 1219 2638 1253
rect 2592 1181 2638 1219
rect 2592 1147 2598 1181
rect 2632 1147 2638 1181
rect 2592 1109 2638 1147
rect 2592 1075 2598 1109
rect 2632 1075 2638 1109
rect 2592 1037 2638 1075
rect 2592 1003 2598 1037
rect 2632 1003 2638 1037
rect 2592 965 2638 1003
rect 2592 931 2598 965
rect 2632 931 2638 965
rect 2592 893 2638 931
rect 2592 859 2598 893
rect 2632 859 2638 893
rect 2592 821 2638 859
rect 2592 787 2598 821
rect 2632 787 2638 821
rect 2592 749 2638 787
rect 2592 715 2598 749
rect 2632 715 2638 749
rect 2592 677 2638 715
rect 2592 643 2598 677
rect 2632 643 2638 677
rect 2592 605 2638 643
rect 2592 571 2598 605
rect 2632 571 2638 605
rect 2592 533 2638 571
rect 2592 499 2598 533
rect 2632 499 2638 533
rect 2592 461 2638 499
rect 2592 427 2598 461
rect 2632 427 2638 461
rect 2592 389 2638 427
rect 2592 355 2598 389
rect 2632 355 2638 389
rect 2592 317 2638 355
rect 2592 283 2598 317
rect 2632 283 2638 317
rect 2592 268 2638 283
rect 2688 1253 2734 1268
rect 2688 1219 2694 1253
rect 2728 1219 2734 1253
rect 2688 1181 2734 1219
rect 2688 1147 2694 1181
rect 2728 1147 2734 1181
rect 2688 1109 2734 1147
rect 2688 1075 2694 1109
rect 2728 1075 2734 1109
rect 2688 1037 2734 1075
rect 2688 1003 2694 1037
rect 2728 1003 2734 1037
rect 2688 965 2734 1003
rect 2688 931 2694 965
rect 2728 931 2734 965
rect 2688 893 2734 931
rect 2688 859 2694 893
rect 2728 859 2734 893
rect 2688 821 2734 859
rect 2688 787 2694 821
rect 2728 787 2734 821
rect 2688 749 2734 787
rect 2688 715 2694 749
rect 2728 715 2734 749
rect 2688 677 2734 715
rect 2688 643 2694 677
rect 2728 643 2734 677
rect 2688 605 2734 643
rect 2688 571 2694 605
rect 2728 571 2734 605
rect 2688 533 2734 571
rect 2688 499 2694 533
rect 2728 499 2734 533
rect 2688 461 2734 499
rect 2688 427 2694 461
rect 2728 427 2734 461
rect 2688 389 2734 427
rect 2688 355 2694 389
rect 2728 355 2734 389
rect 2688 317 2734 355
rect 2688 283 2694 317
rect 2728 283 2734 317
rect 2688 268 2734 283
rect 2784 1253 2830 1268
rect 2784 1219 2790 1253
rect 2824 1219 2830 1253
rect 2784 1181 2830 1219
rect 2784 1147 2790 1181
rect 2824 1147 2830 1181
rect 2784 1109 2830 1147
rect 2784 1075 2790 1109
rect 2824 1075 2830 1109
rect 2784 1037 2830 1075
rect 2784 1003 2790 1037
rect 2824 1003 2830 1037
rect 2784 965 2830 1003
rect 2784 931 2790 965
rect 2824 931 2830 965
rect 2784 893 2830 931
rect 2784 859 2790 893
rect 2824 859 2830 893
rect 2784 821 2830 859
rect 2784 787 2790 821
rect 2824 787 2830 821
rect 2784 749 2830 787
rect 2784 715 2790 749
rect 2824 715 2830 749
rect 2784 677 2830 715
rect 2784 643 2790 677
rect 2824 643 2830 677
rect 2784 605 2830 643
rect 2784 571 2790 605
rect 2824 571 2830 605
rect 2784 533 2830 571
rect 2784 499 2790 533
rect 2824 499 2830 533
rect 2784 461 2830 499
rect 2784 427 2790 461
rect 2824 427 2830 461
rect 2784 389 2830 427
rect 2784 355 2790 389
rect 2824 355 2830 389
rect 2784 317 2830 355
rect 2784 283 2790 317
rect 2824 283 2830 317
rect 2784 268 2830 283
rect 2880 1253 2926 1268
rect 2880 1219 2886 1253
rect 2920 1219 2926 1253
rect 2880 1181 2926 1219
rect 2880 1147 2886 1181
rect 2920 1147 2926 1181
rect 2880 1109 2926 1147
rect 2880 1075 2886 1109
rect 2920 1075 2926 1109
rect 2880 1037 2926 1075
rect 2880 1003 2886 1037
rect 2920 1003 2926 1037
rect 2880 965 2926 1003
rect 2880 931 2886 965
rect 2920 931 2926 965
rect 2880 893 2926 931
rect 2880 859 2886 893
rect 2920 859 2926 893
rect 2880 821 2926 859
rect 2880 787 2886 821
rect 2920 787 2926 821
rect 2880 749 2926 787
rect 2880 715 2886 749
rect 2920 715 2926 749
rect 2880 677 2926 715
rect 2880 643 2886 677
rect 2920 643 2926 677
rect 2880 605 2926 643
rect 2880 571 2886 605
rect 2920 571 2926 605
rect 2880 533 2926 571
rect 2880 499 2886 533
rect 2920 499 2926 533
rect 2880 461 2926 499
rect 2880 427 2886 461
rect 2920 427 2926 461
rect 2880 389 2926 427
rect 2880 355 2886 389
rect 2920 355 2926 389
rect 2880 317 2926 355
rect 2880 283 2886 317
rect 2920 283 2926 317
rect 2880 268 2926 283
rect 2976 1253 3022 1268
rect 2976 1219 2982 1253
rect 3016 1219 3022 1253
rect 15416 1257 15462 1300
rect 2976 1181 3022 1219
rect 2976 1147 2982 1181
rect 3016 1147 3022 1181
rect 2976 1109 3022 1147
rect 2976 1075 2982 1109
rect 3016 1075 3022 1109
rect 2976 1037 3022 1075
rect 2976 1003 2982 1037
rect 3016 1003 3022 1037
rect 2976 965 3022 1003
rect 2976 931 2982 965
rect 3016 931 3022 965
rect 2976 893 3022 931
rect 2976 859 2982 893
rect 3016 859 3022 893
rect 2976 821 3022 859
rect 2976 787 2982 821
rect 3016 787 3022 821
rect 2976 749 3022 787
rect 2976 715 2982 749
rect 3016 715 3022 749
rect 2976 677 3022 715
rect 2976 643 2982 677
rect 3016 643 3022 677
rect 2976 605 3022 643
rect 2976 571 2982 605
rect 3016 571 3022 605
rect 2976 533 3022 571
rect 2976 499 2982 533
rect 3016 499 3022 533
rect 2976 461 3022 499
rect 2976 427 2982 461
rect 3016 427 3022 461
rect 2976 389 3022 427
rect 2976 355 2982 389
rect 3016 355 3022 389
rect 2976 317 3022 355
rect 2976 283 2982 317
rect 3016 283 3022 317
rect 2976 268 3022 283
rect 3108 1237 3154 1252
rect 3108 1203 3114 1237
rect 3148 1203 3154 1237
rect 3108 1165 3154 1203
rect 3108 1131 3114 1165
rect 3148 1131 3154 1165
rect 3108 1093 3154 1131
rect 3108 1059 3114 1093
rect 3148 1059 3154 1093
rect 3108 1021 3154 1059
rect 3108 987 3114 1021
rect 3148 987 3154 1021
rect 3108 949 3154 987
rect 3108 915 3114 949
rect 3148 915 3154 949
rect 3108 877 3154 915
rect 3108 843 3114 877
rect 3148 843 3154 877
rect 3108 805 3154 843
rect 3108 771 3114 805
rect 3148 771 3154 805
rect 3108 733 3154 771
rect 3108 699 3114 733
rect 3148 699 3154 733
rect 3108 661 3154 699
rect 3108 627 3114 661
rect 3148 627 3154 661
rect 3108 589 3154 627
rect 3108 555 3114 589
rect 3148 555 3154 589
rect 3108 517 3154 555
rect 3108 483 3114 517
rect 3148 483 3154 517
rect 3108 445 3154 483
rect 3108 411 3114 445
rect 3148 411 3154 445
rect 3108 373 3154 411
rect 3108 339 3114 373
rect 3148 339 3154 373
rect 3108 301 3154 339
rect 3108 267 3114 301
rect 3148 267 3154 301
rect 3108 252 3154 267
rect 3204 1237 3250 1252
rect 3204 1203 3210 1237
rect 3244 1203 3250 1237
rect 3204 1165 3250 1203
rect 3204 1131 3210 1165
rect 3244 1131 3250 1165
rect 3204 1093 3250 1131
rect 3204 1059 3210 1093
rect 3244 1059 3250 1093
rect 3204 1021 3250 1059
rect 3204 987 3210 1021
rect 3244 987 3250 1021
rect 3204 949 3250 987
rect 3204 915 3210 949
rect 3244 915 3250 949
rect 3204 877 3250 915
rect 3204 843 3210 877
rect 3244 843 3250 877
rect 3204 805 3250 843
rect 3204 771 3210 805
rect 3244 771 3250 805
rect 3204 733 3250 771
rect 3204 699 3210 733
rect 3244 699 3250 733
rect 3204 661 3250 699
rect 3204 627 3210 661
rect 3244 627 3250 661
rect 3204 589 3250 627
rect 3204 555 3210 589
rect 3244 555 3250 589
rect 3204 517 3250 555
rect 3204 483 3210 517
rect 3244 483 3250 517
rect 3204 445 3250 483
rect 3204 411 3210 445
rect 3244 411 3250 445
rect 3204 373 3250 411
rect 3204 339 3210 373
rect 3244 339 3250 373
rect 3204 301 3250 339
rect 3204 267 3210 301
rect 3244 267 3250 301
rect 3204 252 3250 267
rect 3300 1237 3346 1252
rect 3300 1203 3306 1237
rect 3340 1203 3346 1237
rect 3300 1165 3346 1203
rect 3300 1131 3306 1165
rect 3340 1131 3346 1165
rect 3300 1093 3346 1131
rect 3300 1059 3306 1093
rect 3340 1059 3346 1093
rect 3300 1021 3346 1059
rect 3300 987 3306 1021
rect 3340 987 3346 1021
rect 3300 949 3346 987
rect 3300 915 3306 949
rect 3340 915 3346 949
rect 3300 877 3346 915
rect 3300 843 3306 877
rect 3340 843 3346 877
rect 3300 805 3346 843
rect 3300 771 3306 805
rect 3340 771 3346 805
rect 3300 733 3346 771
rect 3300 699 3306 733
rect 3340 699 3346 733
rect 3300 661 3346 699
rect 3300 627 3306 661
rect 3340 627 3346 661
rect 3300 589 3346 627
rect 3300 555 3306 589
rect 3340 555 3346 589
rect 3300 517 3346 555
rect 3300 483 3306 517
rect 3340 483 3346 517
rect 3300 445 3346 483
rect 3300 411 3306 445
rect 3340 411 3346 445
rect 3300 373 3346 411
rect 3300 339 3306 373
rect 3340 339 3346 373
rect 3300 301 3346 339
rect 3300 267 3306 301
rect 3340 267 3346 301
rect 3300 252 3346 267
rect 3396 1237 3442 1252
rect 3396 1203 3402 1237
rect 3436 1203 3442 1237
rect 3396 1165 3442 1203
rect 3396 1131 3402 1165
rect 3436 1131 3442 1165
rect 3396 1093 3442 1131
rect 3396 1059 3402 1093
rect 3436 1059 3442 1093
rect 3396 1021 3442 1059
rect 3396 987 3402 1021
rect 3436 987 3442 1021
rect 3396 949 3442 987
rect 3396 915 3402 949
rect 3436 915 3442 949
rect 3396 877 3442 915
rect 3396 843 3402 877
rect 3436 843 3442 877
rect 3396 805 3442 843
rect 3396 771 3402 805
rect 3436 771 3442 805
rect 3396 733 3442 771
rect 3396 699 3402 733
rect 3436 699 3442 733
rect 3396 661 3442 699
rect 3396 627 3402 661
rect 3436 627 3442 661
rect 3396 589 3442 627
rect 3396 555 3402 589
rect 3436 555 3442 589
rect 3396 517 3442 555
rect 3396 483 3402 517
rect 3436 483 3442 517
rect 3396 445 3442 483
rect 3396 411 3402 445
rect 3436 411 3442 445
rect 3396 373 3442 411
rect 3396 339 3402 373
rect 3436 339 3442 373
rect 3396 301 3442 339
rect 3396 267 3402 301
rect 3436 267 3442 301
rect 3396 252 3442 267
rect 3492 1237 3538 1252
rect 3492 1203 3498 1237
rect 3532 1203 3538 1237
rect 3492 1165 3538 1203
rect 3492 1131 3498 1165
rect 3532 1131 3538 1165
rect 3492 1093 3538 1131
rect 3492 1059 3498 1093
rect 3532 1059 3538 1093
rect 3492 1021 3538 1059
rect 3492 987 3498 1021
rect 3532 987 3538 1021
rect 3492 949 3538 987
rect 3492 915 3498 949
rect 3532 915 3538 949
rect 3492 877 3538 915
rect 3492 843 3498 877
rect 3532 843 3538 877
rect 3492 805 3538 843
rect 3492 771 3498 805
rect 3532 771 3538 805
rect 3492 733 3538 771
rect 3492 699 3498 733
rect 3532 699 3538 733
rect 3492 661 3538 699
rect 3492 627 3498 661
rect 3532 627 3538 661
rect 3492 589 3538 627
rect 3492 555 3498 589
rect 3532 555 3538 589
rect 3492 517 3538 555
rect 3492 483 3498 517
rect 3532 483 3538 517
rect 3492 445 3538 483
rect 3492 411 3498 445
rect 3532 411 3538 445
rect 3492 373 3538 411
rect 3492 339 3498 373
rect 3532 339 3538 373
rect 3492 301 3538 339
rect 3492 267 3498 301
rect 3532 267 3538 301
rect 3492 252 3538 267
rect 3588 1237 3634 1252
rect 3588 1203 3594 1237
rect 3628 1203 3634 1237
rect 3588 1165 3634 1203
rect 3588 1131 3594 1165
rect 3628 1131 3634 1165
rect 3588 1093 3634 1131
rect 3588 1059 3594 1093
rect 3628 1059 3634 1093
rect 3588 1021 3634 1059
rect 3588 987 3594 1021
rect 3628 987 3634 1021
rect 3588 949 3634 987
rect 3588 915 3594 949
rect 3628 915 3634 949
rect 3588 877 3634 915
rect 3588 843 3594 877
rect 3628 843 3634 877
rect 3588 805 3634 843
rect 3588 771 3594 805
rect 3628 771 3634 805
rect 3588 733 3634 771
rect 3588 699 3594 733
rect 3628 699 3634 733
rect 3588 661 3634 699
rect 3588 627 3594 661
rect 3628 627 3634 661
rect 3588 589 3634 627
rect 3588 555 3594 589
rect 3628 555 3634 589
rect 3588 517 3634 555
rect 3588 483 3594 517
rect 3628 483 3634 517
rect 3588 445 3634 483
rect 3588 411 3594 445
rect 3628 411 3634 445
rect 3588 373 3634 411
rect 3588 339 3594 373
rect 3628 339 3634 373
rect 3588 301 3634 339
rect 3588 267 3594 301
rect 3628 267 3634 301
rect 3588 252 3634 267
rect 3684 1237 3730 1252
rect 3684 1203 3690 1237
rect 3724 1203 3730 1237
rect 3684 1165 3730 1203
rect 3684 1131 3690 1165
rect 3724 1131 3730 1165
rect 3684 1093 3730 1131
rect 3684 1059 3690 1093
rect 3724 1059 3730 1093
rect 3684 1021 3730 1059
rect 3684 987 3690 1021
rect 3724 987 3730 1021
rect 3684 949 3730 987
rect 3684 915 3690 949
rect 3724 915 3730 949
rect 3684 877 3730 915
rect 3684 843 3690 877
rect 3724 843 3730 877
rect 3684 805 3730 843
rect 3684 771 3690 805
rect 3724 771 3730 805
rect 3684 733 3730 771
rect 3684 699 3690 733
rect 3724 699 3730 733
rect 3684 661 3730 699
rect 3684 627 3690 661
rect 3724 627 3730 661
rect 3684 589 3730 627
rect 3684 555 3690 589
rect 3724 555 3730 589
rect 3684 517 3730 555
rect 3684 483 3690 517
rect 3724 483 3730 517
rect 3684 445 3730 483
rect 3684 411 3690 445
rect 3724 411 3730 445
rect 3684 373 3730 411
rect 3684 339 3690 373
rect 3724 339 3730 373
rect 3684 301 3730 339
rect 3684 267 3690 301
rect 3724 267 3730 301
rect 3684 252 3730 267
rect 3780 1237 3826 1252
rect 3780 1203 3786 1237
rect 3820 1203 3826 1237
rect 3780 1165 3826 1203
rect 3780 1131 3786 1165
rect 3820 1131 3826 1165
rect 3780 1093 3826 1131
rect 3780 1059 3786 1093
rect 3820 1059 3826 1093
rect 3780 1021 3826 1059
rect 3780 987 3786 1021
rect 3820 987 3826 1021
rect 3780 949 3826 987
rect 3780 915 3786 949
rect 3820 915 3826 949
rect 3780 877 3826 915
rect 3780 843 3786 877
rect 3820 843 3826 877
rect 3780 805 3826 843
rect 3780 771 3786 805
rect 3820 771 3826 805
rect 3780 733 3826 771
rect 3780 699 3786 733
rect 3820 699 3826 733
rect 3780 661 3826 699
rect 3780 627 3786 661
rect 3820 627 3826 661
rect 3780 589 3826 627
rect 3780 555 3786 589
rect 3820 555 3826 589
rect 3780 517 3826 555
rect 3780 483 3786 517
rect 3820 483 3826 517
rect 3780 445 3826 483
rect 3780 411 3786 445
rect 3820 411 3826 445
rect 3780 373 3826 411
rect 3780 339 3786 373
rect 3820 339 3826 373
rect 3780 301 3826 339
rect 3780 267 3786 301
rect 3820 267 3826 301
rect 3780 252 3826 267
rect 3876 1237 3922 1252
rect 3876 1203 3882 1237
rect 3916 1203 3922 1237
rect 3876 1165 3922 1203
rect 3876 1131 3882 1165
rect 3916 1131 3922 1165
rect 3876 1093 3922 1131
rect 3876 1059 3882 1093
rect 3916 1059 3922 1093
rect 3876 1021 3922 1059
rect 3876 987 3882 1021
rect 3916 987 3922 1021
rect 3876 949 3922 987
rect 3876 915 3882 949
rect 3916 915 3922 949
rect 3876 877 3922 915
rect 3876 843 3882 877
rect 3916 843 3922 877
rect 3876 805 3922 843
rect 3876 771 3882 805
rect 3916 771 3922 805
rect 3876 733 3922 771
rect 3876 699 3882 733
rect 3916 699 3922 733
rect 3876 661 3922 699
rect 3876 627 3882 661
rect 3916 627 3922 661
rect 3876 589 3922 627
rect 3876 555 3882 589
rect 3916 555 3922 589
rect 3876 517 3922 555
rect 3876 483 3882 517
rect 3916 483 3922 517
rect 3876 445 3922 483
rect 3876 411 3882 445
rect 3916 411 3922 445
rect 3876 373 3922 411
rect 3876 339 3882 373
rect 3916 339 3922 373
rect 3876 301 3922 339
rect 3876 267 3882 301
rect 3916 267 3922 301
rect 3876 252 3922 267
rect 3972 1237 4018 1252
rect 3972 1203 3978 1237
rect 4012 1203 4018 1237
rect 3972 1165 4018 1203
rect 3972 1131 3978 1165
rect 4012 1131 4018 1165
rect 3972 1093 4018 1131
rect 3972 1059 3978 1093
rect 4012 1059 4018 1093
rect 3972 1021 4018 1059
rect 3972 987 3978 1021
rect 4012 987 4018 1021
rect 3972 949 4018 987
rect 3972 915 3978 949
rect 4012 915 4018 949
rect 3972 877 4018 915
rect 3972 843 3978 877
rect 4012 843 4018 877
rect 3972 805 4018 843
rect 3972 771 3978 805
rect 4012 771 4018 805
rect 3972 733 4018 771
rect 3972 699 3978 733
rect 4012 699 4018 733
rect 3972 661 4018 699
rect 3972 627 3978 661
rect 4012 627 4018 661
rect 3972 589 4018 627
rect 3972 555 3978 589
rect 4012 555 4018 589
rect 3972 517 4018 555
rect 3972 483 3978 517
rect 4012 483 4018 517
rect 3972 445 4018 483
rect 3972 411 3978 445
rect 4012 411 4018 445
rect 3972 373 4018 411
rect 3972 339 3978 373
rect 4012 339 4018 373
rect 3972 301 4018 339
rect 3972 267 3978 301
rect 4012 267 4018 301
rect 3972 252 4018 267
rect 4068 1237 4114 1252
rect 4068 1203 4074 1237
rect 4108 1203 4114 1237
rect 4068 1165 4114 1203
rect 4068 1131 4074 1165
rect 4108 1131 4114 1165
rect 4068 1093 4114 1131
rect 4068 1059 4074 1093
rect 4108 1059 4114 1093
rect 4068 1021 4114 1059
rect 4068 987 4074 1021
rect 4108 987 4114 1021
rect 4068 949 4114 987
rect 4068 915 4074 949
rect 4108 915 4114 949
rect 4068 877 4114 915
rect 4068 843 4074 877
rect 4108 843 4114 877
rect 4068 805 4114 843
rect 4068 771 4074 805
rect 4108 771 4114 805
rect 4068 733 4114 771
rect 4068 699 4074 733
rect 4108 699 4114 733
rect 4068 661 4114 699
rect 4068 627 4074 661
rect 4108 627 4114 661
rect 4068 589 4114 627
rect 4068 555 4074 589
rect 4108 555 4114 589
rect 4068 517 4114 555
rect 4068 483 4074 517
rect 4108 483 4114 517
rect 4068 445 4114 483
rect 4068 411 4074 445
rect 4108 411 4114 445
rect 4068 373 4114 411
rect 4068 339 4074 373
rect 4108 339 4114 373
rect 4068 301 4114 339
rect 4068 267 4074 301
rect 4108 267 4114 301
rect 4068 252 4114 267
rect 4164 1237 4210 1252
rect 4164 1203 4170 1237
rect 4204 1203 4210 1237
rect 4164 1165 4210 1203
rect 4164 1131 4170 1165
rect 4204 1131 4210 1165
rect 4164 1093 4210 1131
rect 4164 1059 4170 1093
rect 4204 1059 4210 1093
rect 4164 1021 4210 1059
rect 4164 987 4170 1021
rect 4204 987 4210 1021
rect 4164 949 4210 987
rect 4164 915 4170 949
rect 4204 915 4210 949
rect 4164 877 4210 915
rect 4164 843 4170 877
rect 4204 843 4210 877
rect 4164 805 4210 843
rect 4164 771 4170 805
rect 4204 771 4210 805
rect 4164 733 4210 771
rect 4164 699 4170 733
rect 4204 699 4210 733
rect 4164 661 4210 699
rect 4164 627 4170 661
rect 4204 627 4210 661
rect 4164 589 4210 627
rect 4164 555 4170 589
rect 4204 555 4210 589
rect 4164 517 4210 555
rect 4164 483 4170 517
rect 4204 483 4210 517
rect 4164 445 4210 483
rect 4164 411 4170 445
rect 4204 411 4210 445
rect 4164 373 4210 411
rect 4164 339 4170 373
rect 4204 339 4210 373
rect 4164 301 4210 339
rect 4164 267 4170 301
rect 4204 267 4210 301
rect 4164 252 4210 267
rect 4260 1237 4306 1252
rect 4260 1203 4266 1237
rect 4300 1203 4306 1237
rect 4260 1165 4306 1203
rect 4260 1131 4266 1165
rect 4300 1131 4306 1165
rect 4260 1093 4306 1131
rect 4260 1059 4266 1093
rect 4300 1059 4306 1093
rect 4260 1021 4306 1059
rect 4260 987 4266 1021
rect 4300 987 4306 1021
rect 4260 949 4306 987
rect 4260 915 4266 949
rect 4300 915 4306 949
rect 4260 877 4306 915
rect 4260 843 4266 877
rect 4300 843 4306 877
rect 4260 805 4306 843
rect 4260 771 4266 805
rect 4300 771 4306 805
rect 4260 733 4306 771
rect 4260 699 4266 733
rect 4300 699 4306 733
rect 4260 661 4306 699
rect 4260 627 4266 661
rect 4300 627 4306 661
rect 4260 589 4306 627
rect 4260 555 4266 589
rect 4300 555 4306 589
rect 4260 517 4306 555
rect 4260 483 4266 517
rect 4300 483 4306 517
rect 4260 445 4306 483
rect 4260 411 4266 445
rect 4300 411 4306 445
rect 4260 373 4306 411
rect 4260 339 4266 373
rect 4300 339 4306 373
rect 4260 301 4306 339
rect 4260 267 4266 301
rect 4300 267 4306 301
rect 4260 252 4306 267
rect 4876 1237 4922 1252
rect 4876 1203 4882 1237
rect 4916 1203 4922 1237
rect 4876 1165 4922 1203
rect 4876 1131 4882 1165
rect 4916 1131 4922 1165
rect 4876 1093 4922 1131
rect 4876 1059 4882 1093
rect 4916 1059 4922 1093
rect 4876 1021 4922 1059
rect 4876 987 4882 1021
rect 4916 987 4922 1021
rect 4876 949 4922 987
rect 4876 915 4882 949
rect 4916 915 4922 949
rect 4876 877 4922 915
rect 4876 843 4882 877
rect 4916 843 4922 877
rect 4876 805 4922 843
rect 4876 771 4882 805
rect 4916 771 4922 805
rect 4876 733 4922 771
rect 4876 699 4882 733
rect 4916 699 4922 733
rect 4876 661 4922 699
rect 4876 627 4882 661
rect 4916 627 4922 661
rect 4876 589 4922 627
rect 4876 555 4882 589
rect 4916 555 4922 589
rect 4876 517 4922 555
rect 4876 483 4882 517
rect 4916 483 4922 517
rect 4876 445 4922 483
rect 4876 411 4882 445
rect 4916 411 4922 445
rect 4876 373 4922 411
rect 4876 339 4882 373
rect 4916 339 4922 373
rect 4876 301 4922 339
rect 4876 267 4882 301
rect 4916 267 4922 301
rect 4876 252 4922 267
rect 4972 1237 5018 1252
rect 4972 1203 4978 1237
rect 5012 1203 5018 1237
rect 4972 1165 5018 1203
rect 4972 1131 4978 1165
rect 5012 1131 5018 1165
rect 4972 1093 5018 1131
rect 4972 1059 4978 1093
rect 5012 1059 5018 1093
rect 4972 1021 5018 1059
rect 4972 987 4978 1021
rect 5012 987 5018 1021
rect 4972 949 5018 987
rect 4972 915 4978 949
rect 5012 915 5018 949
rect 4972 877 5018 915
rect 4972 843 4978 877
rect 5012 843 5018 877
rect 4972 805 5018 843
rect 4972 771 4978 805
rect 5012 771 5018 805
rect 4972 733 5018 771
rect 4972 699 4978 733
rect 5012 699 5018 733
rect 4972 661 5018 699
rect 4972 627 4978 661
rect 5012 627 5018 661
rect 4972 589 5018 627
rect 4972 555 4978 589
rect 5012 555 5018 589
rect 4972 517 5018 555
rect 4972 483 4978 517
rect 5012 483 5018 517
rect 4972 445 5018 483
rect 4972 411 4978 445
rect 5012 411 5018 445
rect 4972 373 5018 411
rect 4972 339 4978 373
rect 5012 339 5018 373
rect 4972 301 5018 339
rect 4972 267 4978 301
rect 5012 267 5018 301
rect 4972 252 5018 267
rect 5068 1237 5114 1252
rect 5068 1203 5074 1237
rect 5108 1203 5114 1237
rect 5068 1165 5114 1203
rect 5068 1131 5074 1165
rect 5108 1131 5114 1165
rect 5068 1093 5114 1131
rect 5068 1059 5074 1093
rect 5108 1059 5114 1093
rect 5068 1021 5114 1059
rect 5068 987 5074 1021
rect 5108 987 5114 1021
rect 5068 949 5114 987
rect 5068 915 5074 949
rect 5108 915 5114 949
rect 5068 877 5114 915
rect 5068 843 5074 877
rect 5108 843 5114 877
rect 5068 805 5114 843
rect 5068 771 5074 805
rect 5108 771 5114 805
rect 5068 733 5114 771
rect 5068 699 5074 733
rect 5108 699 5114 733
rect 5068 661 5114 699
rect 5068 627 5074 661
rect 5108 627 5114 661
rect 5068 589 5114 627
rect 5068 555 5074 589
rect 5108 555 5114 589
rect 5068 517 5114 555
rect 5068 483 5074 517
rect 5108 483 5114 517
rect 5068 445 5114 483
rect 5068 411 5074 445
rect 5108 411 5114 445
rect 5068 373 5114 411
rect 5068 339 5074 373
rect 5108 339 5114 373
rect 5068 301 5114 339
rect 5068 267 5074 301
rect 5108 267 5114 301
rect 5068 252 5114 267
rect 5164 1237 5210 1252
rect 5164 1203 5170 1237
rect 5204 1203 5210 1237
rect 5164 1165 5210 1203
rect 5164 1131 5170 1165
rect 5204 1131 5210 1165
rect 5164 1093 5210 1131
rect 5164 1059 5170 1093
rect 5204 1059 5210 1093
rect 5164 1021 5210 1059
rect 5164 987 5170 1021
rect 5204 987 5210 1021
rect 5164 949 5210 987
rect 5164 915 5170 949
rect 5204 915 5210 949
rect 5164 877 5210 915
rect 5164 843 5170 877
rect 5204 843 5210 877
rect 5164 805 5210 843
rect 5164 771 5170 805
rect 5204 771 5210 805
rect 5164 733 5210 771
rect 5164 699 5170 733
rect 5204 699 5210 733
rect 5164 661 5210 699
rect 5164 627 5170 661
rect 5204 627 5210 661
rect 5164 589 5210 627
rect 5164 555 5170 589
rect 5204 555 5210 589
rect 5164 517 5210 555
rect 5164 483 5170 517
rect 5204 483 5210 517
rect 5164 445 5210 483
rect 5164 411 5170 445
rect 5204 411 5210 445
rect 5164 373 5210 411
rect 5164 339 5170 373
rect 5204 339 5210 373
rect 5164 301 5210 339
rect 5164 267 5170 301
rect 5204 267 5210 301
rect 5164 252 5210 267
rect 5260 1237 5306 1252
rect 5260 1203 5266 1237
rect 5300 1203 5306 1237
rect 5260 1165 5306 1203
rect 5260 1131 5266 1165
rect 5300 1131 5306 1165
rect 5260 1093 5306 1131
rect 5260 1059 5266 1093
rect 5300 1059 5306 1093
rect 5260 1021 5306 1059
rect 5260 987 5266 1021
rect 5300 987 5306 1021
rect 5260 949 5306 987
rect 5260 915 5266 949
rect 5300 915 5306 949
rect 5260 877 5306 915
rect 5260 843 5266 877
rect 5300 843 5306 877
rect 5260 805 5306 843
rect 5260 771 5266 805
rect 5300 771 5306 805
rect 5260 733 5306 771
rect 5260 699 5266 733
rect 5300 699 5306 733
rect 5260 661 5306 699
rect 5260 627 5266 661
rect 5300 627 5306 661
rect 5260 589 5306 627
rect 5260 555 5266 589
rect 5300 555 5306 589
rect 5260 517 5306 555
rect 5260 483 5266 517
rect 5300 483 5306 517
rect 5260 445 5306 483
rect 5260 411 5266 445
rect 5300 411 5306 445
rect 5260 373 5306 411
rect 5260 339 5266 373
rect 5300 339 5306 373
rect 5260 301 5306 339
rect 5260 267 5266 301
rect 5300 267 5306 301
rect 5260 252 5306 267
rect 5356 1237 5402 1252
rect 5356 1203 5362 1237
rect 5396 1203 5402 1237
rect 5356 1165 5402 1203
rect 5356 1131 5362 1165
rect 5396 1131 5402 1165
rect 5356 1093 5402 1131
rect 5356 1059 5362 1093
rect 5396 1059 5402 1093
rect 5356 1021 5402 1059
rect 5356 987 5362 1021
rect 5396 987 5402 1021
rect 5356 949 5402 987
rect 5356 915 5362 949
rect 5396 915 5402 949
rect 5356 877 5402 915
rect 5356 843 5362 877
rect 5396 843 5402 877
rect 5356 805 5402 843
rect 5356 771 5362 805
rect 5396 771 5402 805
rect 5356 733 5402 771
rect 5356 699 5362 733
rect 5396 699 5402 733
rect 5356 661 5402 699
rect 5356 627 5362 661
rect 5396 627 5402 661
rect 5356 589 5402 627
rect 5356 555 5362 589
rect 5396 555 5402 589
rect 5356 517 5402 555
rect 5356 483 5362 517
rect 5396 483 5402 517
rect 5356 445 5402 483
rect 5356 411 5362 445
rect 5396 411 5402 445
rect 5356 373 5402 411
rect 5356 339 5362 373
rect 5396 339 5402 373
rect 5356 301 5402 339
rect 5356 267 5362 301
rect 5396 267 5402 301
rect 5356 252 5402 267
rect 5452 1237 5498 1252
rect 5452 1203 5458 1237
rect 5492 1203 5498 1237
rect 5452 1165 5498 1203
rect 5452 1131 5458 1165
rect 5492 1131 5498 1165
rect 5452 1093 5498 1131
rect 5452 1059 5458 1093
rect 5492 1059 5498 1093
rect 5452 1021 5498 1059
rect 5452 987 5458 1021
rect 5492 987 5498 1021
rect 5452 949 5498 987
rect 5452 915 5458 949
rect 5492 915 5498 949
rect 5452 877 5498 915
rect 5452 843 5458 877
rect 5492 843 5498 877
rect 5452 805 5498 843
rect 5452 771 5458 805
rect 5492 771 5498 805
rect 5452 733 5498 771
rect 5452 699 5458 733
rect 5492 699 5498 733
rect 5452 661 5498 699
rect 5452 627 5458 661
rect 5492 627 5498 661
rect 5452 589 5498 627
rect 5452 555 5458 589
rect 5492 555 5498 589
rect 5452 517 5498 555
rect 5452 483 5458 517
rect 5492 483 5498 517
rect 5452 445 5498 483
rect 5452 411 5458 445
rect 5492 411 5498 445
rect 5452 373 5498 411
rect 5452 339 5458 373
rect 5492 339 5498 373
rect 5452 301 5498 339
rect 5452 267 5458 301
rect 5492 267 5498 301
rect 5452 252 5498 267
rect 5548 1237 5594 1252
rect 5548 1203 5554 1237
rect 5588 1203 5594 1237
rect 5548 1165 5594 1203
rect 5548 1131 5554 1165
rect 5588 1131 5594 1165
rect 5548 1093 5594 1131
rect 5548 1059 5554 1093
rect 5588 1059 5594 1093
rect 5548 1021 5594 1059
rect 5548 987 5554 1021
rect 5588 987 5594 1021
rect 5548 949 5594 987
rect 5548 915 5554 949
rect 5588 915 5594 949
rect 5548 877 5594 915
rect 5548 843 5554 877
rect 5588 843 5594 877
rect 5548 805 5594 843
rect 5548 771 5554 805
rect 5588 771 5594 805
rect 5548 733 5594 771
rect 5548 699 5554 733
rect 5588 699 5594 733
rect 5548 661 5594 699
rect 5548 627 5554 661
rect 5588 627 5594 661
rect 5548 589 5594 627
rect 5548 555 5554 589
rect 5588 555 5594 589
rect 5548 517 5594 555
rect 5548 483 5554 517
rect 5588 483 5594 517
rect 5548 445 5594 483
rect 5548 411 5554 445
rect 5588 411 5594 445
rect 5548 373 5594 411
rect 5548 339 5554 373
rect 5588 339 5594 373
rect 5548 301 5594 339
rect 5548 267 5554 301
rect 5588 267 5594 301
rect 5548 252 5594 267
rect 5644 1237 5690 1252
rect 5644 1203 5650 1237
rect 5684 1203 5690 1237
rect 5644 1165 5690 1203
rect 5644 1131 5650 1165
rect 5684 1131 5690 1165
rect 5644 1093 5690 1131
rect 5644 1059 5650 1093
rect 5684 1059 5690 1093
rect 5644 1021 5690 1059
rect 5644 987 5650 1021
rect 5684 987 5690 1021
rect 5644 949 5690 987
rect 5644 915 5650 949
rect 5684 915 5690 949
rect 5644 877 5690 915
rect 5644 843 5650 877
rect 5684 843 5690 877
rect 5644 805 5690 843
rect 5644 771 5650 805
rect 5684 771 5690 805
rect 5644 733 5690 771
rect 5644 699 5650 733
rect 5684 699 5690 733
rect 5644 661 5690 699
rect 5644 627 5650 661
rect 5684 627 5690 661
rect 5644 589 5690 627
rect 5644 555 5650 589
rect 5684 555 5690 589
rect 5644 517 5690 555
rect 5644 483 5650 517
rect 5684 483 5690 517
rect 5644 445 5690 483
rect 5644 411 5650 445
rect 5684 411 5690 445
rect 5644 373 5690 411
rect 5644 339 5650 373
rect 5684 339 5690 373
rect 5644 301 5690 339
rect 5644 267 5650 301
rect 5684 267 5690 301
rect 5644 252 5690 267
rect 5740 1237 5786 1252
rect 5740 1203 5746 1237
rect 5780 1203 5786 1237
rect 5740 1165 5786 1203
rect 5740 1131 5746 1165
rect 5780 1131 5786 1165
rect 5740 1093 5786 1131
rect 5740 1059 5746 1093
rect 5780 1059 5786 1093
rect 5740 1021 5786 1059
rect 5740 987 5746 1021
rect 5780 987 5786 1021
rect 5740 949 5786 987
rect 5740 915 5746 949
rect 5780 915 5786 949
rect 5740 877 5786 915
rect 5740 843 5746 877
rect 5780 843 5786 877
rect 5740 805 5786 843
rect 5740 771 5746 805
rect 5780 771 5786 805
rect 5740 733 5786 771
rect 5740 699 5746 733
rect 5780 699 5786 733
rect 5740 661 5786 699
rect 5740 627 5746 661
rect 5780 627 5786 661
rect 5740 589 5786 627
rect 5740 555 5746 589
rect 5780 555 5786 589
rect 5740 517 5786 555
rect 5740 483 5746 517
rect 5780 483 5786 517
rect 5740 445 5786 483
rect 5740 411 5746 445
rect 5780 411 5786 445
rect 5740 373 5786 411
rect 5740 339 5746 373
rect 5780 339 5786 373
rect 5740 301 5786 339
rect 5740 267 5746 301
rect 5780 267 5786 301
rect 5740 252 5786 267
rect 5836 1237 5882 1252
rect 5836 1203 5842 1237
rect 5876 1203 5882 1237
rect 5836 1165 5882 1203
rect 5836 1131 5842 1165
rect 5876 1131 5882 1165
rect 5836 1093 5882 1131
rect 5836 1059 5842 1093
rect 5876 1059 5882 1093
rect 5836 1021 5882 1059
rect 5836 987 5842 1021
rect 5876 987 5882 1021
rect 5836 949 5882 987
rect 5836 915 5842 949
rect 5876 915 5882 949
rect 5836 877 5882 915
rect 5836 843 5842 877
rect 5876 843 5882 877
rect 5836 805 5882 843
rect 5836 771 5842 805
rect 5876 771 5882 805
rect 5836 733 5882 771
rect 5836 699 5842 733
rect 5876 699 5882 733
rect 5836 661 5882 699
rect 5836 627 5842 661
rect 5876 627 5882 661
rect 5836 589 5882 627
rect 5836 555 5842 589
rect 5876 555 5882 589
rect 5836 517 5882 555
rect 5836 483 5842 517
rect 5876 483 5882 517
rect 5836 445 5882 483
rect 5836 411 5842 445
rect 5876 411 5882 445
rect 5836 373 5882 411
rect 5836 339 5842 373
rect 5876 339 5882 373
rect 5836 301 5882 339
rect 5836 267 5842 301
rect 5876 267 5882 301
rect 5836 252 5882 267
rect 5932 1237 5978 1252
rect 5932 1203 5938 1237
rect 5972 1203 5978 1237
rect 5932 1165 5978 1203
rect 5932 1131 5938 1165
rect 5972 1131 5978 1165
rect 5932 1093 5978 1131
rect 5932 1059 5938 1093
rect 5972 1059 5978 1093
rect 5932 1021 5978 1059
rect 5932 987 5938 1021
rect 5972 987 5978 1021
rect 5932 949 5978 987
rect 5932 915 5938 949
rect 5972 915 5978 949
rect 5932 877 5978 915
rect 5932 843 5938 877
rect 5972 843 5978 877
rect 5932 805 5978 843
rect 5932 771 5938 805
rect 5972 771 5978 805
rect 5932 733 5978 771
rect 5932 699 5938 733
rect 5972 699 5978 733
rect 5932 661 5978 699
rect 5932 627 5938 661
rect 5972 627 5978 661
rect 5932 589 5978 627
rect 5932 555 5938 589
rect 5972 555 5978 589
rect 5932 517 5978 555
rect 5932 483 5938 517
rect 5972 483 5978 517
rect 5932 445 5978 483
rect 5932 411 5938 445
rect 5972 411 5978 445
rect 5932 373 5978 411
rect 5932 339 5938 373
rect 5972 339 5978 373
rect 5932 301 5978 339
rect 5932 267 5938 301
rect 5972 267 5978 301
rect 5932 252 5978 267
rect 6138 1237 6184 1252
rect 6138 1203 6144 1237
rect 6178 1203 6184 1237
rect 6138 1165 6184 1203
rect 6138 1131 6144 1165
rect 6178 1131 6184 1165
rect 6138 1093 6184 1131
rect 6138 1059 6144 1093
rect 6178 1059 6184 1093
rect 6138 1021 6184 1059
rect 6138 987 6144 1021
rect 6178 987 6184 1021
rect 6138 949 6184 987
rect 6138 915 6144 949
rect 6178 915 6184 949
rect 6138 877 6184 915
rect 6138 843 6144 877
rect 6178 843 6184 877
rect 6138 805 6184 843
rect 6138 771 6144 805
rect 6178 771 6184 805
rect 6138 733 6184 771
rect 6138 699 6144 733
rect 6178 699 6184 733
rect 6138 661 6184 699
rect 6138 627 6144 661
rect 6178 627 6184 661
rect 6138 589 6184 627
rect 6138 555 6144 589
rect 6178 555 6184 589
rect 6138 517 6184 555
rect 6138 483 6144 517
rect 6178 483 6184 517
rect 6138 445 6184 483
rect 6138 411 6144 445
rect 6178 411 6184 445
rect 6138 373 6184 411
rect 6138 339 6144 373
rect 6178 339 6184 373
rect 6138 301 6184 339
rect 6138 267 6144 301
rect 6178 267 6184 301
rect 6138 252 6184 267
rect 6234 1237 6280 1252
rect 6234 1203 6240 1237
rect 6274 1203 6280 1237
rect 6234 1165 6280 1203
rect 6234 1131 6240 1165
rect 6274 1131 6280 1165
rect 6234 1093 6280 1131
rect 6234 1059 6240 1093
rect 6274 1059 6280 1093
rect 6234 1021 6280 1059
rect 6234 987 6240 1021
rect 6274 987 6280 1021
rect 6234 949 6280 987
rect 6234 915 6240 949
rect 6274 915 6280 949
rect 6234 877 6280 915
rect 6234 843 6240 877
rect 6274 843 6280 877
rect 6234 805 6280 843
rect 6234 771 6240 805
rect 6274 771 6280 805
rect 6234 733 6280 771
rect 6234 699 6240 733
rect 6274 699 6280 733
rect 6234 661 6280 699
rect 6234 627 6240 661
rect 6274 627 6280 661
rect 6234 589 6280 627
rect 6234 555 6240 589
rect 6274 555 6280 589
rect 6234 517 6280 555
rect 6234 483 6240 517
rect 6274 483 6280 517
rect 6234 445 6280 483
rect 6234 411 6240 445
rect 6274 411 6280 445
rect 6234 373 6280 411
rect 6234 339 6240 373
rect 6274 339 6280 373
rect 6234 301 6280 339
rect 6234 267 6240 301
rect 6274 267 6280 301
rect 6234 252 6280 267
rect 6330 1237 6376 1252
rect 6330 1203 6336 1237
rect 6370 1203 6376 1237
rect 6330 1165 6376 1203
rect 6330 1131 6336 1165
rect 6370 1131 6376 1165
rect 6330 1093 6376 1131
rect 6330 1059 6336 1093
rect 6370 1059 6376 1093
rect 6330 1021 6376 1059
rect 6330 987 6336 1021
rect 6370 987 6376 1021
rect 6330 949 6376 987
rect 6330 915 6336 949
rect 6370 915 6376 949
rect 6330 877 6376 915
rect 6330 843 6336 877
rect 6370 843 6376 877
rect 6330 805 6376 843
rect 6330 771 6336 805
rect 6370 771 6376 805
rect 6330 733 6376 771
rect 6330 699 6336 733
rect 6370 699 6376 733
rect 6330 661 6376 699
rect 6330 627 6336 661
rect 6370 627 6376 661
rect 6330 589 6376 627
rect 6330 555 6336 589
rect 6370 555 6376 589
rect 6330 517 6376 555
rect 6330 483 6336 517
rect 6370 483 6376 517
rect 6330 445 6376 483
rect 6330 411 6336 445
rect 6370 411 6376 445
rect 6330 373 6376 411
rect 6330 339 6336 373
rect 6370 339 6376 373
rect 6330 301 6376 339
rect 6330 267 6336 301
rect 6370 267 6376 301
rect 6330 252 6376 267
rect 6426 1237 6472 1252
rect 6426 1203 6432 1237
rect 6466 1203 6472 1237
rect 6426 1165 6472 1203
rect 6426 1131 6432 1165
rect 6466 1131 6472 1165
rect 6426 1093 6472 1131
rect 6426 1059 6432 1093
rect 6466 1059 6472 1093
rect 6426 1021 6472 1059
rect 6426 987 6432 1021
rect 6466 987 6472 1021
rect 6426 949 6472 987
rect 6426 915 6432 949
rect 6466 915 6472 949
rect 6426 877 6472 915
rect 6426 843 6432 877
rect 6466 843 6472 877
rect 6426 805 6472 843
rect 6426 771 6432 805
rect 6466 771 6472 805
rect 6426 733 6472 771
rect 6426 699 6432 733
rect 6466 699 6472 733
rect 6426 661 6472 699
rect 6426 627 6432 661
rect 6466 627 6472 661
rect 6426 589 6472 627
rect 6426 555 6432 589
rect 6466 555 6472 589
rect 6426 517 6472 555
rect 6426 483 6432 517
rect 6466 483 6472 517
rect 6426 445 6472 483
rect 6426 411 6432 445
rect 6466 411 6472 445
rect 6426 373 6472 411
rect 6426 339 6432 373
rect 6466 339 6472 373
rect 6426 301 6472 339
rect 6426 267 6432 301
rect 6466 267 6472 301
rect 6426 252 6472 267
rect 6522 1237 6568 1252
rect 6522 1203 6528 1237
rect 6562 1203 6568 1237
rect 6522 1165 6568 1203
rect 6522 1131 6528 1165
rect 6562 1131 6568 1165
rect 6522 1093 6568 1131
rect 6522 1059 6528 1093
rect 6562 1059 6568 1093
rect 6522 1021 6568 1059
rect 6522 987 6528 1021
rect 6562 987 6568 1021
rect 6522 949 6568 987
rect 6522 915 6528 949
rect 6562 915 6568 949
rect 6522 877 6568 915
rect 6522 843 6528 877
rect 6562 843 6568 877
rect 6522 805 6568 843
rect 6522 771 6528 805
rect 6562 771 6568 805
rect 6522 733 6568 771
rect 6522 699 6528 733
rect 6562 699 6568 733
rect 6522 661 6568 699
rect 6522 627 6528 661
rect 6562 627 6568 661
rect 6522 589 6568 627
rect 6522 555 6528 589
rect 6562 555 6568 589
rect 6522 517 6568 555
rect 6522 483 6528 517
rect 6562 483 6568 517
rect 6522 445 6568 483
rect 6522 411 6528 445
rect 6562 411 6568 445
rect 6522 373 6568 411
rect 6522 339 6528 373
rect 6562 339 6568 373
rect 6522 301 6568 339
rect 6522 267 6528 301
rect 6562 267 6568 301
rect 6522 252 6568 267
rect 6618 1237 6664 1252
rect 6618 1203 6624 1237
rect 6658 1203 6664 1237
rect 6618 1165 6664 1203
rect 6618 1131 6624 1165
rect 6658 1131 6664 1165
rect 6618 1093 6664 1131
rect 6618 1059 6624 1093
rect 6658 1059 6664 1093
rect 6618 1021 6664 1059
rect 6618 987 6624 1021
rect 6658 987 6664 1021
rect 6618 949 6664 987
rect 6618 915 6624 949
rect 6658 915 6664 949
rect 6618 877 6664 915
rect 6618 843 6624 877
rect 6658 843 6664 877
rect 6618 805 6664 843
rect 6618 771 6624 805
rect 6658 771 6664 805
rect 6618 733 6664 771
rect 6618 699 6624 733
rect 6658 699 6664 733
rect 6618 661 6664 699
rect 6618 627 6624 661
rect 6658 627 6664 661
rect 6618 589 6664 627
rect 6618 555 6624 589
rect 6658 555 6664 589
rect 6618 517 6664 555
rect 6618 483 6624 517
rect 6658 483 6664 517
rect 6618 445 6664 483
rect 6618 411 6624 445
rect 6658 411 6664 445
rect 6618 373 6664 411
rect 6618 339 6624 373
rect 6658 339 6664 373
rect 6618 301 6664 339
rect 6618 267 6624 301
rect 6658 267 6664 301
rect 6618 252 6664 267
rect 6714 1237 6760 1252
rect 6714 1203 6720 1237
rect 6754 1203 6760 1237
rect 6714 1165 6760 1203
rect 6714 1131 6720 1165
rect 6754 1131 6760 1165
rect 6714 1093 6760 1131
rect 6714 1059 6720 1093
rect 6754 1059 6760 1093
rect 6714 1021 6760 1059
rect 6714 987 6720 1021
rect 6754 987 6760 1021
rect 6714 949 6760 987
rect 6714 915 6720 949
rect 6754 915 6760 949
rect 6714 877 6760 915
rect 6714 843 6720 877
rect 6754 843 6760 877
rect 6714 805 6760 843
rect 6714 771 6720 805
rect 6754 771 6760 805
rect 6714 733 6760 771
rect 6714 699 6720 733
rect 6754 699 6760 733
rect 6714 661 6760 699
rect 6714 627 6720 661
rect 6754 627 6760 661
rect 6714 589 6760 627
rect 6714 555 6720 589
rect 6754 555 6760 589
rect 6714 517 6760 555
rect 6714 483 6720 517
rect 6754 483 6760 517
rect 6714 445 6760 483
rect 6714 411 6720 445
rect 6754 411 6760 445
rect 6714 373 6760 411
rect 6714 339 6720 373
rect 6754 339 6760 373
rect 6714 301 6760 339
rect 6714 267 6720 301
rect 6754 267 6760 301
rect 6714 252 6760 267
rect 6810 1237 6856 1252
rect 6810 1203 6816 1237
rect 6850 1203 6856 1237
rect 6810 1165 6856 1203
rect 6810 1131 6816 1165
rect 6850 1131 6856 1165
rect 6810 1093 6856 1131
rect 6810 1059 6816 1093
rect 6850 1059 6856 1093
rect 6810 1021 6856 1059
rect 6810 987 6816 1021
rect 6850 987 6856 1021
rect 6810 949 6856 987
rect 6810 915 6816 949
rect 6850 915 6856 949
rect 6810 877 6856 915
rect 6810 843 6816 877
rect 6850 843 6856 877
rect 6810 805 6856 843
rect 6810 771 6816 805
rect 6850 771 6856 805
rect 6810 733 6856 771
rect 6810 699 6816 733
rect 6850 699 6856 733
rect 6810 661 6856 699
rect 6810 627 6816 661
rect 6850 627 6856 661
rect 6810 589 6856 627
rect 6810 555 6816 589
rect 6850 555 6856 589
rect 6810 517 6856 555
rect 6810 483 6816 517
rect 6850 483 6856 517
rect 6810 445 6856 483
rect 6810 411 6816 445
rect 6850 411 6856 445
rect 6810 373 6856 411
rect 6810 339 6816 373
rect 6850 339 6856 373
rect 6810 301 6856 339
rect 6810 267 6816 301
rect 6850 267 6856 301
rect 6810 252 6856 267
rect 6906 1237 6952 1252
rect 6906 1203 6912 1237
rect 6946 1203 6952 1237
rect 6906 1165 6952 1203
rect 6906 1131 6912 1165
rect 6946 1131 6952 1165
rect 6906 1093 6952 1131
rect 6906 1059 6912 1093
rect 6946 1059 6952 1093
rect 6906 1021 6952 1059
rect 6906 987 6912 1021
rect 6946 987 6952 1021
rect 6906 949 6952 987
rect 6906 915 6912 949
rect 6946 915 6952 949
rect 6906 877 6952 915
rect 6906 843 6912 877
rect 6946 843 6952 877
rect 6906 805 6952 843
rect 6906 771 6912 805
rect 6946 771 6952 805
rect 6906 733 6952 771
rect 6906 699 6912 733
rect 6946 699 6952 733
rect 6906 661 6952 699
rect 6906 627 6912 661
rect 6946 627 6952 661
rect 6906 589 6952 627
rect 6906 555 6912 589
rect 6946 555 6952 589
rect 6906 517 6952 555
rect 6906 483 6912 517
rect 6946 483 6952 517
rect 6906 445 6952 483
rect 6906 411 6912 445
rect 6946 411 6952 445
rect 6906 373 6952 411
rect 6906 339 6912 373
rect 6946 339 6952 373
rect 6906 301 6952 339
rect 6906 267 6912 301
rect 6946 267 6952 301
rect 6906 252 6952 267
rect 7002 1237 7048 1252
rect 7002 1203 7008 1237
rect 7042 1203 7048 1237
rect 7002 1165 7048 1203
rect 7002 1131 7008 1165
rect 7042 1131 7048 1165
rect 7002 1093 7048 1131
rect 7002 1059 7008 1093
rect 7042 1059 7048 1093
rect 7002 1021 7048 1059
rect 7002 987 7008 1021
rect 7042 987 7048 1021
rect 7002 949 7048 987
rect 7002 915 7008 949
rect 7042 915 7048 949
rect 7002 877 7048 915
rect 7002 843 7008 877
rect 7042 843 7048 877
rect 7002 805 7048 843
rect 7002 771 7008 805
rect 7042 771 7048 805
rect 7002 733 7048 771
rect 7002 699 7008 733
rect 7042 699 7048 733
rect 7002 661 7048 699
rect 7002 627 7008 661
rect 7042 627 7048 661
rect 7002 589 7048 627
rect 7002 555 7008 589
rect 7042 555 7048 589
rect 7002 517 7048 555
rect 7002 483 7008 517
rect 7042 483 7048 517
rect 7002 445 7048 483
rect 7002 411 7008 445
rect 7042 411 7048 445
rect 7002 373 7048 411
rect 7002 339 7008 373
rect 7042 339 7048 373
rect 7002 301 7048 339
rect 7002 267 7008 301
rect 7042 267 7048 301
rect 7002 252 7048 267
rect 7098 1237 7144 1252
rect 7098 1203 7104 1237
rect 7138 1203 7144 1237
rect 7098 1165 7144 1203
rect 7098 1131 7104 1165
rect 7138 1131 7144 1165
rect 7098 1093 7144 1131
rect 7098 1059 7104 1093
rect 7138 1059 7144 1093
rect 7098 1021 7144 1059
rect 7098 987 7104 1021
rect 7138 987 7144 1021
rect 7098 949 7144 987
rect 7098 915 7104 949
rect 7138 915 7144 949
rect 7098 877 7144 915
rect 7098 843 7104 877
rect 7138 843 7144 877
rect 7098 805 7144 843
rect 7098 771 7104 805
rect 7138 771 7144 805
rect 7098 733 7144 771
rect 7098 699 7104 733
rect 7138 699 7144 733
rect 7098 661 7144 699
rect 7098 627 7104 661
rect 7138 627 7144 661
rect 7098 589 7144 627
rect 7098 555 7104 589
rect 7138 555 7144 589
rect 7098 517 7144 555
rect 7098 483 7104 517
rect 7138 483 7144 517
rect 7098 445 7144 483
rect 7098 411 7104 445
rect 7138 411 7144 445
rect 7098 373 7144 411
rect 7098 339 7104 373
rect 7138 339 7144 373
rect 7098 301 7144 339
rect 7098 267 7104 301
rect 7138 267 7144 301
rect 7098 252 7144 267
rect 7194 1237 7240 1252
rect 7194 1203 7200 1237
rect 7234 1203 7240 1237
rect 7194 1165 7240 1203
rect 7194 1131 7200 1165
rect 7234 1131 7240 1165
rect 7194 1093 7240 1131
rect 7194 1059 7200 1093
rect 7234 1059 7240 1093
rect 7194 1021 7240 1059
rect 7194 987 7200 1021
rect 7234 987 7240 1021
rect 7194 949 7240 987
rect 7194 915 7200 949
rect 7234 915 7240 949
rect 7194 877 7240 915
rect 7194 843 7200 877
rect 7234 843 7240 877
rect 7194 805 7240 843
rect 7194 771 7200 805
rect 7234 771 7240 805
rect 7194 733 7240 771
rect 7194 699 7200 733
rect 7234 699 7240 733
rect 7194 661 7240 699
rect 7194 627 7200 661
rect 7234 627 7240 661
rect 7194 589 7240 627
rect 7194 555 7200 589
rect 7234 555 7240 589
rect 7194 517 7240 555
rect 7194 483 7200 517
rect 7234 483 7240 517
rect 7194 445 7240 483
rect 7194 411 7200 445
rect 7234 411 7240 445
rect 7194 373 7240 411
rect 7194 339 7200 373
rect 7234 339 7240 373
rect 7194 301 7240 339
rect 7194 267 7200 301
rect 7234 267 7240 301
rect 7194 252 7240 267
rect 7290 1237 7336 1252
rect 7290 1203 7296 1237
rect 7330 1203 7336 1237
rect 7290 1165 7336 1203
rect 7290 1131 7296 1165
rect 7330 1131 7336 1165
rect 7290 1093 7336 1131
rect 7290 1059 7296 1093
rect 7330 1059 7336 1093
rect 7290 1021 7336 1059
rect 7290 987 7296 1021
rect 7330 987 7336 1021
rect 7290 949 7336 987
rect 7290 915 7296 949
rect 7330 915 7336 949
rect 7290 877 7336 915
rect 7290 843 7296 877
rect 7330 843 7336 877
rect 7290 805 7336 843
rect 7290 771 7296 805
rect 7330 771 7336 805
rect 7290 733 7336 771
rect 7290 699 7296 733
rect 7330 699 7336 733
rect 7290 661 7336 699
rect 7290 627 7296 661
rect 7330 627 7336 661
rect 7290 589 7336 627
rect 7290 555 7296 589
rect 7330 555 7336 589
rect 7290 517 7336 555
rect 7290 483 7296 517
rect 7330 483 7336 517
rect 7290 445 7336 483
rect 7290 411 7296 445
rect 7330 411 7336 445
rect 7290 373 7336 411
rect 7290 339 7296 373
rect 7330 339 7336 373
rect 7290 301 7336 339
rect 7290 267 7296 301
rect 7330 267 7336 301
rect 7290 252 7336 267
rect 7906 1237 7952 1252
rect 7906 1203 7912 1237
rect 7946 1203 7952 1237
rect 7906 1165 7952 1203
rect 7906 1131 7912 1165
rect 7946 1131 7952 1165
rect 7906 1093 7952 1131
rect 7906 1059 7912 1093
rect 7946 1059 7952 1093
rect 7906 1021 7952 1059
rect 7906 987 7912 1021
rect 7946 987 7952 1021
rect 7906 949 7952 987
rect 7906 915 7912 949
rect 7946 915 7952 949
rect 7906 877 7952 915
rect 7906 843 7912 877
rect 7946 843 7952 877
rect 7906 805 7952 843
rect 7906 771 7912 805
rect 7946 771 7952 805
rect 7906 733 7952 771
rect 7906 699 7912 733
rect 7946 699 7952 733
rect 7906 661 7952 699
rect 7906 627 7912 661
rect 7946 627 7952 661
rect 7906 589 7952 627
rect 7906 555 7912 589
rect 7946 555 7952 589
rect 7906 517 7952 555
rect 7906 483 7912 517
rect 7946 483 7952 517
rect 7906 445 7952 483
rect 7906 411 7912 445
rect 7946 411 7952 445
rect 7906 373 7952 411
rect 7906 339 7912 373
rect 7946 339 7952 373
rect 7906 301 7952 339
rect 7906 267 7912 301
rect 7946 267 7952 301
rect 7906 252 7952 267
rect 8002 1237 8048 1252
rect 8002 1203 8008 1237
rect 8042 1203 8048 1237
rect 8002 1165 8048 1203
rect 8002 1131 8008 1165
rect 8042 1131 8048 1165
rect 8002 1093 8048 1131
rect 8002 1059 8008 1093
rect 8042 1059 8048 1093
rect 8002 1021 8048 1059
rect 8002 987 8008 1021
rect 8042 987 8048 1021
rect 8002 949 8048 987
rect 8002 915 8008 949
rect 8042 915 8048 949
rect 8002 877 8048 915
rect 8002 843 8008 877
rect 8042 843 8048 877
rect 8002 805 8048 843
rect 8002 771 8008 805
rect 8042 771 8048 805
rect 8002 733 8048 771
rect 8002 699 8008 733
rect 8042 699 8048 733
rect 8002 661 8048 699
rect 8002 627 8008 661
rect 8042 627 8048 661
rect 8002 589 8048 627
rect 8002 555 8008 589
rect 8042 555 8048 589
rect 8002 517 8048 555
rect 8002 483 8008 517
rect 8042 483 8048 517
rect 8002 445 8048 483
rect 8002 411 8008 445
rect 8042 411 8048 445
rect 8002 373 8048 411
rect 8002 339 8008 373
rect 8042 339 8048 373
rect 8002 301 8048 339
rect 8002 267 8008 301
rect 8042 267 8048 301
rect 8002 252 8048 267
rect 8098 1237 8144 1252
rect 8098 1203 8104 1237
rect 8138 1203 8144 1237
rect 8098 1165 8144 1203
rect 8098 1131 8104 1165
rect 8138 1131 8144 1165
rect 8098 1093 8144 1131
rect 8098 1059 8104 1093
rect 8138 1059 8144 1093
rect 8098 1021 8144 1059
rect 8098 987 8104 1021
rect 8138 987 8144 1021
rect 8098 949 8144 987
rect 8098 915 8104 949
rect 8138 915 8144 949
rect 8098 877 8144 915
rect 8098 843 8104 877
rect 8138 843 8144 877
rect 8098 805 8144 843
rect 8098 771 8104 805
rect 8138 771 8144 805
rect 8098 733 8144 771
rect 8098 699 8104 733
rect 8138 699 8144 733
rect 8098 661 8144 699
rect 8098 627 8104 661
rect 8138 627 8144 661
rect 8098 589 8144 627
rect 8098 555 8104 589
rect 8138 555 8144 589
rect 8098 517 8144 555
rect 8098 483 8104 517
rect 8138 483 8144 517
rect 8098 445 8144 483
rect 8098 411 8104 445
rect 8138 411 8144 445
rect 8098 373 8144 411
rect 8098 339 8104 373
rect 8138 339 8144 373
rect 8098 301 8144 339
rect 8098 267 8104 301
rect 8138 267 8144 301
rect 8098 252 8144 267
rect 8194 1237 8240 1252
rect 8194 1203 8200 1237
rect 8234 1203 8240 1237
rect 8194 1165 8240 1203
rect 8194 1131 8200 1165
rect 8234 1131 8240 1165
rect 8194 1093 8240 1131
rect 8194 1059 8200 1093
rect 8234 1059 8240 1093
rect 8194 1021 8240 1059
rect 8194 987 8200 1021
rect 8234 987 8240 1021
rect 8194 949 8240 987
rect 8194 915 8200 949
rect 8234 915 8240 949
rect 8194 877 8240 915
rect 8194 843 8200 877
rect 8234 843 8240 877
rect 8194 805 8240 843
rect 8194 771 8200 805
rect 8234 771 8240 805
rect 8194 733 8240 771
rect 8194 699 8200 733
rect 8234 699 8240 733
rect 8194 661 8240 699
rect 8194 627 8200 661
rect 8234 627 8240 661
rect 8194 589 8240 627
rect 8194 555 8200 589
rect 8234 555 8240 589
rect 8194 517 8240 555
rect 8194 483 8200 517
rect 8234 483 8240 517
rect 8194 445 8240 483
rect 8194 411 8200 445
rect 8234 411 8240 445
rect 8194 373 8240 411
rect 8194 339 8200 373
rect 8234 339 8240 373
rect 8194 301 8240 339
rect 8194 267 8200 301
rect 8234 267 8240 301
rect 8194 252 8240 267
rect 8290 1237 8336 1252
rect 8290 1203 8296 1237
rect 8330 1203 8336 1237
rect 8290 1165 8336 1203
rect 8290 1131 8296 1165
rect 8330 1131 8336 1165
rect 8290 1093 8336 1131
rect 8290 1059 8296 1093
rect 8330 1059 8336 1093
rect 8290 1021 8336 1059
rect 8290 987 8296 1021
rect 8330 987 8336 1021
rect 8290 949 8336 987
rect 8290 915 8296 949
rect 8330 915 8336 949
rect 8290 877 8336 915
rect 8290 843 8296 877
rect 8330 843 8336 877
rect 8290 805 8336 843
rect 8290 771 8296 805
rect 8330 771 8336 805
rect 8290 733 8336 771
rect 8290 699 8296 733
rect 8330 699 8336 733
rect 8290 661 8336 699
rect 8290 627 8296 661
rect 8330 627 8336 661
rect 8290 589 8336 627
rect 8290 555 8296 589
rect 8330 555 8336 589
rect 8290 517 8336 555
rect 8290 483 8296 517
rect 8330 483 8336 517
rect 8290 445 8336 483
rect 8290 411 8296 445
rect 8330 411 8336 445
rect 8290 373 8336 411
rect 8290 339 8296 373
rect 8330 339 8336 373
rect 8290 301 8336 339
rect 8290 267 8296 301
rect 8330 267 8336 301
rect 8290 252 8336 267
rect 8386 1237 8432 1252
rect 8386 1203 8392 1237
rect 8426 1203 8432 1237
rect 8386 1165 8432 1203
rect 8386 1131 8392 1165
rect 8426 1131 8432 1165
rect 8386 1093 8432 1131
rect 8386 1059 8392 1093
rect 8426 1059 8432 1093
rect 8386 1021 8432 1059
rect 8386 987 8392 1021
rect 8426 987 8432 1021
rect 8386 949 8432 987
rect 8386 915 8392 949
rect 8426 915 8432 949
rect 8386 877 8432 915
rect 8386 843 8392 877
rect 8426 843 8432 877
rect 8386 805 8432 843
rect 8386 771 8392 805
rect 8426 771 8432 805
rect 8386 733 8432 771
rect 8386 699 8392 733
rect 8426 699 8432 733
rect 8386 661 8432 699
rect 8386 627 8392 661
rect 8426 627 8432 661
rect 8386 589 8432 627
rect 8386 555 8392 589
rect 8426 555 8432 589
rect 8386 517 8432 555
rect 8386 483 8392 517
rect 8426 483 8432 517
rect 8386 445 8432 483
rect 8386 411 8392 445
rect 8426 411 8432 445
rect 8386 373 8432 411
rect 8386 339 8392 373
rect 8426 339 8432 373
rect 8386 301 8432 339
rect 8386 267 8392 301
rect 8426 267 8432 301
rect 8386 252 8432 267
rect 8482 1237 8528 1252
rect 8482 1203 8488 1237
rect 8522 1203 8528 1237
rect 8482 1165 8528 1203
rect 8482 1131 8488 1165
rect 8522 1131 8528 1165
rect 8482 1093 8528 1131
rect 8482 1059 8488 1093
rect 8522 1059 8528 1093
rect 8482 1021 8528 1059
rect 8482 987 8488 1021
rect 8522 987 8528 1021
rect 8482 949 8528 987
rect 8482 915 8488 949
rect 8522 915 8528 949
rect 8482 877 8528 915
rect 8482 843 8488 877
rect 8522 843 8528 877
rect 8482 805 8528 843
rect 8482 771 8488 805
rect 8522 771 8528 805
rect 8482 733 8528 771
rect 8482 699 8488 733
rect 8522 699 8528 733
rect 8482 661 8528 699
rect 8482 627 8488 661
rect 8522 627 8528 661
rect 8482 589 8528 627
rect 8482 555 8488 589
rect 8522 555 8528 589
rect 8482 517 8528 555
rect 8482 483 8488 517
rect 8522 483 8528 517
rect 8482 445 8528 483
rect 8482 411 8488 445
rect 8522 411 8528 445
rect 8482 373 8528 411
rect 8482 339 8488 373
rect 8522 339 8528 373
rect 8482 301 8528 339
rect 8482 267 8488 301
rect 8522 267 8528 301
rect 8482 252 8528 267
rect 8578 1237 8624 1252
rect 8578 1203 8584 1237
rect 8618 1203 8624 1237
rect 8578 1165 8624 1203
rect 8578 1131 8584 1165
rect 8618 1131 8624 1165
rect 8578 1093 8624 1131
rect 8578 1059 8584 1093
rect 8618 1059 8624 1093
rect 8578 1021 8624 1059
rect 8578 987 8584 1021
rect 8618 987 8624 1021
rect 8578 949 8624 987
rect 8578 915 8584 949
rect 8618 915 8624 949
rect 8578 877 8624 915
rect 8578 843 8584 877
rect 8618 843 8624 877
rect 8578 805 8624 843
rect 8578 771 8584 805
rect 8618 771 8624 805
rect 8578 733 8624 771
rect 8578 699 8584 733
rect 8618 699 8624 733
rect 8578 661 8624 699
rect 8578 627 8584 661
rect 8618 627 8624 661
rect 8578 589 8624 627
rect 8578 555 8584 589
rect 8618 555 8624 589
rect 8578 517 8624 555
rect 8578 483 8584 517
rect 8618 483 8624 517
rect 8578 445 8624 483
rect 8578 411 8584 445
rect 8618 411 8624 445
rect 8578 373 8624 411
rect 8578 339 8584 373
rect 8618 339 8624 373
rect 8578 301 8624 339
rect 8578 267 8584 301
rect 8618 267 8624 301
rect 8578 252 8624 267
rect 8674 1237 8720 1252
rect 8674 1203 8680 1237
rect 8714 1203 8720 1237
rect 8674 1165 8720 1203
rect 8674 1131 8680 1165
rect 8714 1131 8720 1165
rect 8674 1093 8720 1131
rect 8674 1059 8680 1093
rect 8714 1059 8720 1093
rect 8674 1021 8720 1059
rect 8674 987 8680 1021
rect 8714 987 8720 1021
rect 8674 949 8720 987
rect 8674 915 8680 949
rect 8714 915 8720 949
rect 8674 877 8720 915
rect 8674 843 8680 877
rect 8714 843 8720 877
rect 8674 805 8720 843
rect 8674 771 8680 805
rect 8714 771 8720 805
rect 8674 733 8720 771
rect 8674 699 8680 733
rect 8714 699 8720 733
rect 8674 661 8720 699
rect 8674 627 8680 661
rect 8714 627 8720 661
rect 8674 589 8720 627
rect 8674 555 8680 589
rect 8714 555 8720 589
rect 8674 517 8720 555
rect 8674 483 8680 517
rect 8714 483 8720 517
rect 8674 445 8720 483
rect 8674 411 8680 445
rect 8714 411 8720 445
rect 8674 373 8720 411
rect 8674 339 8680 373
rect 8714 339 8720 373
rect 8674 301 8720 339
rect 8674 267 8680 301
rect 8714 267 8720 301
rect 8674 252 8720 267
rect 8770 1237 8816 1252
rect 8770 1203 8776 1237
rect 8810 1203 8816 1237
rect 8770 1165 8816 1203
rect 8770 1131 8776 1165
rect 8810 1131 8816 1165
rect 8770 1093 8816 1131
rect 8770 1059 8776 1093
rect 8810 1059 8816 1093
rect 8770 1021 8816 1059
rect 8770 987 8776 1021
rect 8810 987 8816 1021
rect 8770 949 8816 987
rect 8770 915 8776 949
rect 8810 915 8816 949
rect 8770 877 8816 915
rect 8770 843 8776 877
rect 8810 843 8816 877
rect 8770 805 8816 843
rect 8770 771 8776 805
rect 8810 771 8816 805
rect 8770 733 8816 771
rect 8770 699 8776 733
rect 8810 699 8816 733
rect 8770 661 8816 699
rect 8770 627 8776 661
rect 8810 627 8816 661
rect 8770 589 8816 627
rect 8770 555 8776 589
rect 8810 555 8816 589
rect 8770 517 8816 555
rect 8770 483 8776 517
rect 8810 483 8816 517
rect 8770 445 8816 483
rect 8770 411 8776 445
rect 8810 411 8816 445
rect 8770 373 8816 411
rect 8770 339 8776 373
rect 8810 339 8816 373
rect 8770 301 8816 339
rect 8770 267 8776 301
rect 8810 267 8816 301
rect 8770 252 8816 267
rect 8866 1237 8912 1252
rect 8866 1203 8872 1237
rect 8906 1203 8912 1237
rect 8866 1165 8912 1203
rect 8866 1131 8872 1165
rect 8906 1131 8912 1165
rect 8866 1093 8912 1131
rect 8866 1059 8872 1093
rect 8906 1059 8912 1093
rect 8866 1021 8912 1059
rect 8866 987 8872 1021
rect 8906 987 8912 1021
rect 8866 949 8912 987
rect 8866 915 8872 949
rect 8906 915 8912 949
rect 8866 877 8912 915
rect 8866 843 8872 877
rect 8906 843 8912 877
rect 8866 805 8912 843
rect 8866 771 8872 805
rect 8906 771 8912 805
rect 8866 733 8912 771
rect 8866 699 8872 733
rect 8906 699 8912 733
rect 8866 661 8912 699
rect 8866 627 8872 661
rect 8906 627 8912 661
rect 8866 589 8912 627
rect 8866 555 8872 589
rect 8906 555 8912 589
rect 8866 517 8912 555
rect 8866 483 8872 517
rect 8906 483 8912 517
rect 8866 445 8912 483
rect 8866 411 8872 445
rect 8906 411 8912 445
rect 8866 373 8912 411
rect 8866 339 8872 373
rect 8906 339 8912 373
rect 8866 301 8912 339
rect 8866 267 8872 301
rect 8906 267 8912 301
rect 8866 252 8912 267
rect 8962 1237 9008 1252
rect 8962 1203 8968 1237
rect 9002 1203 9008 1237
rect 8962 1165 9008 1203
rect 8962 1131 8968 1165
rect 9002 1131 9008 1165
rect 8962 1093 9008 1131
rect 8962 1059 8968 1093
rect 9002 1059 9008 1093
rect 8962 1021 9008 1059
rect 8962 987 8968 1021
rect 9002 987 9008 1021
rect 8962 949 9008 987
rect 8962 915 8968 949
rect 9002 915 9008 949
rect 8962 877 9008 915
rect 8962 843 8968 877
rect 9002 843 9008 877
rect 8962 805 9008 843
rect 8962 771 8968 805
rect 9002 771 9008 805
rect 8962 733 9008 771
rect 8962 699 8968 733
rect 9002 699 9008 733
rect 8962 661 9008 699
rect 8962 627 8968 661
rect 9002 627 9008 661
rect 8962 589 9008 627
rect 8962 555 8968 589
rect 9002 555 9008 589
rect 8962 517 9008 555
rect 8962 483 8968 517
rect 9002 483 9008 517
rect 8962 445 9008 483
rect 8962 411 8968 445
rect 9002 411 9008 445
rect 8962 373 9008 411
rect 8962 339 8968 373
rect 9002 339 9008 373
rect 8962 301 9008 339
rect 8962 267 8968 301
rect 9002 267 9008 301
rect 8962 252 9008 267
rect 9226 1235 9272 1250
rect 9226 1201 9232 1235
rect 9266 1201 9272 1235
rect 9226 1163 9272 1201
rect 9226 1129 9232 1163
rect 9266 1129 9272 1163
rect 9226 1091 9272 1129
rect 9226 1057 9232 1091
rect 9266 1057 9272 1091
rect 9226 1019 9272 1057
rect 9226 985 9232 1019
rect 9266 985 9272 1019
rect 9226 947 9272 985
rect 9226 913 9232 947
rect 9266 913 9272 947
rect 9226 875 9272 913
rect 9226 841 9232 875
rect 9266 841 9272 875
rect 9226 803 9272 841
rect 9226 769 9232 803
rect 9266 769 9272 803
rect 9226 731 9272 769
rect 9226 697 9232 731
rect 9266 697 9272 731
rect 9226 659 9272 697
rect 9226 625 9232 659
rect 9266 625 9272 659
rect 9226 587 9272 625
rect 9226 553 9232 587
rect 9266 553 9272 587
rect 9226 515 9272 553
rect 9226 481 9232 515
rect 9266 481 9272 515
rect 9226 443 9272 481
rect 9226 409 9232 443
rect 9266 409 9272 443
rect 9226 371 9272 409
rect 9226 337 9232 371
rect 9266 337 9272 371
rect 9226 299 9272 337
rect 9226 265 9232 299
rect 9266 265 9272 299
rect 9226 250 9272 265
rect 9322 1235 9368 1250
rect 9322 1201 9328 1235
rect 9362 1201 9368 1235
rect 9322 1163 9368 1201
rect 9322 1129 9328 1163
rect 9362 1129 9368 1163
rect 9322 1091 9368 1129
rect 9322 1057 9328 1091
rect 9362 1057 9368 1091
rect 9322 1019 9368 1057
rect 9322 985 9328 1019
rect 9362 985 9368 1019
rect 9322 947 9368 985
rect 9322 913 9328 947
rect 9362 913 9368 947
rect 9322 875 9368 913
rect 9322 841 9328 875
rect 9362 841 9368 875
rect 9322 803 9368 841
rect 9322 769 9328 803
rect 9362 769 9368 803
rect 9322 731 9368 769
rect 9322 697 9328 731
rect 9362 697 9368 731
rect 9322 659 9368 697
rect 9322 625 9328 659
rect 9362 625 9368 659
rect 9322 587 9368 625
rect 9322 553 9328 587
rect 9362 553 9368 587
rect 9322 515 9368 553
rect 9322 481 9328 515
rect 9362 481 9368 515
rect 9322 443 9368 481
rect 9322 409 9328 443
rect 9362 409 9368 443
rect 9322 371 9368 409
rect 9322 337 9328 371
rect 9362 337 9368 371
rect 9322 299 9368 337
rect 9322 265 9328 299
rect 9362 265 9368 299
rect 9322 250 9368 265
rect 9418 1235 9464 1250
rect 9418 1201 9424 1235
rect 9458 1201 9464 1235
rect 9418 1163 9464 1201
rect 9418 1129 9424 1163
rect 9458 1129 9464 1163
rect 9418 1091 9464 1129
rect 9418 1057 9424 1091
rect 9458 1057 9464 1091
rect 9418 1019 9464 1057
rect 9418 985 9424 1019
rect 9458 985 9464 1019
rect 9418 947 9464 985
rect 9418 913 9424 947
rect 9458 913 9464 947
rect 9418 875 9464 913
rect 9418 841 9424 875
rect 9458 841 9464 875
rect 9418 803 9464 841
rect 9418 769 9424 803
rect 9458 769 9464 803
rect 9418 731 9464 769
rect 9418 697 9424 731
rect 9458 697 9464 731
rect 9418 659 9464 697
rect 9418 625 9424 659
rect 9458 625 9464 659
rect 9418 587 9464 625
rect 9418 553 9424 587
rect 9458 553 9464 587
rect 9418 515 9464 553
rect 9418 481 9424 515
rect 9458 481 9464 515
rect 9418 443 9464 481
rect 9418 409 9424 443
rect 9458 409 9464 443
rect 9418 371 9464 409
rect 9418 337 9424 371
rect 9458 337 9464 371
rect 9418 299 9464 337
rect 9418 265 9424 299
rect 9458 265 9464 299
rect 9418 250 9464 265
rect 9514 1235 9560 1250
rect 9514 1201 9520 1235
rect 9554 1201 9560 1235
rect 9514 1163 9560 1201
rect 9514 1129 9520 1163
rect 9554 1129 9560 1163
rect 9514 1091 9560 1129
rect 9514 1057 9520 1091
rect 9554 1057 9560 1091
rect 9514 1019 9560 1057
rect 9514 985 9520 1019
rect 9554 985 9560 1019
rect 9514 947 9560 985
rect 9514 913 9520 947
rect 9554 913 9560 947
rect 9514 875 9560 913
rect 9514 841 9520 875
rect 9554 841 9560 875
rect 9514 803 9560 841
rect 9514 769 9520 803
rect 9554 769 9560 803
rect 9514 731 9560 769
rect 9514 697 9520 731
rect 9554 697 9560 731
rect 9514 659 9560 697
rect 9514 625 9520 659
rect 9554 625 9560 659
rect 9514 587 9560 625
rect 9514 553 9520 587
rect 9554 553 9560 587
rect 9514 515 9560 553
rect 9514 481 9520 515
rect 9554 481 9560 515
rect 9514 443 9560 481
rect 9514 409 9520 443
rect 9554 409 9560 443
rect 9514 371 9560 409
rect 9514 337 9520 371
rect 9554 337 9560 371
rect 9514 299 9560 337
rect 9514 265 9520 299
rect 9554 265 9560 299
rect 9514 250 9560 265
rect 9610 1235 9656 1250
rect 9610 1201 9616 1235
rect 9650 1201 9656 1235
rect 9610 1163 9656 1201
rect 9610 1129 9616 1163
rect 9650 1129 9656 1163
rect 9610 1091 9656 1129
rect 9610 1057 9616 1091
rect 9650 1057 9656 1091
rect 9610 1019 9656 1057
rect 9610 985 9616 1019
rect 9650 985 9656 1019
rect 9610 947 9656 985
rect 9610 913 9616 947
rect 9650 913 9656 947
rect 9610 875 9656 913
rect 9610 841 9616 875
rect 9650 841 9656 875
rect 9610 803 9656 841
rect 9610 769 9616 803
rect 9650 769 9656 803
rect 9610 731 9656 769
rect 9610 697 9616 731
rect 9650 697 9656 731
rect 9610 659 9656 697
rect 9610 625 9616 659
rect 9650 625 9656 659
rect 9610 587 9656 625
rect 9610 553 9616 587
rect 9650 553 9656 587
rect 9610 515 9656 553
rect 9610 481 9616 515
rect 9650 481 9656 515
rect 9610 443 9656 481
rect 9610 409 9616 443
rect 9650 409 9656 443
rect 9610 371 9656 409
rect 9610 337 9616 371
rect 9650 337 9656 371
rect 9610 299 9656 337
rect 9610 265 9616 299
rect 9650 265 9656 299
rect 9610 250 9656 265
rect 9706 1235 9752 1250
rect 9706 1201 9712 1235
rect 9746 1201 9752 1235
rect 9706 1163 9752 1201
rect 9706 1129 9712 1163
rect 9746 1129 9752 1163
rect 9706 1091 9752 1129
rect 9706 1057 9712 1091
rect 9746 1057 9752 1091
rect 9706 1019 9752 1057
rect 9706 985 9712 1019
rect 9746 985 9752 1019
rect 9706 947 9752 985
rect 9706 913 9712 947
rect 9746 913 9752 947
rect 9706 875 9752 913
rect 9706 841 9712 875
rect 9746 841 9752 875
rect 9706 803 9752 841
rect 9706 769 9712 803
rect 9746 769 9752 803
rect 9706 731 9752 769
rect 9706 697 9712 731
rect 9746 697 9752 731
rect 9706 659 9752 697
rect 9706 625 9712 659
rect 9746 625 9752 659
rect 9706 587 9752 625
rect 9706 553 9712 587
rect 9746 553 9752 587
rect 9706 515 9752 553
rect 9706 481 9712 515
rect 9746 481 9752 515
rect 9706 443 9752 481
rect 9706 409 9712 443
rect 9746 409 9752 443
rect 9706 371 9752 409
rect 9706 337 9712 371
rect 9746 337 9752 371
rect 9706 299 9752 337
rect 9706 265 9712 299
rect 9746 265 9752 299
rect 9706 250 9752 265
rect 9802 1235 9848 1250
rect 9802 1201 9808 1235
rect 9842 1201 9848 1235
rect 9802 1163 9848 1201
rect 9802 1129 9808 1163
rect 9842 1129 9848 1163
rect 9802 1091 9848 1129
rect 9802 1057 9808 1091
rect 9842 1057 9848 1091
rect 9802 1019 9848 1057
rect 9802 985 9808 1019
rect 9842 985 9848 1019
rect 9802 947 9848 985
rect 9802 913 9808 947
rect 9842 913 9848 947
rect 9802 875 9848 913
rect 9802 841 9808 875
rect 9842 841 9848 875
rect 9802 803 9848 841
rect 9802 769 9808 803
rect 9842 769 9848 803
rect 9802 731 9848 769
rect 9802 697 9808 731
rect 9842 697 9848 731
rect 9802 659 9848 697
rect 9802 625 9808 659
rect 9842 625 9848 659
rect 9802 587 9848 625
rect 9802 553 9808 587
rect 9842 553 9848 587
rect 9802 515 9848 553
rect 9802 481 9808 515
rect 9842 481 9848 515
rect 9802 443 9848 481
rect 9802 409 9808 443
rect 9842 409 9848 443
rect 9802 371 9848 409
rect 9802 337 9808 371
rect 9842 337 9848 371
rect 9802 299 9848 337
rect 9802 265 9808 299
rect 9842 265 9848 299
rect 9802 250 9848 265
rect 9898 1235 9944 1250
rect 9898 1201 9904 1235
rect 9938 1201 9944 1235
rect 9898 1163 9944 1201
rect 9898 1129 9904 1163
rect 9938 1129 9944 1163
rect 9898 1091 9944 1129
rect 9898 1057 9904 1091
rect 9938 1057 9944 1091
rect 9898 1019 9944 1057
rect 9898 985 9904 1019
rect 9938 985 9944 1019
rect 9898 947 9944 985
rect 9898 913 9904 947
rect 9938 913 9944 947
rect 9898 875 9944 913
rect 9898 841 9904 875
rect 9938 841 9944 875
rect 9898 803 9944 841
rect 9898 769 9904 803
rect 9938 769 9944 803
rect 9898 731 9944 769
rect 9898 697 9904 731
rect 9938 697 9944 731
rect 9898 659 9944 697
rect 9898 625 9904 659
rect 9938 625 9944 659
rect 9898 587 9944 625
rect 9898 553 9904 587
rect 9938 553 9944 587
rect 9898 515 9944 553
rect 9898 481 9904 515
rect 9938 481 9944 515
rect 9898 443 9944 481
rect 9898 409 9904 443
rect 9938 409 9944 443
rect 9898 371 9944 409
rect 9898 337 9904 371
rect 9938 337 9944 371
rect 9898 299 9944 337
rect 9898 265 9904 299
rect 9938 265 9944 299
rect 9898 250 9944 265
rect 9994 1235 10040 1250
rect 9994 1201 10000 1235
rect 10034 1201 10040 1235
rect 9994 1163 10040 1201
rect 9994 1129 10000 1163
rect 10034 1129 10040 1163
rect 9994 1091 10040 1129
rect 9994 1057 10000 1091
rect 10034 1057 10040 1091
rect 9994 1019 10040 1057
rect 9994 985 10000 1019
rect 10034 985 10040 1019
rect 9994 947 10040 985
rect 9994 913 10000 947
rect 10034 913 10040 947
rect 9994 875 10040 913
rect 9994 841 10000 875
rect 10034 841 10040 875
rect 9994 803 10040 841
rect 9994 769 10000 803
rect 10034 769 10040 803
rect 9994 731 10040 769
rect 9994 697 10000 731
rect 10034 697 10040 731
rect 9994 659 10040 697
rect 9994 625 10000 659
rect 10034 625 10040 659
rect 9994 587 10040 625
rect 9994 553 10000 587
rect 10034 553 10040 587
rect 9994 515 10040 553
rect 9994 481 10000 515
rect 10034 481 10040 515
rect 9994 443 10040 481
rect 9994 409 10000 443
rect 10034 409 10040 443
rect 9994 371 10040 409
rect 9994 337 10000 371
rect 10034 337 10040 371
rect 9994 299 10040 337
rect 9994 265 10000 299
rect 10034 265 10040 299
rect 9994 250 10040 265
rect 10090 1235 10136 1250
rect 10090 1201 10096 1235
rect 10130 1201 10136 1235
rect 10090 1163 10136 1201
rect 10090 1129 10096 1163
rect 10130 1129 10136 1163
rect 10090 1091 10136 1129
rect 10090 1057 10096 1091
rect 10130 1057 10136 1091
rect 10090 1019 10136 1057
rect 10090 985 10096 1019
rect 10130 985 10136 1019
rect 10090 947 10136 985
rect 10090 913 10096 947
rect 10130 913 10136 947
rect 10090 875 10136 913
rect 10090 841 10096 875
rect 10130 841 10136 875
rect 10090 803 10136 841
rect 10090 769 10096 803
rect 10130 769 10136 803
rect 10090 731 10136 769
rect 10090 697 10096 731
rect 10130 697 10136 731
rect 10090 659 10136 697
rect 10090 625 10096 659
rect 10130 625 10136 659
rect 10090 587 10136 625
rect 10090 553 10096 587
rect 10130 553 10136 587
rect 10090 515 10136 553
rect 10090 481 10096 515
rect 10130 481 10136 515
rect 10090 443 10136 481
rect 10090 409 10096 443
rect 10130 409 10136 443
rect 10090 371 10136 409
rect 10090 337 10096 371
rect 10130 337 10136 371
rect 10090 299 10136 337
rect 10090 265 10096 299
rect 10130 265 10136 299
rect 10090 250 10136 265
rect 10186 1235 10232 1250
rect 10186 1201 10192 1235
rect 10226 1201 10232 1235
rect 10186 1163 10232 1201
rect 10186 1129 10192 1163
rect 10226 1129 10232 1163
rect 10186 1091 10232 1129
rect 10186 1057 10192 1091
rect 10226 1057 10232 1091
rect 10186 1019 10232 1057
rect 10186 985 10192 1019
rect 10226 985 10232 1019
rect 10186 947 10232 985
rect 10186 913 10192 947
rect 10226 913 10232 947
rect 10186 875 10232 913
rect 10186 841 10192 875
rect 10226 841 10232 875
rect 10186 803 10232 841
rect 10186 769 10192 803
rect 10226 769 10232 803
rect 10186 731 10232 769
rect 10186 697 10192 731
rect 10226 697 10232 731
rect 10186 659 10232 697
rect 10186 625 10192 659
rect 10226 625 10232 659
rect 10186 587 10232 625
rect 10186 553 10192 587
rect 10226 553 10232 587
rect 10186 515 10232 553
rect 10186 481 10192 515
rect 10226 481 10232 515
rect 10186 443 10232 481
rect 10186 409 10192 443
rect 10226 409 10232 443
rect 10186 371 10232 409
rect 10186 337 10192 371
rect 10226 337 10232 371
rect 10186 299 10232 337
rect 10186 265 10192 299
rect 10226 265 10232 299
rect 10186 250 10232 265
rect 10282 1235 10328 1250
rect 10282 1201 10288 1235
rect 10322 1201 10328 1235
rect 10282 1163 10328 1201
rect 10282 1129 10288 1163
rect 10322 1129 10328 1163
rect 10282 1091 10328 1129
rect 10282 1057 10288 1091
rect 10322 1057 10328 1091
rect 10282 1019 10328 1057
rect 10282 985 10288 1019
rect 10322 985 10328 1019
rect 10282 947 10328 985
rect 10282 913 10288 947
rect 10322 913 10328 947
rect 10282 875 10328 913
rect 10282 841 10288 875
rect 10322 841 10328 875
rect 10282 803 10328 841
rect 10282 769 10288 803
rect 10322 769 10328 803
rect 10282 731 10328 769
rect 10282 697 10288 731
rect 10322 697 10328 731
rect 10282 659 10328 697
rect 10282 625 10288 659
rect 10322 625 10328 659
rect 10282 587 10328 625
rect 10282 553 10288 587
rect 10322 553 10328 587
rect 10282 515 10328 553
rect 10282 481 10288 515
rect 10322 481 10328 515
rect 10282 443 10328 481
rect 10282 409 10288 443
rect 10322 409 10328 443
rect 10282 371 10328 409
rect 10282 337 10288 371
rect 10322 337 10328 371
rect 10282 299 10328 337
rect 10282 265 10288 299
rect 10322 265 10328 299
rect 10282 250 10328 265
rect 10378 1235 10424 1250
rect 10378 1201 10384 1235
rect 10418 1201 10424 1235
rect 10378 1163 10424 1201
rect 10378 1129 10384 1163
rect 10418 1129 10424 1163
rect 10378 1091 10424 1129
rect 10378 1057 10384 1091
rect 10418 1057 10424 1091
rect 10378 1019 10424 1057
rect 10378 985 10384 1019
rect 10418 985 10424 1019
rect 10378 947 10424 985
rect 10378 913 10384 947
rect 10418 913 10424 947
rect 10378 875 10424 913
rect 10378 841 10384 875
rect 10418 841 10424 875
rect 10378 803 10424 841
rect 10378 769 10384 803
rect 10418 769 10424 803
rect 10378 731 10424 769
rect 10378 697 10384 731
rect 10418 697 10424 731
rect 10378 659 10424 697
rect 10378 625 10384 659
rect 10418 625 10424 659
rect 10378 587 10424 625
rect 10378 553 10384 587
rect 10418 553 10424 587
rect 10378 515 10424 553
rect 10378 481 10384 515
rect 10418 481 10424 515
rect 10378 443 10424 481
rect 10378 409 10384 443
rect 10418 409 10424 443
rect 10378 371 10424 409
rect 10378 337 10384 371
rect 10418 337 10424 371
rect 10378 299 10424 337
rect 10378 265 10384 299
rect 10418 265 10424 299
rect 10378 250 10424 265
rect 10994 1235 11040 1250
rect 10994 1201 11000 1235
rect 11034 1201 11040 1235
rect 10994 1163 11040 1201
rect 10994 1129 11000 1163
rect 11034 1129 11040 1163
rect 10994 1091 11040 1129
rect 10994 1057 11000 1091
rect 11034 1057 11040 1091
rect 10994 1019 11040 1057
rect 10994 985 11000 1019
rect 11034 985 11040 1019
rect 10994 947 11040 985
rect 10994 913 11000 947
rect 11034 913 11040 947
rect 10994 875 11040 913
rect 10994 841 11000 875
rect 11034 841 11040 875
rect 10994 803 11040 841
rect 10994 769 11000 803
rect 11034 769 11040 803
rect 10994 731 11040 769
rect 10994 697 11000 731
rect 11034 697 11040 731
rect 10994 659 11040 697
rect 10994 625 11000 659
rect 11034 625 11040 659
rect 10994 587 11040 625
rect 10994 553 11000 587
rect 11034 553 11040 587
rect 10994 515 11040 553
rect 10994 481 11000 515
rect 11034 481 11040 515
rect 10994 443 11040 481
rect 10994 409 11000 443
rect 11034 409 11040 443
rect 10994 371 11040 409
rect 10994 337 11000 371
rect 11034 337 11040 371
rect 10994 299 11040 337
rect 10994 265 11000 299
rect 11034 265 11040 299
rect 10994 250 11040 265
rect 11090 1235 11136 1250
rect 11090 1201 11096 1235
rect 11130 1201 11136 1235
rect 11090 1163 11136 1201
rect 11090 1129 11096 1163
rect 11130 1129 11136 1163
rect 11090 1091 11136 1129
rect 11090 1057 11096 1091
rect 11130 1057 11136 1091
rect 11090 1019 11136 1057
rect 11090 985 11096 1019
rect 11130 985 11136 1019
rect 11090 947 11136 985
rect 11090 913 11096 947
rect 11130 913 11136 947
rect 11090 875 11136 913
rect 11090 841 11096 875
rect 11130 841 11136 875
rect 11090 803 11136 841
rect 11090 769 11096 803
rect 11130 769 11136 803
rect 11090 731 11136 769
rect 11090 697 11096 731
rect 11130 697 11136 731
rect 11090 659 11136 697
rect 11090 625 11096 659
rect 11130 625 11136 659
rect 11090 587 11136 625
rect 11090 553 11096 587
rect 11130 553 11136 587
rect 11090 515 11136 553
rect 11090 481 11096 515
rect 11130 481 11136 515
rect 11090 443 11136 481
rect 11090 409 11096 443
rect 11130 409 11136 443
rect 11090 371 11136 409
rect 11090 337 11096 371
rect 11130 337 11136 371
rect 11090 299 11136 337
rect 11090 265 11096 299
rect 11130 265 11136 299
rect 11090 250 11136 265
rect 11186 1235 11232 1250
rect 11186 1201 11192 1235
rect 11226 1201 11232 1235
rect 11186 1163 11232 1201
rect 11186 1129 11192 1163
rect 11226 1129 11232 1163
rect 11186 1091 11232 1129
rect 11186 1057 11192 1091
rect 11226 1057 11232 1091
rect 11186 1019 11232 1057
rect 11186 985 11192 1019
rect 11226 985 11232 1019
rect 11186 947 11232 985
rect 11186 913 11192 947
rect 11226 913 11232 947
rect 11186 875 11232 913
rect 11186 841 11192 875
rect 11226 841 11232 875
rect 11186 803 11232 841
rect 11186 769 11192 803
rect 11226 769 11232 803
rect 11186 731 11232 769
rect 11186 697 11192 731
rect 11226 697 11232 731
rect 11186 659 11232 697
rect 11186 625 11192 659
rect 11226 625 11232 659
rect 11186 587 11232 625
rect 11186 553 11192 587
rect 11226 553 11232 587
rect 11186 515 11232 553
rect 11186 481 11192 515
rect 11226 481 11232 515
rect 11186 443 11232 481
rect 11186 409 11192 443
rect 11226 409 11232 443
rect 11186 371 11232 409
rect 11186 337 11192 371
rect 11226 337 11232 371
rect 11186 299 11232 337
rect 11186 265 11192 299
rect 11226 265 11232 299
rect 11186 250 11232 265
rect 11282 1235 11328 1250
rect 11282 1201 11288 1235
rect 11322 1201 11328 1235
rect 11282 1163 11328 1201
rect 11282 1129 11288 1163
rect 11322 1129 11328 1163
rect 11282 1091 11328 1129
rect 11282 1057 11288 1091
rect 11322 1057 11328 1091
rect 11282 1019 11328 1057
rect 11282 985 11288 1019
rect 11322 985 11328 1019
rect 11282 947 11328 985
rect 11282 913 11288 947
rect 11322 913 11328 947
rect 11282 875 11328 913
rect 11282 841 11288 875
rect 11322 841 11328 875
rect 11282 803 11328 841
rect 11282 769 11288 803
rect 11322 769 11328 803
rect 11282 731 11328 769
rect 11282 697 11288 731
rect 11322 697 11328 731
rect 11282 659 11328 697
rect 11282 625 11288 659
rect 11322 625 11328 659
rect 11282 587 11328 625
rect 11282 553 11288 587
rect 11322 553 11328 587
rect 11282 515 11328 553
rect 11282 481 11288 515
rect 11322 481 11328 515
rect 11282 443 11328 481
rect 11282 409 11288 443
rect 11322 409 11328 443
rect 11282 371 11328 409
rect 11282 337 11288 371
rect 11322 337 11328 371
rect 11282 299 11328 337
rect 11282 265 11288 299
rect 11322 265 11328 299
rect 11282 250 11328 265
rect 11378 1235 11424 1250
rect 11378 1201 11384 1235
rect 11418 1201 11424 1235
rect 11378 1163 11424 1201
rect 11378 1129 11384 1163
rect 11418 1129 11424 1163
rect 11378 1091 11424 1129
rect 11378 1057 11384 1091
rect 11418 1057 11424 1091
rect 11378 1019 11424 1057
rect 11378 985 11384 1019
rect 11418 985 11424 1019
rect 11378 947 11424 985
rect 11378 913 11384 947
rect 11418 913 11424 947
rect 11378 875 11424 913
rect 11378 841 11384 875
rect 11418 841 11424 875
rect 11378 803 11424 841
rect 11378 769 11384 803
rect 11418 769 11424 803
rect 11378 731 11424 769
rect 11378 697 11384 731
rect 11418 697 11424 731
rect 11378 659 11424 697
rect 11378 625 11384 659
rect 11418 625 11424 659
rect 11378 587 11424 625
rect 11378 553 11384 587
rect 11418 553 11424 587
rect 11378 515 11424 553
rect 11378 481 11384 515
rect 11418 481 11424 515
rect 11378 443 11424 481
rect 11378 409 11384 443
rect 11418 409 11424 443
rect 11378 371 11424 409
rect 11378 337 11384 371
rect 11418 337 11424 371
rect 11378 299 11424 337
rect 11378 265 11384 299
rect 11418 265 11424 299
rect 11378 250 11424 265
rect 11474 1235 11520 1250
rect 11474 1201 11480 1235
rect 11514 1201 11520 1235
rect 11474 1163 11520 1201
rect 11474 1129 11480 1163
rect 11514 1129 11520 1163
rect 11474 1091 11520 1129
rect 11474 1057 11480 1091
rect 11514 1057 11520 1091
rect 11474 1019 11520 1057
rect 11474 985 11480 1019
rect 11514 985 11520 1019
rect 11474 947 11520 985
rect 11474 913 11480 947
rect 11514 913 11520 947
rect 11474 875 11520 913
rect 11474 841 11480 875
rect 11514 841 11520 875
rect 11474 803 11520 841
rect 11474 769 11480 803
rect 11514 769 11520 803
rect 11474 731 11520 769
rect 11474 697 11480 731
rect 11514 697 11520 731
rect 11474 659 11520 697
rect 11474 625 11480 659
rect 11514 625 11520 659
rect 11474 587 11520 625
rect 11474 553 11480 587
rect 11514 553 11520 587
rect 11474 515 11520 553
rect 11474 481 11480 515
rect 11514 481 11520 515
rect 11474 443 11520 481
rect 11474 409 11480 443
rect 11514 409 11520 443
rect 11474 371 11520 409
rect 11474 337 11480 371
rect 11514 337 11520 371
rect 11474 299 11520 337
rect 11474 265 11480 299
rect 11514 265 11520 299
rect 11474 250 11520 265
rect 11570 1235 11616 1250
rect 11570 1201 11576 1235
rect 11610 1201 11616 1235
rect 11570 1163 11616 1201
rect 11570 1129 11576 1163
rect 11610 1129 11616 1163
rect 11570 1091 11616 1129
rect 11570 1057 11576 1091
rect 11610 1057 11616 1091
rect 11570 1019 11616 1057
rect 11570 985 11576 1019
rect 11610 985 11616 1019
rect 11570 947 11616 985
rect 11570 913 11576 947
rect 11610 913 11616 947
rect 11570 875 11616 913
rect 11570 841 11576 875
rect 11610 841 11616 875
rect 11570 803 11616 841
rect 11570 769 11576 803
rect 11610 769 11616 803
rect 11570 731 11616 769
rect 11570 697 11576 731
rect 11610 697 11616 731
rect 11570 659 11616 697
rect 11570 625 11576 659
rect 11610 625 11616 659
rect 11570 587 11616 625
rect 11570 553 11576 587
rect 11610 553 11616 587
rect 11570 515 11616 553
rect 11570 481 11576 515
rect 11610 481 11616 515
rect 11570 443 11616 481
rect 11570 409 11576 443
rect 11610 409 11616 443
rect 11570 371 11616 409
rect 11570 337 11576 371
rect 11610 337 11616 371
rect 11570 299 11616 337
rect 11570 265 11576 299
rect 11610 265 11616 299
rect 11570 250 11616 265
rect 11666 1235 11712 1250
rect 11666 1201 11672 1235
rect 11706 1201 11712 1235
rect 11666 1163 11712 1201
rect 11666 1129 11672 1163
rect 11706 1129 11712 1163
rect 11666 1091 11712 1129
rect 11666 1057 11672 1091
rect 11706 1057 11712 1091
rect 11666 1019 11712 1057
rect 11666 985 11672 1019
rect 11706 985 11712 1019
rect 11666 947 11712 985
rect 11666 913 11672 947
rect 11706 913 11712 947
rect 11666 875 11712 913
rect 11666 841 11672 875
rect 11706 841 11712 875
rect 11666 803 11712 841
rect 11666 769 11672 803
rect 11706 769 11712 803
rect 11666 731 11712 769
rect 11666 697 11672 731
rect 11706 697 11712 731
rect 11666 659 11712 697
rect 11666 625 11672 659
rect 11706 625 11712 659
rect 11666 587 11712 625
rect 11666 553 11672 587
rect 11706 553 11712 587
rect 11666 515 11712 553
rect 11666 481 11672 515
rect 11706 481 11712 515
rect 11666 443 11712 481
rect 11666 409 11672 443
rect 11706 409 11712 443
rect 11666 371 11712 409
rect 11666 337 11672 371
rect 11706 337 11712 371
rect 11666 299 11712 337
rect 11666 265 11672 299
rect 11706 265 11712 299
rect 11666 250 11712 265
rect 11762 1235 11808 1250
rect 11762 1201 11768 1235
rect 11802 1201 11808 1235
rect 11762 1163 11808 1201
rect 11762 1129 11768 1163
rect 11802 1129 11808 1163
rect 11762 1091 11808 1129
rect 11762 1057 11768 1091
rect 11802 1057 11808 1091
rect 11762 1019 11808 1057
rect 11762 985 11768 1019
rect 11802 985 11808 1019
rect 11762 947 11808 985
rect 11762 913 11768 947
rect 11802 913 11808 947
rect 11762 875 11808 913
rect 11762 841 11768 875
rect 11802 841 11808 875
rect 11762 803 11808 841
rect 11762 769 11768 803
rect 11802 769 11808 803
rect 11762 731 11808 769
rect 11762 697 11768 731
rect 11802 697 11808 731
rect 11762 659 11808 697
rect 11762 625 11768 659
rect 11802 625 11808 659
rect 11762 587 11808 625
rect 11762 553 11768 587
rect 11802 553 11808 587
rect 11762 515 11808 553
rect 11762 481 11768 515
rect 11802 481 11808 515
rect 11762 443 11808 481
rect 11762 409 11768 443
rect 11802 409 11808 443
rect 11762 371 11808 409
rect 11762 337 11768 371
rect 11802 337 11808 371
rect 11762 299 11808 337
rect 11762 265 11768 299
rect 11802 265 11808 299
rect 11762 250 11808 265
rect 11858 1235 11904 1250
rect 11858 1201 11864 1235
rect 11898 1201 11904 1235
rect 11858 1163 11904 1201
rect 11858 1129 11864 1163
rect 11898 1129 11904 1163
rect 11858 1091 11904 1129
rect 11858 1057 11864 1091
rect 11898 1057 11904 1091
rect 11858 1019 11904 1057
rect 11858 985 11864 1019
rect 11898 985 11904 1019
rect 11858 947 11904 985
rect 11858 913 11864 947
rect 11898 913 11904 947
rect 11858 875 11904 913
rect 11858 841 11864 875
rect 11898 841 11904 875
rect 11858 803 11904 841
rect 11858 769 11864 803
rect 11898 769 11904 803
rect 11858 731 11904 769
rect 11858 697 11864 731
rect 11898 697 11904 731
rect 11858 659 11904 697
rect 11858 625 11864 659
rect 11898 625 11904 659
rect 11858 587 11904 625
rect 11858 553 11864 587
rect 11898 553 11904 587
rect 11858 515 11904 553
rect 11858 481 11864 515
rect 11898 481 11904 515
rect 11858 443 11904 481
rect 11858 409 11864 443
rect 11898 409 11904 443
rect 11858 371 11904 409
rect 11858 337 11864 371
rect 11898 337 11904 371
rect 11858 299 11904 337
rect 11858 265 11864 299
rect 11898 265 11904 299
rect 11858 250 11904 265
rect 11954 1235 12000 1250
rect 11954 1201 11960 1235
rect 11994 1201 12000 1235
rect 11954 1163 12000 1201
rect 11954 1129 11960 1163
rect 11994 1129 12000 1163
rect 11954 1091 12000 1129
rect 11954 1057 11960 1091
rect 11994 1057 12000 1091
rect 11954 1019 12000 1057
rect 11954 985 11960 1019
rect 11994 985 12000 1019
rect 11954 947 12000 985
rect 11954 913 11960 947
rect 11994 913 12000 947
rect 11954 875 12000 913
rect 11954 841 11960 875
rect 11994 841 12000 875
rect 11954 803 12000 841
rect 11954 769 11960 803
rect 11994 769 12000 803
rect 11954 731 12000 769
rect 11954 697 11960 731
rect 11994 697 12000 731
rect 11954 659 12000 697
rect 11954 625 11960 659
rect 11994 625 12000 659
rect 11954 587 12000 625
rect 11954 553 11960 587
rect 11994 553 12000 587
rect 11954 515 12000 553
rect 11954 481 11960 515
rect 11994 481 12000 515
rect 11954 443 12000 481
rect 11954 409 11960 443
rect 11994 409 12000 443
rect 11954 371 12000 409
rect 11954 337 11960 371
rect 11994 337 12000 371
rect 11954 299 12000 337
rect 11954 265 11960 299
rect 11994 265 12000 299
rect 11954 250 12000 265
rect 12050 1235 12096 1250
rect 12050 1201 12056 1235
rect 12090 1201 12096 1235
rect 12050 1163 12096 1201
rect 12050 1129 12056 1163
rect 12090 1129 12096 1163
rect 12050 1091 12096 1129
rect 12050 1057 12056 1091
rect 12090 1057 12096 1091
rect 12050 1019 12096 1057
rect 12050 985 12056 1019
rect 12090 985 12096 1019
rect 12050 947 12096 985
rect 12050 913 12056 947
rect 12090 913 12096 947
rect 12050 875 12096 913
rect 12050 841 12056 875
rect 12090 841 12096 875
rect 12050 803 12096 841
rect 12050 769 12056 803
rect 12090 769 12096 803
rect 12050 731 12096 769
rect 12050 697 12056 731
rect 12090 697 12096 731
rect 12050 659 12096 697
rect 12050 625 12056 659
rect 12090 625 12096 659
rect 12050 587 12096 625
rect 12050 553 12056 587
rect 12090 553 12096 587
rect 12050 515 12096 553
rect 12050 481 12056 515
rect 12090 481 12096 515
rect 12050 443 12096 481
rect 12050 409 12056 443
rect 12090 409 12096 443
rect 12050 371 12096 409
rect 12050 337 12056 371
rect 12090 337 12096 371
rect 12050 299 12096 337
rect 12050 265 12056 299
rect 12090 265 12096 299
rect 12050 250 12096 265
rect 12382 1209 12428 1224
rect 12382 1175 12388 1209
rect 12422 1175 12428 1209
rect 12382 1137 12428 1175
rect 12382 1103 12388 1137
rect 12422 1103 12428 1137
rect 12382 1065 12428 1103
rect 12382 1031 12388 1065
rect 12422 1031 12428 1065
rect 12382 993 12428 1031
rect 12382 959 12388 993
rect 12422 959 12428 993
rect 12382 921 12428 959
rect 12382 887 12388 921
rect 12422 887 12428 921
rect 12382 849 12428 887
rect 12382 815 12388 849
rect 12422 815 12428 849
rect 12382 777 12428 815
rect 12382 743 12388 777
rect 12422 743 12428 777
rect 12382 705 12428 743
rect 12382 671 12388 705
rect 12422 671 12428 705
rect 12382 633 12428 671
rect 12382 599 12388 633
rect 12422 599 12428 633
rect 12382 561 12428 599
rect 12382 527 12388 561
rect 12422 527 12428 561
rect 12382 489 12428 527
rect 12382 455 12388 489
rect 12422 455 12428 489
rect 12382 417 12428 455
rect 12382 383 12388 417
rect 12422 383 12428 417
rect 12382 345 12428 383
rect 12382 311 12388 345
rect 12422 311 12428 345
rect 12382 273 12428 311
rect 12382 239 12388 273
rect 12422 239 12428 273
rect 12382 224 12428 239
rect 12478 1209 12524 1224
rect 12478 1175 12484 1209
rect 12518 1175 12524 1209
rect 12478 1137 12524 1175
rect 12478 1103 12484 1137
rect 12518 1103 12524 1137
rect 12478 1065 12524 1103
rect 12478 1031 12484 1065
rect 12518 1031 12524 1065
rect 12478 993 12524 1031
rect 12478 959 12484 993
rect 12518 959 12524 993
rect 12478 921 12524 959
rect 12478 887 12484 921
rect 12518 887 12524 921
rect 12478 849 12524 887
rect 12478 815 12484 849
rect 12518 815 12524 849
rect 12478 777 12524 815
rect 12478 743 12484 777
rect 12518 743 12524 777
rect 12478 705 12524 743
rect 12478 671 12484 705
rect 12518 671 12524 705
rect 12478 633 12524 671
rect 12478 599 12484 633
rect 12518 599 12524 633
rect 12478 561 12524 599
rect 12478 527 12484 561
rect 12518 527 12524 561
rect 12478 489 12524 527
rect 12478 455 12484 489
rect 12518 455 12524 489
rect 12478 417 12524 455
rect 12478 383 12484 417
rect 12518 383 12524 417
rect 12478 345 12524 383
rect 12478 311 12484 345
rect 12518 311 12524 345
rect 12478 273 12524 311
rect 12478 239 12484 273
rect 12518 239 12524 273
rect 12478 224 12524 239
rect 12574 1209 12620 1224
rect 12574 1175 12580 1209
rect 12614 1175 12620 1209
rect 12574 1137 12620 1175
rect 12574 1103 12580 1137
rect 12614 1103 12620 1137
rect 12574 1065 12620 1103
rect 12574 1031 12580 1065
rect 12614 1031 12620 1065
rect 12574 993 12620 1031
rect 12574 959 12580 993
rect 12614 959 12620 993
rect 12574 921 12620 959
rect 12574 887 12580 921
rect 12614 887 12620 921
rect 12574 849 12620 887
rect 12574 815 12580 849
rect 12614 815 12620 849
rect 12574 777 12620 815
rect 12574 743 12580 777
rect 12614 743 12620 777
rect 12574 705 12620 743
rect 12574 671 12580 705
rect 12614 671 12620 705
rect 12574 633 12620 671
rect 12574 599 12580 633
rect 12614 599 12620 633
rect 12574 561 12620 599
rect 12574 527 12580 561
rect 12614 527 12620 561
rect 12574 489 12620 527
rect 12574 455 12580 489
rect 12614 455 12620 489
rect 12574 417 12620 455
rect 12574 383 12580 417
rect 12614 383 12620 417
rect 12574 345 12620 383
rect 12574 311 12580 345
rect 12614 311 12620 345
rect 12574 273 12620 311
rect 12574 239 12580 273
rect 12614 239 12620 273
rect 12574 224 12620 239
rect 12670 1209 12716 1224
rect 12670 1175 12676 1209
rect 12710 1175 12716 1209
rect 12670 1137 12716 1175
rect 12670 1103 12676 1137
rect 12710 1103 12716 1137
rect 12670 1065 12716 1103
rect 12670 1031 12676 1065
rect 12710 1031 12716 1065
rect 12670 993 12716 1031
rect 12670 959 12676 993
rect 12710 959 12716 993
rect 12670 921 12716 959
rect 12670 887 12676 921
rect 12710 887 12716 921
rect 12670 849 12716 887
rect 12670 815 12676 849
rect 12710 815 12716 849
rect 12670 777 12716 815
rect 12670 743 12676 777
rect 12710 743 12716 777
rect 12670 705 12716 743
rect 12670 671 12676 705
rect 12710 671 12716 705
rect 12670 633 12716 671
rect 12670 599 12676 633
rect 12710 599 12716 633
rect 12670 561 12716 599
rect 12670 527 12676 561
rect 12710 527 12716 561
rect 12670 489 12716 527
rect 12670 455 12676 489
rect 12710 455 12716 489
rect 12670 417 12716 455
rect 12670 383 12676 417
rect 12710 383 12716 417
rect 12670 345 12716 383
rect 12670 311 12676 345
rect 12710 311 12716 345
rect 12670 273 12716 311
rect 12670 239 12676 273
rect 12710 239 12716 273
rect 12670 224 12716 239
rect 12766 1209 12812 1224
rect 12766 1175 12772 1209
rect 12806 1175 12812 1209
rect 12766 1137 12812 1175
rect 12766 1103 12772 1137
rect 12806 1103 12812 1137
rect 12766 1065 12812 1103
rect 12766 1031 12772 1065
rect 12806 1031 12812 1065
rect 12766 993 12812 1031
rect 12766 959 12772 993
rect 12806 959 12812 993
rect 12766 921 12812 959
rect 12766 887 12772 921
rect 12806 887 12812 921
rect 12766 849 12812 887
rect 12766 815 12772 849
rect 12806 815 12812 849
rect 12766 777 12812 815
rect 12766 743 12772 777
rect 12806 743 12812 777
rect 12766 705 12812 743
rect 12766 671 12772 705
rect 12806 671 12812 705
rect 12766 633 12812 671
rect 12766 599 12772 633
rect 12806 599 12812 633
rect 12766 561 12812 599
rect 12766 527 12772 561
rect 12806 527 12812 561
rect 12766 489 12812 527
rect 12766 455 12772 489
rect 12806 455 12812 489
rect 12766 417 12812 455
rect 12766 383 12772 417
rect 12806 383 12812 417
rect 12766 345 12812 383
rect 12766 311 12772 345
rect 12806 311 12812 345
rect 12766 273 12812 311
rect 12766 239 12772 273
rect 12806 239 12812 273
rect 12766 224 12812 239
rect 12862 1209 12908 1224
rect 12862 1175 12868 1209
rect 12902 1175 12908 1209
rect 12862 1137 12908 1175
rect 12862 1103 12868 1137
rect 12902 1103 12908 1137
rect 12862 1065 12908 1103
rect 12862 1031 12868 1065
rect 12902 1031 12908 1065
rect 12862 993 12908 1031
rect 12862 959 12868 993
rect 12902 959 12908 993
rect 12862 921 12908 959
rect 12862 887 12868 921
rect 12902 887 12908 921
rect 12862 849 12908 887
rect 12862 815 12868 849
rect 12902 815 12908 849
rect 12862 777 12908 815
rect 12862 743 12868 777
rect 12902 743 12908 777
rect 12862 705 12908 743
rect 12862 671 12868 705
rect 12902 671 12908 705
rect 12862 633 12908 671
rect 12862 599 12868 633
rect 12902 599 12908 633
rect 12862 561 12908 599
rect 12862 527 12868 561
rect 12902 527 12908 561
rect 12862 489 12908 527
rect 12862 455 12868 489
rect 12902 455 12908 489
rect 12862 417 12908 455
rect 12862 383 12868 417
rect 12902 383 12908 417
rect 12862 345 12908 383
rect 12862 311 12868 345
rect 12902 311 12908 345
rect 12862 273 12908 311
rect 12862 239 12868 273
rect 12902 239 12908 273
rect 12862 224 12908 239
rect 12958 1209 13004 1224
rect 12958 1175 12964 1209
rect 12998 1175 13004 1209
rect 12958 1137 13004 1175
rect 12958 1103 12964 1137
rect 12998 1103 13004 1137
rect 12958 1065 13004 1103
rect 12958 1031 12964 1065
rect 12998 1031 13004 1065
rect 12958 993 13004 1031
rect 12958 959 12964 993
rect 12998 959 13004 993
rect 12958 921 13004 959
rect 12958 887 12964 921
rect 12998 887 13004 921
rect 12958 849 13004 887
rect 12958 815 12964 849
rect 12998 815 13004 849
rect 12958 777 13004 815
rect 12958 743 12964 777
rect 12998 743 13004 777
rect 12958 705 13004 743
rect 12958 671 12964 705
rect 12998 671 13004 705
rect 12958 633 13004 671
rect 12958 599 12964 633
rect 12998 599 13004 633
rect 12958 561 13004 599
rect 12958 527 12964 561
rect 12998 527 13004 561
rect 12958 489 13004 527
rect 12958 455 12964 489
rect 12998 455 13004 489
rect 12958 417 13004 455
rect 12958 383 12964 417
rect 12998 383 13004 417
rect 12958 345 13004 383
rect 12958 311 12964 345
rect 12998 311 13004 345
rect 12958 273 13004 311
rect 12958 239 12964 273
rect 12998 239 13004 273
rect 12958 224 13004 239
rect 13054 1209 13100 1224
rect 13054 1175 13060 1209
rect 13094 1175 13100 1209
rect 13054 1137 13100 1175
rect 13054 1103 13060 1137
rect 13094 1103 13100 1137
rect 13054 1065 13100 1103
rect 13054 1031 13060 1065
rect 13094 1031 13100 1065
rect 13054 993 13100 1031
rect 13054 959 13060 993
rect 13094 959 13100 993
rect 13054 921 13100 959
rect 13054 887 13060 921
rect 13094 887 13100 921
rect 13054 849 13100 887
rect 13054 815 13060 849
rect 13094 815 13100 849
rect 13054 777 13100 815
rect 13054 743 13060 777
rect 13094 743 13100 777
rect 13054 705 13100 743
rect 13054 671 13060 705
rect 13094 671 13100 705
rect 13054 633 13100 671
rect 13054 599 13060 633
rect 13094 599 13100 633
rect 13054 561 13100 599
rect 13054 527 13060 561
rect 13094 527 13100 561
rect 13054 489 13100 527
rect 13054 455 13060 489
rect 13094 455 13100 489
rect 13054 417 13100 455
rect 13054 383 13060 417
rect 13094 383 13100 417
rect 13054 345 13100 383
rect 13054 311 13060 345
rect 13094 311 13100 345
rect 13054 273 13100 311
rect 13054 239 13060 273
rect 13094 239 13100 273
rect 13054 224 13100 239
rect 13150 1209 13196 1224
rect 13150 1175 13156 1209
rect 13190 1175 13196 1209
rect 13150 1137 13196 1175
rect 13150 1103 13156 1137
rect 13190 1103 13196 1137
rect 13150 1065 13196 1103
rect 13150 1031 13156 1065
rect 13190 1031 13196 1065
rect 13150 993 13196 1031
rect 13150 959 13156 993
rect 13190 959 13196 993
rect 13150 921 13196 959
rect 13150 887 13156 921
rect 13190 887 13196 921
rect 13150 849 13196 887
rect 13150 815 13156 849
rect 13190 815 13196 849
rect 13150 777 13196 815
rect 13150 743 13156 777
rect 13190 743 13196 777
rect 13150 705 13196 743
rect 13150 671 13156 705
rect 13190 671 13196 705
rect 13150 633 13196 671
rect 13150 599 13156 633
rect 13190 599 13196 633
rect 13150 561 13196 599
rect 13150 527 13156 561
rect 13190 527 13196 561
rect 13150 489 13196 527
rect 13150 455 13156 489
rect 13190 455 13196 489
rect 13150 417 13196 455
rect 13150 383 13156 417
rect 13190 383 13196 417
rect 13150 345 13196 383
rect 13150 311 13156 345
rect 13190 311 13196 345
rect 13150 273 13196 311
rect 13150 239 13156 273
rect 13190 239 13196 273
rect 13150 224 13196 239
rect 13246 1209 13292 1224
rect 13246 1175 13252 1209
rect 13286 1175 13292 1209
rect 13246 1137 13292 1175
rect 13246 1103 13252 1137
rect 13286 1103 13292 1137
rect 13246 1065 13292 1103
rect 13246 1031 13252 1065
rect 13286 1031 13292 1065
rect 13246 993 13292 1031
rect 13246 959 13252 993
rect 13286 959 13292 993
rect 13246 921 13292 959
rect 13246 887 13252 921
rect 13286 887 13292 921
rect 13246 849 13292 887
rect 13246 815 13252 849
rect 13286 815 13292 849
rect 13246 777 13292 815
rect 13246 743 13252 777
rect 13286 743 13292 777
rect 13246 705 13292 743
rect 13246 671 13252 705
rect 13286 671 13292 705
rect 13246 633 13292 671
rect 13246 599 13252 633
rect 13286 599 13292 633
rect 13246 561 13292 599
rect 13246 527 13252 561
rect 13286 527 13292 561
rect 13246 489 13292 527
rect 13246 455 13252 489
rect 13286 455 13292 489
rect 13246 417 13292 455
rect 13246 383 13252 417
rect 13286 383 13292 417
rect 13246 345 13292 383
rect 13246 311 13252 345
rect 13286 311 13292 345
rect 13246 273 13292 311
rect 13246 239 13252 273
rect 13286 239 13292 273
rect 13246 224 13292 239
rect 13342 1209 13388 1224
rect 13342 1175 13348 1209
rect 13382 1175 13388 1209
rect 13342 1137 13388 1175
rect 13342 1103 13348 1137
rect 13382 1103 13388 1137
rect 13342 1065 13388 1103
rect 13342 1031 13348 1065
rect 13382 1031 13388 1065
rect 13342 993 13388 1031
rect 13342 959 13348 993
rect 13382 959 13388 993
rect 13342 921 13388 959
rect 13342 887 13348 921
rect 13382 887 13388 921
rect 13342 849 13388 887
rect 13342 815 13348 849
rect 13382 815 13388 849
rect 13342 777 13388 815
rect 13342 743 13348 777
rect 13382 743 13388 777
rect 13342 705 13388 743
rect 13342 671 13348 705
rect 13382 671 13388 705
rect 13342 633 13388 671
rect 13342 599 13348 633
rect 13382 599 13388 633
rect 13342 561 13388 599
rect 13342 527 13348 561
rect 13382 527 13388 561
rect 13342 489 13388 527
rect 13342 455 13348 489
rect 13382 455 13388 489
rect 13342 417 13388 455
rect 13342 383 13348 417
rect 13382 383 13388 417
rect 13342 345 13388 383
rect 13342 311 13348 345
rect 13382 311 13388 345
rect 13342 273 13388 311
rect 13342 239 13348 273
rect 13382 239 13388 273
rect 13342 224 13388 239
rect 13438 1209 13484 1224
rect 13438 1175 13444 1209
rect 13478 1175 13484 1209
rect 13438 1137 13484 1175
rect 13438 1103 13444 1137
rect 13478 1103 13484 1137
rect 13438 1065 13484 1103
rect 13438 1031 13444 1065
rect 13478 1031 13484 1065
rect 13438 993 13484 1031
rect 13438 959 13444 993
rect 13478 959 13484 993
rect 13438 921 13484 959
rect 13438 887 13444 921
rect 13478 887 13484 921
rect 13438 849 13484 887
rect 13438 815 13444 849
rect 13478 815 13484 849
rect 13438 777 13484 815
rect 13438 743 13444 777
rect 13478 743 13484 777
rect 13438 705 13484 743
rect 13438 671 13444 705
rect 13478 671 13484 705
rect 13438 633 13484 671
rect 13438 599 13444 633
rect 13478 599 13484 633
rect 13438 561 13484 599
rect 13438 527 13444 561
rect 13478 527 13484 561
rect 13438 489 13484 527
rect 13438 455 13444 489
rect 13478 455 13484 489
rect 13438 417 13484 455
rect 13438 383 13444 417
rect 13478 383 13484 417
rect 13438 345 13484 383
rect 13438 311 13444 345
rect 13478 311 13484 345
rect 13438 273 13484 311
rect 13438 239 13444 273
rect 13478 239 13484 273
rect 13438 224 13484 239
rect 13534 1209 13580 1224
rect 13534 1175 13540 1209
rect 13574 1175 13580 1209
rect 13534 1137 13580 1175
rect 13534 1103 13540 1137
rect 13574 1103 13580 1137
rect 13534 1065 13580 1103
rect 13534 1031 13540 1065
rect 13574 1031 13580 1065
rect 13534 993 13580 1031
rect 13534 959 13540 993
rect 13574 959 13580 993
rect 13534 921 13580 959
rect 13534 887 13540 921
rect 13574 887 13580 921
rect 13534 849 13580 887
rect 13534 815 13540 849
rect 13574 815 13580 849
rect 13534 777 13580 815
rect 13534 743 13540 777
rect 13574 743 13580 777
rect 13534 705 13580 743
rect 13534 671 13540 705
rect 13574 671 13580 705
rect 13534 633 13580 671
rect 13534 599 13540 633
rect 13574 599 13580 633
rect 13534 561 13580 599
rect 13534 527 13540 561
rect 13574 527 13580 561
rect 13534 489 13580 527
rect 13534 455 13540 489
rect 13574 455 13580 489
rect 13534 417 13580 455
rect 13534 383 13540 417
rect 13574 383 13580 417
rect 13534 345 13580 383
rect 13534 311 13540 345
rect 13574 311 13580 345
rect 13534 273 13580 311
rect 13534 239 13540 273
rect 13574 239 13580 273
rect 13534 224 13580 239
rect 14150 1209 14196 1224
rect 14150 1175 14156 1209
rect 14190 1175 14196 1209
rect 14150 1137 14196 1175
rect 14150 1103 14156 1137
rect 14190 1103 14196 1137
rect 14150 1065 14196 1103
rect 14150 1031 14156 1065
rect 14190 1031 14196 1065
rect 14150 993 14196 1031
rect 14150 959 14156 993
rect 14190 959 14196 993
rect 14150 921 14196 959
rect 14150 887 14156 921
rect 14190 887 14196 921
rect 14150 849 14196 887
rect 14150 815 14156 849
rect 14190 815 14196 849
rect 14150 777 14196 815
rect 14150 743 14156 777
rect 14190 743 14196 777
rect 14150 705 14196 743
rect 14150 671 14156 705
rect 14190 671 14196 705
rect 14150 633 14196 671
rect 14150 599 14156 633
rect 14190 599 14196 633
rect 14150 561 14196 599
rect 14150 527 14156 561
rect 14190 527 14196 561
rect 14150 489 14196 527
rect 14150 455 14156 489
rect 14190 455 14196 489
rect 14150 417 14196 455
rect 14150 383 14156 417
rect 14190 383 14196 417
rect 14150 345 14196 383
rect 14150 311 14156 345
rect 14190 311 14196 345
rect 14150 273 14196 311
rect 14150 239 14156 273
rect 14190 239 14196 273
rect 14150 224 14196 239
rect 14246 1209 14292 1224
rect 14246 1175 14252 1209
rect 14286 1175 14292 1209
rect 14246 1137 14292 1175
rect 14246 1103 14252 1137
rect 14286 1103 14292 1137
rect 14246 1065 14292 1103
rect 14246 1031 14252 1065
rect 14286 1031 14292 1065
rect 14246 993 14292 1031
rect 14246 959 14252 993
rect 14286 959 14292 993
rect 14246 921 14292 959
rect 14246 887 14252 921
rect 14286 887 14292 921
rect 14246 849 14292 887
rect 14246 815 14252 849
rect 14286 815 14292 849
rect 14246 777 14292 815
rect 14246 743 14252 777
rect 14286 743 14292 777
rect 14246 705 14292 743
rect 14246 671 14252 705
rect 14286 671 14292 705
rect 14246 633 14292 671
rect 14246 599 14252 633
rect 14286 599 14292 633
rect 14246 561 14292 599
rect 14246 527 14252 561
rect 14286 527 14292 561
rect 14246 489 14292 527
rect 14246 455 14252 489
rect 14286 455 14292 489
rect 14246 417 14292 455
rect 14246 383 14252 417
rect 14286 383 14292 417
rect 14246 345 14292 383
rect 14246 311 14252 345
rect 14286 311 14292 345
rect 14246 273 14292 311
rect 14246 239 14252 273
rect 14286 239 14292 273
rect 14246 224 14292 239
rect 14342 1209 14388 1224
rect 14342 1175 14348 1209
rect 14382 1175 14388 1209
rect 14342 1137 14388 1175
rect 14342 1103 14348 1137
rect 14382 1103 14388 1137
rect 14342 1065 14388 1103
rect 14342 1031 14348 1065
rect 14382 1031 14388 1065
rect 14342 993 14388 1031
rect 14342 959 14348 993
rect 14382 959 14388 993
rect 14342 921 14388 959
rect 14342 887 14348 921
rect 14382 887 14388 921
rect 14342 849 14388 887
rect 14342 815 14348 849
rect 14382 815 14388 849
rect 14342 777 14388 815
rect 14342 743 14348 777
rect 14382 743 14388 777
rect 14342 705 14388 743
rect 14342 671 14348 705
rect 14382 671 14388 705
rect 14342 633 14388 671
rect 14342 599 14348 633
rect 14382 599 14388 633
rect 14342 561 14388 599
rect 14342 527 14348 561
rect 14382 527 14388 561
rect 14342 489 14388 527
rect 14342 455 14348 489
rect 14382 455 14388 489
rect 14342 417 14388 455
rect 14342 383 14348 417
rect 14382 383 14388 417
rect 14342 345 14388 383
rect 14342 311 14348 345
rect 14382 311 14388 345
rect 14342 273 14388 311
rect 14342 239 14348 273
rect 14382 239 14388 273
rect 14342 224 14388 239
rect 14438 1209 14484 1224
rect 14438 1175 14444 1209
rect 14478 1175 14484 1209
rect 14438 1137 14484 1175
rect 14438 1103 14444 1137
rect 14478 1103 14484 1137
rect 14438 1065 14484 1103
rect 14438 1031 14444 1065
rect 14478 1031 14484 1065
rect 14438 993 14484 1031
rect 14438 959 14444 993
rect 14478 959 14484 993
rect 14438 921 14484 959
rect 14438 887 14444 921
rect 14478 887 14484 921
rect 14438 849 14484 887
rect 14438 815 14444 849
rect 14478 815 14484 849
rect 14438 777 14484 815
rect 14438 743 14444 777
rect 14478 743 14484 777
rect 14438 705 14484 743
rect 14438 671 14444 705
rect 14478 671 14484 705
rect 14438 633 14484 671
rect 14438 599 14444 633
rect 14478 599 14484 633
rect 14438 561 14484 599
rect 14438 527 14444 561
rect 14478 527 14484 561
rect 14438 489 14484 527
rect 14438 455 14444 489
rect 14478 455 14484 489
rect 14438 417 14484 455
rect 14438 383 14444 417
rect 14478 383 14484 417
rect 14438 345 14484 383
rect 14438 311 14444 345
rect 14478 311 14484 345
rect 14438 273 14484 311
rect 14438 239 14444 273
rect 14478 239 14484 273
rect 14438 224 14484 239
rect 14534 1209 14580 1224
rect 14534 1175 14540 1209
rect 14574 1175 14580 1209
rect 14534 1137 14580 1175
rect 14534 1103 14540 1137
rect 14574 1103 14580 1137
rect 14534 1065 14580 1103
rect 14534 1031 14540 1065
rect 14574 1031 14580 1065
rect 14534 993 14580 1031
rect 14534 959 14540 993
rect 14574 959 14580 993
rect 14534 921 14580 959
rect 14534 887 14540 921
rect 14574 887 14580 921
rect 14534 849 14580 887
rect 14534 815 14540 849
rect 14574 815 14580 849
rect 14534 777 14580 815
rect 14534 743 14540 777
rect 14574 743 14580 777
rect 14534 705 14580 743
rect 14534 671 14540 705
rect 14574 671 14580 705
rect 14534 633 14580 671
rect 14534 599 14540 633
rect 14574 599 14580 633
rect 14534 561 14580 599
rect 14534 527 14540 561
rect 14574 527 14580 561
rect 14534 489 14580 527
rect 14534 455 14540 489
rect 14574 455 14580 489
rect 14534 417 14580 455
rect 14534 383 14540 417
rect 14574 383 14580 417
rect 14534 345 14580 383
rect 14534 311 14540 345
rect 14574 311 14580 345
rect 14534 273 14580 311
rect 14534 239 14540 273
rect 14574 239 14580 273
rect 14534 224 14580 239
rect 14630 1209 14676 1224
rect 14630 1175 14636 1209
rect 14670 1175 14676 1209
rect 14630 1137 14676 1175
rect 14630 1103 14636 1137
rect 14670 1103 14676 1137
rect 14630 1065 14676 1103
rect 14630 1031 14636 1065
rect 14670 1031 14676 1065
rect 14630 993 14676 1031
rect 14630 959 14636 993
rect 14670 959 14676 993
rect 14630 921 14676 959
rect 14630 887 14636 921
rect 14670 887 14676 921
rect 14630 849 14676 887
rect 14630 815 14636 849
rect 14670 815 14676 849
rect 14630 777 14676 815
rect 14630 743 14636 777
rect 14670 743 14676 777
rect 14630 705 14676 743
rect 14630 671 14636 705
rect 14670 671 14676 705
rect 14630 633 14676 671
rect 14630 599 14636 633
rect 14670 599 14676 633
rect 14630 561 14676 599
rect 14630 527 14636 561
rect 14670 527 14676 561
rect 14630 489 14676 527
rect 14630 455 14636 489
rect 14670 455 14676 489
rect 14630 417 14676 455
rect 14630 383 14636 417
rect 14670 383 14676 417
rect 14630 345 14676 383
rect 14630 311 14636 345
rect 14670 311 14676 345
rect 14630 273 14676 311
rect 14630 239 14636 273
rect 14670 239 14676 273
rect 14630 224 14676 239
rect 14726 1209 14772 1224
rect 14726 1175 14732 1209
rect 14766 1175 14772 1209
rect 14726 1137 14772 1175
rect 14726 1103 14732 1137
rect 14766 1103 14772 1137
rect 14726 1065 14772 1103
rect 14726 1031 14732 1065
rect 14766 1031 14772 1065
rect 14726 993 14772 1031
rect 14726 959 14732 993
rect 14766 959 14772 993
rect 14726 921 14772 959
rect 14726 887 14732 921
rect 14766 887 14772 921
rect 14726 849 14772 887
rect 14726 815 14732 849
rect 14766 815 14772 849
rect 14726 777 14772 815
rect 14726 743 14732 777
rect 14766 743 14772 777
rect 14726 705 14772 743
rect 14726 671 14732 705
rect 14766 671 14772 705
rect 14726 633 14772 671
rect 14726 599 14732 633
rect 14766 599 14772 633
rect 14726 561 14772 599
rect 14726 527 14732 561
rect 14766 527 14772 561
rect 14726 489 14772 527
rect 14726 455 14732 489
rect 14766 455 14772 489
rect 14726 417 14772 455
rect 14726 383 14732 417
rect 14766 383 14772 417
rect 14726 345 14772 383
rect 14726 311 14732 345
rect 14766 311 14772 345
rect 14726 273 14772 311
rect 14726 239 14732 273
rect 14766 239 14772 273
rect 14726 224 14772 239
rect 14822 1209 14868 1224
rect 14822 1175 14828 1209
rect 14862 1175 14868 1209
rect 14822 1137 14868 1175
rect 14822 1103 14828 1137
rect 14862 1103 14868 1137
rect 14822 1065 14868 1103
rect 14822 1031 14828 1065
rect 14862 1031 14868 1065
rect 14822 993 14868 1031
rect 14822 959 14828 993
rect 14862 959 14868 993
rect 14822 921 14868 959
rect 14822 887 14828 921
rect 14862 887 14868 921
rect 14822 849 14868 887
rect 14822 815 14828 849
rect 14862 815 14868 849
rect 14822 777 14868 815
rect 14822 743 14828 777
rect 14862 743 14868 777
rect 14822 705 14868 743
rect 14822 671 14828 705
rect 14862 671 14868 705
rect 14822 633 14868 671
rect 14822 599 14828 633
rect 14862 599 14868 633
rect 14822 561 14868 599
rect 14822 527 14828 561
rect 14862 527 14868 561
rect 14822 489 14868 527
rect 14822 455 14828 489
rect 14862 455 14868 489
rect 14822 417 14868 455
rect 14822 383 14828 417
rect 14862 383 14868 417
rect 14822 345 14868 383
rect 14822 311 14828 345
rect 14862 311 14868 345
rect 14822 273 14868 311
rect 14822 239 14828 273
rect 14862 239 14868 273
rect 14822 224 14868 239
rect 14918 1209 14964 1224
rect 14918 1175 14924 1209
rect 14958 1175 14964 1209
rect 14918 1137 14964 1175
rect 14918 1103 14924 1137
rect 14958 1103 14964 1137
rect 14918 1065 14964 1103
rect 14918 1031 14924 1065
rect 14958 1031 14964 1065
rect 14918 993 14964 1031
rect 14918 959 14924 993
rect 14958 959 14964 993
rect 14918 921 14964 959
rect 14918 887 14924 921
rect 14958 887 14964 921
rect 14918 849 14964 887
rect 14918 815 14924 849
rect 14958 815 14964 849
rect 14918 777 14964 815
rect 14918 743 14924 777
rect 14958 743 14964 777
rect 14918 705 14964 743
rect 14918 671 14924 705
rect 14958 671 14964 705
rect 14918 633 14964 671
rect 14918 599 14924 633
rect 14958 599 14964 633
rect 14918 561 14964 599
rect 14918 527 14924 561
rect 14958 527 14964 561
rect 14918 489 14964 527
rect 14918 455 14924 489
rect 14958 455 14964 489
rect 14918 417 14964 455
rect 14918 383 14924 417
rect 14958 383 14964 417
rect 14918 345 14964 383
rect 14918 311 14924 345
rect 14958 311 14964 345
rect 14918 273 14964 311
rect 14918 239 14924 273
rect 14958 239 14964 273
rect 14918 224 14964 239
rect 15014 1209 15060 1224
rect 15014 1175 15020 1209
rect 15054 1175 15060 1209
rect 15014 1137 15060 1175
rect 15014 1103 15020 1137
rect 15054 1103 15060 1137
rect 15014 1065 15060 1103
rect 15014 1031 15020 1065
rect 15054 1031 15060 1065
rect 15014 993 15060 1031
rect 15014 959 15020 993
rect 15054 959 15060 993
rect 15014 921 15060 959
rect 15014 887 15020 921
rect 15054 887 15060 921
rect 15014 849 15060 887
rect 15014 815 15020 849
rect 15054 815 15060 849
rect 15014 777 15060 815
rect 15014 743 15020 777
rect 15054 743 15060 777
rect 15014 705 15060 743
rect 15014 671 15020 705
rect 15054 671 15060 705
rect 15014 633 15060 671
rect 15014 599 15020 633
rect 15054 599 15060 633
rect 15014 561 15060 599
rect 15014 527 15020 561
rect 15054 527 15060 561
rect 15014 489 15060 527
rect 15014 455 15020 489
rect 15054 455 15060 489
rect 15014 417 15060 455
rect 15014 383 15020 417
rect 15054 383 15060 417
rect 15014 345 15060 383
rect 15014 311 15020 345
rect 15054 311 15060 345
rect 15014 273 15060 311
rect 15014 239 15020 273
rect 15054 239 15060 273
rect 15014 224 15060 239
rect 15110 1209 15156 1224
rect 15110 1175 15116 1209
rect 15150 1175 15156 1209
rect 15110 1137 15156 1175
rect 15110 1103 15116 1137
rect 15150 1103 15156 1137
rect 15110 1065 15156 1103
rect 15110 1031 15116 1065
rect 15150 1031 15156 1065
rect 15110 993 15156 1031
rect 15110 959 15116 993
rect 15150 959 15156 993
rect 15110 921 15156 959
rect 15110 887 15116 921
rect 15150 887 15156 921
rect 15110 849 15156 887
rect 15110 815 15116 849
rect 15150 815 15156 849
rect 15110 777 15156 815
rect 15110 743 15116 777
rect 15150 743 15156 777
rect 15110 705 15156 743
rect 15110 671 15116 705
rect 15150 671 15156 705
rect 15110 633 15156 671
rect 15110 599 15116 633
rect 15150 599 15156 633
rect 15110 561 15156 599
rect 15110 527 15116 561
rect 15150 527 15156 561
rect 15110 489 15156 527
rect 15110 455 15116 489
rect 15150 455 15156 489
rect 15110 417 15156 455
rect 15110 383 15116 417
rect 15150 383 15156 417
rect 15110 345 15156 383
rect 15110 311 15116 345
rect 15150 311 15156 345
rect 15110 273 15156 311
rect 15110 239 15116 273
rect 15150 239 15156 273
rect 15110 224 15156 239
rect 15206 1209 15252 1224
rect 15206 1175 15212 1209
rect 15246 1175 15252 1209
rect 15206 1137 15252 1175
rect 15206 1103 15212 1137
rect 15246 1103 15252 1137
rect 15206 1065 15252 1103
rect 15206 1031 15212 1065
rect 15246 1031 15252 1065
rect 15206 993 15252 1031
rect 15206 959 15212 993
rect 15246 959 15252 993
rect 15206 921 15252 959
rect 15206 887 15212 921
rect 15246 887 15252 921
rect 15206 849 15252 887
rect 15206 815 15212 849
rect 15246 815 15252 849
rect 15206 777 15252 815
rect 15206 743 15212 777
rect 15246 743 15252 777
rect 15206 705 15252 743
rect 15206 671 15212 705
rect 15246 671 15252 705
rect 15206 633 15252 671
rect 15206 599 15212 633
rect 15246 599 15252 633
rect 15206 561 15252 599
rect 15206 527 15212 561
rect 15246 527 15252 561
rect 15206 489 15252 527
rect 15206 455 15212 489
rect 15246 455 15252 489
rect 15206 417 15252 455
rect 15206 383 15212 417
rect 15246 383 15252 417
rect 15206 345 15252 383
rect 15206 311 15212 345
rect 15246 311 15252 345
rect 15206 273 15252 311
rect 15206 239 15212 273
rect 15246 239 15252 273
rect 15206 224 15252 239
rect 15416 1223 15422 1257
rect 15456 1223 15462 1257
rect 15416 1185 15462 1223
rect 15416 1151 15422 1185
rect 15456 1151 15462 1185
rect 15416 1113 15462 1151
rect 15416 1079 15422 1113
rect 15456 1079 15462 1113
rect 15416 1041 15462 1079
rect 15416 1007 15422 1041
rect 15456 1007 15462 1041
rect 15416 969 15462 1007
rect 15416 935 15422 969
rect 15456 935 15462 969
rect 15416 897 15462 935
rect 15416 863 15422 897
rect 15456 863 15462 897
rect 15416 825 15462 863
rect 15416 791 15422 825
rect 15456 791 15462 825
rect 15416 753 15462 791
rect 15416 719 15422 753
rect 15456 719 15462 753
rect 15416 681 15462 719
rect 15416 647 15422 681
rect 15456 647 15462 681
rect 15416 609 15462 647
rect 15416 575 15422 609
rect 15456 575 15462 609
rect 15416 537 15462 575
rect 15416 503 15422 537
rect 15456 503 15462 537
rect 15416 465 15462 503
rect 15416 431 15422 465
rect 15456 431 15462 465
rect 15416 393 15462 431
rect 15416 359 15422 393
rect 15456 359 15462 393
rect 15416 321 15462 359
rect 15416 287 15422 321
rect 15456 287 15462 321
rect 15416 249 15462 287
rect 15416 215 15422 249
rect 15456 215 15462 249
rect 15416 177 15462 215
rect 2482 146 2540 160
rect 142 130 204 144
rect 142 96 156 130
rect 190 96 204 130
rect 142 -76 204 96
rect 818 120 876 130
rect 818 86 830 120
rect 864 86 876 120
rect 818 40 876 86
rect 2482 112 2494 146
rect 2528 112 2540 146
rect 2482 40 2540 112
rect 2774 130 2836 144
rect 2774 96 2788 130
rect 2822 96 2836 130
rect 5438 130 5496 144
rect 818 24 2544 40
rect 818 -10 1664 24
rect 1698 -10 2544 24
rect 818 -20 2544 -10
rect 2774 -15 2836 96
rect 1700 -45 1774 -20
rect 142 -126 206 -76
rect 1700 -97 1711 -45
rect 1763 -97 1774 -45
rect 2774 -67 2779 -15
rect 2831 -67 2836 -15
rect 2774 -82 2836 -67
rect 3098 114 3160 128
rect 3098 80 3112 114
rect 3146 80 3160 114
rect 3098 -76 3160 80
rect 3774 104 3832 114
rect 3774 70 3786 104
rect 3820 70 3832 104
rect 3774 24 3832 70
rect 5438 96 5450 130
rect 5484 96 5496 130
rect 8468 130 8526 144
rect 15416 143 15422 177
rect 15456 143 15462 177
rect 5438 24 5496 96
rect 5730 122 5790 124
rect 5730 114 5792 122
rect 5730 80 5744 114
rect 5778 80 5792 114
rect 3774 13 5500 24
rect 3774 -21 4665 13
rect 4699 -21 5500 13
rect 3774 -23 5500 -21
rect 3774 -36 4871 -23
rect 4856 -75 4871 -36
rect 4923 -36 5500 -23
rect 5730 -11 5792 80
rect 4923 -75 4938 -36
rect 1700 -98 1774 -97
rect 3098 -126 3162 -76
rect 4856 -80 4938 -75
rect 5730 -63 5735 -11
rect 5787 -63 5792 -11
rect 5730 -78 5792 -63
rect 6128 114 6190 126
rect 6128 80 6142 114
rect 6176 80 6190 114
rect 6128 -78 6190 80
rect 6804 104 6862 114
rect 6804 70 6816 104
rect 6850 70 6862 104
rect 6804 24 6862 70
rect 8468 96 8480 130
rect 8514 96 8526 130
rect 11556 128 11614 142
rect 8468 24 8526 96
rect 8760 122 8820 124
rect 8760 114 8822 122
rect 8760 80 8774 114
rect 8808 80 8822 114
rect 6804 15 8530 24
rect 6804 -19 7665 15
rect 7699 -13 8530 15
rect 7699 -19 7837 -13
rect 6804 -36 7837 -19
rect 7822 -65 7837 -36
rect 7889 -36 8530 -13
rect 8760 -25 8822 80
rect 7889 -65 7904 -36
rect 7822 -70 7904 -65
rect 6126 -126 6190 -78
rect 8760 -77 8765 -25
rect 8817 -77 8822 -25
rect 8760 -92 8822 -77
rect 9214 112 9276 128
rect 9214 78 9230 112
rect 9264 78 9276 112
rect 9214 -76 9276 78
rect 9892 102 9950 112
rect 9892 68 9904 102
rect 9938 68 9950 102
rect 9892 22 9950 68
rect 11556 94 11568 128
rect 11602 94 11614 128
rect 11556 22 11614 94
rect 11848 112 11910 122
rect 11848 78 11862 112
rect 11896 78 11910 112
rect 9892 11 11618 22
rect 9892 -23 10663 11
rect 10697 -23 11618 11
rect 9892 -34 11618 -23
rect 9892 -38 10945 -34
rect 9214 -126 9278 -76
rect 10930 -86 10945 -38
rect 10997 -38 11618 -34
rect 11848 -25 11910 78
rect 10997 -86 11012 -38
rect 10930 -96 11012 -86
rect 11848 -77 11853 -25
rect 11905 -77 11910 -25
rect 11848 -92 11910 -77
rect 12346 86 12464 104
rect 14712 102 14770 116
rect 12346 52 12386 86
rect 12420 52 12464 86
rect 12346 -126 12464 52
rect 13048 76 13106 86
rect 13048 42 13060 76
rect 13094 42 13106 76
rect 13048 -4 13106 42
rect 14712 68 14724 102
rect 14758 68 14770 102
rect 15416 100 15462 143
rect 15504 1257 15550 1300
rect 15504 1223 15510 1257
rect 15544 1223 15550 1257
rect 15504 1185 15550 1223
rect 15504 1151 15510 1185
rect 15544 1151 15550 1185
rect 15504 1113 15550 1151
rect 15504 1079 15510 1113
rect 15544 1079 15550 1113
rect 15504 1041 15550 1079
rect 15504 1007 15510 1041
rect 15544 1007 15550 1041
rect 15504 969 15550 1007
rect 15504 935 15510 969
rect 15544 935 15550 969
rect 15504 897 15550 935
rect 15504 863 15510 897
rect 15544 863 15550 897
rect 15504 825 15550 863
rect 15504 791 15510 825
rect 15544 791 15550 825
rect 15504 753 15550 791
rect 15504 719 15510 753
rect 15544 719 15550 753
rect 15504 681 15550 719
rect 15504 647 15510 681
rect 15544 647 15550 681
rect 15504 609 15550 647
rect 15504 575 15510 609
rect 15544 575 15550 609
rect 15504 537 15550 575
rect 15504 503 15510 537
rect 15544 503 15550 537
rect 15504 465 15550 503
rect 15504 431 15510 465
rect 15544 431 15550 465
rect 15504 393 15550 431
rect 15504 359 15510 393
rect 15544 359 15550 393
rect 15504 321 15550 359
rect 15504 287 15510 321
rect 15544 287 15550 321
rect 15504 249 15550 287
rect 15504 215 15510 249
rect 15544 215 15550 249
rect 15504 177 15550 215
rect 15504 143 15510 177
rect 15544 143 15550 177
rect 15504 100 15550 143
rect 14712 -4 14770 68
rect 15002 86 15064 98
rect 15002 52 15018 86
rect 15052 52 15064 86
rect 13048 -15 14774 -4
rect 13048 -49 13965 -15
rect 13999 -45 14774 -15
rect 13999 -49 14121 -45
rect 13048 -64 14121 -49
rect 14106 -97 14121 -64
rect 14173 -64 14774 -45
rect 14173 -97 14188 -64
rect 14106 -104 14188 -97
rect 15002 -66 15064 52
rect 15322 52 15554 64
rect 15322 18 15510 52
rect 15544 18 15554 52
rect 15322 2 15554 18
rect 15322 -66 15384 2
rect -564 -280 12464 -126
rect 15002 -128 15384 -66
rect 15320 -258 15384 -128
rect 15698 -258 15760 3726
rect 15320 -320 15760 -258
rect 15320 -400 15384 -320
rect 2794 -442 15384 -400
rect 2794 -456 11746 -442
rect 2794 -458 5634 -456
rect 2794 -518 2884 -458
rect 2946 -516 5634 -458
rect 5696 -460 11746 -456
rect 5696 -512 8672 -460
rect 8734 -502 11746 -460
rect 11808 -502 15384 -442
rect 8734 -512 15384 -502
rect 5696 -516 15384 -512
rect 2946 -518 15384 -516
rect 2794 -570 15384 -518
<< via1 >>
rect 1748 7820 1840 7926
rect 1770 6895 1822 6947
rect 2893 6757 2945 6809
rect 4688 6875 4740 6927
rect 5923 6751 5975 6803
rect 7688 6882 7740 6934
rect 8905 6747 8957 6799
rect 10758 6870 10810 6922
rect 12055 6749 12107 6801
rect 13953 6847 14005 6899
rect 14855 6717 14907 6769
rect 15603 6293 15655 6345
rect -1896 3354 -1782 3462
rect 2101 3735 2153 3787
rect 4933 3717 4985 3769
rect 3663 3253 3715 3305
rect 1409 2961 1461 3013
rect 10023 3715 10075 3767
rect 7127 3427 7179 3479
rect 5605 3163 5657 3215
rect 7286 3092 7374 3158
rect 2570 2540 2622 2592
rect 11064 3706 11150 3780
rect 8682 3592 8752 3676
rect 10409 3419 10461 3471
rect 8746 3352 8850 3408
rect 13081 3419 13133 3471
rect 13436 3412 13498 3464
rect 15336 3732 15398 3794
rect 5570 2540 5622 2592
rect 8571 2545 8623 2597
rect 11570 2516 11622 2568
rect 15456 1596 15538 1692
rect 1711 -97 1763 -45
rect 2779 -67 2831 -15
rect 4871 -75 4923 -23
rect 5735 -63 5787 -11
rect 7837 -65 7889 -13
rect 8765 -77 8817 -25
rect 10945 -86 10997 -34
rect 11853 -77 11905 -25
rect 14121 -97 14173 -45
rect 2884 -518 2946 -458
rect 5634 -516 5696 -456
rect 8672 -512 8734 -460
rect 11746 -502 11808 -442
<< metal2 >>
rect 1768 7936 1826 7944
rect 1748 7926 1840 7936
rect 1748 7810 1840 7820
rect 1768 7040 1826 7810
rect 2814 7344 15262 7564
rect 1768 6947 1824 7040
rect 1768 6895 1770 6947
rect 1822 6895 1824 6947
rect 1768 6882 1824 6895
rect 2888 6809 2950 7344
rect 4678 7173 4750 7190
rect 4678 7117 4686 7173
rect 4742 7117 4750 7173
rect 4678 6927 4750 7117
rect 4678 6875 4688 6927
rect 4740 6875 4750 6927
rect 4678 6858 4750 6875
rect 2888 6757 2893 6809
rect 2945 6757 2950 6809
rect 2888 6742 2950 6757
rect 5918 6803 5980 7344
rect 7672 7238 7756 7264
rect 7672 7182 7686 7238
rect 7742 7182 7756 7238
rect 7672 6934 7756 7182
rect 7672 6882 7688 6934
rect 7740 6882 7756 6934
rect 7672 6854 7756 6882
rect 5918 6751 5923 6803
rect 5975 6751 5980 6803
rect 5918 6738 5980 6751
rect 8900 6799 8962 7344
rect 10740 7202 10828 7228
rect 10740 7146 10756 7202
rect 10812 7146 10828 7202
rect 10740 6922 10828 7146
rect 10740 6870 10758 6922
rect 10810 6870 10828 6922
rect 10740 6842 10828 6870
rect 8900 6747 8905 6799
rect 8957 6747 8962 6799
rect 8900 6732 8962 6747
rect 12050 6801 12112 7344
rect 13932 7135 14026 7164
rect 13932 7079 13951 7135
rect 14007 7079 14026 7135
rect 13932 6899 14026 7079
rect 13932 6847 13953 6899
rect 14005 6847 14026 6899
rect 13932 6816 14026 6847
rect 12050 6749 12055 6801
rect 12107 6749 12112 6801
rect 12050 6734 12112 6749
rect 14850 6769 14912 7344
rect 14850 6717 14855 6769
rect 14907 6717 14912 6769
rect 14850 6702 14912 6717
rect 2096 3787 2158 3802
rect 2096 3735 2101 3787
rect 2153 3735 2158 3787
rect 2096 3484 2158 3735
rect 4928 3769 4990 3784
rect 4928 3717 4933 3769
rect 4985 3717 4990 3769
rect 4928 3666 4990 3717
rect 10018 3767 10080 3782
rect 10018 3715 10023 3767
rect 10075 3715 10080 3767
rect 8682 3676 8752 3686
rect 4928 3664 5082 3666
rect 5484 3664 8682 3666
rect 4928 3646 8682 3664
rect 4928 3604 5364 3646
rect 5458 3604 8682 3646
rect 8682 3582 8752 3592
rect 5364 3556 5458 3566
rect 2720 3490 2824 3500
rect -1896 3462 -1782 3472
rect 2096 3422 2720 3484
rect 2824 3479 7194 3484
rect 2824 3427 7127 3479
rect 7179 3427 7194 3479
rect 2824 3422 7194 3427
rect 2720 3408 2824 3418
rect 8746 3408 8850 3418
rect -1896 3344 -1782 3354
rect 8746 3342 8850 3352
rect 10018 3310 10080 3715
rect 11064 3780 11150 3790
rect 11064 3696 11150 3706
rect 10394 3471 13148 3476
rect 10394 3419 10409 3471
rect 10461 3419 13081 3471
rect 13133 3419 13148 3471
rect 10394 3414 13148 3419
rect 13436 3464 13498 3474
rect 3648 3305 10080 3310
rect 3648 3253 3663 3305
rect 3715 3253 10080 3305
rect 3648 3248 10080 3253
rect 1404 3215 5680 3220
rect 1404 3163 5605 3215
rect 5657 3163 5680 3215
rect 1404 3158 5680 3163
rect 7286 3158 7374 3168
rect 1404 3013 1466 3158
rect 13436 3156 13498 3412
rect 7374 3094 13498 3156
rect 7286 3082 7374 3092
rect 1404 2961 1409 3013
rect 1461 2961 1466 3013
rect 1404 2946 1466 2961
rect 2540 2594 2828 2612
rect 2540 2592 2744 2594
rect 2540 2540 2570 2592
rect 2622 2540 2744 2592
rect 2540 2538 2744 2540
rect 2800 2538 2828 2594
rect 2540 2520 2828 2538
rect 5356 2594 5652 2612
rect 5356 2538 5384 2594
rect 5440 2592 5652 2594
rect 5440 2540 5570 2592
rect 5622 2540 5652 2592
rect 5440 2538 5652 2540
rect 5356 2520 5652 2538
rect 8540 2599 8856 2618
rect 8540 2597 8771 2599
rect 8540 2545 8571 2597
rect 8623 2545 8771 2597
rect 8540 2543 8771 2545
rect 8827 2543 8856 2599
rect 8540 2524 8856 2543
rect 11540 2570 11836 2588
rect 11540 2568 11752 2570
rect 11540 2516 11570 2568
rect 11622 2516 11752 2568
rect 11540 2514 11752 2516
rect 11808 2514 11836 2570
rect 11540 2496 11836 2514
rect 15056 1746 15262 7344
rect 15592 6653 15666 6672
rect 15592 6597 15601 6653
rect 15657 6597 15666 6653
rect 15592 6345 15666 6597
rect 15592 6293 15603 6345
rect 15655 6293 15666 6345
rect 15592 6272 15666 6293
rect 15336 3794 15398 3804
rect 15336 3676 15398 3732
rect 15336 3614 15946 3676
rect 15056 1692 15548 1746
rect 15056 1596 15456 1692
rect 15538 1596 15548 1692
rect 15056 1574 15548 1596
rect 2764 -15 2946 -10
rect 1706 -45 1768 -30
rect 1706 -97 1711 -45
rect 1763 -97 1768 -45
rect 2764 -67 2779 -15
rect 2831 -67 2946 -15
rect 2764 -72 2946 -67
rect 1706 -223 1768 -97
rect 1706 -279 1709 -223
rect 1765 -279 1768 -223
rect 1706 -292 1768 -279
rect 2884 -458 2946 -72
rect 4866 -23 4928 -8
rect 4866 -75 4871 -23
rect 4923 -75 4928 -23
rect 4866 -237 4928 -75
rect 4866 -293 4869 -237
rect 4925 -293 4928 -237
rect 4866 -306 4928 -293
rect 5634 -11 5802 -6
rect 5634 -63 5735 -11
rect 5787 -63 5802 -11
rect 5634 -68 5802 -63
rect 7832 -13 7894 2
rect 7832 -65 7837 -13
rect 7889 -65 7894 -13
rect 2884 -528 2946 -518
rect 5634 -456 5696 -68
rect 7832 -225 7894 -65
rect 7832 -281 7835 -225
rect 7891 -281 7894 -225
rect 7832 -294 7894 -281
rect 8672 -25 8832 -20
rect 8672 -77 8765 -25
rect 8817 -77 8832 -25
rect 8672 -82 8832 -77
rect 10940 -34 11002 -14
rect 5634 -526 5696 -516
rect 8672 -460 8734 -82
rect 10940 -86 10945 -34
rect 10997 -86 11002 -34
rect 10940 -238 11002 -86
rect 10940 -294 10943 -238
rect 10999 -294 11002 -238
rect 10940 -312 11002 -294
rect 11746 -25 11920 -20
rect 11746 -77 11853 -25
rect 11905 -77 11920 -25
rect 11746 -82 11920 -77
rect 14116 -45 14178 -28
rect 11746 -442 11808 -82
rect 14116 -97 14121 -45
rect 14173 -97 14178 -45
rect 15882 -60 15946 3614
rect 14116 -177 14178 -97
rect 14116 -233 14119 -177
rect 14175 -233 14178 -177
rect 15576 -116 15946 -60
rect 15576 -184 15626 -116
rect 14116 -248 14178 -233
rect 15572 -194 15630 -184
rect 15572 -250 15573 -194
rect 15629 -250 15630 -194
rect 15572 -260 15630 -250
rect 11746 -512 11808 -502
rect 8672 -522 8734 -512
<< via2 >>
rect 1748 7820 1840 7926
rect 4686 7117 4742 7173
rect 7686 7182 7742 7238
rect 10756 7146 10812 7202
rect 13951 7079 14007 7135
rect 5364 3566 5458 3646
rect -1896 3354 -1782 3462
rect 2720 3418 2824 3490
rect 8746 3352 8850 3408
rect 11064 3706 11150 3780
rect 2744 2538 2800 2594
rect 5384 2538 5440 2594
rect 8771 2543 8827 2599
rect 11752 2514 11808 2570
rect 15601 6597 15657 6653
rect 15456 1596 15538 1692
rect 1709 -279 1765 -223
rect 4869 -293 4925 -237
rect 7835 -281 7891 -225
rect 10943 -294 10999 -238
rect 14119 -233 14175 -177
rect 15573 -250 15629 -194
<< metal3 >>
rect 1738 7926 1850 7931
rect 1738 7820 1748 7926
rect 1840 7820 1850 7926
rect 1738 7815 1850 7820
rect 4862 7632 4968 7642
rect 4862 7568 4883 7632
rect 4947 7568 4968 7632
rect 4862 7558 4968 7568
rect 7910 7601 8028 7618
rect 4872 7188 4958 7558
rect 7910 7537 7937 7601
rect 8001 7537 8028 7601
rect 14298 7604 14422 7624
rect 7910 7520 8028 7537
rect 11076 7580 11196 7598
rect 7920 7260 8018 7520
rect 11076 7516 11104 7580
rect 11168 7516 11196 7580
rect 14298 7540 14328 7604
rect 14392 7540 14422 7604
rect 14298 7520 14422 7540
rect 11076 7498 11196 7516
rect 7746 7259 8018 7260
rect 4660 7173 4958 7188
rect 4660 7117 4686 7173
rect 4742 7117 4958 7173
rect 7662 7238 8018 7259
rect 7662 7182 7686 7238
rect 7742 7182 8018 7238
rect 11086 7224 11186 7498
rect 10830 7223 11186 7224
rect 7662 7162 8018 7182
rect 10730 7202 11186 7223
rect 7662 7161 7766 7162
rect 10730 7146 10756 7202
rect 10812 7146 11186 7202
rect 14308 7160 14412 7520
rect 13932 7159 14412 7160
rect 10730 7125 11186 7146
rect 10830 7124 11186 7125
rect 13922 7135 14412 7159
rect 4660 7102 4958 7117
rect 13922 7079 13951 7135
rect 14007 7079 14412 7135
rect 13922 7056 14412 7079
rect 13922 7055 14036 7056
rect 14308 7054 14412 7056
rect 15570 7063 15688 7080
rect 15570 6999 15597 7063
rect 15661 6999 15688 7063
rect 15570 6982 15688 6999
rect 15580 6653 15678 6982
rect 15580 6597 15601 6653
rect 15657 6597 15678 6653
rect 15580 6576 15678 6597
rect 11054 3780 11160 3785
rect 11726 3780 11832 3782
rect 11054 3706 11064 3780
rect 11150 3706 11832 3780
rect 11054 3701 11160 3706
rect 5360 3651 5464 3672
rect 5354 3646 5468 3651
rect 5354 3566 5364 3646
rect 5458 3566 5468 3646
rect 5354 3561 5468 3566
rect 2710 3490 2834 3495
rect -1906 3462 -1772 3467
rect -1906 3354 -1896 3462
rect -1782 3354 -1772 3462
rect 2710 3418 2720 3490
rect 2824 3418 2834 3490
rect 2710 3413 2834 3418
rect -1906 3349 -1772 3354
rect 2720 2616 2824 3413
rect 2721 2594 2823 2616
rect 2721 2538 2744 2594
rect 2800 2538 2823 2594
rect 5360 2594 5464 3561
rect 8746 3413 8852 3414
rect 8736 3408 8860 3413
rect 8736 3352 8746 3408
rect 8850 3352 8860 3408
rect 8736 3347 8860 3352
rect 8746 2624 8852 3347
rect 5360 2582 5384 2594
rect 2721 2510 2823 2538
rect 5361 2538 5384 2582
rect 5440 2582 5464 2594
rect 8747 2599 8851 2624
rect 5440 2538 5463 2582
rect 5361 2510 5463 2538
rect 8747 2543 8771 2599
rect 8827 2543 8851 2599
rect 11728 2590 11832 3706
rect 8747 2514 8851 2543
rect 11729 2570 11831 2590
rect 11729 2514 11752 2570
rect 11808 2514 11831 2570
rect 11729 2486 11831 2514
rect 15446 1694 15548 1697
rect 15444 1692 15884 1694
rect 15444 1596 15456 1692
rect 15538 1677 15884 1692
rect 15538 1613 15793 1677
rect 15857 1613 15884 1677
rect 15538 1596 15884 1613
rect 15446 1591 15548 1596
rect 14102 -177 14366 -162
rect 1688 -223 1916 -202
rect 1688 -279 1709 -223
rect 1765 -279 1916 -223
rect 1688 -296 1916 -279
rect 1822 -361 1916 -296
rect 4852 -237 5070 -224
rect 4852 -293 4869 -237
rect 4925 -293 5070 -237
rect 4852 -312 5070 -293
rect 7806 -225 8070 -210
rect 7806 -281 7835 -225
rect 7891 -281 8070 -225
rect 7806 -302 8070 -281
rect 1821 -368 1916 -361
rect 1821 -386 1915 -368
rect 1821 -450 1836 -386
rect 1900 -450 1915 -386
rect 1821 -475 1915 -450
rect 4982 -643 5070 -312
rect 7978 -583 8070 -302
rect 10924 -238 11126 -222
rect 10924 -294 10943 -238
rect 10999 -294 11126 -238
rect 14102 -233 14119 -177
rect 14175 -233 14366 -177
rect 14102 -248 14366 -233
rect 10924 -318 11126 -294
rect 4981 -644 5070 -643
rect 7969 -607 8073 -583
rect 4981 -665 5069 -644
rect 4981 -729 4993 -665
rect 5057 -729 5069 -665
rect 7969 -671 7989 -607
rect 8053 -671 8073 -607
rect 11032 -607 11126 -318
rect 14282 -598 14366 -248
rect 15542 -194 15654 -178
rect 15542 -250 15573 -194
rect 15629 -250 15654 -194
rect 15542 -330 15654 -250
rect 15532 -345 15664 -330
rect 15532 -409 15566 -345
rect 15630 -409 15664 -345
rect 15532 -424 15664 -409
rect 11032 -608 11127 -607
rect 7969 -695 8073 -671
rect 11033 -632 11127 -608
rect 11033 -696 11048 -632
rect 11112 -696 11127 -632
rect 14283 -613 14363 -598
rect 14283 -677 14291 -613
rect 14355 -677 14363 -613
rect 14283 -695 14363 -677
rect 11033 -721 11127 -696
rect 4981 -751 5069 -729
<< via3 >>
rect 1748 7820 1840 7926
rect 4883 7568 4947 7632
rect 7937 7537 8001 7601
rect 11104 7516 11168 7580
rect 14328 7540 14392 7604
rect 15597 6999 15661 7063
rect -1896 3354 -1782 3462
rect 15793 1613 15857 1677
rect 1836 -450 1900 -386
rect 4993 -729 5057 -665
rect 7989 -671 8053 -607
rect 15566 -409 15630 -345
rect 11048 -696 11112 -632
rect 14291 -677 14355 -613
<< metal4 >>
rect 1684 7926 15998 8098
rect 1684 7820 1748 7926
rect 1840 7820 15998 7926
rect 1684 7792 15998 7820
rect 1684 7790 1812 7792
rect 2002 7790 15998 7792
rect 4864 7632 4964 7790
rect 7916 7706 8020 7790
rect 4864 7568 4883 7632
rect 4947 7568 4964 7632
rect 4864 7552 4964 7568
rect 7918 7601 8020 7706
rect 7918 7537 7937 7601
rect 8001 7537 8020 7601
rect 7918 7518 8020 7537
rect 11084 7580 11188 7790
rect 11084 7516 11104 7580
rect 11168 7516 11188 7580
rect 14306 7604 14414 7790
rect 14306 7540 14328 7604
rect 14392 7540 14414 7604
rect 14306 7518 14414 7540
rect 11084 7496 11188 7516
rect 15578 7063 15680 7790
rect 15578 6999 15597 7063
rect 15661 6999 15680 7063
rect 15578 6980 15680 6999
rect -2630 3526 -1690 3576
rect -2630 3462 -1688 3526
rect -2630 3354 -1896 3462
rect -1782 3354 -1688 3462
rect -2630 3302 -1688 3354
rect -2630 3278 -1690 3302
rect 16036 1764 16284 1770
rect 16036 1696 16042 1764
rect 15774 1677 16042 1696
rect 15774 1613 15793 1677
rect 15857 1613 16042 1677
rect 15774 1596 16042 1613
rect 15775 1595 15875 1596
rect 16036 1528 16042 1596
rect 16278 1528 16284 1764
rect 16036 1522 16284 1528
rect 15541 -345 15655 -329
rect 1812 -386 2086 -366
rect 1812 -450 1836 -386
rect 1900 -450 2086 -386
rect 15541 -409 15566 -345
rect 15630 -409 15655 -345
rect 15541 -425 15655 -409
rect 1812 -470 2086 -450
rect 1982 -826 2086 -470
rect 7968 -607 8232 -592
rect 4976 -665 5228 -648
rect 4976 -729 4993 -665
rect 5057 -729 5228 -665
rect 7968 -671 7989 -607
rect 8053 -671 8232 -607
rect 7968 -686 8232 -671
rect 4976 -748 5228 -729
rect 5128 -826 5228 -748
rect 8126 -826 8232 -686
rect 11028 -632 11290 -612
rect 11028 -696 11048 -632
rect 11112 -696 11290 -632
rect 14280 -613 14520 -602
rect 14280 -677 14291 -613
rect 14355 -677 14520 -613
rect 14280 -688 14520 -677
rect 11028 -714 11290 -696
rect 11196 -826 11290 -714
rect 14436 -826 14520 -688
rect 15542 -826 15654 -425
rect 1900 -1158 15656 -826
<< via4 >>
rect 16042 1528 16278 1764
<< metal5 >>
rect 15972 1764 16782 1860
rect 15972 1528 16042 1764
rect 16278 1528 16782 1764
rect 15972 1432 16782 1528
<< labels >>
rlabel metal4 7152 7932 7152 7932 1 VP
port 3 n
rlabel metal4 11374 -976 11374 -976 1 VN
port 5 n
rlabel metal5 16574 1566 16574 1566 1 VCT
port 4 n
rlabel metal1 13934 3282 13934 3282 1 OUT
port 2 n
rlabel metal4 -2578 3420 -2578 3420 1 VB
port 1 n
<< end >>
