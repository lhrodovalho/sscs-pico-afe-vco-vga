magic
tech sky130A
timestamp 1638390070
<< psubdiff >>
rect -6440 1800 -6360 1840
rect 7360 1800 7440 1840
rect -6440 1760 -6400 1800
rect -6440 720 -6400 760
rect 7400 1760 7440 1800
rect 7400 720 7440 760
rect -6440 680 -6360 720
rect 7360 680 7440 720
<< psubdiffcont >>
rect -6360 1800 7360 1840
rect -6440 760 -6400 1760
rect 7400 760 7440 1760
rect -6360 680 7360 720
<< locali >>
rect -6440 1800 -6360 1840
rect 7360 1800 7440 1840
rect -6440 1760 -6400 1800
rect -6440 720 -6400 760
rect 7400 1760 7440 1800
rect 7400 720 7440 760
rect -6440 680 -6360 720
rect 7360 680 7440 720
<< metal3 >>
rect -6360 1756 -6160 1760
rect -6360 1724 -6356 1756
rect -6324 1724 -6276 1756
rect -6244 1724 -6196 1756
rect -6164 1724 -6160 1756
rect -6360 1596 -6160 1724
rect 7160 1756 7360 1760
rect 7160 1724 7164 1756
rect 7196 1724 7244 1756
rect 7276 1724 7324 1756
rect 7356 1724 7360 1756
rect -6360 1564 -6356 1596
rect -6324 1564 -6276 1596
rect -6244 1564 -6196 1596
rect -6164 1564 -6160 1596
rect -6360 1436 -6160 1564
rect -5520 1676 -5480 1680
rect -5520 1644 -5516 1676
rect -5484 1644 -5480 1676
rect -6360 1404 -6356 1436
rect -6324 1404 -6276 1436
rect -6244 1404 -6196 1436
rect -6164 1404 -6160 1436
rect -6360 1116 -6160 1404
rect -6360 1084 -6356 1116
rect -6324 1084 -6276 1116
rect -6244 1084 -6196 1116
rect -6164 1084 -6160 1116
rect -6360 956 -6160 1084
rect -6120 1436 -6080 1440
rect -6120 1404 -6116 1436
rect -6084 1404 -6080 1436
rect -6120 1116 -6080 1404
rect -5520 1360 -5480 1644
rect -4320 1676 -4280 1680
rect -4320 1644 -4316 1676
rect -4284 1644 -4280 1676
rect -4920 1436 -4880 1440
rect -4920 1404 -4916 1436
rect -4884 1404 -4880 1436
rect -6040 1160 -4960 1360
rect -6120 1084 -6116 1116
rect -6084 1084 -6080 1116
rect -6120 1080 -6080 1084
rect -6360 924 -6356 956
rect -6324 924 -6276 956
rect -6244 924 -6196 956
rect -6164 924 -6160 956
rect -6360 796 -6160 924
rect -5520 876 -5480 1160
rect -4920 1116 -4880 1404
rect -4320 1360 -4280 1644
rect -3120 1676 -3080 1680
rect -3120 1644 -3116 1676
rect -3084 1644 -3080 1676
rect -3720 1436 -3680 1440
rect -3720 1404 -3716 1436
rect -3684 1404 -3680 1436
rect -4840 1160 -3760 1360
rect -4920 1084 -4916 1116
rect -4884 1084 -4880 1116
rect -4920 1080 -4880 1084
rect -5520 844 -5516 876
rect -5484 844 -5480 876
rect -5520 840 -5480 844
rect -4320 876 -4280 1160
rect -3720 1116 -3680 1404
rect -3120 1360 -3080 1644
rect -1920 1676 -1880 1680
rect -1920 1644 -1916 1676
rect -1884 1644 -1880 1676
rect -2520 1436 -2480 1440
rect -2520 1404 -2516 1436
rect -2484 1404 -2480 1436
rect -3640 1160 -2560 1360
rect -3720 1084 -3716 1116
rect -3684 1084 -3680 1116
rect -3720 1080 -3680 1084
rect -4320 844 -4316 876
rect -4284 844 -4280 876
rect -4320 840 -4280 844
rect -3120 876 -3080 1160
rect -2520 1116 -2480 1404
rect -1920 1360 -1880 1644
rect -720 1676 -680 1680
rect -720 1644 -716 1676
rect -684 1644 -680 1676
rect -1320 1436 -1280 1440
rect -1320 1404 -1316 1436
rect -1284 1404 -1280 1436
rect -2440 1160 -1360 1360
rect -2520 1084 -2516 1116
rect -2484 1084 -2480 1116
rect -2520 1080 -2480 1084
rect -3120 844 -3116 876
rect -3084 844 -3080 876
rect -3120 840 -3080 844
rect -1920 876 -1880 1160
rect -1320 1116 -1280 1404
rect -720 1360 -680 1644
rect 1680 1676 1720 1680
rect 1680 1644 1684 1676
rect 1716 1644 1720 1676
rect 480 1516 520 1520
rect 480 1484 484 1516
rect 516 1484 520 1516
rect -120 1436 -80 1440
rect -120 1404 -116 1436
rect -84 1404 -80 1436
rect -1240 1160 -160 1360
rect -1320 1084 -1316 1116
rect -1284 1084 -1280 1116
rect -1320 1080 -1280 1084
rect -1920 844 -1916 876
rect -1884 844 -1880 876
rect -1920 840 -1880 844
rect -720 876 -680 1160
rect -120 1116 -80 1404
rect 480 1360 520 1484
rect 1080 1436 1120 1440
rect 1080 1404 1084 1436
rect 1116 1404 1120 1436
rect -40 1160 1040 1360
rect -120 1084 -116 1116
rect -84 1084 -80 1116
rect -120 1080 -80 1084
rect 480 1036 520 1160
rect 1080 1116 1120 1404
rect 1680 1360 1720 1644
rect 2880 1676 2920 1680
rect 2880 1644 2884 1676
rect 2916 1644 2920 1676
rect 2280 1436 2320 1440
rect 2280 1404 2284 1436
rect 2316 1404 2320 1436
rect 1160 1160 2240 1360
rect 1080 1084 1084 1116
rect 1116 1084 1120 1116
rect 1080 1080 1120 1084
rect 480 1004 484 1036
rect 516 1004 520 1036
rect 480 1000 520 1004
rect -720 844 -716 876
rect -684 844 -680 876
rect -720 840 -680 844
rect 1680 876 1720 1160
rect 2280 1116 2320 1404
rect 2880 1360 2920 1644
rect 4080 1676 4120 1680
rect 4080 1644 4084 1676
rect 4116 1644 4120 1676
rect 3480 1436 3520 1440
rect 3480 1404 3484 1436
rect 3516 1404 3520 1436
rect 2360 1160 3440 1360
rect 2280 1084 2284 1116
rect 2316 1084 2320 1116
rect 2280 1080 2320 1084
rect 1680 844 1684 876
rect 1716 844 1720 876
rect 1680 840 1720 844
rect 2880 876 2920 1160
rect 3480 1116 3520 1404
rect 4080 1360 4120 1644
rect 5280 1676 5320 1680
rect 5280 1644 5284 1676
rect 5316 1644 5320 1676
rect 4680 1436 4720 1440
rect 4680 1404 4684 1436
rect 4716 1404 4720 1436
rect 3560 1160 4640 1360
rect 3480 1084 3484 1116
rect 3516 1084 3520 1116
rect 3480 1080 3520 1084
rect 2880 844 2884 876
rect 2916 844 2920 876
rect 2880 840 2920 844
rect 4080 876 4120 1160
rect 4680 1116 4720 1404
rect 5280 1360 5320 1644
rect 6480 1676 6520 1680
rect 6480 1644 6484 1676
rect 6516 1644 6520 1676
rect 5880 1436 5920 1440
rect 5880 1404 5884 1436
rect 5916 1404 5920 1436
rect 4760 1160 5840 1360
rect 4680 1084 4684 1116
rect 4716 1084 4720 1116
rect 4680 1080 4720 1084
rect 4080 844 4084 876
rect 4116 844 4120 876
rect 4080 840 4120 844
rect 5280 876 5320 1160
rect 5880 1116 5920 1404
rect 6480 1360 6520 1644
rect 7160 1676 7360 1724
rect 7160 1644 7164 1676
rect 7196 1644 7244 1676
rect 7276 1644 7324 1676
rect 7356 1644 7360 1676
rect 7160 1596 7360 1644
rect 7160 1564 7164 1596
rect 7196 1564 7244 1596
rect 7276 1564 7324 1596
rect 7356 1564 7360 1596
rect 7160 1516 7360 1564
rect 7160 1484 7164 1516
rect 7196 1484 7244 1516
rect 7276 1484 7324 1516
rect 7356 1484 7360 1516
rect 7080 1436 7120 1440
rect 7080 1404 7084 1436
rect 7116 1404 7120 1436
rect 5960 1160 7040 1360
rect 5880 1084 5884 1116
rect 5916 1084 5920 1116
rect 5880 1080 5920 1084
rect 5280 844 5284 876
rect 5316 844 5320 876
rect 5280 840 5320 844
rect 6480 876 6520 1160
rect 7080 1116 7120 1404
rect 7080 1084 7084 1116
rect 7116 1084 7120 1116
rect 7080 1080 7120 1084
rect 7160 1436 7360 1484
rect 7160 1404 7164 1436
rect 7196 1404 7244 1436
rect 7276 1404 7324 1436
rect 7356 1404 7360 1436
rect 7160 1116 7360 1404
rect 7160 1084 7164 1116
rect 7196 1084 7244 1116
rect 7276 1084 7324 1116
rect 7356 1084 7360 1116
rect 6480 844 6484 876
rect 6516 844 6520 876
rect 6480 840 6520 844
rect 7160 1036 7360 1084
rect 7160 1004 7164 1036
rect 7196 1004 7244 1036
rect 7276 1004 7324 1036
rect 7356 1004 7360 1036
rect 7160 956 7360 1004
rect 7160 924 7164 956
rect 7196 924 7244 956
rect 7276 924 7324 956
rect 7356 924 7360 956
rect 7160 876 7360 924
rect 7160 844 7164 876
rect 7196 844 7244 876
rect 7276 844 7324 876
rect 7356 844 7360 876
rect -6360 764 -6356 796
rect -6324 764 -6276 796
rect -6244 764 -6196 796
rect -6164 764 -6160 796
rect -6360 760 -6160 764
rect 7160 796 7360 844
rect 7160 764 7164 796
rect 7196 764 7244 796
rect 7276 764 7324 796
rect 7356 764 7360 796
rect 7160 760 7360 764
<< via3 >>
rect -6356 1724 -6324 1756
rect -6276 1724 -6244 1756
rect -6196 1724 -6164 1756
rect 7164 1724 7196 1756
rect 7244 1724 7276 1756
rect 7324 1724 7356 1756
rect -6356 1564 -6324 1596
rect -6276 1564 -6244 1596
rect -6196 1564 -6164 1596
rect -5516 1644 -5484 1676
rect -6356 1404 -6324 1436
rect -6276 1404 -6244 1436
rect -6196 1404 -6164 1436
rect -6356 1084 -6324 1116
rect -6276 1084 -6244 1116
rect -6196 1084 -6164 1116
rect -6116 1404 -6084 1436
rect -4316 1644 -4284 1676
rect -4916 1404 -4884 1436
rect -6116 1084 -6084 1116
rect -6356 924 -6324 956
rect -6276 924 -6244 956
rect -6196 924 -6164 956
rect -3116 1644 -3084 1676
rect -3716 1404 -3684 1436
rect -4916 1084 -4884 1116
rect -5516 844 -5484 876
rect -1916 1644 -1884 1676
rect -2516 1404 -2484 1436
rect -3716 1084 -3684 1116
rect -4316 844 -4284 876
rect -716 1644 -684 1676
rect -1316 1404 -1284 1436
rect -2516 1084 -2484 1116
rect -3116 844 -3084 876
rect 1684 1644 1716 1676
rect 484 1484 516 1516
rect -116 1404 -84 1436
rect -1316 1084 -1284 1116
rect -1916 844 -1884 876
rect 1084 1404 1116 1436
rect -116 1084 -84 1116
rect 2884 1644 2916 1676
rect 2284 1404 2316 1436
rect 1084 1084 1116 1116
rect 484 1004 516 1036
rect -716 844 -684 876
rect 4084 1644 4116 1676
rect 3484 1404 3516 1436
rect 2284 1084 2316 1116
rect 1684 844 1716 876
rect 5284 1644 5316 1676
rect 4684 1404 4716 1436
rect 3484 1084 3516 1116
rect 2884 844 2916 876
rect 6484 1644 6516 1676
rect 5884 1404 5916 1436
rect 4684 1084 4716 1116
rect 4084 844 4116 876
rect 7164 1644 7196 1676
rect 7244 1644 7276 1676
rect 7324 1644 7356 1676
rect 7164 1564 7196 1596
rect 7244 1564 7276 1596
rect 7324 1564 7356 1596
rect 7164 1484 7196 1516
rect 7244 1484 7276 1516
rect 7324 1484 7356 1516
rect 7084 1404 7116 1436
rect 5884 1084 5916 1116
rect 5284 844 5316 876
rect 7084 1084 7116 1116
rect 7164 1404 7196 1436
rect 7244 1404 7276 1436
rect 7324 1404 7356 1436
rect 7164 1084 7196 1116
rect 7244 1084 7276 1116
rect 7324 1084 7356 1116
rect 6484 844 6516 876
rect 7164 1004 7196 1036
rect 7244 1004 7276 1036
rect 7324 1004 7356 1036
rect 7164 924 7196 956
rect 7244 924 7276 956
rect 7324 924 7356 956
rect 7164 844 7196 876
rect 7244 844 7276 876
rect 7324 844 7356 876
rect -6356 764 -6324 796
rect -6276 764 -6244 796
rect -6196 764 -6164 796
rect 7164 764 7196 796
rect 7244 764 7276 796
rect 7324 764 7356 796
<< mimcap >>
rect -6320 1280 -6200 1320
rect -6320 1240 -6280 1280
rect -6240 1240 -6200 1280
rect -6320 1200 -6200 1240
rect -6000 1280 -5000 1320
rect -6000 1240 -5960 1280
rect -5040 1240 -5000 1280
rect -6000 1200 -5000 1240
rect -4800 1280 -3800 1320
rect -4800 1240 -4760 1280
rect -3840 1240 -3800 1280
rect -4800 1200 -3800 1240
rect -3600 1280 -2600 1320
rect -3600 1240 -3560 1280
rect -2640 1240 -2600 1280
rect -3600 1200 -2600 1240
rect -2400 1280 -1400 1320
rect -2400 1240 -2360 1280
rect -1440 1240 -1400 1280
rect -2400 1200 -1400 1240
rect -1200 1280 -200 1320
rect -1200 1240 -1160 1280
rect -240 1240 -200 1280
rect -1200 1200 -200 1240
rect 0 1280 1000 1320
rect 0 1240 40 1280
rect 960 1240 1000 1280
rect 0 1200 1000 1240
rect 1200 1280 2200 1320
rect 1200 1240 1240 1280
rect 2160 1240 2200 1280
rect 1200 1200 2200 1240
rect 2400 1280 3400 1320
rect 2400 1240 2440 1280
rect 3360 1240 3400 1280
rect 2400 1200 3400 1240
rect 3600 1280 4600 1320
rect 3600 1240 3640 1280
rect 4560 1240 4600 1280
rect 3600 1200 4600 1240
rect 4800 1280 5800 1320
rect 4800 1240 4840 1280
rect 5760 1240 5800 1280
rect 4800 1200 5800 1240
rect 6000 1280 7000 1320
rect 6000 1240 6040 1280
rect 6960 1240 7000 1280
rect 6000 1200 7000 1240
rect 7200 1280 7320 1320
rect 7200 1240 7240 1280
rect 7280 1240 7320 1280
rect 7200 1200 7320 1240
<< mimcapcontact >>
rect -6280 1240 -6240 1280
rect -5960 1240 -5040 1280
rect -4760 1240 -3840 1280
rect -3560 1240 -2640 1280
rect -2360 1240 -1440 1280
rect -1160 1240 -240 1280
rect 40 1240 960 1280
rect 1240 1240 2160 1280
rect 2440 1240 3360 1280
rect 3640 1240 4560 1280
rect 4840 1240 5760 1280
rect 6040 1240 6960 1280
rect 7240 1240 7280 1280
<< metal4 >>
rect -6360 1756 7440 1760
rect -6360 1724 -6356 1756
rect -6324 1724 -6276 1756
rect -6244 1724 -6196 1756
rect -6164 1724 7164 1756
rect 7196 1724 7244 1756
rect 7276 1724 7324 1756
rect 7356 1724 7440 1756
rect -6360 1720 7440 1724
rect -6360 1676 7440 1680
rect -6360 1644 -5516 1676
rect -5484 1644 -4316 1676
rect -4284 1644 -3116 1676
rect -3084 1644 -1916 1676
rect -1884 1644 -716 1676
rect -684 1644 1684 1676
rect 1716 1644 2884 1676
rect 2916 1644 4084 1676
rect 4116 1644 5284 1676
rect 5316 1644 6484 1676
rect 6516 1644 7164 1676
rect 7196 1644 7244 1676
rect 7276 1644 7324 1676
rect 7356 1644 7440 1676
rect -6360 1640 7440 1644
rect -5520 1600 -5480 1640
rect -4320 1600 -4280 1640
rect -3120 1600 -3080 1640
rect -1920 1600 -1880 1640
rect -720 1600 -680 1640
rect 1680 1600 1720 1640
rect 2880 1600 2920 1640
rect 4080 1600 4120 1640
rect 5280 1600 5320 1640
rect 6480 1600 6520 1640
rect -6360 1596 7440 1600
rect -6360 1564 -6356 1596
rect -6324 1564 -6276 1596
rect -6244 1564 -6196 1596
rect -6164 1564 7164 1596
rect 7196 1564 7244 1596
rect 7276 1564 7324 1596
rect 7356 1564 7440 1596
rect -6360 1560 7440 1564
rect -5520 1520 -5480 1560
rect -4320 1520 -4280 1560
rect -3120 1520 -3080 1560
rect -1920 1520 -1880 1560
rect -720 1520 -680 1560
rect 1680 1520 1720 1560
rect 2880 1520 2920 1560
rect 4080 1520 4120 1560
rect 5280 1520 5320 1560
rect 6480 1520 6520 1560
rect -6360 1516 7440 1520
rect -6360 1484 484 1516
rect 516 1484 7164 1516
rect 7196 1484 7244 1516
rect 7276 1484 7324 1516
rect 7356 1484 7440 1516
rect -6360 1480 7440 1484
rect -5520 1440 -5480 1480
rect -4320 1440 -4280 1480
rect -3120 1440 -3080 1480
rect -1920 1440 -1880 1480
rect -720 1440 -680 1480
rect 480 1440 520 1480
rect 1680 1440 1720 1480
rect 2880 1440 2920 1480
rect 4080 1440 4120 1480
rect 5280 1440 5320 1480
rect 6480 1440 6520 1480
rect -6360 1436 7440 1440
rect -6360 1404 -6356 1436
rect -6324 1404 -6276 1436
rect -6244 1404 -6196 1436
rect -6164 1404 -6116 1436
rect -6084 1404 -4916 1436
rect -4884 1404 -3716 1436
rect -3684 1404 -2516 1436
rect -2484 1404 -1316 1436
rect -1284 1404 -116 1436
rect -84 1404 1084 1436
rect 1116 1404 2284 1436
rect 2316 1404 3484 1436
rect 3516 1404 4684 1436
rect 4716 1404 5884 1436
rect 5916 1404 7084 1436
rect 7116 1404 7164 1436
rect 7196 1404 7244 1436
rect 7276 1404 7324 1436
rect 7356 1404 7440 1436
rect -6360 1400 7440 1404
rect -6360 1360 -6320 1400
rect -6280 1360 -6240 1400
rect -6200 1360 -6160 1400
rect -6360 1280 -6160 1360
rect -6360 1240 -6280 1280
rect -6240 1240 -6160 1280
rect -6360 1160 -6160 1240
rect -6360 1120 -6320 1160
rect -6280 1120 -6240 1160
rect -6200 1120 -6160 1160
rect -6120 1120 -6080 1400
rect -5520 1360 -5480 1400
rect -6040 1280 -4960 1360
rect -6040 1240 -5960 1280
rect -5040 1240 -4960 1280
rect -6040 1160 -4960 1240
rect -5520 1120 -5480 1160
rect -4920 1120 -4880 1400
rect -4320 1360 -4280 1400
rect -4840 1280 -3760 1360
rect -4840 1240 -4760 1280
rect -3840 1240 -3760 1280
rect -4840 1160 -3760 1240
rect -4320 1120 -4280 1160
rect -3720 1120 -3680 1400
rect -3120 1360 -3080 1400
rect -3640 1280 -2560 1360
rect -3640 1240 -3560 1280
rect -2640 1240 -2560 1280
rect -3640 1160 -2560 1240
rect -3120 1120 -3080 1160
rect -2520 1120 -2480 1400
rect -1920 1360 -1880 1400
rect -2440 1280 -1360 1360
rect -2440 1240 -2360 1280
rect -1440 1240 -1360 1280
rect -2440 1160 -1360 1240
rect -1920 1120 -1880 1160
rect -1320 1120 -1280 1400
rect -720 1360 -680 1400
rect -1240 1280 -160 1360
rect -1240 1240 -1160 1280
rect -240 1240 -160 1280
rect -1240 1160 -160 1240
rect -720 1120 -680 1160
rect -120 1120 -80 1400
rect 480 1360 520 1400
rect -40 1280 1040 1360
rect -40 1240 40 1280
rect 960 1240 1040 1280
rect -40 1160 1040 1240
rect 480 1120 520 1160
rect 1080 1120 1120 1400
rect 1680 1360 1720 1400
rect 1160 1280 2240 1360
rect 1160 1240 1240 1280
rect 2160 1240 2240 1280
rect 1160 1160 2240 1240
rect 1680 1120 1720 1160
rect 2280 1120 2320 1400
rect 2880 1360 2920 1400
rect 2360 1280 3440 1360
rect 2360 1240 2440 1280
rect 3360 1240 3440 1280
rect 2360 1160 3440 1240
rect 2880 1120 2920 1160
rect 3480 1120 3520 1400
rect 4080 1360 4120 1400
rect 3560 1280 4640 1360
rect 3560 1240 3640 1280
rect 4560 1240 4640 1280
rect 3560 1160 4640 1240
rect 4080 1120 4120 1160
rect 4680 1120 4720 1400
rect 5280 1360 5320 1400
rect 4760 1280 5840 1360
rect 4760 1240 4840 1280
rect 5760 1240 5840 1280
rect 4760 1160 5840 1240
rect 5280 1120 5320 1160
rect 5880 1120 5920 1400
rect 6480 1360 6520 1400
rect 5960 1280 7040 1360
rect 5960 1240 6040 1280
rect 6960 1240 7040 1280
rect 5960 1160 7040 1240
rect 6480 1120 6520 1160
rect 7080 1120 7120 1400
rect 7160 1360 7200 1400
rect 7240 1360 7280 1400
rect 7320 1360 7360 1400
rect 7160 1280 7360 1360
rect 7160 1240 7240 1280
rect 7280 1240 7360 1280
rect 7160 1160 7360 1240
rect 7160 1120 7200 1160
rect 7240 1120 7280 1160
rect 7320 1120 7360 1160
rect -6400 1116 7440 1120
rect -6400 1084 -6356 1116
rect -6324 1084 -6276 1116
rect -6244 1084 -6196 1116
rect -6164 1084 -6116 1116
rect -6084 1084 -4916 1116
rect -4884 1084 -3716 1116
rect -3684 1084 -2516 1116
rect -2484 1084 -1316 1116
rect -1284 1084 -116 1116
rect -84 1084 1084 1116
rect 1116 1084 2284 1116
rect 2316 1084 3484 1116
rect 3516 1084 4684 1116
rect 4716 1084 5884 1116
rect 5916 1084 7084 1116
rect 7116 1084 7164 1116
rect 7196 1084 7244 1116
rect 7276 1084 7324 1116
rect 7356 1084 7440 1116
rect -6400 1080 7440 1084
rect -5520 1040 -5480 1080
rect -4320 1040 -4280 1080
rect -3120 1040 -3080 1080
rect -1920 1040 -1880 1080
rect -720 1040 -680 1080
rect 480 1040 520 1080
rect 1680 1040 1720 1080
rect 2880 1040 2920 1080
rect 4080 1040 4120 1080
rect 5280 1040 5320 1080
rect 6480 1040 6520 1080
rect -6400 1036 7440 1040
rect -6400 1004 484 1036
rect 516 1004 7164 1036
rect 7196 1004 7244 1036
rect 7276 1004 7324 1036
rect 7356 1004 7440 1036
rect -6400 1000 7440 1004
rect -5520 960 -5480 1000
rect -4320 960 -4280 1000
rect -3120 960 -3080 1000
rect -1920 960 -1880 1000
rect -720 960 -680 1000
rect 1680 960 1720 1000
rect 2880 960 2920 1000
rect 4080 960 4120 1000
rect 5280 960 5320 1000
rect 6480 960 6520 1000
rect -6400 956 7440 960
rect -6400 924 -6356 956
rect -6324 924 -6276 956
rect -6244 924 -6196 956
rect -6164 924 7164 956
rect 7196 924 7244 956
rect 7276 924 7324 956
rect 7356 924 7440 956
rect -6400 920 7440 924
rect -5520 880 -5480 920
rect -4320 880 -4280 920
rect -3120 880 -3080 920
rect -1920 880 -1880 920
rect -720 880 -680 920
rect 1680 880 1720 920
rect 2880 880 2920 920
rect 4080 880 4120 920
rect 5280 880 5320 920
rect 6480 880 6520 920
rect -6400 876 7440 880
rect -6400 844 -5516 876
rect -5484 844 -4316 876
rect -4284 844 -3116 876
rect -3084 844 -1916 876
rect -1884 844 -716 876
rect -684 844 1684 876
rect 1716 844 2884 876
rect 2916 844 4084 876
rect 4116 844 5284 876
rect 5316 844 6484 876
rect 6516 844 7164 876
rect 7196 844 7244 876
rect 7276 844 7324 876
rect 7356 844 7440 876
rect -6400 840 7440 844
rect -6400 796 7440 800
rect -6400 764 -6356 796
rect -6324 764 -6276 796
rect -6244 764 -6196 796
rect -6164 764 7164 796
rect 7196 764 7244 796
rect 7276 764 7324 796
rect 7356 764 7440 796
rect -6400 760 7440 764
<< labels >>
rlabel metal4 7400 1720 7440 1760 0 gnda
port 12 nsew
rlabel locali 7400 1800 7440 1840 0 vssa
port 13 nsew
<< end >>
