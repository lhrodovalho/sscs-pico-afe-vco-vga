magic
tech sky130A
timestamp 1638398216
<< locali >>
rect -14960 21430 -14920 21440
rect -14960 21410 -14950 21430
rect -14930 21410 -14920 21430
rect -14960 21270 -14920 21410
rect -14960 21250 -14950 21270
rect -14930 21250 -14920 21270
rect -14960 21110 -14920 21250
rect -14960 21090 -14950 21110
rect -14930 21090 -14920 21110
rect -14960 20950 -14920 21090
rect -14960 20930 -14950 20950
rect -14930 20930 -14920 20950
rect -14960 20920 -14920 20930
rect -14880 21430 -14840 21440
rect -14880 21410 -14870 21430
rect -14850 21410 -14840 21430
rect -14880 21270 -14840 21410
rect -14880 21250 -14870 21270
rect -14850 21250 -14840 21270
rect -14880 21110 -14840 21250
rect -14880 21090 -14870 21110
rect -14850 21090 -14840 21110
rect -14880 20950 -14840 21090
rect -14880 20930 -14870 20950
rect -14850 20930 -14840 20950
rect -14880 20920 -14840 20930
rect -14800 21430 -14760 21440
rect -14800 21410 -14790 21430
rect -14770 21410 -14760 21430
rect -14800 21270 -14760 21410
rect -14800 21250 -14790 21270
rect -14770 21250 -14760 21270
rect -14800 21110 -14760 21250
rect -14800 21090 -14790 21110
rect -14770 21090 -14760 21110
rect -14800 20950 -14760 21090
rect -14800 20930 -14790 20950
rect -14770 20930 -14760 20950
rect -14800 20920 -14760 20930
rect -14720 21430 -14680 21440
rect -14720 21410 -14710 21430
rect -14690 21410 -14680 21430
rect -14720 21270 -14680 21410
rect -14720 21250 -14710 21270
rect -14690 21250 -14680 21270
rect -14720 21110 -14680 21250
rect -14720 21090 -14710 21110
rect -14690 21090 -14680 21110
rect -14720 20950 -14680 21090
rect -14720 20930 -14710 20950
rect -14690 20930 -14680 20950
rect -14720 20920 -14680 20930
rect -14640 21430 -14600 21440
rect -14640 21410 -14630 21430
rect -14610 21410 -14600 21430
rect -14640 21270 -14600 21410
rect -14640 21250 -14630 21270
rect -14610 21250 -14600 21270
rect -14640 21110 -14600 21250
rect -14640 21090 -14630 21110
rect -14610 21090 -14600 21110
rect -14640 20950 -14600 21090
rect -14640 20930 -14630 20950
rect -14610 20930 -14600 20950
rect -14640 20920 -14600 20930
rect -14560 21430 -14520 21440
rect -14560 21410 -14550 21430
rect -14530 21410 -14520 21430
rect -14560 21270 -14520 21410
rect -14560 21250 -14550 21270
rect -14530 21250 -14520 21270
rect -14560 21110 -14520 21250
rect -14560 21090 -14550 21110
rect -14530 21090 -14520 21110
rect -14560 20950 -14520 21090
rect -14560 20930 -14550 20950
rect -14530 20930 -14520 20950
rect -14560 20920 -14520 20930
rect -14480 21430 -14440 21440
rect -14480 21410 -14470 21430
rect -14450 21410 -14440 21430
rect -14480 21270 -14440 21410
rect -14480 21250 -14470 21270
rect -14450 21250 -14440 21270
rect -14480 21110 -14440 21250
rect -14480 21090 -14470 21110
rect -14450 21090 -14440 21110
rect -14480 20950 -14440 21090
rect -14480 20930 -14470 20950
rect -14450 20930 -14440 20950
rect -14480 20920 -14440 20930
rect -14400 21430 -14360 21440
rect -14400 21410 -14390 21430
rect -14370 21410 -14360 21430
rect -14400 21270 -14360 21410
rect -14400 21250 -14390 21270
rect -14370 21250 -14360 21270
rect -14400 21110 -14360 21250
rect -14400 21090 -14390 21110
rect -14370 21090 -14360 21110
rect -14400 20950 -14360 21090
rect -14400 20930 -14390 20950
rect -14370 20930 -14360 20950
rect -14400 20920 -14360 20930
rect -14320 21430 -14280 21440
rect -14320 21410 -14310 21430
rect -14290 21410 -14280 21430
rect -14320 21270 -14280 21410
rect -14320 21250 -14310 21270
rect -14290 21250 -14280 21270
rect -14320 21110 -14280 21250
rect -14320 21090 -14310 21110
rect -14290 21090 -14280 21110
rect -14320 20950 -14280 21090
rect -14320 20930 -14310 20950
rect -14290 20930 -14280 20950
rect -14320 20920 -14280 20930
rect -14240 21430 -14200 21440
rect -14240 21410 -14230 21430
rect -14210 21410 -14200 21430
rect -14240 21270 -14200 21410
rect -14240 21250 -14230 21270
rect -14210 21250 -14200 21270
rect -14240 21110 -14200 21250
rect -14240 21090 -14230 21110
rect -14210 21090 -14200 21110
rect -14240 20950 -14200 21090
rect -14240 20930 -14230 20950
rect -14210 20930 -14200 20950
rect -14240 20920 -14200 20930
rect -14160 21430 -14120 21440
rect -14160 21410 -14150 21430
rect -14130 21410 -14120 21430
rect -14160 21270 -14120 21410
rect -14160 21250 -14150 21270
rect -14130 21250 -14120 21270
rect -14160 21110 -14120 21250
rect -14160 21090 -14150 21110
rect -14130 21090 -14120 21110
rect -14160 20950 -14120 21090
rect -14160 20930 -14150 20950
rect -14130 20930 -14120 20950
rect -14160 20920 -14120 20930
rect -14080 21430 -14040 21440
rect -14080 21410 -14070 21430
rect -14050 21410 -14040 21430
rect -14080 21270 -14040 21410
rect -14080 21250 -14070 21270
rect -14050 21250 -14040 21270
rect -14080 21110 -14040 21250
rect -14080 21090 -14070 21110
rect -14050 21090 -14040 21110
rect -14080 20950 -14040 21090
rect -14080 20930 -14070 20950
rect -14050 20930 -14040 20950
rect -14080 20920 -14040 20930
rect -14000 21430 -13960 21440
rect -14000 21410 -13990 21430
rect -13970 21410 -13960 21430
rect -14000 21270 -13960 21410
rect -14000 21250 -13990 21270
rect -13970 21250 -13960 21270
rect -14000 21110 -13960 21250
rect -14000 21090 -13990 21110
rect -13970 21090 -13960 21110
rect -14000 20950 -13960 21090
rect -14000 20930 -13990 20950
rect -13970 20930 -13960 20950
rect -14000 20920 -13960 20930
rect -13920 21430 -13880 21440
rect -13920 21410 -13910 21430
rect -13890 21410 -13880 21430
rect -13920 21270 -13880 21410
rect -13920 21250 -13910 21270
rect -13890 21250 -13880 21270
rect -13920 21110 -13880 21250
rect -13920 21090 -13910 21110
rect -13890 21090 -13880 21110
rect -13920 20950 -13880 21090
rect -13920 20930 -13910 20950
rect -13890 20930 -13880 20950
rect -13920 20920 -13880 20930
rect -13840 21430 -13800 21440
rect -13840 21410 -13830 21430
rect -13810 21410 -13800 21430
rect -13840 21270 -13800 21410
rect -13840 21250 -13830 21270
rect -13810 21250 -13800 21270
rect -13840 21110 -13800 21250
rect -13840 21090 -13830 21110
rect -13810 21090 -13800 21110
rect -13840 20950 -13800 21090
rect -13840 20930 -13830 20950
rect -13810 20930 -13800 20950
rect -13840 20920 -13800 20930
rect -13760 21430 -13720 21440
rect -13760 21410 -13750 21430
rect -13730 21410 -13720 21430
rect -13760 21270 -13720 21410
rect -13760 21250 -13750 21270
rect -13730 21250 -13720 21270
rect -13760 21110 -13720 21250
rect -13760 21090 -13750 21110
rect -13730 21090 -13720 21110
rect -13760 20950 -13720 21090
rect -13760 20930 -13750 20950
rect -13730 20930 -13720 20950
rect -13760 20920 -13720 20930
rect -13680 21430 -13640 21440
rect -13680 21410 -13670 21430
rect -13650 21410 -13640 21430
rect -13680 21270 -13640 21410
rect -13680 21250 -13670 21270
rect -13650 21250 -13640 21270
rect -13680 21110 -13640 21250
rect -13680 21090 -13670 21110
rect -13650 21090 -13640 21110
rect -13680 20950 -13640 21090
rect -13680 20930 -13670 20950
rect -13650 20930 -13640 20950
rect -13680 20920 -13640 20930
rect -13600 21430 -13560 21440
rect -13600 21410 -13590 21430
rect -13570 21410 -13560 21430
rect -13600 21270 -13560 21410
rect -13600 21250 -13590 21270
rect -13570 21250 -13560 21270
rect -13600 21110 -13560 21250
rect -13600 21090 -13590 21110
rect -13570 21090 -13560 21110
rect -13600 20950 -13560 21090
rect -13600 20930 -13590 20950
rect -13570 20930 -13560 20950
rect -13600 20920 -13560 20930
rect -13520 21430 -13480 21440
rect -13520 21410 -13510 21430
rect -13490 21410 -13480 21430
rect -13520 21270 -13480 21410
rect -13520 21250 -13510 21270
rect -13490 21250 -13480 21270
rect -13520 21110 -13480 21250
rect -13520 21090 -13510 21110
rect -13490 21090 -13480 21110
rect -13520 20950 -13480 21090
rect -13520 20930 -13510 20950
rect -13490 20930 -13480 20950
rect -13520 20920 -13480 20930
rect -13440 21430 -13400 21440
rect -13440 21410 -13430 21430
rect -13410 21410 -13400 21430
rect -13440 21270 -13400 21410
rect -13440 21250 -13430 21270
rect -13410 21250 -13400 21270
rect -13440 21110 -13400 21250
rect -13440 21090 -13430 21110
rect -13410 21090 -13400 21110
rect -13440 20950 -13400 21090
rect -13440 20930 -13430 20950
rect -13410 20930 -13400 20950
rect -13440 20920 -13400 20930
rect -13360 21430 -13320 21440
rect -13360 21410 -13350 21430
rect -13330 21410 -13320 21430
rect -13360 21270 -13320 21410
rect -13360 21250 -13350 21270
rect -13330 21250 -13320 21270
rect -13360 21110 -13320 21250
rect -13360 21090 -13350 21110
rect -13330 21090 -13320 21110
rect -13360 20950 -13320 21090
rect -13360 20930 -13350 20950
rect -13330 20930 -13320 20950
rect -13360 20920 -13320 20930
rect -13280 21430 -13240 21440
rect -13280 21410 -13270 21430
rect -13250 21410 -13240 21430
rect -13280 21270 -13240 21410
rect -13280 21250 -13270 21270
rect -13250 21250 -13240 21270
rect -13280 21110 -13240 21250
rect -13280 21090 -13270 21110
rect -13250 21090 -13240 21110
rect -13280 20950 -13240 21090
rect -13280 20930 -13270 20950
rect -13250 20930 -13240 20950
rect -13280 20920 -13240 20930
rect -13200 21430 -13160 21440
rect -13200 21410 -13190 21430
rect -13170 21410 -13160 21430
rect -13200 21270 -13160 21410
rect -13200 21250 -13190 21270
rect -13170 21250 -13160 21270
rect -13200 21110 -13160 21250
rect -13200 21090 -13190 21110
rect -13170 21090 -13160 21110
rect -13200 20950 -13160 21090
rect -13200 20930 -13190 20950
rect -13170 20930 -13160 20950
rect -13200 20920 -13160 20930
rect -13120 21430 -13080 21440
rect -13120 21410 -13110 21430
rect -13090 21410 -13080 21430
rect -13120 21270 -13080 21410
rect -13120 21250 -13110 21270
rect -13090 21250 -13080 21270
rect -13120 21110 -13080 21250
rect -13120 21090 -13110 21110
rect -13090 21090 -13080 21110
rect -13120 20950 -13080 21090
rect -13120 20930 -13110 20950
rect -13090 20930 -13080 20950
rect -13120 20920 -13080 20930
rect -13040 21430 -13000 21440
rect -13040 21410 -13030 21430
rect -13010 21410 -13000 21430
rect -13040 21270 -13000 21410
rect -13040 21250 -13030 21270
rect -13010 21250 -13000 21270
rect -13040 21110 -13000 21250
rect -13040 21090 -13030 21110
rect -13010 21090 -13000 21110
rect -13040 20950 -13000 21090
rect -13040 20930 -13030 20950
rect -13010 20930 -13000 20950
rect -13040 20920 -13000 20930
rect -12960 21430 -12920 21440
rect -12960 21410 -12950 21430
rect -12930 21410 -12920 21430
rect -12960 21270 -12920 21410
rect -12960 21250 -12950 21270
rect -12930 21250 -12920 21270
rect -12960 21110 -12920 21250
rect -12960 21090 -12950 21110
rect -12930 21090 -12920 21110
rect -12960 20950 -12920 21090
rect -12960 20930 -12950 20950
rect -12930 20930 -12920 20950
rect -12960 20920 -12920 20930
rect -12880 21430 -12840 21440
rect -12880 21410 -12870 21430
rect -12850 21410 -12840 21430
rect -12880 21270 -12840 21410
rect -12880 21250 -12870 21270
rect -12850 21250 -12840 21270
rect -12880 21110 -12840 21250
rect -12880 21090 -12870 21110
rect -12850 21090 -12840 21110
rect -12880 20950 -12840 21090
rect -12880 20930 -12870 20950
rect -12850 20930 -12840 20950
rect -12880 20920 -12840 20930
rect -12800 21430 -12760 21440
rect -12800 21410 -12790 21430
rect -12770 21410 -12760 21430
rect -12800 21270 -12760 21410
rect -12800 21250 -12790 21270
rect -12770 21250 -12760 21270
rect -12800 21110 -12760 21250
rect -12800 21090 -12790 21110
rect -12770 21090 -12760 21110
rect -12800 20950 -12760 21090
rect -12800 20930 -12790 20950
rect -12770 20930 -12760 20950
rect -12800 20920 -12760 20930
rect -12720 21430 -12680 21440
rect -12720 21410 -12710 21430
rect -12690 21410 -12680 21430
rect -12720 21270 -12680 21410
rect -12720 21250 -12710 21270
rect -12690 21250 -12680 21270
rect -12720 21110 -12680 21250
rect -12720 21090 -12710 21110
rect -12690 21090 -12680 21110
rect -12720 20950 -12680 21090
rect -12720 20930 -12710 20950
rect -12690 20930 -12680 20950
rect -12720 20920 -12680 20930
rect -12640 21430 -12600 21440
rect -12640 21410 -12630 21430
rect -12610 21410 -12600 21430
rect -12640 21270 -12600 21410
rect -12640 21250 -12630 21270
rect -12610 21250 -12600 21270
rect -12640 21110 -12600 21250
rect -12640 21090 -12630 21110
rect -12610 21090 -12600 21110
rect -12640 20950 -12600 21090
rect -12640 20930 -12630 20950
rect -12610 20930 -12600 20950
rect -12640 20920 -12600 20930
rect -12560 21430 -12520 21440
rect -12560 21410 -12550 21430
rect -12530 21410 -12520 21430
rect -12560 21270 -12520 21410
rect -12560 21250 -12550 21270
rect -12530 21250 -12520 21270
rect -12560 21110 -12520 21250
rect -12560 21090 -12550 21110
rect -12530 21090 -12520 21110
rect -12560 20950 -12520 21090
rect -12560 20930 -12550 20950
rect -12530 20930 -12520 20950
rect -12560 20920 -12520 20930
rect -12480 21430 -12440 21440
rect -12480 21410 -12470 21430
rect -12450 21410 -12440 21430
rect -12480 21270 -12440 21410
rect -12480 21250 -12470 21270
rect -12450 21250 -12440 21270
rect -12480 21110 -12440 21250
rect -12480 21090 -12470 21110
rect -12450 21090 -12440 21110
rect -12480 20950 -12440 21090
rect -12480 20930 -12470 20950
rect -12450 20930 -12440 20950
rect -12480 20920 -12440 20930
rect -12400 21430 -12360 21440
rect -12400 21410 -12390 21430
rect -12370 21410 -12360 21430
rect -12400 21270 -12360 21410
rect -12400 21250 -12390 21270
rect -12370 21250 -12360 21270
rect -12400 21110 -12360 21250
rect -12400 21090 -12390 21110
rect -12370 21090 -12360 21110
rect -12400 20950 -12360 21090
rect -12400 20930 -12390 20950
rect -12370 20930 -12360 20950
rect -12400 20920 -12360 20930
rect -12320 21430 -12280 21440
rect -12320 21410 -12310 21430
rect -12290 21410 -12280 21430
rect -12320 21270 -12280 21410
rect -12320 21250 -12310 21270
rect -12290 21250 -12280 21270
rect -12320 21110 -12280 21250
rect -12320 21090 -12310 21110
rect -12290 21090 -12280 21110
rect -12320 20950 -12280 21090
rect -12320 20930 -12310 20950
rect -12290 20930 -12280 20950
rect -12320 20920 -12280 20930
rect -12240 21430 -12200 21440
rect -12240 21410 -12230 21430
rect -12210 21410 -12200 21430
rect -12240 21270 -12200 21410
rect -12240 21250 -12230 21270
rect -12210 21250 -12200 21270
rect -12240 21110 -12200 21250
rect -12240 21090 -12230 21110
rect -12210 21090 -12200 21110
rect -12240 20950 -12200 21090
rect -12240 20930 -12230 20950
rect -12210 20930 -12200 20950
rect -12240 20920 -12200 20930
rect -12160 21430 -12120 21440
rect -12160 21410 -12150 21430
rect -12130 21410 -12120 21430
rect -12160 21270 -12120 21410
rect -12160 21250 -12150 21270
rect -12130 21250 -12120 21270
rect -12160 21110 -12120 21250
rect -12160 21090 -12150 21110
rect -12130 21090 -12120 21110
rect -12160 20950 -12120 21090
rect -12160 20930 -12150 20950
rect -12130 20930 -12120 20950
rect -12160 20920 -12120 20930
rect -12080 21430 -12040 21440
rect -12080 21410 -12070 21430
rect -12050 21410 -12040 21430
rect -12080 21270 -12040 21410
rect -12080 21250 -12070 21270
rect -12050 21250 -12040 21270
rect -12080 21110 -12040 21250
rect -12080 21090 -12070 21110
rect -12050 21090 -12040 21110
rect -12080 20950 -12040 21090
rect -12080 20930 -12070 20950
rect -12050 20930 -12040 20950
rect -12080 20920 -12040 20930
rect -12000 21430 -11960 21440
rect -12000 21410 -11990 21430
rect -11970 21410 -11960 21430
rect -12000 21270 -11960 21410
rect -12000 21250 -11990 21270
rect -11970 21250 -11960 21270
rect -12000 21110 -11960 21250
rect -12000 21090 -11990 21110
rect -11970 21090 -11960 21110
rect -12000 20950 -11960 21090
rect -12000 20930 -11990 20950
rect -11970 20930 -11960 20950
rect -12000 20920 -11960 20930
rect -11920 21430 -11880 21440
rect -11920 21410 -11910 21430
rect -11890 21410 -11880 21430
rect -11920 21270 -11880 21410
rect -11920 21250 -11910 21270
rect -11890 21250 -11880 21270
rect -11920 21110 -11880 21250
rect -11920 21090 -11910 21110
rect -11890 21090 -11880 21110
rect -11920 20950 -11880 21090
rect -11920 20930 -11910 20950
rect -11890 20930 -11880 20950
rect -11920 20920 -11880 20930
rect -11840 21430 -11800 21440
rect -11840 21410 -11830 21430
rect -11810 21410 -11800 21430
rect -11840 21270 -11800 21410
rect -11840 21250 -11830 21270
rect -11810 21250 -11800 21270
rect -11840 21110 -11800 21250
rect -11840 21090 -11830 21110
rect -11810 21090 -11800 21110
rect -11840 20950 -11800 21090
rect -11840 20930 -11830 20950
rect -11810 20930 -11800 20950
rect -11840 20920 -11800 20930
rect -11760 21430 -11720 21440
rect -11760 21410 -11750 21430
rect -11730 21410 -11720 21430
rect -11760 21270 -11720 21410
rect -11760 21250 -11750 21270
rect -11730 21250 -11720 21270
rect -11760 21110 -11720 21250
rect -11760 21090 -11750 21110
rect -11730 21090 -11720 21110
rect -11760 20950 -11720 21090
rect -11760 20930 -11750 20950
rect -11730 20930 -11720 20950
rect -11760 20920 -11720 20930
rect -11680 21430 -11640 21440
rect -11680 21410 -11670 21430
rect -11650 21410 -11640 21430
rect -11680 21270 -11640 21410
rect -11680 21250 -11670 21270
rect -11650 21250 -11640 21270
rect -11680 21110 -11640 21250
rect -11680 21090 -11670 21110
rect -11650 21090 -11640 21110
rect -11680 20950 -11640 21090
rect -11680 20930 -11670 20950
rect -11650 20930 -11640 20950
rect -11680 20920 -11640 20930
rect -11600 21430 -11560 21440
rect -11600 21410 -11590 21430
rect -11570 21410 -11560 21430
rect -11600 21270 -11560 21410
rect -11600 21250 -11590 21270
rect -11570 21250 -11560 21270
rect -11600 21110 -11560 21250
rect -11600 21090 -11590 21110
rect -11570 21090 -11560 21110
rect -11600 20950 -11560 21090
rect -11600 20930 -11590 20950
rect -11570 20930 -11560 20950
rect -11600 20920 -11560 20930
rect -11520 21430 -11480 21440
rect -11520 21410 -11510 21430
rect -11490 21410 -11480 21430
rect -11520 21270 -11480 21410
rect -11520 21250 -11510 21270
rect -11490 21250 -11480 21270
rect -11520 21110 -11480 21250
rect -11520 21090 -11510 21110
rect -11490 21090 -11480 21110
rect -11520 20950 -11480 21090
rect -11520 20930 -11510 20950
rect -11490 20930 -11480 20950
rect -11520 20920 -11480 20930
rect -11440 21430 -11400 21440
rect -11440 21410 -11430 21430
rect -11410 21410 -11400 21430
rect -11440 21270 -11400 21410
rect -11440 21250 -11430 21270
rect -11410 21250 -11400 21270
rect -11440 21110 -11400 21250
rect -11440 21090 -11430 21110
rect -11410 21090 -11400 21110
rect -11440 20950 -11400 21090
rect -11440 20930 -11430 20950
rect -11410 20930 -11400 20950
rect -11440 20920 -11400 20930
rect -11360 21430 -11320 21440
rect -11360 21410 -11350 21430
rect -11330 21410 -11320 21430
rect -11360 21270 -11320 21410
rect -11360 21250 -11350 21270
rect -11330 21250 -11320 21270
rect -11360 21110 -11320 21250
rect -11360 21090 -11350 21110
rect -11330 21090 -11320 21110
rect -11360 20950 -11320 21090
rect -11360 20930 -11350 20950
rect -11330 20930 -11320 20950
rect -11360 20920 -11320 20930
rect -11280 21430 -11240 21440
rect -11280 21410 -11270 21430
rect -11250 21410 -11240 21430
rect -11280 21270 -11240 21410
rect -11280 21250 -11270 21270
rect -11250 21250 -11240 21270
rect -11280 21110 -11240 21250
rect -11280 21090 -11270 21110
rect -11250 21090 -11240 21110
rect -11280 20950 -11240 21090
rect -11280 20930 -11270 20950
rect -11250 20930 -11240 20950
rect -11280 20920 -11240 20930
rect -11200 21430 -11160 21440
rect -11200 21410 -11190 21430
rect -11170 21410 -11160 21430
rect -11200 21270 -11160 21410
rect -11200 21250 -11190 21270
rect -11170 21250 -11160 21270
rect -11200 21110 -11160 21250
rect -11200 21090 -11190 21110
rect -11170 21090 -11160 21110
rect -11200 20950 -11160 21090
rect -11200 20930 -11190 20950
rect -11170 20930 -11160 20950
rect -11200 20920 -11160 20930
rect -11120 21430 -11080 21440
rect -11120 21410 -11110 21430
rect -11090 21410 -11080 21430
rect -11120 21270 -11080 21410
rect -11120 21250 -11110 21270
rect -11090 21250 -11080 21270
rect -11120 21110 -11080 21250
rect -11120 21090 -11110 21110
rect -11090 21090 -11080 21110
rect -11120 20950 -11080 21090
rect -11120 20930 -11110 20950
rect -11090 20930 -11080 20950
rect -11120 20920 -11080 20930
rect -11040 21430 -11000 21440
rect -11040 21410 -11030 21430
rect -11010 21410 -11000 21430
rect -11040 21270 -11000 21410
rect -11040 21250 -11030 21270
rect -11010 21250 -11000 21270
rect -11040 21110 -11000 21250
rect -11040 21090 -11030 21110
rect -11010 21090 -11000 21110
rect -11040 20950 -11000 21090
rect -11040 20930 -11030 20950
rect -11010 20930 -11000 20950
rect -11040 20920 -11000 20930
rect -10960 21430 -10920 21440
rect -10960 21410 -10950 21430
rect -10930 21410 -10920 21430
rect -10960 21270 -10920 21410
rect -10960 21250 -10950 21270
rect -10930 21250 -10920 21270
rect -10960 21110 -10920 21250
rect -10960 21090 -10950 21110
rect -10930 21090 -10920 21110
rect -10960 20950 -10920 21090
rect -10960 20930 -10950 20950
rect -10930 20930 -10920 20950
rect -10960 20920 -10920 20930
rect -10880 21430 -10840 21440
rect -10880 21410 -10870 21430
rect -10850 21410 -10840 21430
rect -10880 21270 -10840 21410
rect -10880 21250 -10870 21270
rect -10850 21250 -10840 21270
rect -10880 21110 -10840 21250
rect -10880 21090 -10870 21110
rect -10850 21090 -10840 21110
rect -10880 20950 -10840 21090
rect -10880 20930 -10870 20950
rect -10850 20930 -10840 20950
rect -10880 20920 -10840 20930
rect -10800 21430 -10760 21440
rect -10800 21410 -10790 21430
rect -10770 21410 -10760 21430
rect -10800 21270 -10760 21410
rect -10800 21250 -10790 21270
rect -10770 21250 -10760 21270
rect -10800 21110 -10760 21250
rect -10800 21090 -10790 21110
rect -10770 21090 -10760 21110
rect -10800 20950 -10760 21090
rect -10800 20930 -10790 20950
rect -10770 20930 -10760 20950
rect -10800 20920 -10760 20930
rect -10720 21430 -10680 21440
rect -10720 21410 -10710 21430
rect -10690 21410 -10680 21430
rect -10720 21270 -10680 21410
rect -10720 21250 -10710 21270
rect -10690 21250 -10680 21270
rect -10720 21110 -10680 21250
rect -10720 21090 -10710 21110
rect -10690 21090 -10680 21110
rect -10720 20950 -10680 21090
rect -10720 20930 -10710 20950
rect -10690 20930 -10680 20950
rect -10720 20920 -10680 20930
rect -10640 21430 -10600 21440
rect -10640 21410 -10630 21430
rect -10610 21410 -10600 21430
rect -10640 21270 -10600 21410
rect -10640 21250 -10630 21270
rect -10610 21250 -10600 21270
rect -10640 21110 -10600 21250
rect -10640 21090 -10630 21110
rect -10610 21090 -10600 21110
rect -10640 20950 -10600 21090
rect -10640 20930 -10630 20950
rect -10610 20930 -10600 20950
rect -10640 20920 -10600 20930
rect -10560 21430 -10520 21440
rect -10560 21410 -10550 21430
rect -10530 21410 -10520 21430
rect -10560 21270 -10520 21410
rect -10560 21250 -10550 21270
rect -10530 21250 -10520 21270
rect -10560 21110 -10520 21250
rect -10560 21090 -10550 21110
rect -10530 21090 -10520 21110
rect -10560 20950 -10520 21090
rect -10560 20930 -10550 20950
rect -10530 20930 -10520 20950
rect -10560 20920 -10520 20930
rect -10480 21430 -10440 21440
rect -10480 21410 -10470 21430
rect -10450 21410 -10440 21430
rect -10480 21270 -10440 21410
rect -10480 21250 -10470 21270
rect -10450 21250 -10440 21270
rect -10480 21110 -10440 21250
rect -10480 21090 -10470 21110
rect -10450 21090 -10440 21110
rect -10480 20950 -10440 21090
rect -10480 20930 -10470 20950
rect -10450 20930 -10440 20950
rect -10480 20920 -10440 20930
rect -10400 21430 -10360 21440
rect -10400 21410 -10390 21430
rect -10370 21410 -10360 21430
rect -10400 21270 -10360 21410
rect -10400 21250 -10390 21270
rect -10370 21250 -10360 21270
rect -10400 21110 -10360 21250
rect -10400 21090 -10390 21110
rect -10370 21090 -10360 21110
rect -10400 20950 -10360 21090
rect -10400 20930 -10390 20950
rect -10370 20930 -10360 20950
rect -10400 20920 -10360 20930
rect -10320 21430 -10280 21440
rect -10320 21410 -10310 21430
rect -10290 21410 -10280 21430
rect -10320 21270 -10280 21410
rect -10320 21250 -10310 21270
rect -10290 21250 -10280 21270
rect -10320 21110 -10280 21250
rect -10320 21090 -10310 21110
rect -10290 21090 -10280 21110
rect -10320 20950 -10280 21090
rect -10320 20930 -10310 20950
rect -10290 20930 -10280 20950
rect -10320 20920 -10280 20930
rect -10240 21430 -10200 21440
rect -10240 21410 -10230 21430
rect -10210 21410 -10200 21430
rect -10240 21270 -10200 21410
rect -10240 21250 -10230 21270
rect -10210 21250 -10200 21270
rect -10240 21110 -10200 21250
rect -10240 21090 -10230 21110
rect -10210 21090 -10200 21110
rect -10240 20950 -10200 21090
rect -10240 20930 -10230 20950
rect -10210 20930 -10200 20950
rect -10240 20920 -10200 20930
rect -10160 21430 -10120 21440
rect -10160 21410 -10150 21430
rect -10130 21410 -10120 21430
rect -10160 21270 -10120 21410
rect -10160 21250 -10150 21270
rect -10130 21250 -10120 21270
rect -10160 21110 -10120 21250
rect -10160 21090 -10150 21110
rect -10130 21090 -10120 21110
rect -10160 20950 -10120 21090
rect -10160 20930 -10150 20950
rect -10130 20930 -10120 20950
rect -10160 20920 -10120 20930
rect -10080 21430 -10040 21440
rect -10080 21410 -10070 21430
rect -10050 21410 -10040 21430
rect -10080 21270 -10040 21410
rect -10080 21250 -10070 21270
rect -10050 21250 -10040 21270
rect -10080 21110 -10040 21250
rect -10080 21090 -10070 21110
rect -10050 21090 -10040 21110
rect -10080 20950 -10040 21090
rect -10080 20930 -10070 20950
rect -10050 20930 -10040 20950
rect -10080 20920 -10040 20930
rect -10000 21430 -9960 21440
rect -10000 21410 -9990 21430
rect -9970 21410 -9960 21430
rect -10000 21270 -9960 21410
rect -10000 21250 -9990 21270
rect -9970 21250 -9960 21270
rect -10000 21110 -9960 21250
rect -10000 21090 -9990 21110
rect -9970 21090 -9960 21110
rect -10000 20950 -9960 21090
rect -10000 20930 -9990 20950
rect -9970 20930 -9960 20950
rect -10000 20920 -9960 20930
rect -9920 21430 -9880 21440
rect -9920 21410 -9910 21430
rect -9890 21410 -9880 21430
rect -9920 21270 -9880 21410
rect -9920 21250 -9910 21270
rect -9890 21250 -9880 21270
rect -9920 21110 -9880 21250
rect -9920 21090 -9910 21110
rect -9890 21090 -9880 21110
rect -9920 20950 -9880 21090
rect -9920 20930 -9910 20950
rect -9890 20930 -9880 20950
rect -9920 20920 -9880 20930
rect -9840 21430 -9800 21440
rect -9840 21410 -9830 21430
rect -9810 21410 -9800 21430
rect -9840 21270 -9800 21410
rect -9840 21250 -9830 21270
rect -9810 21250 -9800 21270
rect -9840 21110 -9800 21250
rect -9840 21090 -9830 21110
rect -9810 21090 -9800 21110
rect -9840 20950 -9800 21090
rect -9840 20930 -9830 20950
rect -9810 20930 -9800 20950
rect -9840 20920 -9800 20930
rect -9760 21430 -9720 21440
rect -9760 21410 -9750 21430
rect -9730 21410 -9720 21430
rect -9760 21270 -9720 21410
rect -9760 21250 -9750 21270
rect -9730 21250 -9720 21270
rect -9760 21110 -9720 21250
rect -9760 21090 -9750 21110
rect -9730 21090 -9720 21110
rect -9760 20950 -9720 21090
rect -9760 20930 -9750 20950
rect -9730 20930 -9720 20950
rect -9760 20920 -9720 20930
rect -9680 21430 -9640 21440
rect -9680 21410 -9670 21430
rect -9650 21410 -9640 21430
rect -9680 21270 -9640 21410
rect -9680 21250 -9670 21270
rect -9650 21250 -9640 21270
rect -9680 21110 -9640 21250
rect -9680 21090 -9670 21110
rect -9650 21090 -9640 21110
rect -9680 20950 -9640 21090
rect -9680 20930 -9670 20950
rect -9650 20930 -9640 20950
rect -9680 20920 -9640 20930
rect -9600 21430 -9560 21440
rect -9600 21410 -9590 21430
rect -9570 21410 -9560 21430
rect -9600 21270 -9560 21410
rect -9600 21250 -9590 21270
rect -9570 21250 -9560 21270
rect -9600 21110 -9560 21250
rect -9600 21090 -9590 21110
rect -9570 21090 -9560 21110
rect -9600 20950 -9560 21090
rect -9600 20930 -9590 20950
rect -9570 20930 -9560 20950
rect -9600 20920 -9560 20930
rect -9520 21430 -9480 21440
rect -9520 21410 -9510 21430
rect -9490 21410 -9480 21430
rect -9520 21270 -9480 21410
rect -9520 21250 -9510 21270
rect -9490 21250 -9480 21270
rect -9520 21110 -9480 21250
rect -9520 21090 -9510 21110
rect -9490 21090 -9480 21110
rect -9520 20950 -9480 21090
rect -9520 20930 -9510 20950
rect -9490 20930 -9480 20950
rect -9520 20920 -9480 20930
rect -9440 21430 -9400 21440
rect -9440 21410 -9430 21430
rect -9410 21410 -9400 21430
rect -9440 21270 -9400 21410
rect -9440 21250 -9430 21270
rect -9410 21250 -9400 21270
rect -9440 21110 -9400 21250
rect -9440 21090 -9430 21110
rect -9410 21090 -9400 21110
rect -9440 20950 -9400 21090
rect -9440 20930 -9430 20950
rect -9410 20930 -9400 20950
rect -9440 20920 -9400 20930
rect -9360 21430 -9320 21440
rect -9360 21410 -9350 21430
rect -9330 21410 -9320 21430
rect -9360 21270 -9320 21410
rect -9360 21250 -9350 21270
rect -9330 21250 -9320 21270
rect -9360 21110 -9320 21250
rect -9360 21090 -9350 21110
rect -9330 21090 -9320 21110
rect -9360 20950 -9320 21090
rect -9360 20930 -9350 20950
rect -9330 20930 -9320 20950
rect -9360 20920 -9320 20930
rect -9280 21430 -9240 21440
rect -9280 21410 -9270 21430
rect -9250 21410 -9240 21430
rect -9280 21270 -9240 21410
rect -9280 21250 -9270 21270
rect -9250 21250 -9240 21270
rect -9280 21110 -9240 21250
rect -9280 21090 -9270 21110
rect -9250 21090 -9240 21110
rect -9280 20950 -9240 21090
rect -9280 20930 -9270 20950
rect -9250 20930 -9240 20950
rect -9280 20920 -9240 20930
rect -9200 21430 -9160 21440
rect -9200 21410 -9190 21430
rect -9170 21410 -9160 21430
rect -9200 21270 -9160 21410
rect -9200 21250 -9190 21270
rect -9170 21250 -9160 21270
rect -9200 21110 -9160 21250
rect -9200 21090 -9190 21110
rect -9170 21090 -9160 21110
rect -9200 20950 -9160 21090
rect -9200 20930 -9190 20950
rect -9170 20930 -9160 20950
rect -9200 20920 -9160 20930
rect -9120 21430 -9080 21440
rect -9120 21410 -9110 21430
rect -9090 21410 -9080 21430
rect -9120 21270 -9080 21410
rect -9120 21250 -9110 21270
rect -9090 21250 -9080 21270
rect -9120 21110 -9080 21250
rect -9120 21090 -9110 21110
rect -9090 21090 -9080 21110
rect -9120 20950 -9080 21090
rect -9120 20930 -9110 20950
rect -9090 20930 -9080 20950
rect -9120 20920 -9080 20930
rect -9040 21430 -9000 21440
rect -9040 21410 -9030 21430
rect -9010 21410 -9000 21430
rect -9040 21270 -9000 21410
rect -9040 21250 -9030 21270
rect -9010 21250 -9000 21270
rect -9040 21110 -9000 21250
rect -9040 21090 -9030 21110
rect -9010 21090 -9000 21110
rect -9040 20950 -9000 21090
rect -9040 20930 -9030 20950
rect -9010 20930 -9000 20950
rect -9040 20920 -9000 20930
rect -8960 21430 -8920 21440
rect -8960 21410 -8950 21430
rect -8930 21410 -8920 21430
rect -8960 21270 -8920 21410
rect -8960 21250 -8950 21270
rect -8930 21250 -8920 21270
rect -8960 21110 -8920 21250
rect -8960 21090 -8950 21110
rect -8930 21090 -8920 21110
rect -8960 20950 -8920 21090
rect -8960 20930 -8950 20950
rect -8930 20930 -8920 20950
rect -8960 20920 -8920 20930
rect -8880 21430 -8840 21440
rect -8880 21410 -8870 21430
rect -8850 21410 -8840 21430
rect -8880 21270 -8840 21410
rect -8880 21250 -8870 21270
rect -8850 21250 -8840 21270
rect -8880 21110 -8840 21250
rect -8880 21090 -8870 21110
rect -8850 21090 -8840 21110
rect -8880 20950 -8840 21090
rect -8880 20930 -8870 20950
rect -8850 20930 -8840 20950
rect -8880 20920 -8840 20930
rect -8800 21430 -8760 21440
rect -8800 21410 -8790 21430
rect -8770 21410 -8760 21430
rect -8800 21270 -8760 21410
rect -8800 21250 -8790 21270
rect -8770 21250 -8760 21270
rect -8800 21110 -8760 21250
rect -8800 21090 -8790 21110
rect -8770 21090 -8760 21110
rect -8800 20950 -8760 21090
rect -8800 20930 -8790 20950
rect -8770 20930 -8760 20950
rect -8800 20920 -8760 20930
rect -8720 21430 -8680 21440
rect -8720 21410 -8710 21430
rect -8690 21410 -8680 21430
rect -8720 21270 -8680 21410
rect -8720 21250 -8710 21270
rect -8690 21250 -8680 21270
rect -8720 21110 -8680 21250
rect -8720 21090 -8710 21110
rect -8690 21090 -8680 21110
rect -8720 20950 -8680 21090
rect -8720 20930 -8710 20950
rect -8690 20930 -8680 20950
rect -8720 20920 -8680 20930
rect -8640 21430 -8600 21440
rect -8640 21410 -8630 21430
rect -8610 21410 -8600 21430
rect -8640 21270 -8600 21410
rect -8640 21250 -8630 21270
rect -8610 21250 -8600 21270
rect -8640 21110 -8600 21250
rect -8640 21090 -8630 21110
rect -8610 21090 -8600 21110
rect -8640 20950 -8600 21090
rect -8640 20930 -8630 20950
rect -8610 20930 -8600 20950
rect -8640 20920 -8600 20930
rect -8560 21430 -8520 21440
rect -8560 21410 -8550 21430
rect -8530 21410 -8520 21430
rect -8560 21270 -8520 21410
rect -8560 21250 -8550 21270
rect -8530 21250 -8520 21270
rect -8560 21110 -8520 21250
rect -8560 21090 -8550 21110
rect -8530 21090 -8520 21110
rect -8560 20950 -8520 21090
rect -8560 20930 -8550 20950
rect -8530 20930 -8520 20950
rect -8560 20920 -8520 20930
rect -8480 21430 -8440 21440
rect -8480 21410 -8470 21430
rect -8450 21410 -8440 21430
rect -8480 21270 -8440 21410
rect -8480 21250 -8470 21270
rect -8450 21250 -8440 21270
rect -8480 21110 -8440 21250
rect -8480 21090 -8470 21110
rect -8450 21090 -8440 21110
rect -8480 20950 -8440 21090
rect -8480 20930 -8470 20950
rect -8450 20930 -8440 20950
rect -8480 20920 -8440 20930
rect -8400 21430 -8360 21440
rect -8400 21410 -8390 21430
rect -8370 21410 -8360 21430
rect -8400 21270 -8360 21410
rect -8400 21250 -8390 21270
rect -8370 21250 -8360 21270
rect -8400 21110 -8360 21250
rect -8400 21090 -8390 21110
rect -8370 21090 -8360 21110
rect -8400 20950 -8360 21090
rect -8400 20930 -8390 20950
rect -8370 20930 -8360 20950
rect -8400 20920 -8360 20930
rect -8320 21430 -8280 21440
rect -8320 21410 -8310 21430
rect -8290 21410 -8280 21430
rect -8320 21270 -8280 21410
rect -8320 21250 -8310 21270
rect -8290 21250 -8280 21270
rect -8320 21110 -8280 21250
rect -8320 21090 -8310 21110
rect -8290 21090 -8280 21110
rect -8320 20950 -8280 21090
rect -8320 20930 -8310 20950
rect -8290 20930 -8280 20950
rect -8320 20920 -8280 20930
rect -8240 21430 -8200 21440
rect -8240 21410 -8230 21430
rect -8210 21410 -8200 21430
rect -8240 21270 -8200 21410
rect -8240 21250 -8230 21270
rect -8210 21250 -8200 21270
rect -8240 21110 -8200 21250
rect -8240 21090 -8230 21110
rect -8210 21090 -8200 21110
rect -8240 20950 -8200 21090
rect -8240 20930 -8230 20950
rect -8210 20930 -8200 20950
rect -8240 20920 -8200 20930
rect -8160 21430 -8120 21440
rect -8160 21410 -8150 21430
rect -8130 21410 -8120 21430
rect -8160 21270 -8120 21410
rect -8160 21250 -8150 21270
rect -8130 21250 -8120 21270
rect -8160 21110 -8120 21250
rect -8160 21090 -8150 21110
rect -8130 21090 -8120 21110
rect -8160 20950 -8120 21090
rect -8160 20930 -8150 20950
rect -8130 20930 -8120 20950
rect -8160 20920 -8120 20930
rect -8080 21430 -8040 21440
rect -8080 21410 -8070 21430
rect -8050 21410 -8040 21430
rect -8080 21270 -8040 21410
rect -8080 21250 -8070 21270
rect -8050 21250 -8040 21270
rect -8080 21110 -8040 21250
rect -8080 21090 -8070 21110
rect -8050 21090 -8040 21110
rect -8080 20950 -8040 21090
rect -8080 20930 -8070 20950
rect -8050 20930 -8040 20950
rect -8080 20920 -8040 20930
rect -8000 21430 -7960 21440
rect -8000 21410 -7990 21430
rect -7970 21410 -7960 21430
rect -8000 21270 -7960 21410
rect -8000 21250 -7990 21270
rect -7970 21250 -7960 21270
rect -8000 21110 -7960 21250
rect -8000 21090 -7990 21110
rect -7970 21090 -7960 21110
rect -8000 20950 -7960 21090
rect -8000 20930 -7990 20950
rect -7970 20930 -7960 20950
rect -8000 20920 -7960 20930
rect -7920 21430 -7880 21440
rect -7920 21410 -7910 21430
rect -7890 21410 -7880 21430
rect -7920 21270 -7880 21410
rect -7920 21250 -7910 21270
rect -7890 21250 -7880 21270
rect -7920 21110 -7880 21250
rect -7920 21090 -7910 21110
rect -7890 21090 -7880 21110
rect -7920 20950 -7880 21090
rect -7920 20930 -7910 20950
rect -7890 20930 -7880 20950
rect -7920 20920 -7880 20930
rect -7840 21430 -7800 21440
rect -7840 21410 -7830 21430
rect -7810 21410 -7800 21430
rect -7840 21270 -7800 21410
rect -7840 21250 -7830 21270
rect -7810 21250 -7800 21270
rect -7840 21110 -7800 21250
rect -7840 21090 -7830 21110
rect -7810 21090 -7800 21110
rect -7840 20950 -7800 21090
rect -7840 20930 -7830 20950
rect -7810 20930 -7800 20950
rect -7840 20920 -7800 20930
rect -7760 21430 -7720 21440
rect -7760 21410 -7750 21430
rect -7730 21410 -7720 21430
rect -7760 21270 -7720 21410
rect -7760 21250 -7750 21270
rect -7730 21250 -7720 21270
rect -7760 21110 -7720 21250
rect -7760 21090 -7750 21110
rect -7730 21090 -7720 21110
rect -7760 20950 -7720 21090
rect -7760 20930 -7750 20950
rect -7730 20930 -7720 20950
rect -7760 20920 -7720 20930
rect -7680 21430 -7640 21440
rect -7680 21410 -7670 21430
rect -7650 21410 -7640 21430
rect -7680 21270 -7640 21410
rect -7680 21250 -7670 21270
rect -7650 21250 -7640 21270
rect -7680 21110 -7640 21250
rect -7680 21090 -7670 21110
rect -7650 21090 -7640 21110
rect -7680 20950 -7640 21090
rect -7680 20930 -7670 20950
rect -7650 20930 -7640 20950
rect -7680 20920 -7640 20930
rect -7600 21430 -7560 21440
rect -7600 21410 -7590 21430
rect -7570 21410 -7560 21430
rect -7600 21270 -7560 21410
rect -7600 21250 -7590 21270
rect -7570 21250 -7560 21270
rect -7600 21110 -7560 21250
rect -7600 21090 -7590 21110
rect -7570 21090 -7560 21110
rect -7600 20950 -7560 21090
rect -7600 20930 -7590 20950
rect -7570 20930 -7560 20950
rect -7600 20920 -7560 20930
rect -7520 21430 -7480 21440
rect -7520 21410 -7510 21430
rect -7490 21410 -7480 21430
rect -7520 21270 -7480 21410
rect -7520 21250 -7510 21270
rect -7490 21250 -7480 21270
rect -7520 21110 -7480 21250
rect -7520 21090 -7510 21110
rect -7490 21090 -7480 21110
rect -7520 20950 -7480 21090
rect -7520 20930 -7510 20950
rect -7490 20930 -7480 20950
rect -7520 20920 -7480 20930
rect -7440 21430 -7400 21440
rect -7440 21410 -7430 21430
rect -7410 21410 -7400 21430
rect -7440 21270 -7400 21410
rect -7440 21250 -7430 21270
rect -7410 21250 -7400 21270
rect -7440 21110 -7400 21250
rect -7440 21090 -7430 21110
rect -7410 21090 -7400 21110
rect -7440 20950 -7400 21090
rect -7440 20930 -7430 20950
rect -7410 20930 -7400 20950
rect -7440 20920 -7400 20930
rect -7360 21430 -7320 21440
rect -7360 21410 -7350 21430
rect -7330 21410 -7320 21430
rect -7360 21270 -7320 21410
rect -7360 21250 -7350 21270
rect -7330 21250 -7320 21270
rect -7360 21110 -7320 21250
rect -7360 21090 -7350 21110
rect -7330 21090 -7320 21110
rect -7360 20950 -7320 21090
rect -7360 20930 -7350 20950
rect -7330 20930 -7320 20950
rect -7360 20920 -7320 20930
rect -7280 21430 -7240 21440
rect -7280 21410 -7270 21430
rect -7250 21410 -7240 21430
rect -7280 21270 -7240 21410
rect -7280 21250 -7270 21270
rect -7250 21250 -7240 21270
rect -7280 21110 -7240 21250
rect -7280 21090 -7270 21110
rect -7250 21090 -7240 21110
rect -7280 20950 -7240 21090
rect -7280 20930 -7270 20950
rect -7250 20930 -7240 20950
rect -7280 20920 -7240 20930
rect -7200 21430 -7160 21440
rect -7200 21410 -7190 21430
rect -7170 21410 -7160 21430
rect -7200 21270 -7160 21410
rect -7200 21250 -7190 21270
rect -7170 21250 -7160 21270
rect -7200 21110 -7160 21250
rect -7200 21090 -7190 21110
rect -7170 21090 -7160 21110
rect -7200 20950 -7160 21090
rect -7200 20930 -7190 20950
rect -7170 20930 -7160 20950
rect -7200 20920 -7160 20930
rect -7120 21430 -7080 21440
rect -7120 21410 -7110 21430
rect -7090 21410 -7080 21430
rect -7120 21270 -7080 21410
rect -7120 21250 -7110 21270
rect -7090 21250 -7080 21270
rect -7120 21110 -7080 21250
rect -7120 21090 -7110 21110
rect -7090 21090 -7080 21110
rect -7120 20950 -7080 21090
rect -7120 20930 -7110 20950
rect -7090 20930 -7080 20950
rect -7120 20920 -7080 20930
rect -7040 21430 -7000 21440
rect -7040 21410 -7030 21430
rect -7010 21410 -7000 21430
rect -7040 21270 -7000 21410
rect -7040 21250 -7030 21270
rect -7010 21250 -7000 21270
rect -7040 21110 -7000 21250
rect -7040 21090 -7030 21110
rect -7010 21090 -7000 21110
rect -7040 20950 -7000 21090
rect -7040 20930 -7030 20950
rect -7010 20930 -7000 20950
rect -7040 20920 -7000 20930
rect -6960 21430 -6920 21440
rect -6960 21410 -6950 21430
rect -6930 21410 -6920 21430
rect -6960 21270 -6920 21410
rect -6960 21250 -6950 21270
rect -6930 21250 -6920 21270
rect -6960 21110 -6920 21250
rect -6960 21090 -6950 21110
rect -6930 21090 -6920 21110
rect -6960 20950 -6920 21090
rect -6960 20930 -6950 20950
rect -6930 20930 -6920 20950
rect -6960 20920 -6920 20930
rect -6880 21430 -6840 21440
rect -6880 21410 -6870 21430
rect -6850 21410 -6840 21430
rect -6880 21270 -6840 21410
rect -6880 21250 -6870 21270
rect -6850 21250 -6840 21270
rect -6880 21110 -6840 21250
rect -6880 21090 -6870 21110
rect -6850 21090 -6840 21110
rect -6880 20950 -6840 21090
rect -6880 20930 -6870 20950
rect -6850 20930 -6840 20950
rect -6880 20920 -6840 20930
rect -6800 21430 -6760 21440
rect -6800 21410 -6790 21430
rect -6770 21410 -6760 21430
rect -6800 21270 -6760 21410
rect -6800 21250 -6790 21270
rect -6770 21250 -6760 21270
rect -6800 21110 -6760 21250
rect -6800 21090 -6790 21110
rect -6770 21090 -6760 21110
rect -6800 20950 -6760 21090
rect -6800 20930 -6790 20950
rect -6770 20930 -6760 20950
rect -6800 20920 -6760 20930
rect -6720 21430 -6680 21440
rect -6720 21410 -6710 21430
rect -6690 21410 -6680 21430
rect -6720 21270 -6680 21410
rect -6720 21250 -6710 21270
rect -6690 21250 -6680 21270
rect -6720 21110 -6680 21250
rect -6720 21090 -6710 21110
rect -6690 21090 -6680 21110
rect -6720 20950 -6680 21090
rect -6720 20930 -6710 20950
rect -6690 20930 -6680 20950
rect -6720 20920 -6680 20930
rect -6640 21430 -6600 21440
rect -6640 21410 -6630 21430
rect -6610 21410 -6600 21430
rect -6640 21270 -6600 21410
rect -6640 21250 -6630 21270
rect -6610 21250 -6600 21270
rect -6640 21110 -6600 21250
rect -6640 21090 -6630 21110
rect -6610 21090 -6600 21110
rect -6640 20950 -6600 21090
rect -6640 20930 -6630 20950
rect -6610 20930 -6600 20950
rect -6640 20920 -6600 20930
rect -6560 21430 -6520 21440
rect -6560 21410 -6550 21430
rect -6530 21410 -6520 21430
rect -6560 21270 -6520 21410
rect -6560 21250 -6550 21270
rect -6530 21250 -6520 21270
rect -6560 21110 -6520 21250
rect -6560 21090 -6550 21110
rect -6530 21090 -6520 21110
rect -6560 20950 -6520 21090
rect -6560 20930 -6550 20950
rect -6530 20930 -6520 20950
rect -6560 20920 -6520 20930
rect -6480 21430 -6440 21440
rect -6480 21410 -6470 21430
rect -6450 21410 -6440 21430
rect -6480 21270 -6440 21410
rect -6480 21250 -6470 21270
rect -6450 21250 -6440 21270
rect -6480 21110 -6440 21250
rect -6480 21090 -6470 21110
rect -6450 21090 -6440 21110
rect -6480 20950 -6440 21090
rect -6480 20930 -6470 20950
rect -6450 20930 -6440 20950
rect -6480 20920 -6440 20930
rect -6400 21430 -6360 21440
rect -6400 21410 -6390 21430
rect -6370 21410 -6360 21430
rect -6400 21270 -6360 21410
rect -6400 21250 -6390 21270
rect -6370 21250 -6360 21270
rect -6400 21110 -6360 21250
rect -6400 21090 -6390 21110
rect -6370 21090 -6360 21110
rect -6400 20950 -6360 21090
rect -6400 20930 -6390 20950
rect -6370 20930 -6360 20950
rect -6400 20920 -6360 20930
rect -6320 21430 -6280 21440
rect -6320 21410 -6310 21430
rect -6290 21410 -6280 21430
rect -6320 21270 -6280 21410
rect -6320 21250 -6310 21270
rect -6290 21250 -6280 21270
rect -6320 21110 -6280 21250
rect -6320 21090 -6310 21110
rect -6290 21090 -6280 21110
rect -6320 20950 -6280 21090
rect -6320 20930 -6310 20950
rect -6290 20930 -6280 20950
rect -6320 20920 -6280 20930
rect -6240 21430 -6200 21440
rect -6240 21410 -6230 21430
rect -6210 21410 -6200 21430
rect -6240 21270 -6200 21410
rect -6240 21250 -6230 21270
rect -6210 21250 -6200 21270
rect -6240 21110 -6200 21250
rect -6240 21090 -6230 21110
rect -6210 21090 -6200 21110
rect -6240 20950 -6200 21090
rect -6240 20930 -6230 20950
rect -6210 20930 -6200 20950
rect -6240 20920 -6200 20930
rect -6160 21430 -6120 21440
rect -6160 21410 -6150 21430
rect -6130 21410 -6120 21430
rect -6160 21270 -6120 21410
rect -6160 21250 -6150 21270
rect -6130 21250 -6120 21270
rect -6160 21110 -6120 21250
rect -6160 21090 -6150 21110
rect -6130 21090 -6120 21110
rect -6160 20950 -6120 21090
rect -6160 20930 -6150 20950
rect -6130 20930 -6120 20950
rect -6160 20920 -6120 20930
rect -5680 21430 -5640 21440
rect -5680 21410 -5670 21430
rect -5650 21410 -5640 21430
rect -5680 21270 -5640 21410
rect -5680 21250 -5670 21270
rect -5650 21250 -5640 21270
rect -5680 21110 -5640 21250
rect -5680 21090 -5670 21110
rect -5650 21090 -5640 21110
rect -5680 20950 -5640 21090
rect -5680 20930 -5670 20950
rect -5650 20930 -5640 20950
rect -5680 20920 -5640 20930
rect -5600 21430 -5560 21440
rect -5600 21410 -5590 21430
rect -5570 21410 -5560 21430
rect -5600 21270 -5560 21410
rect -5600 21250 -5590 21270
rect -5570 21250 -5560 21270
rect -5600 21110 -5560 21250
rect -5600 21090 -5590 21110
rect -5570 21090 -5560 21110
rect -5600 20950 -5560 21090
rect -5600 20930 -5590 20950
rect -5570 20930 -5560 20950
rect -5600 20920 -5560 20930
rect -5520 21430 -5480 21440
rect -5520 21410 -5510 21430
rect -5490 21410 -5480 21430
rect -5520 21270 -5480 21410
rect -5520 21250 -5510 21270
rect -5490 21250 -5480 21270
rect -5520 21110 -5480 21250
rect -5520 21090 -5510 21110
rect -5490 21090 -5480 21110
rect -5520 20950 -5480 21090
rect -5520 20930 -5510 20950
rect -5490 20930 -5480 20950
rect -5520 20920 -5480 20930
rect -5440 21430 -5400 21440
rect -5440 21410 -5430 21430
rect -5410 21410 -5400 21430
rect -5440 21270 -5400 21410
rect -5440 21250 -5430 21270
rect -5410 21250 -5400 21270
rect -5440 21110 -5400 21250
rect -5440 21090 -5430 21110
rect -5410 21090 -5400 21110
rect -5440 20950 -5400 21090
rect -5440 20930 -5430 20950
rect -5410 20930 -5400 20950
rect -5440 20920 -5400 20930
rect -5360 21430 -5320 21440
rect -5360 21410 -5350 21430
rect -5330 21410 -5320 21430
rect -5360 21270 -5320 21410
rect -5360 21250 -5350 21270
rect -5330 21250 -5320 21270
rect -5360 21110 -5320 21250
rect -5360 21090 -5350 21110
rect -5330 21090 -5320 21110
rect -5360 20950 -5320 21090
rect -5360 20930 -5350 20950
rect -5330 20930 -5320 20950
rect -5360 20920 -5320 20930
rect -5280 21430 -5240 21440
rect -5280 21410 -5270 21430
rect -5250 21410 -5240 21430
rect -5280 21270 -5240 21410
rect -5280 21250 -5270 21270
rect -5250 21250 -5240 21270
rect -5280 21110 -5240 21250
rect -5280 21090 -5270 21110
rect -5250 21090 -5240 21110
rect -5280 20950 -5240 21090
rect -5280 20930 -5270 20950
rect -5250 20930 -5240 20950
rect -5280 20920 -5240 20930
rect -5200 21430 -5160 21440
rect -5200 21410 -5190 21430
rect -5170 21410 -5160 21430
rect -5200 21270 -5160 21410
rect -5200 21250 -5190 21270
rect -5170 21250 -5160 21270
rect -5200 21110 -5160 21250
rect -5200 21090 -5190 21110
rect -5170 21090 -5160 21110
rect -5200 20950 -5160 21090
rect -5200 20930 -5190 20950
rect -5170 20930 -5160 20950
rect -5200 20920 -5160 20930
rect -5120 21430 -5080 21440
rect -5120 21410 -5110 21430
rect -5090 21410 -5080 21430
rect -5120 21270 -5080 21410
rect -5120 21250 -5110 21270
rect -5090 21250 -5080 21270
rect -5120 21110 -5080 21250
rect -5120 21090 -5110 21110
rect -5090 21090 -5080 21110
rect -5120 20950 -5080 21090
rect -5120 20930 -5110 20950
rect -5090 20930 -5080 20950
rect -5120 20920 -5080 20930
rect -5040 21430 -5000 21440
rect -5040 21410 -5030 21430
rect -5010 21410 -5000 21430
rect -5040 21270 -5000 21410
rect -5040 21250 -5030 21270
rect -5010 21250 -5000 21270
rect -5040 21110 -5000 21250
rect -5040 21090 -5030 21110
rect -5010 21090 -5000 21110
rect -5040 20950 -5000 21090
rect -5040 20930 -5030 20950
rect -5010 20930 -5000 20950
rect -5040 20920 -5000 20930
rect -4960 21430 -4920 21440
rect -4960 21410 -4950 21430
rect -4930 21410 -4920 21430
rect -4960 21270 -4920 21410
rect -4960 21250 -4950 21270
rect -4930 21250 -4920 21270
rect -4960 21110 -4920 21250
rect -4960 21090 -4950 21110
rect -4930 21090 -4920 21110
rect -4960 20950 -4920 21090
rect -4960 20930 -4950 20950
rect -4930 20930 -4920 20950
rect -4960 20920 -4920 20930
rect -4880 21430 -4840 21440
rect -4880 21410 -4870 21430
rect -4850 21410 -4840 21430
rect -4880 21270 -4840 21410
rect -4880 21250 -4870 21270
rect -4850 21250 -4840 21270
rect -4880 21110 -4840 21250
rect -4880 21090 -4870 21110
rect -4850 21090 -4840 21110
rect -4880 20950 -4840 21090
rect -4880 20930 -4870 20950
rect -4850 20930 -4840 20950
rect -4880 20920 -4840 20930
rect -4800 21430 -4760 21440
rect -4800 21410 -4790 21430
rect -4770 21410 -4760 21430
rect -4800 21270 -4760 21410
rect -4800 21250 -4790 21270
rect -4770 21250 -4760 21270
rect -4800 21110 -4760 21250
rect -4800 21090 -4790 21110
rect -4770 21090 -4760 21110
rect -4800 20950 -4760 21090
rect -4800 20930 -4790 20950
rect -4770 20930 -4760 20950
rect -4800 20920 -4760 20930
rect -4720 21430 -4680 21440
rect -4720 21410 -4710 21430
rect -4690 21410 -4680 21430
rect -4720 21270 -4680 21410
rect -4720 21250 -4710 21270
rect -4690 21250 -4680 21270
rect -4720 21110 -4680 21250
rect -4720 21090 -4710 21110
rect -4690 21090 -4680 21110
rect -4720 20950 -4680 21090
rect -4720 20930 -4710 20950
rect -4690 20930 -4680 20950
rect -4720 20920 -4680 20930
rect -4640 21430 -4600 21440
rect -4640 21410 -4630 21430
rect -4610 21410 -4600 21430
rect -4640 21270 -4600 21410
rect -4640 21250 -4630 21270
rect -4610 21250 -4600 21270
rect -4640 21110 -4600 21250
rect -4640 21090 -4630 21110
rect -4610 21090 -4600 21110
rect -4640 20950 -4600 21090
rect -4640 20930 -4630 20950
rect -4610 20930 -4600 20950
rect -4640 20920 -4600 20930
rect -4560 21430 -4520 21440
rect -4560 21410 -4550 21430
rect -4530 21410 -4520 21430
rect -4560 21270 -4520 21410
rect -4560 21250 -4550 21270
rect -4530 21250 -4520 21270
rect -4560 21110 -4520 21250
rect -4560 21090 -4550 21110
rect -4530 21090 -4520 21110
rect -4560 20950 -4520 21090
rect -4560 20930 -4550 20950
rect -4530 20930 -4520 20950
rect -4560 20920 -4520 20930
rect -4480 21430 -4440 21440
rect -4480 21410 -4470 21430
rect -4450 21410 -4440 21430
rect -4480 21270 -4440 21410
rect -4480 21250 -4470 21270
rect -4450 21250 -4440 21270
rect -4480 21110 -4440 21250
rect -4480 21090 -4470 21110
rect -4450 21090 -4440 21110
rect -4480 20950 -4440 21090
rect -4480 20930 -4470 20950
rect -4450 20930 -4440 20950
rect -4480 20920 -4440 20930
rect -4400 21430 -4360 21440
rect -4400 21410 -4390 21430
rect -4370 21410 -4360 21430
rect -4400 21270 -4360 21410
rect -4400 21250 -4390 21270
rect -4370 21250 -4360 21270
rect -4400 21110 -4360 21250
rect -4400 21090 -4390 21110
rect -4370 21090 -4360 21110
rect -4400 20950 -4360 21090
rect -4400 20930 -4390 20950
rect -4370 20930 -4360 20950
rect -4400 20920 -4360 20930
rect -4320 21430 -4280 21440
rect -4320 21410 -4310 21430
rect -4290 21410 -4280 21430
rect -4320 21270 -4280 21410
rect -4320 21250 -4310 21270
rect -4290 21250 -4280 21270
rect -4320 21110 -4280 21250
rect -4320 21090 -4310 21110
rect -4290 21090 -4280 21110
rect -4320 20950 -4280 21090
rect -4320 20930 -4310 20950
rect -4290 20930 -4280 20950
rect -4320 20920 -4280 20930
rect -4240 21430 -4200 21440
rect -4240 21410 -4230 21430
rect -4210 21410 -4200 21430
rect -4240 21270 -4200 21410
rect -4240 21250 -4230 21270
rect -4210 21250 -4200 21270
rect -4240 21110 -4200 21250
rect -4240 21090 -4230 21110
rect -4210 21090 -4200 21110
rect -4240 20950 -4200 21090
rect -4240 20930 -4230 20950
rect -4210 20930 -4200 20950
rect -4240 20920 -4200 20930
rect -4160 21430 -4120 21440
rect -4160 21410 -4150 21430
rect -4130 21410 -4120 21430
rect -4160 21270 -4120 21410
rect -4160 21250 -4150 21270
rect -4130 21250 -4120 21270
rect -4160 21110 -4120 21250
rect -4160 21090 -4150 21110
rect -4130 21090 -4120 21110
rect -4160 20950 -4120 21090
rect -4160 20930 -4150 20950
rect -4130 20930 -4120 20950
rect -4160 20920 -4120 20930
rect -4080 21430 -4040 21440
rect -4080 21410 -4070 21430
rect -4050 21410 -4040 21430
rect -4080 21270 -4040 21410
rect -4080 21250 -4070 21270
rect -4050 21250 -4040 21270
rect -4080 21110 -4040 21250
rect -4080 21090 -4070 21110
rect -4050 21090 -4040 21110
rect -4080 20950 -4040 21090
rect -4080 20930 -4070 20950
rect -4050 20930 -4040 20950
rect -4080 20920 -4040 20930
rect -4000 21430 -3960 21440
rect -4000 21410 -3990 21430
rect -3970 21410 -3960 21430
rect -4000 21270 -3960 21410
rect -4000 21250 -3990 21270
rect -3970 21250 -3960 21270
rect -4000 21110 -3960 21250
rect -4000 21090 -3990 21110
rect -3970 21090 -3960 21110
rect -4000 20950 -3960 21090
rect -4000 20930 -3990 20950
rect -3970 20930 -3960 20950
rect -4000 20920 -3960 20930
rect -3920 21430 -3880 21440
rect -3920 21410 -3910 21430
rect -3890 21410 -3880 21430
rect -3920 21270 -3880 21410
rect -3920 21250 -3910 21270
rect -3890 21250 -3880 21270
rect -3920 21110 -3880 21250
rect -3920 21090 -3910 21110
rect -3890 21090 -3880 21110
rect -3920 20950 -3880 21090
rect -3920 20930 -3910 20950
rect -3890 20930 -3880 20950
rect -3920 20920 -3880 20930
rect -3840 21430 -3800 21440
rect -3840 21410 -3830 21430
rect -3810 21410 -3800 21430
rect -3840 21270 -3800 21410
rect -3840 21250 -3830 21270
rect -3810 21250 -3800 21270
rect -3840 21110 -3800 21250
rect -3840 21090 -3830 21110
rect -3810 21090 -3800 21110
rect -3840 20950 -3800 21090
rect -3840 20930 -3830 20950
rect -3810 20930 -3800 20950
rect -3840 20920 -3800 20930
rect -3760 21430 -3720 21440
rect -3760 21410 -3750 21430
rect -3730 21410 -3720 21430
rect -3760 21270 -3720 21410
rect -3760 21250 -3750 21270
rect -3730 21250 -3720 21270
rect -3760 21110 -3720 21250
rect -3760 21090 -3750 21110
rect -3730 21090 -3720 21110
rect -3760 20950 -3720 21090
rect -3760 20930 -3750 20950
rect -3730 20930 -3720 20950
rect -3760 20920 -3720 20930
rect -3680 21430 -3640 21440
rect -3680 21410 -3670 21430
rect -3650 21410 -3640 21430
rect -3680 21270 -3640 21410
rect -3680 21250 -3670 21270
rect -3650 21250 -3640 21270
rect -3680 21110 -3640 21250
rect -3680 21090 -3670 21110
rect -3650 21090 -3640 21110
rect -3680 20950 -3640 21090
rect -3680 20930 -3670 20950
rect -3650 20930 -3640 20950
rect -3680 20920 -3640 20930
rect -3600 21430 -3560 21440
rect -3600 21410 -3590 21430
rect -3570 21410 -3560 21430
rect -3600 21270 -3560 21410
rect -3600 21250 -3590 21270
rect -3570 21250 -3560 21270
rect -3600 21110 -3560 21250
rect -3600 21090 -3590 21110
rect -3570 21090 -3560 21110
rect -3600 20950 -3560 21090
rect -3600 20930 -3590 20950
rect -3570 20930 -3560 20950
rect -3600 20920 -3560 20930
rect -3520 21430 -3480 21440
rect -3520 21410 -3510 21430
rect -3490 21410 -3480 21430
rect -3520 21270 -3480 21410
rect -3520 21250 -3510 21270
rect -3490 21250 -3480 21270
rect -3520 21110 -3480 21250
rect -3520 21090 -3510 21110
rect -3490 21090 -3480 21110
rect -3520 20950 -3480 21090
rect -3520 20930 -3510 20950
rect -3490 20930 -3480 20950
rect -3520 20920 -3480 20930
rect -3440 21430 -3400 21440
rect -3440 21410 -3430 21430
rect -3410 21410 -3400 21430
rect -3440 21270 -3400 21410
rect -3440 21250 -3430 21270
rect -3410 21250 -3400 21270
rect -3440 21110 -3400 21250
rect -3440 21090 -3430 21110
rect -3410 21090 -3400 21110
rect -3440 20950 -3400 21090
rect -3440 20930 -3430 20950
rect -3410 20930 -3400 20950
rect -3440 20920 -3400 20930
rect -3360 21430 -3320 21440
rect -3360 21410 -3350 21430
rect -3330 21410 -3320 21430
rect -3360 21270 -3320 21410
rect -3360 21250 -3350 21270
rect -3330 21250 -3320 21270
rect -3360 21110 -3320 21250
rect -3360 21090 -3350 21110
rect -3330 21090 -3320 21110
rect -3360 20950 -3320 21090
rect -3360 20930 -3350 20950
rect -3330 20930 -3320 20950
rect -3360 20920 -3320 20930
rect -3280 21430 -3240 21440
rect -3280 21410 -3270 21430
rect -3250 21410 -3240 21430
rect -3280 21270 -3240 21410
rect -3280 21250 -3270 21270
rect -3250 21250 -3240 21270
rect -3280 21110 -3240 21250
rect -3280 21090 -3270 21110
rect -3250 21090 -3240 21110
rect -3280 20950 -3240 21090
rect -3280 20930 -3270 20950
rect -3250 20930 -3240 20950
rect -3280 20920 -3240 20930
rect -3200 21430 -3160 21440
rect -3200 21410 -3190 21430
rect -3170 21410 -3160 21430
rect -3200 21270 -3160 21410
rect -3200 21250 -3190 21270
rect -3170 21250 -3160 21270
rect -3200 21110 -3160 21250
rect -3200 21090 -3190 21110
rect -3170 21090 -3160 21110
rect -3200 20950 -3160 21090
rect -3200 20930 -3190 20950
rect -3170 20930 -3160 20950
rect -3200 20920 -3160 20930
rect -3120 21430 -3080 21440
rect -3120 21410 -3110 21430
rect -3090 21410 -3080 21430
rect -3120 21270 -3080 21410
rect -3120 21250 -3110 21270
rect -3090 21250 -3080 21270
rect -3120 21110 -3080 21250
rect -3120 21090 -3110 21110
rect -3090 21090 -3080 21110
rect -3120 20950 -3080 21090
rect -3120 20930 -3110 20950
rect -3090 20930 -3080 20950
rect -3120 20920 -3080 20930
rect -3040 21430 -3000 21440
rect -3040 21410 -3030 21430
rect -3010 21410 -3000 21430
rect -3040 21270 -3000 21410
rect -3040 21250 -3030 21270
rect -3010 21250 -3000 21270
rect -3040 21110 -3000 21250
rect -3040 21090 -3030 21110
rect -3010 21090 -3000 21110
rect -3040 20950 -3000 21090
rect -3040 20930 -3030 20950
rect -3010 20930 -3000 20950
rect -3040 20920 -3000 20930
rect -2960 21430 -2920 21440
rect -2960 21410 -2950 21430
rect -2930 21410 -2920 21430
rect -2960 21270 -2920 21410
rect -2960 21250 -2950 21270
rect -2930 21250 -2920 21270
rect -2960 21110 -2920 21250
rect -2960 21090 -2950 21110
rect -2930 21090 -2920 21110
rect -2960 20950 -2920 21090
rect -2960 20930 -2950 20950
rect -2930 20930 -2920 20950
rect -2960 20920 -2920 20930
rect -2880 21430 -2840 21440
rect -2880 21410 -2870 21430
rect -2850 21410 -2840 21430
rect -2880 21270 -2840 21410
rect -2880 21250 -2870 21270
rect -2850 21250 -2840 21270
rect -2880 21110 -2840 21250
rect -2880 21090 -2870 21110
rect -2850 21090 -2840 21110
rect -2880 20950 -2840 21090
rect -2880 20930 -2870 20950
rect -2850 20930 -2840 20950
rect -2880 20920 -2840 20930
rect -2800 21430 -2760 21440
rect -2800 21410 -2790 21430
rect -2770 21410 -2760 21430
rect -2800 21270 -2760 21410
rect -2800 21250 -2790 21270
rect -2770 21250 -2760 21270
rect -2800 21110 -2760 21250
rect -2800 21090 -2790 21110
rect -2770 21090 -2760 21110
rect -2800 20950 -2760 21090
rect -2800 20930 -2790 20950
rect -2770 20930 -2760 20950
rect -2800 20920 -2760 20930
rect -2720 21430 -2680 21440
rect -2720 21410 -2710 21430
rect -2690 21410 -2680 21430
rect -2720 21270 -2680 21410
rect -2720 21250 -2710 21270
rect -2690 21250 -2680 21270
rect -2720 21110 -2680 21250
rect -2720 21090 -2710 21110
rect -2690 21090 -2680 21110
rect -2720 20950 -2680 21090
rect -2720 20930 -2710 20950
rect -2690 20930 -2680 20950
rect -2720 20920 -2680 20930
rect -2640 21430 -2600 21440
rect -2640 21410 -2630 21430
rect -2610 21410 -2600 21430
rect -2640 21270 -2600 21410
rect -2640 21250 -2630 21270
rect -2610 21250 -2600 21270
rect -2640 21110 -2600 21250
rect -2640 21090 -2630 21110
rect -2610 21090 -2600 21110
rect -2640 20950 -2600 21090
rect -2640 20930 -2630 20950
rect -2610 20930 -2600 20950
rect -2640 20920 -2600 20930
rect -2560 21430 -2520 21440
rect -2560 21410 -2550 21430
rect -2530 21410 -2520 21430
rect -2560 21270 -2520 21410
rect -2560 21250 -2550 21270
rect -2530 21250 -2520 21270
rect -2560 21110 -2520 21250
rect -2560 21090 -2550 21110
rect -2530 21090 -2520 21110
rect -2560 20950 -2520 21090
rect -2560 20930 -2550 20950
rect -2530 20930 -2520 20950
rect -2560 20920 -2520 20930
rect -2480 21430 -2440 21440
rect -2480 21410 -2470 21430
rect -2450 21410 -2440 21430
rect -2480 21270 -2440 21410
rect -2480 21250 -2470 21270
rect -2450 21250 -2440 21270
rect -2480 21110 -2440 21250
rect -2480 21090 -2470 21110
rect -2450 21090 -2440 21110
rect -2480 20950 -2440 21090
rect -2480 20930 -2470 20950
rect -2450 20930 -2440 20950
rect -2480 20920 -2440 20930
rect -2400 21430 -2360 21440
rect -2400 21410 -2390 21430
rect -2370 21410 -2360 21430
rect -2400 21270 -2360 21410
rect -2400 21250 -2390 21270
rect -2370 21250 -2360 21270
rect -2400 21110 -2360 21250
rect -2400 21090 -2390 21110
rect -2370 21090 -2360 21110
rect -2400 20950 -2360 21090
rect -2400 20930 -2390 20950
rect -2370 20930 -2360 20950
rect -2400 20920 -2360 20930
rect -2320 21430 -2280 21440
rect -2320 21410 -2310 21430
rect -2290 21410 -2280 21430
rect -2320 21270 -2280 21410
rect -2320 21250 -2310 21270
rect -2290 21250 -2280 21270
rect -2320 21110 -2280 21250
rect -2320 21090 -2310 21110
rect -2290 21090 -2280 21110
rect -2320 20950 -2280 21090
rect -2320 20930 -2310 20950
rect -2290 20930 -2280 20950
rect -2320 20920 -2280 20930
rect -2240 21430 -2200 21440
rect -2240 21410 -2230 21430
rect -2210 21410 -2200 21430
rect -2240 21270 -2200 21410
rect -2240 21250 -2230 21270
rect -2210 21250 -2200 21270
rect -2240 21110 -2200 21250
rect -2240 21090 -2230 21110
rect -2210 21090 -2200 21110
rect -2240 20950 -2200 21090
rect -2240 20930 -2230 20950
rect -2210 20930 -2200 20950
rect -2240 20920 -2200 20930
rect -2160 21430 -2120 21440
rect -2160 21410 -2150 21430
rect -2130 21410 -2120 21430
rect -2160 21270 -2120 21410
rect -2160 21250 -2150 21270
rect -2130 21250 -2120 21270
rect -2160 21110 -2120 21250
rect -2160 21090 -2150 21110
rect -2130 21090 -2120 21110
rect -2160 20950 -2120 21090
rect -2160 20930 -2150 20950
rect -2130 20930 -2120 20950
rect -2160 20920 -2120 20930
rect -2080 21430 -2040 21440
rect -2080 21410 -2070 21430
rect -2050 21410 -2040 21430
rect -2080 21270 -2040 21410
rect -2080 21250 -2070 21270
rect -2050 21250 -2040 21270
rect -2080 21110 -2040 21250
rect -2080 21090 -2070 21110
rect -2050 21090 -2040 21110
rect -2080 20950 -2040 21090
rect -2080 20930 -2070 20950
rect -2050 20930 -2040 20950
rect -2080 20920 -2040 20930
rect -2000 21430 -1960 21440
rect -2000 21410 -1990 21430
rect -1970 21410 -1960 21430
rect -2000 21270 -1960 21410
rect -2000 21250 -1990 21270
rect -1970 21250 -1960 21270
rect -2000 21110 -1960 21250
rect -2000 21090 -1990 21110
rect -1970 21090 -1960 21110
rect -2000 20950 -1960 21090
rect -2000 20930 -1990 20950
rect -1970 20930 -1960 20950
rect -2000 20920 -1960 20930
rect -16560 20670 -16520 20680
rect -16560 20650 -16550 20670
rect -16530 20650 -16520 20670
rect -16560 20510 -16520 20650
rect -16560 20490 -16550 20510
rect -16530 20490 -16520 20510
rect -16560 20480 -16520 20490
rect -16480 20670 -16440 20680
rect -16480 20650 -16470 20670
rect -16450 20650 -16440 20670
rect -16480 20510 -16440 20650
rect -16480 20490 -16470 20510
rect -16450 20490 -16440 20510
rect -16480 20480 -16440 20490
rect -16400 20670 -16360 20680
rect -16400 20650 -16390 20670
rect -16370 20650 -16360 20670
rect -16400 20510 -16360 20650
rect -16400 20490 -16390 20510
rect -16370 20490 -16360 20510
rect -16400 20480 -16360 20490
rect -16320 20670 -16280 20680
rect -16320 20650 -16310 20670
rect -16290 20650 -16280 20670
rect -16320 20510 -16280 20650
rect -16320 20490 -16310 20510
rect -16290 20490 -16280 20510
rect -16320 20480 -16280 20490
rect -16240 20670 -16200 20680
rect -16240 20650 -16230 20670
rect -16210 20650 -16200 20670
rect -16240 20510 -16200 20650
rect -16240 20490 -16230 20510
rect -16210 20490 -16200 20510
rect -16240 20480 -16200 20490
rect -16160 20670 -16120 20680
rect -16160 20650 -16150 20670
rect -16130 20650 -16120 20670
rect -16160 20510 -16120 20650
rect -16160 20490 -16150 20510
rect -16130 20490 -16120 20510
rect -16160 20480 -16120 20490
rect -16080 20670 -16040 20680
rect -16080 20650 -16070 20670
rect -16050 20650 -16040 20670
rect -16080 20510 -16040 20650
rect -16080 20490 -16070 20510
rect -16050 20490 -16040 20510
rect -16080 20480 -16040 20490
rect -16000 20670 -15960 20680
rect -16000 20650 -15990 20670
rect -15970 20650 -15960 20670
rect -16000 20510 -15960 20650
rect -16000 20490 -15990 20510
rect -15970 20490 -15960 20510
rect -16000 20480 -15960 20490
rect -15920 20670 -15880 20680
rect -15920 20650 -15910 20670
rect -15890 20650 -15880 20670
rect -15920 20510 -15880 20650
rect -15920 20490 -15910 20510
rect -15890 20490 -15880 20510
rect -15920 20480 -15880 20490
rect -15840 20670 -15800 20680
rect -15840 20650 -15830 20670
rect -15810 20650 -15800 20670
rect -15840 20510 -15800 20650
rect -15840 20490 -15830 20510
rect -15810 20490 -15800 20510
rect -15840 20480 -15800 20490
rect -15760 20670 -15720 20680
rect -15760 20650 -15750 20670
rect -15730 20650 -15720 20670
rect -15760 20510 -15720 20650
rect -15760 20490 -15750 20510
rect -15730 20490 -15720 20510
rect -15760 20480 -15720 20490
rect -15680 20670 -15640 20680
rect -15680 20650 -15670 20670
rect -15650 20650 -15640 20670
rect -15680 20510 -15640 20650
rect -15680 20490 -15670 20510
rect -15650 20490 -15640 20510
rect -15680 20480 -15640 20490
rect -15600 20670 -15560 20680
rect -15600 20650 -15590 20670
rect -15570 20650 -15560 20670
rect -15600 20510 -15560 20650
rect -15600 20490 -15590 20510
rect -15570 20490 -15560 20510
rect -15600 20480 -15560 20490
rect -14960 20670 -14920 20680
rect -14960 20650 -14950 20670
rect -14930 20650 -14920 20670
rect -14960 20510 -14920 20650
rect -14960 20490 -14950 20510
rect -14930 20490 -14920 20510
rect -14960 20480 -14920 20490
rect -14880 20670 -14840 20680
rect -14880 20650 -14870 20670
rect -14850 20650 -14840 20670
rect -14880 20510 -14840 20650
rect -14880 20490 -14870 20510
rect -14850 20490 -14840 20510
rect -14880 20480 -14840 20490
rect -14800 20670 -14760 20680
rect -14800 20650 -14790 20670
rect -14770 20650 -14760 20670
rect -14800 20510 -14760 20650
rect -14800 20490 -14790 20510
rect -14770 20490 -14760 20510
rect -14800 20480 -14760 20490
rect -14720 20670 -14680 20680
rect -14720 20650 -14710 20670
rect -14690 20650 -14680 20670
rect -14720 20510 -14680 20650
rect -14720 20490 -14710 20510
rect -14690 20490 -14680 20510
rect -14720 20480 -14680 20490
rect -14640 20670 -14600 20680
rect -14640 20650 -14630 20670
rect -14610 20650 -14600 20670
rect -14640 20510 -14600 20650
rect -14640 20490 -14630 20510
rect -14610 20490 -14600 20510
rect -14640 20480 -14600 20490
rect -14560 20670 -14520 20680
rect -14560 20650 -14550 20670
rect -14530 20650 -14520 20670
rect -14560 20510 -14520 20650
rect -14560 20490 -14550 20510
rect -14530 20490 -14520 20510
rect -14560 20480 -14520 20490
rect -14480 20670 -14440 20680
rect -14480 20650 -14470 20670
rect -14450 20650 -14440 20670
rect -14480 20510 -14440 20650
rect -14480 20490 -14470 20510
rect -14450 20490 -14440 20510
rect -14480 20480 -14440 20490
rect -14400 20670 -14360 20680
rect -14400 20650 -14390 20670
rect -14370 20650 -14360 20670
rect -14400 20510 -14360 20650
rect -14400 20490 -14390 20510
rect -14370 20490 -14360 20510
rect -14400 20480 -14360 20490
rect -14320 20670 -14280 20680
rect -14320 20650 -14310 20670
rect -14290 20650 -14280 20670
rect -14320 20510 -14280 20650
rect -14320 20490 -14310 20510
rect -14290 20490 -14280 20510
rect -14320 20480 -14280 20490
rect -14240 20670 -14200 20680
rect -14240 20650 -14230 20670
rect -14210 20650 -14200 20670
rect -14240 20510 -14200 20650
rect -14240 20490 -14230 20510
rect -14210 20490 -14200 20510
rect -14240 20480 -14200 20490
rect -14160 20670 -14120 20680
rect -14160 20650 -14150 20670
rect -14130 20650 -14120 20670
rect -14160 20510 -14120 20650
rect -14160 20490 -14150 20510
rect -14130 20490 -14120 20510
rect -14160 20480 -14120 20490
rect -14080 20670 -14040 20680
rect -14080 20650 -14070 20670
rect -14050 20650 -14040 20670
rect -14080 20510 -14040 20650
rect -14080 20490 -14070 20510
rect -14050 20490 -14040 20510
rect -14080 20480 -14040 20490
rect -14000 20670 -13960 20680
rect -14000 20650 -13990 20670
rect -13970 20650 -13960 20670
rect -14000 20510 -13960 20650
rect -14000 20490 -13990 20510
rect -13970 20490 -13960 20510
rect -14000 20480 -13960 20490
rect -13920 20670 -13880 20680
rect -13920 20650 -13910 20670
rect -13890 20650 -13880 20670
rect -13920 20510 -13880 20650
rect -13920 20490 -13910 20510
rect -13890 20490 -13880 20510
rect -13920 20480 -13880 20490
rect -13840 20670 -13800 20680
rect -13840 20650 -13830 20670
rect -13810 20650 -13800 20670
rect -13840 20510 -13800 20650
rect -13840 20490 -13830 20510
rect -13810 20490 -13800 20510
rect -13840 20480 -13800 20490
rect -13760 20670 -13720 20680
rect -13760 20650 -13750 20670
rect -13730 20650 -13720 20670
rect -13760 20510 -13720 20650
rect -13760 20490 -13750 20510
rect -13730 20490 -13720 20510
rect -13760 20480 -13720 20490
rect -13680 20670 -13640 20680
rect -13680 20650 -13670 20670
rect -13650 20650 -13640 20670
rect -13680 20510 -13640 20650
rect -13680 20490 -13670 20510
rect -13650 20490 -13640 20510
rect -13680 20480 -13640 20490
rect -13600 20670 -13560 20680
rect -13600 20650 -13590 20670
rect -13570 20650 -13560 20670
rect -13600 20510 -13560 20650
rect -13600 20490 -13590 20510
rect -13570 20490 -13560 20510
rect -13600 20480 -13560 20490
rect -13520 20670 -13480 20680
rect -13520 20650 -13510 20670
rect -13490 20650 -13480 20670
rect -13520 20510 -13480 20650
rect -13520 20490 -13510 20510
rect -13490 20490 -13480 20510
rect -13520 20480 -13480 20490
rect -13440 20670 -13400 20680
rect -13440 20650 -13430 20670
rect -13410 20650 -13400 20670
rect -13440 20510 -13400 20650
rect -13440 20490 -13430 20510
rect -13410 20490 -13400 20510
rect -13440 20480 -13400 20490
rect -13360 20670 -13320 20680
rect -13360 20650 -13350 20670
rect -13330 20650 -13320 20670
rect -13360 20510 -13320 20650
rect -13360 20490 -13350 20510
rect -13330 20490 -13320 20510
rect -13360 20480 -13320 20490
rect -13280 20670 -13240 20680
rect -13280 20650 -13270 20670
rect -13250 20650 -13240 20670
rect -13280 20510 -13240 20650
rect -13280 20490 -13270 20510
rect -13250 20490 -13240 20510
rect -13280 20480 -13240 20490
rect -13200 20670 -13160 20680
rect -13200 20650 -13190 20670
rect -13170 20650 -13160 20670
rect -13200 20510 -13160 20650
rect -13200 20490 -13190 20510
rect -13170 20490 -13160 20510
rect -13200 20480 -13160 20490
rect -13120 20670 -13080 20680
rect -13120 20650 -13110 20670
rect -13090 20650 -13080 20670
rect -13120 20510 -13080 20650
rect -13120 20490 -13110 20510
rect -13090 20490 -13080 20510
rect -13120 20480 -13080 20490
rect -13040 20670 -13000 20680
rect -13040 20650 -13030 20670
rect -13010 20650 -13000 20670
rect -13040 20510 -13000 20650
rect -13040 20490 -13030 20510
rect -13010 20490 -13000 20510
rect -13040 20480 -13000 20490
rect -12960 20670 -12920 20680
rect -12960 20650 -12950 20670
rect -12930 20650 -12920 20670
rect -12960 20510 -12920 20650
rect -12960 20490 -12950 20510
rect -12930 20490 -12920 20510
rect -12960 20480 -12920 20490
rect -12880 20670 -12840 20680
rect -12880 20650 -12870 20670
rect -12850 20650 -12840 20670
rect -12880 20510 -12840 20650
rect -12880 20490 -12870 20510
rect -12850 20490 -12840 20510
rect -12880 20480 -12840 20490
rect -12800 20670 -12760 20680
rect -12800 20650 -12790 20670
rect -12770 20650 -12760 20670
rect -12800 20510 -12760 20650
rect -12800 20490 -12790 20510
rect -12770 20490 -12760 20510
rect -12800 20480 -12760 20490
rect -12720 20670 -12680 20680
rect -12720 20650 -12710 20670
rect -12690 20650 -12680 20670
rect -12720 20510 -12680 20650
rect -12720 20490 -12710 20510
rect -12690 20490 -12680 20510
rect -12720 20480 -12680 20490
rect -12640 20670 -12600 20680
rect -12640 20650 -12630 20670
rect -12610 20650 -12600 20670
rect -12640 20510 -12600 20650
rect -12640 20490 -12630 20510
rect -12610 20490 -12600 20510
rect -12640 20480 -12600 20490
rect -12560 20670 -12520 20680
rect -12560 20650 -12550 20670
rect -12530 20650 -12520 20670
rect -12560 20510 -12520 20650
rect -12560 20490 -12550 20510
rect -12530 20490 -12520 20510
rect -12560 20480 -12520 20490
rect -12480 20670 -12440 20680
rect -12480 20650 -12470 20670
rect -12450 20650 -12440 20670
rect -12480 20510 -12440 20650
rect -12480 20490 -12470 20510
rect -12450 20490 -12440 20510
rect -12480 20480 -12440 20490
rect -12400 20670 -12360 20680
rect -12400 20650 -12390 20670
rect -12370 20650 -12360 20670
rect -12400 20510 -12360 20650
rect -12400 20490 -12390 20510
rect -12370 20490 -12360 20510
rect -12400 20480 -12360 20490
rect -12320 20670 -12280 20680
rect -12320 20650 -12310 20670
rect -12290 20650 -12280 20670
rect -12320 20510 -12280 20650
rect -12320 20490 -12310 20510
rect -12290 20490 -12280 20510
rect -12320 20480 -12280 20490
rect -12240 20670 -12200 20680
rect -12240 20650 -12230 20670
rect -12210 20650 -12200 20670
rect -12240 20510 -12200 20650
rect -12240 20490 -12230 20510
rect -12210 20490 -12200 20510
rect -12240 20480 -12200 20490
rect -12160 20670 -12120 20680
rect -12160 20650 -12150 20670
rect -12130 20650 -12120 20670
rect -12160 20510 -12120 20650
rect -12160 20490 -12150 20510
rect -12130 20490 -12120 20510
rect -12160 20480 -12120 20490
rect -12080 20670 -12040 20680
rect -12080 20650 -12070 20670
rect -12050 20650 -12040 20670
rect -12080 20510 -12040 20650
rect -12080 20490 -12070 20510
rect -12050 20490 -12040 20510
rect -12080 20480 -12040 20490
rect -12000 20670 -11960 20680
rect -12000 20650 -11990 20670
rect -11970 20650 -11960 20670
rect -12000 20510 -11960 20650
rect -12000 20490 -11990 20510
rect -11970 20490 -11960 20510
rect -12000 20480 -11960 20490
rect -11920 20670 -11880 20680
rect -11920 20650 -11910 20670
rect -11890 20650 -11880 20670
rect -11920 20510 -11880 20650
rect -11920 20490 -11910 20510
rect -11890 20490 -11880 20510
rect -11920 20480 -11880 20490
rect -11840 20670 -11800 20680
rect -11840 20650 -11830 20670
rect -11810 20650 -11800 20670
rect -11840 20510 -11800 20650
rect -11840 20490 -11830 20510
rect -11810 20490 -11800 20510
rect -11840 20480 -11800 20490
rect -11760 20670 -11720 20680
rect -11760 20650 -11750 20670
rect -11730 20650 -11720 20670
rect -11760 20510 -11720 20650
rect -11760 20490 -11750 20510
rect -11730 20490 -11720 20510
rect -11760 20480 -11720 20490
rect -11680 20670 -11640 20680
rect -11680 20650 -11670 20670
rect -11650 20650 -11640 20670
rect -11680 20510 -11640 20650
rect -11680 20490 -11670 20510
rect -11650 20490 -11640 20510
rect -11680 20480 -11640 20490
rect -11600 20670 -11560 20680
rect -11600 20650 -11590 20670
rect -11570 20650 -11560 20670
rect -11600 20510 -11560 20650
rect -11600 20490 -11590 20510
rect -11570 20490 -11560 20510
rect -11600 20480 -11560 20490
rect -11520 20670 -11480 20680
rect -11520 20650 -11510 20670
rect -11490 20650 -11480 20670
rect -11520 20510 -11480 20650
rect -11520 20490 -11510 20510
rect -11490 20490 -11480 20510
rect -11520 20480 -11480 20490
rect -11440 20670 -11400 20680
rect -11440 20650 -11430 20670
rect -11410 20650 -11400 20670
rect -11440 20510 -11400 20650
rect -11440 20490 -11430 20510
rect -11410 20490 -11400 20510
rect -11440 20480 -11400 20490
rect -11360 20670 -11320 20680
rect -11360 20650 -11350 20670
rect -11330 20650 -11320 20670
rect -11360 20510 -11320 20650
rect -11360 20490 -11350 20510
rect -11330 20490 -11320 20510
rect -11360 20480 -11320 20490
rect -11280 20670 -11240 20680
rect -11280 20650 -11270 20670
rect -11250 20650 -11240 20670
rect -11280 20510 -11240 20650
rect -11280 20490 -11270 20510
rect -11250 20490 -11240 20510
rect -11280 20480 -11240 20490
rect -11200 20670 -11160 20680
rect -11200 20650 -11190 20670
rect -11170 20650 -11160 20670
rect -11200 20510 -11160 20650
rect -11200 20490 -11190 20510
rect -11170 20490 -11160 20510
rect -11200 20480 -11160 20490
rect -11120 20670 -11080 20680
rect -11120 20650 -11110 20670
rect -11090 20650 -11080 20670
rect -11120 20510 -11080 20650
rect -11120 20490 -11110 20510
rect -11090 20490 -11080 20510
rect -11120 20480 -11080 20490
rect -11040 20670 -11000 20680
rect -11040 20650 -11030 20670
rect -11010 20650 -11000 20670
rect -11040 20510 -11000 20650
rect -11040 20490 -11030 20510
rect -11010 20490 -11000 20510
rect -11040 20480 -11000 20490
rect -10960 20670 -10920 20680
rect -10960 20650 -10950 20670
rect -10930 20650 -10920 20670
rect -10960 20510 -10920 20650
rect -10960 20490 -10950 20510
rect -10930 20490 -10920 20510
rect -10960 20480 -10920 20490
rect -10880 20670 -10840 20680
rect -10880 20650 -10870 20670
rect -10850 20650 -10840 20670
rect -10880 20510 -10840 20650
rect -10880 20490 -10870 20510
rect -10850 20490 -10840 20510
rect -10880 20480 -10840 20490
rect -10800 20670 -10760 20680
rect -10800 20650 -10790 20670
rect -10770 20650 -10760 20670
rect -10800 20510 -10760 20650
rect -10800 20490 -10790 20510
rect -10770 20490 -10760 20510
rect -10800 20480 -10760 20490
rect -10720 20670 -10680 20680
rect -10720 20650 -10710 20670
rect -10690 20650 -10680 20670
rect -10720 20510 -10680 20650
rect -10720 20490 -10710 20510
rect -10690 20490 -10680 20510
rect -10720 20480 -10680 20490
rect -10640 20670 -10600 20680
rect -10640 20650 -10630 20670
rect -10610 20650 -10600 20670
rect -10640 20510 -10600 20650
rect -10640 20490 -10630 20510
rect -10610 20490 -10600 20510
rect -10640 20480 -10600 20490
rect -10560 20670 -10520 20680
rect -10560 20650 -10550 20670
rect -10530 20650 -10520 20670
rect -10560 20510 -10520 20650
rect -10560 20490 -10550 20510
rect -10530 20490 -10520 20510
rect -10560 20480 -10520 20490
rect -10480 20670 -10440 20680
rect -10480 20650 -10470 20670
rect -10450 20650 -10440 20670
rect -10480 20510 -10440 20650
rect -10480 20490 -10470 20510
rect -10450 20490 -10440 20510
rect -10480 20480 -10440 20490
rect -10400 20670 -10360 20680
rect -10400 20650 -10390 20670
rect -10370 20650 -10360 20670
rect -10400 20510 -10360 20650
rect -10400 20490 -10390 20510
rect -10370 20490 -10360 20510
rect -10400 20480 -10360 20490
rect -10320 20670 -10280 20680
rect -10320 20650 -10310 20670
rect -10290 20650 -10280 20670
rect -10320 20510 -10280 20650
rect -10320 20490 -10310 20510
rect -10290 20490 -10280 20510
rect -10320 20480 -10280 20490
rect -10240 20670 -10200 20680
rect -10240 20650 -10230 20670
rect -10210 20650 -10200 20670
rect -10240 20510 -10200 20650
rect -10240 20490 -10230 20510
rect -10210 20490 -10200 20510
rect -10240 20480 -10200 20490
rect -10160 20670 -10120 20680
rect -10160 20650 -10150 20670
rect -10130 20650 -10120 20670
rect -10160 20510 -10120 20650
rect -10160 20490 -10150 20510
rect -10130 20490 -10120 20510
rect -10160 20480 -10120 20490
rect -10080 20670 -10040 20680
rect -10080 20650 -10070 20670
rect -10050 20650 -10040 20670
rect -10080 20510 -10040 20650
rect -10080 20490 -10070 20510
rect -10050 20490 -10040 20510
rect -10080 20480 -10040 20490
rect -10000 20670 -9960 20680
rect -10000 20650 -9990 20670
rect -9970 20650 -9960 20670
rect -10000 20510 -9960 20650
rect -10000 20490 -9990 20510
rect -9970 20490 -9960 20510
rect -10000 20480 -9960 20490
rect -9920 20670 -9880 20680
rect -9920 20650 -9910 20670
rect -9890 20650 -9880 20670
rect -9920 20510 -9880 20650
rect -9920 20490 -9910 20510
rect -9890 20490 -9880 20510
rect -9920 20480 -9880 20490
rect -9840 20670 -9800 20680
rect -9840 20650 -9830 20670
rect -9810 20650 -9800 20670
rect -9840 20510 -9800 20650
rect -9840 20490 -9830 20510
rect -9810 20490 -9800 20510
rect -9840 20480 -9800 20490
rect -9760 20670 -9720 20680
rect -9760 20650 -9750 20670
rect -9730 20650 -9720 20670
rect -9760 20510 -9720 20650
rect -9760 20490 -9750 20510
rect -9730 20490 -9720 20510
rect -9760 20480 -9720 20490
rect -9680 20670 -9640 20680
rect -9680 20650 -9670 20670
rect -9650 20650 -9640 20670
rect -9680 20510 -9640 20650
rect -9680 20490 -9670 20510
rect -9650 20490 -9640 20510
rect -9680 20480 -9640 20490
rect -9600 20670 -9560 20680
rect -9600 20650 -9590 20670
rect -9570 20650 -9560 20670
rect -9600 20510 -9560 20650
rect -9600 20490 -9590 20510
rect -9570 20490 -9560 20510
rect -9600 20480 -9560 20490
rect -9520 20670 -9480 20680
rect -9520 20650 -9510 20670
rect -9490 20650 -9480 20670
rect -9520 20510 -9480 20650
rect -9520 20490 -9510 20510
rect -9490 20490 -9480 20510
rect -9520 20480 -9480 20490
rect -9440 20670 -9400 20680
rect -9440 20650 -9430 20670
rect -9410 20650 -9400 20670
rect -9440 20510 -9400 20650
rect -9440 20490 -9430 20510
rect -9410 20490 -9400 20510
rect -9440 20480 -9400 20490
rect -9360 20670 -9320 20680
rect -9360 20650 -9350 20670
rect -9330 20650 -9320 20670
rect -9360 20510 -9320 20650
rect -9360 20490 -9350 20510
rect -9330 20490 -9320 20510
rect -9360 20480 -9320 20490
rect -9280 20670 -9240 20680
rect -9280 20650 -9270 20670
rect -9250 20650 -9240 20670
rect -9280 20510 -9240 20650
rect -9280 20490 -9270 20510
rect -9250 20490 -9240 20510
rect -9280 20480 -9240 20490
rect -9200 20670 -9160 20680
rect -9200 20650 -9190 20670
rect -9170 20650 -9160 20670
rect -9200 20510 -9160 20650
rect -9200 20490 -9190 20510
rect -9170 20490 -9160 20510
rect -9200 20480 -9160 20490
rect -9120 20670 -9080 20680
rect -9120 20650 -9110 20670
rect -9090 20650 -9080 20670
rect -9120 20510 -9080 20650
rect -9120 20490 -9110 20510
rect -9090 20490 -9080 20510
rect -9120 20480 -9080 20490
rect -9040 20670 -9000 20680
rect -9040 20650 -9030 20670
rect -9010 20650 -9000 20670
rect -9040 20510 -9000 20650
rect -9040 20490 -9030 20510
rect -9010 20490 -9000 20510
rect -9040 20480 -9000 20490
rect -8960 20670 -8920 20680
rect -8960 20650 -8950 20670
rect -8930 20650 -8920 20670
rect -8960 20510 -8920 20650
rect -8960 20490 -8950 20510
rect -8930 20490 -8920 20510
rect -8960 20480 -8920 20490
rect -8880 20670 -8840 20680
rect -8880 20650 -8870 20670
rect -8850 20650 -8840 20670
rect -8880 20510 -8840 20650
rect -8880 20490 -8870 20510
rect -8850 20490 -8840 20510
rect -8880 20480 -8840 20490
rect -8800 20670 -8760 20680
rect -8800 20650 -8790 20670
rect -8770 20650 -8760 20670
rect -8800 20510 -8760 20650
rect -8800 20490 -8790 20510
rect -8770 20490 -8760 20510
rect -8800 20480 -8760 20490
rect -8720 20670 -8680 20680
rect -8720 20650 -8710 20670
rect -8690 20650 -8680 20670
rect -8720 20510 -8680 20650
rect -8720 20490 -8710 20510
rect -8690 20490 -8680 20510
rect -8720 20480 -8680 20490
rect -8640 20670 -8600 20680
rect -8640 20650 -8630 20670
rect -8610 20650 -8600 20670
rect -8640 20510 -8600 20650
rect -8640 20490 -8630 20510
rect -8610 20490 -8600 20510
rect -8640 20480 -8600 20490
rect -8560 20670 -8520 20680
rect -8560 20650 -8550 20670
rect -8530 20650 -8520 20670
rect -8560 20510 -8520 20650
rect -8560 20490 -8550 20510
rect -8530 20490 -8520 20510
rect -8560 20480 -8520 20490
rect -8480 20670 -8440 20680
rect -8480 20650 -8470 20670
rect -8450 20650 -8440 20670
rect -8480 20510 -8440 20650
rect -8480 20490 -8470 20510
rect -8450 20490 -8440 20510
rect -8480 20480 -8440 20490
rect -8400 20670 -8360 20680
rect -8400 20650 -8390 20670
rect -8370 20650 -8360 20670
rect -8400 20510 -8360 20650
rect -8400 20490 -8390 20510
rect -8370 20490 -8360 20510
rect -8400 20480 -8360 20490
rect -8320 20670 -8280 20680
rect -8320 20650 -8310 20670
rect -8290 20650 -8280 20670
rect -8320 20510 -8280 20650
rect -8320 20490 -8310 20510
rect -8290 20490 -8280 20510
rect -8320 20480 -8280 20490
rect -8240 20670 -8200 20680
rect -8240 20650 -8230 20670
rect -8210 20650 -8200 20670
rect -8240 20510 -8200 20650
rect -8240 20490 -8230 20510
rect -8210 20490 -8200 20510
rect -8240 20480 -8200 20490
rect -8160 20670 -8120 20680
rect -8160 20650 -8150 20670
rect -8130 20650 -8120 20670
rect -8160 20510 -8120 20650
rect -8160 20490 -8150 20510
rect -8130 20490 -8120 20510
rect -8160 20480 -8120 20490
rect -8080 20670 -8040 20680
rect -8080 20650 -8070 20670
rect -8050 20650 -8040 20670
rect -8080 20510 -8040 20650
rect -8080 20490 -8070 20510
rect -8050 20490 -8040 20510
rect -8080 20480 -8040 20490
rect -8000 20670 -7960 20680
rect -8000 20650 -7990 20670
rect -7970 20650 -7960 20670
rect -8000 20510 -7960 20650
rect -8000 20490 -7990 20510
rect -7970 20490 -7960 20510
rect -8000 20480 -7960 20490
rect -7920 20670 -7880 20680
rect -7920 20650 -7910 20670
rect -7890 20650 -7880 20670
rect -7920 20510 -7880 20650
rect -7920 20490 -7910 20510
rect -7890 20490 -7880 20510
rect -7920 20480 -7880 20490
rect -7840 20670 -7800 20680
rect -7840 20650 -7830 20670
rect -7810 20650 -7800 20670
rect -7840 20510 -7800 20650
rect -7840 20490 -7830 20510
rect -7810 20490 -7800 20510
rect -7840 20480 -7800 20490
rect -7760 20670 -7720 20680
rect -7760 20650 -7750 20670
rect -7730 20650 -7720 20670
rect -7760 20510 -7720 20650
rect -7760 20490 -7750 20510
rect -7730 20490 -7720 20510
rect -7760 20480 -7720 20490
rect -7680 20670 -7640 20680
rect -7680 20650 -7670 20670
rect -7650 20650 -7640 20670
rect -7680 20510 -7640 20650
rect -7680 20490 -7670 20510
rect -7650 20490 -7640 20510
rect -7680 20480 -7640 20490
rect -7600 20670 -7560 20680
rect -7600 20650 -7590 20670
rect -7570 20650 -7560 20670
rect -7600 20510 -7560 20650
rect -7600 20490 -7590 20510
rect -7570 20490 -7560 20510
rect -7600 20480 -7560 20490
rect -7520 20670 -7480 20680
rect -7520 20650 -7510 20670
rect -7490 20650 -7480 20670
rect -7520 20510 -7480 20650
rect -7520 20490 -7510 20510
rect -7490 20490 -7480 20510
rect -7520 20480 -7480 20490
rect -7440 20670 -7400 20680
rect -7440 20650 -7430 20670
rect -7410 20650 -7400 20670
rect -7440 20510 -7400 20650
rect -7440 20490 -7430 20510
rect -7410 20490 -7400 20510
rect -7440 20480 -7400 20490
rect -7360 20670 -7320 20680
rect -7360 20650 -7350 20670
rect -7330 20650 -7320 20670
rect -7360 20510 -7320 20650
rect -7360 20490 -7350 20510
rect -7330 20490 -7320 20510
rect -7360 20480 -7320 20490
rect -7280 20670 -7240 20680
rect -7280 20650 -7270 20670
rect -7250 20650 -7240 20670
rect -7280 20510 -7240 20650
rect -7280 20490 -7270 20510
rect -7250 20490 -7240 20510
rect -7280 20480 -7240 20490
rect -7200 20670 -7160 20680
rect -7200 20650 -7190 20670
rect -7170 20650 -7160 20670
rect -7200 20510 -7160 20650
rect -7200 20490 -7190 20510
rect -7170 20490 -7160 20510
rect -7200 20480 -7160 20490
rect -7120 20670 -7080 20680
rect -7120 20650 -7110 20670
rect -7090 20650 -7080 20670
rect -7120 20510 -7080 20650
rect -7120 20490 -7110 20510
rect -7090 20490 -7080 20510
rect -7120 20480 -7080 20490
rect -7040 20670 -7000 20680
rect -7040 20650 -7030 20670
rect -7010 20650 -7000 20670
rect -7040 20510 -7000 20650
rect -7040 20490 -7030 20510
rect -7010 20490 -7000 20510
rect -7040 20480 -7000 20490
rect -6960 20670 -6920 20680
rect -6960 20650 -6950 20670
rect -6930 20650 -6920 20670
rect -6960 20510 -6920 20650
rect -6960 20490 -6950 20510
rect -6930 20490 -6920 20510
rect -6960 20480 -6920 20490
rect -6880 20670 -6840 20680
rect -6880 20650 -6870 20670
rect -6850 20650 -6840 20670
rect -6880 20510 -6840 20650
rect -6880 20490 -6870 20510
rect -6850 20490 -6840 20510
rect -6880 20480 -6840 20490
rect -6800 20670 -6760 20680
rect -6800 20650 -6790 20670
rect -6770 20650 -6760 20670
rect -6800 20510 -6760 20650
rect -6800 20490 -6790 20510
rect -6770 20490 -6760 20510
rect -6800 20480 -6760 20490
rect -6720 20670 -6680 20680
rect -6720 20650 -6710 20670
rect -6690 20650 -6680 20670
rect -6720 20510 -6680 20650
rect -6720 20490 -6710 20510
rect -6690 20490 -6680 20510
rect -6720 20480 -6680 20490
rect -6640 20670 -6600 20680
rect -6640 20650 -6630 20670
rect -6610 20650 -6600 20670
rect -6640 20510 -6600 20650
rect -6640 20490 -6630 20510
rect -6610 20490 -6600 20510
rect -6640 20480 -6600 20490
rect -6560 20670 -6520 20680
rect -6560 20650 -6550 20670
rect -6530 20650 -6520 20670
rect -6560 20510 -6520 20650
rect -6560 20490 -6550 20510
rect -6530 20490 -6520 20510
rect -6560 20480 -6520 20490
rect -6480 20670 -6440 20680
rect -6480 20650 -6470 20670
rect -6450 20650 -6440 20670
rect -6480 20510 -6440 20650
rect -6480 20490 -6470 20510
rect -6450 20490 -6440 20510
rect -6480 20480 -6440 20490
rect -6400 20670 -6360 20680
rect -6400 20650 -6390 20670
rect -6370 20650 -6360 20670
rect -6400 20510 -6360 20650
rect -6400 20490 -6390 20510
rect -6370 20490 -6360 20510
rect -6400 20480 -6360 20490
rect -6320 20670 -6280 20680
rect -6320 20650 -6310 20670
rect -6290 20650 -6280 20670
rect -6320 20510 -6280 20650
rect -6320 20490 -6310 20510
rect -6290 20490 -6280 20510
rect -6320 20480 -6280 20490
rect -6240 20670 -6200 20680
rect -6240 20650 -6230 20670
rect -6210 20650 -6200 20670
rect -6240 20510 -6200 20650
rect -6240 20490 -6230 20510
rect -6210 20490 -6200 20510
rect -6240 20480 -6200 20490
rect -6160 20670 -6120 20680
rect -6160 20650 -6150 20670
rect -6130 20650 -6120 20670
rect -6160 20510 -6120 20650
rect -6160 20490 -6150 20510
rect -6130 20490 -6120 20510
rect -6160 20480 -6120 20490
rect -5680 20670 -5640 20680
rect -5680 20650 -5670 20670
rect -5650 20650 -5640 20670
rect -5680 20510 -5640 20650
rect -5680 20490 -5670 20510
rect -5650 20490 -5640 20510
rect -5680 20480 -5640 20490
rect -5600 20670 -5560 20680
rect -5600 20650 -5590 20670
rect -5570 20650 -5560 20670
rect -5600 20510 -5560 20650
rect -5600 20490 -5590 20510
rect -5570 20490 -5560 20510
rect -5600 20480 -5560 20490
rect -5520 20670 -5480 20680
rect -5520 20650 -5510 20670
rect -5490 20650 -5480 20670
rect -5520 20510 -5480 20650
rect -5520 20490 -5510 20510
rect -5490 20490 -5480 20510
rect -5520 20480 -5480 20490
rect -5440 20670 -5400 20680
rect -5440 20650 -5430 20670
rect -5410 20650 -5400 20670
rect -5440 20510 -5400 20650
rect -5440 20490 -5430 20510
rect -5410 20490 -5400 20510
rect -5440 20480 -5400 20490
rect -5360 20670 -5320 20680
rect -5360 20650 -5350 20670
rect -5330 20650 -5320 20670
rect -5360 20510 -5320 20650
rect -5360 20490 -5350 20510
rect -5330 20490 -5320 20510
rect -5360 20480 -5320 20490
rect -5280 20670 -5240 20680
rect -5280 20650 -5270 20670
rect -5250 20650 -5240 20670
rect -5280 20510 -5240 20650
rect -5280 20490 -5270 20510
rect -5250 20490 -5240 20510
rect -5280 20480 -5240 20490
rect -5200 20670 -5160 20680
rect -5200 20650 -5190 20670
rect -5170 20650 -5160 20670
rect -5200 20510 -5160 20650
rect -5200 20490 -5190 20510
rect -5170 20490 -5160 20510
rect -5200 20480 -5160 20490
rect -5120 20670 -5080 20680
rect -5120 20650 -5110 20670
rect -5090 20650 -5080 20670
rect -5120 20510 -5080 20650
rect -5120 20490 -5110 20510
rect -5090 20490 -5080 20510
rect -5120 20480 -5080 20490
rect -5040 20670 -5000 20680
rect -5040 20650 -5030 20670
rect -5010 20650 -5000 20670
rect -5040 20510 -5000 20650
rect -5040 20490 -5030 20510
rect -5010 20490 -5000 20510
rect -5040 20480 -5000 20490
rect -4960 20670 -4920 20680
rect -4960 20650 -4950 20670
rect -4930 20650 -4920 20670
rect -4960 20510 -4920 20650
rect -4960 20490 -4950 20510
rect -4930 20490 -4920 20510
rect -4960 20480 -4920 20490
rect -4880 20670 -4840 20680
rect -4880 20650 -4870 20670
rect -4850 20650 -4840 20670
rect -4880 20510 -4840 20650
rect -4880 20490 -4870 20510
rect -4850 20490 -4840 20510
rect -4880 20480 -4840 20490
rect -4800 20670 -4760 20680
rect -4800 20650 -4790 20670
rect -4770 20650 -4760 20670
rect -4800 20510 -4760 20650
rect -4800 20490 -4790 20510
rect -4770 20490 -4760 20510
rect -4800 20480 -4760 20490
rect -4720 20670 -4680 20680
rect -4720 20650 -4710 20670
rect -4690 20650 -4680 20670
rect -4720 20510 -4680 20650
rect -4720 20490 -4710 20510
rect -4690 20490 -4680 20510
rect -4720 20480 -4680 20490
rect -4640 20670 -4600 20680
rect -4640 20650 -4630 20670
rect -4610 20650 -4600 20670
rect -4640 20510 -4600 20650
rect -4640 20490 -4630 20510
rect -4610 20490 -4600 20510
rect -4640 20480 -4600 20490
rect -4560 20670 -4520 20680
rect -4560 20650 -4550 20670
rect -4530 20650 -4520 20670
rect -4560 20510 -4520 20650
rect -4560 20490 -4550 20510
rect -4530 20490 -4520 20510
rect -4560 20480 -4520 20490
rect -4480 20670 -4440 20680
rect -4480 20650 -4470 20670
rect -4450 20650 -4440 20670
rect -4480 20510 -4440 20650
rect -4480 20490 -4470 20510
rect -4450 20490 -4440 20510
rect -4480 20480 -4440 20490
rect -4400 20670 -4360 20680
rect -4400 20650 -4390 20670
rect -4370 20650 -4360 20670
rect -4400 20510 -4360 20650
rect -4400 20490 -4390 20510
rect -4370 20490 -4360 20510
rect -4400 20480 -4360 20490
rect -4320 20670 -4280 20680
rect -4320 20650 -4310 20670
rect -4290 20650 -4280 20670
rect -4320 20510 -4280 20650
rect -4320 20490 -4310 20510
rect -4290 20490 -4280 20510
rect -4320 20480 -4280 20490
rect -4240 20670 -4200 20680
rect -4240 20650 -4230 20670
rect -4210 20650 -4200 20670
rect -4240 20510 -4200 20650
rect -4240 20490 -4230 20510
rect -4210 20490 -4200 20510
rect -4240 20480 -4200 20490
rect -4160 20670 -4120 20680
rect -4160 20650 -4150 20670
rect -4130 20650 -4120 20670
rect -4160 20510 -4120 20650
rect -4160 20490 -4150 20510
rect -4130 20490 -4120 20510
rect -4160 20480 -4120 20490
rect -4080 20670 -4040 20680
rect -4080 20650 -4070 20670
rect -4050 20650 -4040 20670
rect -4080 20510 -4040 20650
rect -4080 20490 -4070 20510
rect -4050 20490 -4040 20510
rect -4080 20480 -4040 20490
rect -4000 20670 -3960 20680
rect -4000 20650 -3990 20670
rect -3970 20650 -3960 20670
rect -4000 20510 -3960 20650
rect -4000 20490 -3990 20510
rect -3970 20490 -3960 20510
rect -4000 20480 -3960 20490
rect -3920 20670 -3880 20680
rect -3920 20650 -3910 20670
rect -3890 20650 -3880 20670
rect -3920 20510 -3880 20650
rect -3920 20490 -3910 20510
rect -3890 20490 -3880 20510
rect -3920 20480 -3880 20490
rect -3840 20670 -3800 20680
rect -3840 20650 -3830 20670
rect -3810 20650 -3800 20670
rect -3840 20510 -3800 20650
rect -3840 20490 -3830 20510
rect -3810 20490 -3800 20510
rect -3840 20480 -3800 20490
rect -3760 20670 -3720 20680
rect -3760 20650 -3750 20670
rect -3730 20650 -3720 20670
rect -3760 20510 -3720 20650
rect -3760 20490 -3750 20510
rect -3730 20490 -3720 20510
rect -3760 20480 -3720 20490
rect -3680 20670 -3640 20680
rect -3680 20650 -3670 20670
rect -3650 20650 -3640 20670
rect -3680 20510 -3640 20650
rect -3680 20490 -3670 20510
rect -3650 20490 -3640 20510
rect -3680 20480 -3640 20490
rect -3600 20670 -3560 20680
rect -3600 20650 -3590 20670
rect -3570 20650 -3560 20670
rect -3600 20510 -3560 20650
rect -3600 20490 -3590 20510
rect -3570 20490 -3560 20510
rect -3600 20480 -3560 20490
rect -3520 20670 -3480 20680
rect -3520 20650 -3510 20670
rect -3490 20650 -3480 20670
rect -3520 20510 -3480 20650
rect -3520 20490 -3510 20510
rect -3490 20490 -3480 20510
rect -3520 20480 -3480 20490
rect -3440 20670 -3400 20680
rect -3440 20650 -3430 20670
rect -3410 20650 -3400 20670
rect -3440 20510 -3400 20650
rect -3440 20490 -3430 20510
rect -3410 20490 -3400 20510
rect -3440 20480 -3400 20490
rect -3360 20670 -3320 20680
rect -3360 20650 -3350 20670
rect -3330 20650 -3320 20670
rect -3360 20510 -3320 20650
rect -3360 20490 -3350 20510
rect -3330 20490 -3320 20510
rect -3360 20480 -3320 20490
rect -3280 20670 -3240 20680
rect -3280 20650 -3270 20670
rect -3250 20650 -3240 20670
rect -3280 20510 -3240 20650
rect -3280 20490 -3270 20510
rect -3250 20490 -3240 20510
rect -3280 20480 -3240 20490
rect -3200 20670 -3160 20680
rect -3200 20650 -3190 20670
rect -3170 20650 -3160 20670
rect -3200 20510 -3160 20650
rect -3200 20490 -3190 20510
rect -3170 20490 -3160 20510
rect -3200 20480 -3160 20490
rect -3120 20670 -3080 20680
rect -3120 20650 -3110 20670
rect -3090 20650 -3080 20670
rect -3120 20510 -3080 20650
rect -3120 20490 -3110 20510
rect -3090 20490 -3080 20510
rect -3120 20480 -3080 20490
rect -3040 20670 -3000 20680
rect -3040 20650 -3030 20670
rect -3010 20650 -3000 20670
rect -3040 20510 -3000 20650
rect -3040 20490 -3030 20510
rect -3010 20490 -3000 20510
rect -3040 20480 -3000 20490
rect -2960 20670 -2920 20680
rect -2960 20650 -2950 20670
rect -2930 20650 -2920 20670
rect -2960 20510 -2920 20650
rect -2960 20490 -2950 20510
rect -2930 20490 -2920 20510
rect -2960 20480 -2920 20490
rect -2880 20670 -2840 20680
rect -2880 20650 -2870 20670
rect -2850 20650 -2840 20670
rect -2880 20510 -2840 20650
rect -2880 20490 -2870 20510
rect -2850 20490 -2840 20510
rect -2880 20480 -2840 20490
rect -2800 20670 -2760 20680
rect -2800 20650 -2790 20670
rect -2770 20650 -2760 20670
rect -2800 20510 -2760 20650
rect -2800 20490 -2790 20510
rect -2770 20490 -2760 20510
rect -2800 20480 -2760 20490
rect -2720 20670 -2680 20680
rect -2720 20650 -2710 20670
rect -2690 20650 -2680 20670
rect -2720 20510 -2680 20650
rect -2720 20490 -2710 20510
rect -2690 20490 -2680 20510
rect -2720 20480 -2680 20490
rect -2640 20670 -2600 20680
rect -2640 20650 -2630 20670
rect -2610 20650 -2600 20670
rect -2640 20510 -2600 20650
rect -2640 20490 -2630 20510
rect -2610 20490 -2600 20510
rect -2640 20480 -2600 20490
rect -2560 20670 -2520 20680
rect -2560 20650 -2550 20670
rect -2530 20650 -2520 20670
rect -2560 20510 -2520 20650
rect -2560 20490 -2550 20510
rect -2530 20490 -2520 20510
rect -2560 20480 -2520 20490
rect -2480 20670 -2440 20680
rect -2480 20650 -2470 20670
rect -2450 20650 -2440 20670
rect -2480 20510 -2440 20650
rect -2480 20490 -2470 20510
rect -2450 20490 -2440 20510
rect -2480 20480 -2440 20490
rect -2400 20670 -2360 20680
rect -2400 20650 -2390 20670
rect -2370 20650 -2360 20670
rect -2400 20510 -2360 20650
rect -2400 20490 -2390 20510
rect -2370 20490 -2360 20510
rect -2400 20480 -2360 20490
rect -2320 20670 -2280 20680
rect -2320 20650 -2310 20670
rect -2290 20650 -2280 20670
rect -2320 20510 -2280 20650
rect -2320 20490 -2310 20510
rect -2290 20490 -2280 20510
rect -2320 20480 -2280 20490
rect -2240 20670 -2200 20680
rect -2240 20650 -2230 20670
rect -2210 20650 -2200 20670
rect -2240 20510 -2200 20650
rect -2240 20490 -2230 20510
rect -2210 20490 -2200 20510
rect -2240 20480 -2200 20490
rect -2160 20670 -2120 20680
rect -2160 20650 -2150 20670
rect -2130 20650 -2120 20670
rect -2160 20510 -2120 20650
rect -2160 20490 -2150 20510
rect -2130 20490 -2120 20510
rect -2160 20480 -2120 20490
rect -2080 20670 -2040 20680
rect -2080 20650 -2070 20670
rect -2050 20650 -2040 20670
rect -2080 20510 -2040 20650
rect -2080 20490 -2070 20510
rect -2050 20490 -2040 20510
rect -2080 20480 -2040 20490
rect -2000 20670 -1960 20680
rect -2000 20650 -1990 20670
rect -1970 20650 -1960 20670
rect -2000 20510 -1960 20650
rect -2000 20490 -1990 20510
rect -1970 20490 -1960 20510
rect -2000 20480 -1960 20490
rect -1920 20670 -1880 21480
rect -1840 21430 -1800 21440
rect -1840 21410 -1830 21430
rect -1810 21410 -1800 21430
rect -1840 21270 -1800 21410
rect -1840 21250 -1830 21270
rect -1810 21250 -1800 21270
rect -1840 21110 -1800 21250
rect -1840 21090 -1830 21110
rect -1810 21090 -1800 21110
rect -1840 20950 -1800 21090
rect -1840 20930 -1830 20950
rect -1810 20930 -1800 20950
rect -1840 20920 -1800 20930
rect -1760 21430 -1720 21440
rect -1760 21410 -1750 21430
rect -1730 21410 -1720 21430
rect -1760 21270 -1720 21410
rect -1760 21250 -1750 21270
rect -1730 21250 -1720 21270
rect -1760 21110 -1720 21250
rect -1760 21090 -1750 21110
rect -1730 21090 -1720 21110
rect -1760 20950 -1720 21090
rect -1760 20930 -1750 20950
rect -1730 20930 -1720 20950
rect -1760 20920 -1720 20930
rect -1680 21430 -1640 21440
rect -1680 21410 -1670 21430
rect -1650 21410 -1640 21430
rect -1680 21270 -1640 21410
rect -1680 21250 -1670 21270
rect -1650 21250 -1640 21270
rect -1680 21110 -1640 21250
rect -1680 21090 -1670 21110
rect -1650 21090 -1640 21110
rect -1680 20950 -1640 21090
rect -1680 20930 -1670 20950
rect -1650 20930 -1640 20950
rect -1680 20920 -1640 20930
rect -1520 21430 -1480 21440
rect -1520 21410 -1510 21430
rect -1490 21410 -1480 21430
rect -1520 21270 -1480 21410
rect -1520 21250 -1510 21270
rect -1490 21250 -1480 21270
rect -1520 21110 -1480 21250
rect -1520 21090 -1510 21110
rect -1490 21090 -1480 21110
rect -1520 20950 -1480 21090
rect -1520 20930 -1510 20950
rect -1490 20930 -1480 20950
rect -1520 20920 -1480 20930
rect -1360 21430 -1320 21440
rect -1360 21410 -1350 21430
rect -1330 21410 -1320 21430
rect -1360 21270 -1320 21410
rect -1360 21250 -1350 21270
rect -1330 21250 -1320 21270
rect -1360 21110 -1320 21250
rect -1360 21090 -1350 21110
rect -1330 21090 -1320 21110
rect -1360 20950 -1320 21090
rect -1360 20930 -1350 20950
rect -1330 20930 -1320 20950
rect -1360 20920 -1320 20930
rect -1280 21430 -1240 21440
rect -1280 21410 -1270 21430
rect -1250 21410 -1240 21430
rect -1280 21270 -1240 21410
rect -1280 21250 -1270 21270
rect -1250 21250 -1240 21270
rect -1280 21110 -1240 21250
rect -1280 21090 -1270 21110
rect -1250 21090 -1240 21110
rect -1280 20950 -1240 21090
rect -1280 20930 -1270 20950
rect -1250 20930 -1240 20950
rect -1280 20920 -1240 20930
rect -1200 21430 -1160 21440
rect -1200 21410 -1190 21430
rect -1170 21410 -1160 21430
rect -1200 21270 -1160 21410
rect -1200 21250 -1190 21270
rect -1170 21250 -1160 21270
rect -1200 21110 -1160 21250
rect -1200 21090 -1190 21110
rect -1170 21090 -1160 21110
rect -1200 20950 -1160 21090
rect -1200 20930 -1190 20950
rect -1170 20930 -1160 20950
rect -1200 20920 -1160 20930
rect -1120 21430 -1080 21440
rect -1120 21410 -1110 21430
rect -1090 21410 -1080 21430
rect -1120 21270 -1080 21410
rect -1120 21250 -1110 21270
rect -1090 21250 -1080 21270
rect -1120 21110 -1080 21250
rect -1120 21090 -1110 21110
rect -1090 21090 -1080 21110
rect -1120 20950 -1080 21090
rect -1120 20930 -1110 20950
rect -1090 20930 -1080 20950
rect -1120 20920 -1080 20930
rect -1040 21430 -1000 21440
rect -1040 21410 -1030 21430
rect -1010 21410 -1000 21430
rect -1040 21270 -1000 21410
rect -1040 21250 -1030 21270
rect -1010 21250 -1000 21270
rect -1040 21110 -1000 21250
rect -1040 21090 -1030 21110
rect -1010 21090 -1000 21110
rect -1040 20950 -1000 21090
rect -1040 20930 -1030 20950
rect -1010 20930 -1000 20950
rect -1040 20920 -1000 20930
rect -880 21430 -840 21440
rect -880 21410 -870 21430
rect -850 21410 -840 21430
rect -880 21270 -840 21410
rect -880 21250 -870 21270
rect -850 21250 -840 21270
rect -880 21110 -840 21250
rect -880 21090 -870 21110
rect -850 21090 -840 21110
rect -880 20950 -840 21090
rect -880 20930 -870 20950
rect -850 20930 -840 20950
rect -880 20920 -840 20930
rect -720 21430 -680 21440
rect -720 21410 -710 21430
rect -690 21410 -680 21430
rect -720 21270 -680 21410
rect -720 21250 -710 21270
rect -690 21250 -680 21270
rect -720 21110 -680 21250
rect -720 21090 -710 21110
rect -690 21090 -680 21110
rect -720 20950 -680 21090
rect -720 20930 -710 20950
rect -690 20930 -680 20950
rect -720 20920 -680 20930
rect -560 21430 -520 21440
rect -560 21410 -550 21430
rect -530 21410 -520 21430
rect -560 21270 -520 21410
rect -560 21250 -550 21270
rect -530 21250 -520 21270
rect -560 21110 -520 21250
rect -560 21090 -550 21110
rect -530 21090 -520 21110
rect -560 20950 -520 21090
rect -560 20930 -550 20950
rect -530 20930 -520 20950
rect -560 20920 -520 20930
rect -1920 20650 -1910 20670
rect -1890 20650 -1880 20670
rect -1920 20510 -1880 20650
rect -1920 20490 -1910 20510
rect -1890 20490 -1880 20510
rect -5280 20350 -5240 20360
rect -5280 20330 -5270 20350
rect -5250 20330 -5240 20350
rect -5280 20190 -5240 20330
rect -5280 20170 -5270 20190
rect -5250 20170 -5240 20190
rect -5280 20160 -5240 20170
rect -5120 20350 -5080 20360
rect -5120 20330 -5110 20350
rect -5090 20330 -5080 20350
rect -5120 20190 -5080 20330
rect -5120 20170 -5110 20190
rect -5090 20170 -5080 20190
rect -5120 20160 -5080 20170
rect -5040 20350 -5000 20360
rect -5040 20330 -5030 20350
rect -5010 20330 -5000 20350
rect -5040 20190 -5000 20330
rect -5040 20170 -5030 20190
rect -5010 20170 -5000 20190
rect -5040 20160 -5000 20170
rect -4960 20350 -4920 20360
rect -4960 20330 -4950 20350
rect -4930 20330 -4920 20350
rect -4960 20190 -4920 20330
rect -4960 20170 -4950 20190
rect -4930 20170 -4920 20190
rect -4960 20160 -4920 20170
rect -4880 20350 -4840 20360
rect -4880 20330 -4870 20350
rect -4850 20330 -4840 20350
rect -4880 20190 -4840 20330
rect -4880 20170 -4870 20190
rect -4850 20170 -4840 20190
rect -4880 20160 -4840 20170
rect -4800 20350 -4760 20360
rect -4800 20330 -4790 20350
rect -4770 20330 -4760 20350
rect -4800 20190 -4760 20330
rect -4800 20170 -4790 20190
rect -4770 20170 -4760 20190
rect -4800 20160 -4760 20170
rect -4720 20350 -4680 20360
rect -4720 20330 -4710 20350
rect -4690 20330 -4680 20350
rect -4720 20190 -4680 20330
rect -4720 20170 -4710 20190
rect -4690 20170 -4680 20190
rect -4720 20160 -4680 20170
rect -4640 20350 -4600 20360
rect -4640 20330 -4630 20350
rect -4610 20330 -4600 20350
rect -4640 20190 -4600 20330
rect -4640 20170 -4630 20190
rect -4610 20170 -4600 20190
rect -4640 20160 -4600 20170
rect -4560 20350 -4520 20360
rect -4560 20330 -4550 20350
rect -4530 20330 -4520 20350
rect -4560 20190 -4520 20330
rect -4560 20170 -4550 20190
rect -4530 20170 -4520 20190
rect -4560 20160 -4520 20170
rect -4480 20350 -4440 20360
rect -4480 20330 -4470 20350
rect -4450 20330 -4440 20350
rect -4480 20190 -4440 20330
rect -4480 20170 -4470 20190
rect -4450 20170 -4440 20190
rect -4480 20160 -4440 20170
rect -4400 20350 -4360 20360
rect -4400 20330 -4390 20350
rect -4370 20330 -4360 20350
rect -4400 20190 -4360 20330
rect -4400 20170 -4390 20190
rect -4370 20170 -4360 20190
rect -4400 20160 -4360 20170
rect -4320 20350 -4280 20360
rect -4320 20330 -4310 20350
rect -4290 20330 -4280 20350
rect -4320 20190 -4280 20330
rect -4320 20170 -4310 20190
rect -4290 20170 -4280 20190
rect -4320 20160 -4280 20170
rect -4240 20350 -4200 20360
rect -4240 20330 -4230 20350
rect -4210 20330 -4200 20350
rect -4240 20190 -4200 20330
rect -4240 20170 -4230 20190
rect -4210 20170 -4200 20190
rect -4240 20160 -4200 20170
rect -4160 20350 -4120 20360
rect -4160 20330 -4150 20350
rect -4130 20330 -4120 20350
rect -4160 20190 -4120 20330
rect -4160 20170 -4150 20190
rect -4130 20170 -4120 20190
rect -4160 20160 -4120 20170
rect -4080 20350 -4040 20360
rect -4080 20330 -4070 20350
rect -4050 20330 -4040 20350
rect -4080 20190 -4040 20330
rect -4080 20170 -4070 20190
rect -4050 20170 -4040 20190
rect -4080 20160 -4040 20170
rect -4000 20350 -3960 20360
rect -4000 20330 -3990 20350
rect -3970 20330 -3960 20350
rect -4000 20190 -3960 20330
rect -4000 20170 -3990 20190
rect -3970 20170 -3960 20190
rect -4000 20160 -3960 20170
rect -3920 20350 -3880 20360
rect -3920 20330 -3910 20350
rect -3890 20330 -3880 20350
rect -3920 20190 -3880 20330
rect -3920 20170 -3910 20190
rect -3890 20170 -3880 20190
rect -3920 20160 -3880 20170
rect -3840 20350 -3800 20360
rect -3840 20330 -3830 20350
rect -3810 20330 -3800 20350
rect -3840 20190 -3800 20330
rect -3840 20170 -3830 20190
rect -3810 20170 -3800 20190
rect -3840 20160 -3800 20170
rect -3760 20350 -3720 20360
rect -3760 20330 -3750 20350
rect -3730 20330 -3720 20350
rect -3760 20190 -3720 20330
rect -3760 20170 -3750 20190
rect -3730 20170 -3720 20190
rect -3760 20160 -3720 20170
rect -3680 20350 -3640 20360
rect -3680 20330 -3670 20350
rect -3650 20330 -3640 20350
rect -3680 20190 -3640 20330
rect -3680 20170 -3670 20190
rect -3650 20170 -3640 20190
rect -3680 20160 -3640 20170
rect -3600 20350 -3560 20360
rect -3600 20330 -3590 20350
rect -3570 20330 -3560 20350
rect -3600 20190 -3560 20330
rect -3600 20170 -3590 20190
rect -3570 20170 -3560 20190
rect -3600 20160 -3560 20170
rect -3520 20350 -3480 20360
rect -3520 20330 -3510 20350
rect -3490 20330 -3480 20350
rect -3520 20190 -3480 20330
rect -3520 20170 -3510 20190
rect -3490 20170 -3480 20190
rect -3520 20160 -3480 20170
rect -3440 20350 -3400 20360
rect -3440 20330 -3430 20350
rect -3410 20330 -3400 20350
rect -3440 20190 -3400 20330
rect -3440 20170 -3430 20190
rect -3410 20170 -3400 20190
rect -3440 20160 -3400 20170
rect -3360 20350 -3320 20360
rect -3360 20330 -3350 20350
rect -3330 20330 -3320 20350
rect -3360 20190 -3320 20330
rect -3360 20170 -3350 20190
rect -3330 20170 -3320 20190
rect -3360 20160 -3320 20170
rect -3280 20350 -3240 20360
rect -3280 20330 -3270 20350
rect -3250 20330 -3240 20350
rect -3280 20190 -3240 20330
rect -3280 20170 -3270 20190
rect -3250 20170 -3240 20190
rect -3280 20160 -3240 20170
rect -3200 20350 -3160 20360
rect -3200 20330 -3190 20350
rect -3170 20330 -3160 20350
rect -3200 20190 -3160 20330
rect -3200 20170 -3190 20190
rect -3170 20170 -3160 20190
rect -3200 20160 -3160 20170
rect -3120 20350 -3080 20360
rect -3120 20330 -3110 20350
rect -3090 20330 -3080 20350
rect -3120 20190 -3080 20330
rect -3120 20170 -3110 20190
rect -3090 20170 -3080 20190
rect -3120 20160 -3080 20170
rect -3040 20350 -3000 20360
rect -3040 20330 -3030 20350
rect -3010 20330 -3000 20350
rect -3040 20190 -3000 20330
rect -3040 20170 -3030 20190
rect -3010 20170 -3000 20190
rect -3040 20160 -3000 20170
rect -2960 20350 -2920 20360
rect -2960 20330 -2950 20350
rect -2930 20330 -2920 20350
rect -2960 20190 -2920 20330
rect -2960 20170 -2950 20190
rect -2930 20170 -2920 20190
rect -2960 20160 -2920 20170
rect -2880 20350 -2840 20360
rect -2880 20330 -2870 20350
rect -2850 20330 -2840 20350
rect -2880 20190 -2840 20330
rect -2880 20170 -2870 20190
rect -2850 20170 -2840 20190
rect -2880 20160 -2840 20170
rect -2800 20350 -2760 20360
rect -2800 20330 -2790 20350
rect -2770 20330 -2760 20350
rect -2800 20190 -2760 20330
rect -2800 20170 -2790 20190
rect -2770 20170 -2760 20190
rect -2800 20160 -2760 20170
rect -2720 20350 -2680 20360
rect -2720 20330 -2710 20350
rect -2690 20330 -2680 20350
rect -2720 20190 -2680 20330
rect -2720 20170 -2710 20190
rect -2690 20170 -2680 20190
rect -2720 20160 -2680 20170
rect -2640 20350 -2600 20360
rect -2640 20330 -2630 20350
rect -2610 20330 -2600 20350
rect -2640 20190 -2600 20330
rect -2640 20170 -2630 20190
rect -2610 20170 -2600 20190
rect -2640 20160 -2600 20170
rect -2560 20350 -2520 20360
rect -2560 20330 -2550 20350
rect -2530 20330 -2520 20350
rect -2560 20190 -2520 20330
rect -2560 20170 -2550 20190
rect -2530 20170 -2520 20190
rect -2560 20160 -2520 20170
rect -2480 20350 -2440 20360
rect -2480 20330 -2470 20350
rect -2450 20330 -2440 20350
rect -2480 20190 -2440 20330
rect -2480 20170 -2470 20190
rect -2450 20170 -2440 20190
rect -2480 20160 -2440 20170
rect -2400 20350 -2360 20360
rect -2400 20330 -2390 20350
rect -2370 20330 -2360 20350
rect -2400 20190 -2360 20330
rect -2400 20170 -2390 20190
rect -2370 20170 -2360 20190
rect -2400 20160 -2360 20170
rect -2320 20350 -2280 20360
rect -2320 20330 -2310 20350
rect -2290 20330 -2280 20350
rect -2320 20190 -2280 20330
rect -2320 20170 -2310 20190
rect -2290 20170 -2280 20190
rect -2320 20160 -2280 20170
rect -2240 20350 -2200 20360
rect -2240 20330 -2230 20350
rect -2210 20330 -2200 20350
rect -2240 20190 -2200 20330
rect -2240 20170 -2230 20190
rect -2210 20170 -2200 20190
rect -2240 20160 -2200 20170
rect -2160 20350 -2120 20360
rect -2160 20330 -2150 20350
rect -2130 20330 -2120 20350
rect -2160 20190 -2120 20330
rect -2160 20170 -2150 20190
rect -2130 20170 -2120 20190
rect -2160 20160 -2120 20170
rect -2080 20350 -2040 20360
rect -2080 20330 -2070 20350
rect -2050 20330 -2040 20350
rect -2080 20190 -2040 20330
rect -2080 20170 -2070 20190
rect -2050 20170 -2040 20190
rect -2080 20160 -2040 20170
rect -2000 20350 -1960 20360
rect -2000 20330 -1990 20350
rect -1970 20330 -1960 20350
rect -2000 20190 -1960 20330
rect -2000 20170 -1990 20190
rect -1970 20170 -1960 20190
rect -2000 20160 -1960 20170
rect -1920 19960 -1880 20490
rect -1840 20670 -1800 20680
rect -1840 20650 -1830 20670
rect -1810 20650 -1800 20670
rect -1840 20510 -1800 20650
rect -1840 20490 -1830 20510
rect -1810 20490 -1800 20510
rect -1840 20480 -1800 20490
rect -1760 20670 -1720 20680
rect -1760 20650 -1750 20670
rect -1730 20650 -1720 20670
rect -1760 20510 -1720 20650
rect -1760 20490 -1750 20510
rect -1730 20490 -1720 20510
rect -1760 20480 -1720 20490
rect 20520 20670 20560 20680
rect 20520 20650 20530 20670
rect 20550 20650 20560 20670
rect 20520 20510 20560 20650
rect 20520 20490 20530 20510
rect 20550 20490 20560 20510
rect 20520 20480 20560 20490
rect 20600 20670 20640 20680
rect 20600 20650 20610 20670
rect 20630 20650 20640 20670
rect 20600 20510 20640 20650
rect 20600 20490 20610 20510
rect 20630 20490 20640 20510
rect 20600 20480 20640 20490
rect 20680 20670 20720 20680
rect 20680 20650 20690 20670
rect 20710 20650 20720 20670
rect 20680 20510 20720 20650
rect 20680 20490 20690 20510
rect 20710 20490 20720 20510
rect 20680 20480 20720 20490
rect 20760 20670 20800 20680
rect 20760 20650 20770 20670
rect 20790 20650 20800 20670
rect 20760 20510 20800 20650
rect 20760 20490 20770 20510
rect 20790 20490 20800 20510
rect 20760 20480 20800 20490
rect 20840 20670 20880 20680
rect 20840 20650 20850 20670
rect 20870 20650 20880 20670
rect 20840 20510 20880 20650
rect 20840 20490 20850 20510
rect 20870 20490 20880 20510
rect 20840 20480 20880 20490
rect 20920 20670 20960 20680
rect 20920 20650 20930 20670
rect 20950 20650 20960 20670
rect 20920 20510 20960 20650
rect 20920 20490 20930 20510
rect 20950 20490 20960 20510
rect 20920 20480 20960 20490
rect 21000 20670 21040 20680
rect 21000 20650 21010 20670
rect 21030 20650 21040 20670
rect 21000 20510 21040 20650
rect 21000 20490 21010 20510
rect 21030 20490 21040 20510
rect 21000 20480 21040 20490
rect 21080 20670 21120 20680
rect 21080 20650 21090 20670
rect 21110 20650 21120 20670
rect 21080 20510 21120 20650
rect 21080 20490 21090 20510
rect 21110 20490 21120 20510
rect 21080 20480 21120 20490
rect 21160 20670 21200 20680
rect 21160 20650 21170 20670
rect 21190 20650 21200 20670
rect 21160 20510 21200 20650
rect 21160 20490 21170 20510
rect 21190 20490 21200 20510
rect 21160 20480 21200 20490
rect 21240 20670 21280 20680
rect 21240 20650 21250 20670
rect 21270 20650 21280 20670
rect 21240 20510 21280 20650
rect 21240 20490 21250 20510
rect 21270 20490 21280 20510
rect 21240 20480 21280 20490
rect 21320 20670 21360 20680
rect 21320 20650 21330 20670
rect 21350 20650 21360 20670
rect 21320 20510 21360 20650
rect 21320 20490 21330 20510
rect 21350 20490 21360 20510
rect 21320 20480 21360 20490
rect 21400 20670 21440 20680
rect 21400 20650 21410 20670
rect 21430 20650 21440 20670
rect 21400 20510 21440 20650
rect 21400 20490 21410 20510
rect 21430 20490 21440 20510
rect 21400 20480 21440 20490
rect 21480 20670 21520 20680
rect 21480 20650 21490 20670
rect 21510 20650 21520 20670
rect 21480 20510 21520 20650
rect 21480 20490 21490 20510
rect 21510 20490 21520 20510
rect 21480 20480 21520 20490
rect 21560 20670 21600 20680
rect 21560 20650 21570 20670
rect 21590 20650 21600 20670
rect 21560 20510 21600 20650
rect 21560 20490 21570 20510
rect 21590 20490 21600 20510
rect 21560 20480 21600 20490
rect -1840 20350 -1800 20360
rect -1840 20330 -1830 20350
rect -1810 20330 -1800 20350
rect -1840 20190 -1800 20330
rect -1840 20170 -1830 20190
rect -1810 20170 -1800 20190
rect -1840 20160 -1800 20170
rect -1760 20350 -1720 20360
rect -1760 20330 -1750 20350
rect -1730 20330 -1720 20350
rect -1760 20190 -1720 20330
rect -1760 20170 -1750 20190
rect -1730 20170 -1720 20190
rect -1760 20160 -1720 20170
rect 20520 20030 20560 20040
rect 20520 20010 20530 20030
rect 20550 20010 20560 20030
rect 20520 19870 20560 20010
rect 20520 19850 20530 19870
rect 20550 19850 20560 19870
rect 20520 19840 20560 19850
rect 20600 20030 20640 20040
rect 20600 20010 20610 20030
rect 20630 20010 20640 20030
rect 20600 19870 20640 20010
rect 20600 19850 20610 19870
rect 20630 19850 20640 19870
rect 20600 19840 20640 19850
rect 20680 20030 20720 20040
rect 20680 20010 20690 20030
rect 20710 20010 20720 20030
rect 20680 19870 20720 20010
rect 20680 19850 20690 19870
rect 20710 19850 20720 19870
rect 20680 19840 20720 19850
rect 20760 20030 20800 20040
rect 20760 20010 20770 20030
rect 20790 20010 20800 20030
rect 20760 19870 20800 20010
rect 20760 19850 20770 19870
rect 20790 19850 20800 19870
rect 20760 19840 20800 19850
rect 20840 20030 20880 20040
rect 20840 20010 20850 20030
rect 20870 20010 20880 20030
rect 20840 19870 20880 20010
rect 20840 19850 20850 19870
rect 20870 19850 20880 19870
rect 20840 19840 20880 19850
rect 20920 20030 20960 20040
rect 20920 20010 20930 20030
rect 20950 20010 20960 20030
rect 20920 19870 20960 20010
rect 20920 19850 20930 19870
rect 20950 19850 20960 19870
rect 20920 19840 20960 19850
rect 21000 20030 21040 20040
rect 21000 20010 21010 20030
rect 21030 20010 21040 20030
rect 21000 19870 21040 20010
rect 21000 19850 21010 19870
rect 21030 19850 21040 19870
rect 21000 19840 21040 19850
rect 21080 20030 21120 20040
rect 21080 20010 21090 20030
rect 21110 20010 21120 20030
rect 21080 19870 21120 20010
rect 21080 19850 21090 19870
rect 21110 19850 21120 19870
rect 21080 19840 21120 19850
rect 21160 20030 21200 20040
rect 21160 20010 21170 20030
rect 21190 20010 21200 20030
rect 21160 19870 21200 20010
rect 21160 19850 21170 19870
rect 21190 19850 21200 19870
rect 21160 19840 21200 19850
rect 21240 20030 21280 20040
rect 21240 20010 21250 20030
rect 21270 20010 21280 20030
rect 21240 19870 21280 20010
rect 21240 19850 21250 19870
rect 21270 19850 21280 19870
rect 21240 19840 21280 19850
rect 21320 20030 21360 20040
rect 21320 20010 21330 20030
rect 21350 20010 21360 20030
rect 21320 19870 21360 20010
rect 21320 19850 21330 19870
rect 21350 19850 21360 19870
rect 21320 19840 21360 19850
rect 21400 20030 21440 20040
rect 21400 20010 21410 20030
rect 21430 20010 21440 20030
rect 21400 19870 21440 20010
rect 21400 19850 21410 19870
rect 21430 19850 21440 19870
rect 21400 19840 21440 19850
rect 21480 20030 21520 20040
rect 21480 20010 21490 20030
rect 21510 20010 21520 20030
rect 21480 19870 21520 20010
rect 21480 19850 21490 19870
rect 21510 19850 21520 19870
rect 21480 19840 21520 19850
rect 21560 20030 21600 20040
rect 21560 20010 21570 20030
rect 21590 20010 21600 20030
rect 21560 19870 21600 20010
rect 21560 19850 21570 19870
rect 21590 19850 21600 19870
rect 21560 19840 21600 19850
rect -16560 18870 -16520 18880
rect -16560 18850 -16550 18870
rect -16530 18850 -16520 18870
rect -16560 18710 -16520 18850
rect -16560 18690 -16550 18710
rect -16530 18690 -16520 18710
rect -16560 18550 -16520 18690
rect -16560 18530 -16550 18550
rect -16530 18530 -16520 18550
rect -16560 18520 -16520 18530
rect -16480 18870 -16440 18880
rect -16480 18850 -16470 18870
rect -16450 18850 -16440 18870
rect -16480 18710 -16440 18850
rect -16480 18690 -16470 18710
rect -16450 18690 -16440 18710
rect -16480 18550 -16440 18690
rect -16480 18530 -16470 18550
rect -16450 18530 -16440 18550
rect -16480 18520 -16440 18530
rect -16400 18870 -16360 18880
rect -16400 18850 -16390 18870
rect -16370 18850 -16360 18870
rect -16400 18710 -16360 18850
rect -16400 18690 -16390 18710
rect -16370 18690 -16360 18710
rect -16400 18550 -16360 18690
rect -16400 18530 -16390 18550
rect -16370 18530 -16360 18550
rect -16400 18520 -16360 18530
rect -16320 18870 -16280 18880
rect -16320 18850 -16310 18870
rect -16290 18850 -16280 18870
rect -16320 18710 -16280 18850
rect -16320 18690 -16310 18710
rect -16290 18690 -16280 18710
rect -16320 18550 -16280 18690
rect -16320 18530 -16310 18550
rect -16290 18530 -16280 18550
rect -16320 18520 -16280 18530
rect -16240 18870 -16200 18880
rect -16240 18850 -16230 18870
rect -16210 18850 -16200 18870
rect -16240 18710 -16200 18850
rect -16240 18690 -16230 18710
rect -16210 18690 -16200 18710
rect -16240 18550 -16200 18690
rect -16240 18530 -16230 18550
rect -16210 18530 -16200 18550
rect -16240 18520 -16200 18530
rect -16160 18870 -16120 18880
rect -16160 18850 -16150 18870
rect -16130 18850 -16120 18870
rect -16160 18710 -16120 18850
rect -16160 18690 -16150 18710
rect -16130 18690 -16120 18710
rect -16160 18550 -16120 18690
rect -16160 18530 -16150 18550
rect -16130 18530 -16120 18550
rect -16160 18520 -16120 18530
rect -16080 18870 -16040 18880
rect -16080 18850 -16070 18870
rect -16050 18850 -16040 18870
rect -16080 18710 -16040 18850
rect -16080 18690 -16070 18710
rect -16050 18690 -16040 18710
rect -16080 18550 -16040 18690
rect -16080 18530 -16070 18550
rect -16050 18530 -16040 18550
rect -16080 18520 -16040 18530
rect -16000 18870 -15960 18880
rect -16000 18850 -15990 18870
rect -15970 18850 -15960 18870
rect -16000 18710 -15960 18850
rect -16000 18690 -15990 18710
rect -15970 18690 -15960 18710
rect -16000 18550 -15960 18690
rect -16000 18530 -15990 18550
rect -15970 18530 -15960 18550
rect -16000 18520 -15960 18530
rect -15920 18870 -15880 18880
rect -15920 18850 -15910 18870
rect -15890 18850 -15880 18870
rect -15920 18710 -15880 18850
rect -15920 18690 -15910 18710
rect -15890 18690 -15880 18710
rect -15920 18550 -15880 18690
rect -15920 18530 -15910 18550
rect -15890 18530 -15880 18550
rect -15920 18520 -15880 18530
rect -15840 18870 -15800 18880
rect -15840 18850 -15830 18870
rect -15810 18850 -15800 18870
rect -15840 18710 -15800 18850
rect -15840 18690 -15830 18710
rect -15810 18690 -15800 18710
rect -15840 18550 -15800 18690
rect -15840 18530 -15830 18550
rect -15810 18530 -15800 18550
rect -15840 18520 -15800 18530
rect -15760 18870 -15720 18880
rect -15760 18850 -15750 18870
rect -15730 18850 -15720 18870
rect -15760 18710 -15720 18850
rect -15760 18690 -15750 18710
rect -15730 18690 -15720 18710
rect -15760 18550 -15720 18690
rect -15760 18530 -15750 18550
rect -15730 18530 -15720 18550
rect -15760 18520 -15720 18530
rect -15680 18870 -15640 18880
rect -15680 18850 -15670 18870
rect -15650 18850 -15640 18870
rect -15680 18710 -15640 18850
rect -15680 18690 -15670 18710
rect -15650 18690 -15640 18710
rect -15680 18550 -15640 18690
rect -15680 18530 -15670 18550
rect -15650 18530 -15640 18550
rect -15680 18520 -15640 18530
rect -15600 18870 -15560 18880
rect -15600 18850 -15590 18870
rect -15570 18850 -15560 18870
rect -15600 18710 -15560 18850
rect -15600 18690 -15590 18710
rect -15570 18690 -15560 18710
rect -15600 18550 -15560 18690
rect -15600 18530 -15590 18550
rect -15570 18530 -15560 18550
rect -15600 18520 -15560 18530
rect 20520 18030 20560 18040
rect 20520 18010 20530 18030
rect 20550 18010 20560 18030
rect 20520 17870 20560 18010
rect 20520 17850 20530 17870
rect 20550 17850 20560 17870
rect 20520 17840 20560 17850
rect 20600 18030 20640 18040
rect 20600 18010 20610 18030
rect 20630 18010 20640 18030
rect 20600 17870 20640 18010
rect 20600 17850 20610 17870
rect 20630 17850 20640 17870
rect 20600 17840 20640 17850
rect 20680 18030 20720 18040
rect 20680 18010 20690 18030
rect 20710 18010 20720 18030
rect 20680 17870 20720 18010
rect 20680 17850 20690 17870
rect 20710 17850 20720 17870
rect 20680 17840 20720 17850
rect 20760 18030 20800 18040
rect 20760 18010 20770 18030
rect 20790 18010 20800 18030
rect 20760 17870 20800 18010
rect 20760 17850 20770 17870
rect 20790 17850 20800 17870
rect 20760 17840 20800 17850
rect 20840 18030 20880 18040
rect 20840 18010 20850 18030
rect 20870 18010 20880 18030
rect 20840 17870 20880 18010
rect 20840 17850 20850 17870
rect 20870 17850 20880 17870
rect 20840 17840 20880 17850
rect 20920 18030 20960 18040
rect 20920 18010 20930 18030
rect 20950 18010 20960 18030
rect 20920 17870 20960 18010
rect 20920 17850 20930 17870
rect 20950 17850 20960 17870
rect 20920 17840 20960 17850
rect 21000 18030 21040 18040
rect 21000 18010 21010 18030
rect 21030 18010 21040 18030
rect 21000 17870 21040 18010
rect 21000 17850 21010 17870
rect 21030 17850 21040 17870
rect 21000 17840 21040 17850
rect 21080 18030 21120 18040
rect 21080 18010 21090 18030
rect 21110 18010 21120 18030
rect 21080 17870 21120 18010
rect 21080 17850 21090 17870
rect 21110 17850 21120 17870
rect 21080 17840 21120 17850
rect 21160 18030 21200 18040
rect 21160 18010 21170 18030
rect 21190 18010 21200 18030
rect 21160 17870 21200 18010
rect 21160 17850 21170 17870
rect 21190 17850 21200 17870
rect 21160 17840 21200 17850
rect 21240 18030 21280 18040
rect 21240 18010 21250 18030
rect 21270 18010 21280 18030
rect 21240 17870 21280 18010
rect 21240 17850 21250 17870
rect 21270 17850 21280 17870
rect 21240 17840 21280 17850
rect 21320 18030 21360 18040
rect 21320 18010 21330 18030
rect 21350 18010 21360 18030
rect 21320 17870 21360 18010
rect 21320 17850 21330 17870
rect 21350 17850 21360 17870
rect 21320 17840 21360 17850
rect 21400 18030 21440 18040
rect 21400 18010 21410 18030
rect 21430 18010 21440 18030
rect 21400 17870 21440 18010
rect 21400 17850 21410 17870
rect 21430 17850 21440 17870
rect 21400 17840 21440 17850
rect 21480 18030 21520 18040
rect 21480 18010 21490 18030
rect 21510 18010 21520 18030
rect 21480 17870 21520 18010
rect 21480 17850 21490 17870
rect 21510 17850 21520 17870
rect 21480 17840 21520 17850
rect 21560 18030 21600 18040
rect 21560 18010 21570 18030
rect 21590 18010 21600 18030
rect 21560 17870 21600 18010
rect 21560 17850 21570 17870
rect 21590 17850 21600 17870
rect 21560 17840 21600 17850
rect -16560 17350 -16520 17360
rect -16560 17330 -16550 17350
rect -16530 17330 -16520 17350
rect -16560 17190 -16520 17330
rect -16560 17170 -16550 17190
rect -16530 17170 -16520 17190
rect -16560 17160 -16520 17170
rect -16480 17350 -16440 17360
rect -16480 17330 -16470 17350
rect -16450 17330 -16440 17350
rect -16480 17190 -16440 17330
rect -16480 17170 -16470 17190
rect -16450 17170 -16440 17190
rect -16480 17160 -16440 17170
rect -16400 17350 -16360 17360
rect -16400 17330 -16390 17350
rect -16370 17330 -16360 17350
rect -16400 17190 -16360 17330
rect -16400 17170 -16390 17190
rect -16370 17170 -16360 17190
rect -16400 17160 -16360 17170
rect -16320 17350 -16280 17360
rect -16320 17330 -16310 17350
rect -16290 17330 -16280 17350
rect -16320 17190 -16280 17330
rect -16320 17170 -16310 17190
rect -16290 17170 -16280 17190
rect -16320 17160 -16280 17170
rect -16240 17350 -16200 17360
rect -16240 17330 -16230 17350
rect -16210 17330 -16200 17350
rect -16240 17190 -16200 17330
rect -16240 17170 -16230 17190
rect -16210 17170 -16200 17190
rect -16240 17160 -16200 17170
rect -16160 17350 -16120 17360
rect -16160 17330 -16150 17350
rect -16130 17330 -16120 17350
rect -16160 17190 -16120 17330
rect -16160 17170 -16150 17190
rect -16130 17170 -16120 17190
rect -16160 17160 -16120 17170
rect -16080 17350 -16040 17360
rect -16080 17330 -16070 17350
rect -16050 17330 -16040 17350
rect -16080 17190 -16040 17330
rect -16080 17170 -16070 17190
rect -16050 17170 -16040 17190
rect -16080 17160 -16040 17170
rect -16000 17350 -15960 17360
rect -16000 17330 -15990 17350
rect -15970 17330 -15960 17350
rect -16000 17190 -15960 17330
rect -16000 17170 -15990 17190
rect -15970 17170 -15960 17190
rect -16000 17160 -15960 17170
rect -15920 17350 -15880 17360
rect -15920 17330 -15910 17350
rect -15890 17330 -15880 17350
rect -15920 17190 -15880 17330
rect -15920 17170 -15910 17190
rect -15890 17170 -15880 17190
rect -15920 17160 -15880 17170
rect -15840 17350 -15800 17360
rect -15840 17330 -15830 17350
rect -15810 17330 -15800 17350
rect -15840 17190 -15800 17330
rect -15840 17170 -15830 17190
rect -15810 17170 -15800 17190
rect -15840 17160 -15800 17170
rect -15760 17350 -15720 17360
rect -15760 17330 -15750 17350
rect -15730 17330 -15720 17350
rect -15760 17190 -15720 17330
rect -15760 17170 -15750 17190
rect -15730 17170 -15720 17190
rect -15760 17160 -15720 17170
rect -15680 17350 -15640 17360
rect -15680 17330 -15670 17350
rect -15650 17330 -15640 17350
rect -15680 17190 -15640 17330
rect -15680 17170 -15670 17190
rect -15650 17170 -15640 17190
rect -15680 17160 -15640 17170
rect -15600 17350 -15560 17360
rect -15600 17330 -15590 17350
rect -15570 17330 -15560 17350
rect -15600 17190 -15560 17330
rect -15600 17170 -15590 17190
rect -15570 17170 -15560 17190
rect -15600 17160 -15560 17170
rect -14960 17350 -14920 17360
rect -14960 17330 -14950 17350
rect -14930 17330 -14920 17350
rect -14960 17190 -14920 17330
rect -14960 17170 -14950 17190
rect -14930 17170 -14920 17190
rect -14960 17160 -14920 17170
rect -14880 17350 -14840 17360
rect -14880 17330 -14870 17350
rect -14850 17330 -14840 17350
rect -14880 17190 -14840 17330
rect -14880 17170 -14870 17190
rect -14850 17170 -14840 17190
rect -14880 17160 -14840 17170
rect -14800 17350 -14760 17360
rect -14800 17330 -14790 17350
rect -14770 17330 -14760 17350
rect -14800 17190 -14760 17330
rect -14800 17170 -14790 17190
rect -14770 17170 -14760 17190
rect -14800 17160 -14760 17170
rect -14720 17350 -14680 17360
rect -14720 17330 -14710 17350
rect -14690 17330 -14680 17350
rect -14720 17190 -14680 17330
rect -14720 17170 -14710 17190
rect -14690 17170 -14680 17190
rect -14720 17160 -14680 17170
rect -14640 17350 -14600 17360
rect -14640 17330 -14630 17350
rect -14610 17330 -14600 17350
rect -14640 17190 -14600 17330
rect -14640 17170 -14630 17190
rect -14610 17170 -14600 17190
rect -14640 17160 -14600 17170
rect -14560 17350 -14520 17360
rect -14560 17330 -14550 17350
rect -14530 17330 -14520 17350
rect -14560 17190 -14520 17330
rect -14560 17170 -14550 17190
rect -14530 17170 -14520 17190
rect -14560 17160 -14520 17170
rect -14480 17350 -14440 17360
rect -14480 17330 -14470 17350
rect -14450 17330 -14440 17350
rect -14480 17190 -14440 17330
rect -14480 17170 -14470 17190
rect -14450 17170 -14440 17190
rect -14480 17160 -14440 17170
rect -14400 17350 -14360 17360
rect -14400 17330 -14390 17350
rect -14370 17330 -14360 17350
rect -14400 17190 -14360 17330
rect -14400 17170 -14390 17190
rect -14370 17170 -14360 17190
rect -14400 17160 -14360 17170
rect -14320 17350 -14280 17360
rect -14320 17330 -14310 17350
rect -14290 17330 -14280 17350
rect -14320 17190 -14280 17330
rect -14320 17170 -14310 17190
rect -14290 17170 -14280 17190
rect -14320 17160 -14280 17170
rect -14240 17350 -14200 17360
rect -14240 17330 -14230 17350
rect -14210 17330 -14200 17350
rect -14240 17190 -14200 17330
rect -14240 17170 -14230 17190
rect -14210 17170 -14200 17190
rect -14240 17160 -14200 17170
rect -14160 17350 -14120 17360
rect -14160 17330 -14150 17350
rect -14130 17330 -14120 17350
rect -14160 17190 -14120 17330
rect -14160 17170 -14150 17190
rect -14130 17170 -14120 17190
rect -14160 17160 -14120 17170
rect -14080 17350 -14040 17360
rect -14080 17330 -14070 17350
rect -14050 17330 -14040 17350
rect -14080 17190 -14040 17330
rect -14080 17170 -14070 17190
rect -14050 17170 -14040 17190
rect -14080 17160 -14040 17170
rect -14000 17350 -13960 17360
rect -14000 17330 -13990 17350
rect -13970 17330 -13960 17350
rect -14000 17190 -13960 17330
rect -14000 17170 -13990 17190
rect -13970 17170 -13960 17190
rect -14000 17160 -13960 17170
rect -13920 17350 -13880 17360
rect -13920 17330 -13910 17350
rect -13890 17330 -13880 17350
rect -13920 17190 -13880 17330
rect -13920 17170 -13910 17190
rect -13890 17170 -13880 17190
rect -13920 17160 -13880 17170
rect -13840 17350 -13800 17360
rect -13840 17330 -13830 17350
rect -13810 17330 -13800 17350
rect -13840 17190 -13800 17330
rect -13840 17170 -13830 17190
rect -13810 17170 -13800 17190
rect -13840 17160 -13800 17170
rect -13760 17350 -13720 17360
rect -13760 17330 -13750 17350
rect -13730 17330 -13720 17350
rect -13760 17190 -13720 17330
rect -13760 17170 -13750 17190
rect -13730 17170 -13720 17190
rect -13760 17160 -13720 17170
rect -13680 17350 -13640 17360
rect -13680 17330 -13670 17350
rect -13650 17330 -13640 17350
rect -13680 17190 -13640 17330
rect -13680 17170 -13670 17190
rect -13650 17170 -13640 17190
rect -13680 17160 -13640 17170
rect -13600 17350 -13560 17360
rect -13600 17330 -13590 17350
rect -13570 17330 -13560 17350
rect -13600 17190 -13560 17330
rect -13600 17170 -13590 17190
rect -13570 17170 -13560 17190
rect -13600 17160 -13560 17170
rect -13520 17350 -13480 17360
rect -13520 17330 -13510 17350
rect -13490 17330 -13480 17350
rect -13520 17190 -13480 17330
rect -13520 17170 -13510 17190
rect -13490 17170 -13480 17190
rect -13520 17160 -13480 17170
rect -13440 17350 -13400 17360
rect -13440 17330 -13430 17350
rect -13410 17330 -13400 17350
rect -13440 17190 -13400 17330
rect -13440 17170 -13430 17190
rect -13410 17170 -13400 17190
rect -13440 17160 -13400 17170
rect -13360 17350 -13320 17360
rect -13360 17330 -13350 17350
rect -13330 17330 -13320 17350
rect -13360 17190 -13320 17330
rect -13360 17170 -13350 17190
rect -13330 17170 -13320 17190
rect -13360 17160 -13320 17170
rect -13280 17350 -13240 17360
rect -13280 17330 -13270 17350
rect -13250 17330 -13240 17350
rect -13280 17190 -13240 17330
rect -13280 17170 -13270 17190
rect -13250 17170 -13240 17190
rect -13280 17160 -13240 17170
rect -13200 17350 -13160 17360
rect -13200 17330 -13190 17350
rect -13170 17330 -13160 17350
rect -13200 17190 -13160 17330
rect -13200 17170 -13190 17190
rect -13170 17170 -13160 17190
rect -13200 17160 -13160 17170
rect -13120 17350 -13080 17360
rect -13120 17330 -13110 17350
rect -13090 17330 -13080 17350
rect -13120 17190 -13080 17330
rect -13120 17170 -13110 17190
rect -13090 17170 -13080 17190
rect -13120 17160 -13080 17170
rect -13040 17350 -13000 17360
rect -13040 17330 -13030 17350
rect -13010 17330 -13000 17350
rect -13040 17190 -13000 17330
rect -13040 17170 -13030 17190
rect -13010 17170 -13000 17190
rect -13040 17160 -13000 17170
rect -12960 17350 -12920 17360
rect -12960 17330 -12950 17350
rect -12930 17330 -12920 17350
rect -12960 17190 -12920 17330
rect -12960 17170 -12950 17190
rect -12930 17170 -12920 17190
rect -12960 17160 -12920 17170
rect -12880 17350 -12840 17360
rect -12880 17330 -12870 17350
rect -12850 17330 -12840 17350
rect -12880 17190 -12840 17330
rect -12880 17170 -12870 17190
rect -12850 17170 -12840 17190
rect -12880 17160 -12840 17170
rect -12800 17350 -12760 17360
rect -12800 17330 -12790 17350
rect -12770 17330 -12760 17350
rect -12800 17190 -12760 17330
rect -12800 17170 -12790 17190
rect -12770 17170 -12760 17190
rect -12800 17160 -12760 17170
rect -12720 17350 -12680 17360
rect -12720 17330 -12710 17350
rect -12690 17330 -12680 17350
rect -12720 17190 -12680 17330
rect -12720 17170 -12710 17190
rect -12690 17170 -12680 17190
rect -12720 17160 -12680 17170
rect -12640 17350 -12600 17360
rect -12640 17330 -12630 17350
rect -12610 17330 -12600 17350
rect -12640 17190 -12600 17330
rect -12640 17170 -12630 17190
rect -12610 17170 -12600 17190
rect -12640 17160 -12600 17170
rect -12560 17350 -12520 17360
rect -12560 17330 -12550 17350
rect -12530 17330 -12520 17350
rect -12560 17190 -12520 17330
rect -12560 17170 -12550 17190
rect -12530 17170 -12520 17190
rect -12560 17160 -12520 17170
rect -12480 17350 -12440 17360
rect -12480 17330 -12470 17350
rect -12450 17330 -12440 17350
rect -12480 17190 -12440 17330
rect -12480 17170 -12470 17190
rect -12450 17170 -12440 17190
rect -12480 17160 -12440 17170
rect -12400 17350 -12360 17360
rect -12400 17330 -12390 17350
rect -12370 17330 -12360 17350
rect -12400 17190 -12360 17330
rect -12400 17170 -12390 17190
rect -12370 17170 -12360 17190
rect -12400 17160 -12360 17170
rect -12320 17350 -12280 17360
rect -12320 17330 -12310 17350
rect -12290 17330 -12280 17350
rect -12320 17190 -12280 17330
rect -12320 17170 -12310 17190
rect -12290 17170 -12280 17190
rect -12320 17160 -12280 17170
rect -12240 17350 -12200 17360
rect -12240 17330 -12230 17350
rect -12210 17330 -12200 17350
rect -12240 17190 -12200 17330
rect -12240 17170 -12230 17190
rect -12210 17170 -12200 17190
rect -12240 17160 -12200 17170
rect -12160 17350 -12120 17360
rect -12160 17330 -12150 17350
rect -12130 17330 -12120 17350
rect -12160 17190 -12120 17330
rect -12160 17170 -12150 17190
rect -12130 17170 -12120 17190
rect -12160 17160 -12120 17170
rect -12080 17350 -12040 17360
rect -12080 17330 -12070 17350
rect -12050 17330 -12040 17350
rect -12080 17190 -12040 17330
rect -12080 17170 -12070 17190
rect -12050 17170 -12040 17190
rect -12080 17160 -12040 17170
rect -12000 17350 -11960 17360
rect -12000 17330 -11990 17350
rect -11970 17330 -11960 17350
rect -12000 17190 -11960 17330
rect -12000 17170 -11990 17190
rect -11970 17170 -11960 17190
rect -12000 17160 -11960 17170
rect -11920 17350 -11880 17360
rect -11920 17330 -11910 17350
rect -11890 17330 -11880 17350
rect -11920 17190 -11880 17330
rect -11920 17170 -11910 17190
rect -11890 17170 -11880 17190
rect -11920 17160 -11880 17170
rect -11840 17350 -11800 17360
rect -11840 17330 -11830 17350
rect -11810 17330 -11800 17350
rect -11840 17190 -11800 17330
rect -11840 17170 -11830 17190
rect -11810 17170 -11800 17190
rect -11840 17160 -11800 17170
rect -11760 17350 -11720 17360
rect -11760 17330 -11750 17350
rect -11730 17330 -11720 17350
rect -11760 17190 -11720 17330
rect -11760 17170 -11750 17190
rect -11730 17170 -11720 17190
rect -11760 17160 -11720 17170
rect -11680 17350 -11640 17360
rect -11680 17330 -11670 17350
rect -11650 17330 -11640 17350
rect -11680 17190 -11640 17330
rect -11680 17170 -11670 17190
rect -11650 17170 -11640 17190
rect -11680 17160 -11640 17170
rect -11600 17350 -11560 17360
rect -11600 17330 -11590 17350
rect -11570 17330 -11560 17350
rect -11600 17190 -11560 17330
rect -11600 17170 -11590 17190
rect -11570 17170 -11560 17190
rect -11600 17160 -11560 17170
rect -11520 17350 -11480 17360
rect -11520 17330 -11510 17350
rect -11490 17330 -11480 17350
rect -11520 17190 -11480 17330
rect -11520 17170 -11510 17190
rect -11490 17170 -11480 17190
rect -11520 17160 -11480 17170
rect -11440 17350 -11400 17360
rect -11440 17330 -11430 17350
rect -11410 17330 -11400 17350
rect -11440 17190 -11400 17330
rect -11440 17170 -11430 17190
rect -11410 17170 -11400 17190
rect -11440 17160 -11400 17170
rect -11360 17350 -11320 17360
rect -11360 17330 -11350 17350
rect -11330 17330 -11320 17350
rect -11360 17190 -11320 17330
rect -11360 17170 -11350 17190
rect -11330 17170 -11320 17190
rect -11360 17160 -11320 17170
rect -11280 17350 -11240 17360
rect -11280 17330 -11270 17350
rect -11250 17330 -11240 17350
rect -11280 17190 -11240 17330
rect -11280 17170 -11270 17190
rect -11250 17170 -11240 17190
rect -11280 17160 -11240 17170
rect -11200 17350 -11160 17360
rect -11200 17330 -11190 17350
rect -11170 17330 -11160 17350
rect -11200 17190 -11160 17330
rect -11200 17170 -11190 17190
rect -11170 17170 -11160 17190
rect -11200 17160 -11160 17170
rect -11120 17350 -11080 17360
rect -11120 17330 -11110 17350
rect -11090 17330 -11080 17350
rect -11120 17190 -11080 17330
rect -11120 17170 -11110 17190
rect -11090 17170 -11080 17190
rect -11120 17160 -11080 17170
rect -11040 17350 -11000 17360
rect -11040 17330 -11030 17350
rect -11010 17330 -11000 17350
rect -11040 17190 -11000 17330
rect -11040 17170 -11030 17190
rect -11010 17170 -11000 17190
rect -11040 17160 -11000 17170
rect -10960 17350 -10920 17360
rect -10960 17330 -10950 17350
rect -10930 17330 -10920 17350
rect -10960 17190 -10920 17330
rect -10960 17170 -10950 17190
rect -10930 17170 -10920 17190
rect -10960 17160 -10920 17170
rect -10880 17350 -10840 17360
rect -10880 17330 -10870 17350
rect -10850 17330 -10840 17350
rect -10880 17190 -10840 17330
rect -10880 17170 -10870 17190
rect -10850 17170 -10840 17190
rect -10880 17160 -10840 17170
rect -10800 17350 -10760 17360
rect -10800 17330 -10790 17350
rect -10770 17330 -10760 17350
rect -10800 17190 -10760 17330
rect -10800 17170 -10790 17190
rect -10770 17170 -10760 17190
rect -10800 17160 -10760 17170
rect -10720 17350 -10680 17360
rect -10720 17330 -10710 17350
rect -10690 17330 -10680 17350
rect -10720 17190 -10680 17330
rect -10720 17170 -10710 17190
rect -10690 17170 -10680 17190
rect -10720 17160 -10680 17170
rect -10640 17350 -10600 17360
rect -10640 17330 -10630 17350
rect -10610 17330 -10600 17350
rect -10640 17190 -10600 17330
rect -10640 17170 -10630 17190
rect -10610 17170 -10600 17190
rect -10640 17160 -10600 17170
rect -10560 17350 -10520 17360
rect -10560 17330 -10550 17350
rect -10530 17330 -10520 17350
rect -10560 17190 -10520 17330
rect -10560 17170 -10550 17190
rect -10530 17170 -10520 17190
rect -10560 17160 -10520 17170
rect -10480 17350 -10440 17360
rect -10480 17330 -10470 17350
rect -10450 17330 -10440 17350
rect -10480 17190 -10440 17330
rect -10480 17170 -10470 17190
rect -10450 17170 -10440 17190
rect -10480 17160 -10440 17170
rect -10400 17350 -10360 17360
rect -10400 17330 -10390 17350
rect -10370 17330 -10360 17350
rect -10400 17190 -10360 17330
rect -10400 17170 -10390 17190
rect -10370 17170 -10360 17190
rect -10400 17160 -10360 17170
rect -10320 17350 -10280 17360
rect -10320 17330 -10310 17350
rect -10290 17330 -10280 17350
rect -10320 17190 -10280 17330
rect -10320 17170 -10310 17190
rect -10290 17170 -10280 17190
rect -10320 17160 -10280 17170
rect -10240 17350 -10200 17360
rect -10240 17330 -10230 17350
rect -10210 17330 -10200 17350
rect -10240 17190 -10200 17330
rect -10240 17170 -10230 17190
rect -10210 17170 -10200 17190
rect -10240 17160 -10200 17170
rect -10160 17350 -10120 17360
rect -10160 17330 -10150 17350
rect -10130 17330 -10120 17350
rect -10160 17190 -10120 17330
rect -10160 17170 -10150 17190
rect -10130 17170 -10120 17190
rect -10160 17160 -10120 17170
rect -10080 17350 -10040 17360
rect -10080 17330 -10070 17350
rect -10050 17330 -10040 17350
rect -10080 17190 -10040 17330
rect -10080 17170 -10070 17190
rect -10050 17170 -10040 17190
rect -10080 17160 -10040 17170
rect -10000 17350 -9960 17360
rect -10000 17330 -9990 17350
rect -9970 17330 -9960 17350
rect -10000 17190 -9960 17330
rect -10000 17170 -9990 17190
rect -9970 17170 -9960 17190
rect -10000 17160 -9960 17170
rect -9920 17350 -9880 17360
rect -9920 17330 -9910 17350
rect -9890 17330 -9880 17350
rect -9920 17190 -9880 17330
rect -9920 17170 -9910 17190
rect -9890 17170 -9880 17190
rect -9920 17160 -9880 17170
rect -9840 17350 -9800 17360
rect -9840 17330 -9830 17350
rect -9810 17330 -9800 17350
rect -9840 17190 -9800 17330
rect -9840 17170 -9830 17190
rect -9810 17170 -9800 17190
rect -9840 17160 -9800 17170
rect -9760 17350 -9720 17360
rect -9760 17330 -9750 17350
rect -9730 17330 -9720 17350
rect -9760 17190 -9720 17330
rect -9760 17170 -9750 17190
rect -9730 17170 -9720 17190
rect -9760 17160 -9720 17170
rect -9680 17350 -9640 17360
rect -9680 17330 -9670 17350
rect -9650 17330 -9640 17350
rect -9680 17190 -9640 17330
rect -9680 17170 -9670 17190
rect -9650 17170 -9640 17190
rect -9680 17160 -9640 17170
rect -9600 17350 -9560 17360
rect -9600 17330 -9590 17350
rect -9570 17330 -9560 17350
rect -9600 17190 -9560 17330
rect -9600 17170 -9590 17190
rect -9570 17170 -9560 17190
rect -9600 17160 -9560 17170
rect -9520 17350 -9480 17360
rect -9520 17330 -9510 17350
rect -9490 17330 -9480 17350
rect -9520 17190 -9480 17330
rect -9520 17170 -9510 17190
rect -9490 17170 -9480 17190
rect -9520 17160 -9480 17170
rect -9440 17350 -9400 17360
rect -9440 17330 -9430 17350
rect -9410 17330 -9400 17350
rect -9440 17190 -9400 17330
rect -9440 17170 -9430 17190
rect -9410 17170 -9400 17190
rect -9440 17160 -9400 17170
rect -9360 17350 -9320 17360
rect -9360 17330 -9350 17350
rect -9330 17330 -9320 17350
rect -9360 17190 -9320 17330
rect -9360 17170 -9350 17190
rect -9330 17170 -9320 17190
rect -9360 17160 -9320 17170
rect -9280 17350 -9240 17360
rect -9280 17330 -9270 17350
rect -9250 17330 -9240 17350
rect -9280 17190 -9240 17330
rect -9280 17170 -9270 17190
rect -9250 17170 -9240 17190
rect -9280 17160 -9240 17170
rect -9200 17350 -9160 17360
rect -9200 17330 -9190 17350
rect -9170 17330 -9160 17350
rect -9200 17190 -9160 17330
rect -9200 17170 -9190 17190
rect -9170 17170 -9160 17190
rect -9200 17160 -9160 17170
rect -9120 17350 -9080 17360
rect -9120 17330 -9110 17350
rect -9090 17330 -9080 17350
rect -9120 17190 -9080 17330
rect -9120 17170 -9110 17190
rect -9090 17170 -9080 17190
rect -9120 17160 -9080 17170
rect -9040 17350 -9000 17360
rect -9040 17330 -9030 17350
rect -9010 17330 -9000 17350
rect -9040 17190 -9000 17330
rect -9040 17170 -9030 17190
rect -9010 17170 -9000 17190
rect -9040 17160 -9000 17170
rect -8960 17350 -8920 17360
rect -8960 17330 -8950 17350
rect -8930 17330 -8920 17350
rect -8960 17190 -8920 17330
rect -8960 17170 -8950 17190
rect -8930 17170 -8920 17190
rect -8960 17160 -8920 17170
rect -8880 17350 -8840 17360
rect -8880 17330 -8870 17350
rect -8850 17330 -8840 17350
rect -8880 17190 -8840 17330
rect -8880 17170 -8870 17190
rect -8850 17170 -8840 17190
rect -8880 17160 -8840 17170
rect -8800 17350 -8760 17360
rect -8800 17330 -8790 17350
rect -8770 17330 -8760 17350
rect -8800 17190 -8760 17330
rect -8800 17170 -8790 17190
rect -8770 17170 -8760 17190
rect -8800 17160 -8760 17170
rect -8720 17350 -8680 17360
rect -8720 17330 -8710 17350
rect -8690 17330 -8680 17350
rect -8720 17190 -8680 17330
rect -8720 17170 -8710 17190
rect -8690 17170 -8680 17190
rect -8720 17160 -8680 17170
rect -8640 17350 -8600 17360
rect -8640 17330 -8630 17350
rect -8610 17330 -8600 17350
rect -8640 17190 -8600 17330
rect -8640 17170 -8630 17190
rect -8610 17170 -8600 17190
rect -8640 17160 -8600 17170
rect -8560 17350 -8520 17360
rect -8560 17330 -8550 17350
rect -8530 17330 -8520 17350
rect -8560 17190 -8520 17330
rect -8560 17170 -8550 17190
rect -8530 17170 -8520 17190
rect -8560 17160 -8520 17170
rect -8480 17350 -8440 17360
rect -8480 17330 -8470 17350
rect -8450 17330 -8440 17350
rect -8480 17190 -8440 17330
rect -8480 17170 -8470 17190
rect -8450 17170 -8440 17190
rect -8480 17160 -8440 17170
rect -8400 17350 -8360 17360
rect -8400 17330 -8390 17350
rect -8370 17330 -8360 17350
rect -8400 17190 -8360 17330
rect -8400 17170 -8390 17190
rect -8370 17170 -8360 17190
rect -8400 17160 -8360 17170
rect -8320 17350 -8280 17360
rect -8320 17330 -8310 17350
rect -8290 17330 -8280 17350
rect -8320 17190 -8280 17330
rect -8320 17170 -8310 17190
rect -8290 17170 -8280 17190
rect -8320 17160 -8280 17170
rect -8240 17350 -8200 17360
rect -8240 17330 -8230 17350
rect -8210 17330 -8200 17350
rect -8240 17190 -8200 17330
rect -8240 17170 -8230 17190
rect -8210 17170 -8200 17190
rect -8240 17160 -8200 17170
rect -8160 17350 -8120 17360
rect -8160 17330 -8150 17350
rect -8130 17330 -8120 17350
rect -8160 17190 -8120 17330
rect -8160 17170 -8150 17190
rect -8130 17170 -8120 17190
rect -8160 17160 -8120 17170
rect -8080 17350 -8040 17360
rect -8080 17330 -8070 17350
rect -8050 17330 -8040 17350
rect -8080 17190 -8040 17330
rect -8080 17170 -8070 17190
rect -8050 17170 -8040 17190
rect -8080 17160 -8040 17170
rect -8000 17350 -7960 17360
rect -8000 17330 -7990 17350
rect -7970 17330 -7960 17350
rect -8000 17190 -7960 17330
rect -8000 17170 -7990 17190
rect -7970 17170 -7960 17190
rect -8000 17160 -7960 17170
rect -7920 17350 -7880 17360
rect -7920 17330 -7910 17350
rect -7890 17330 -7880 17350
rect -7920 17190 -7880 17330
rect -7920 17170 -7910 17190
rect -7890 17170 -7880 17190
rect -7920 17160 -7880 17170
rect -7840 17350 -7800 17360
rect -7840 17330 -7830 17350
rect -7810 17330 -7800 17350
rect -7840 17190 -7800 17330
rect -7840 17170 -7830 17190
rect -7810 17170 -7800 17190
rect -7840 17160 -7800 17170
rect -7760 17350 -7720 17360
rect -7760 17330 -7750 17350
rect -7730 17330 -7720 17350
rect -7760 17190 -7720 17330
rect -7760 17170 -7750 17190
rect -7730 17170 -7720 17190
rect -7760 17160 -7720 17170
rect -7680 17350 -7640 17360
rect -7680 17330 -7670 17350
rect -7650 17330 -7640 17350
rect -7680 17190 -7640 17330
rect -7680 17170 -7670 17190
rect -7650 17170 -7640 17190
rect -7680 17160 -7640 17170
rect -7600 17350 -7560 17360
rect -7600 17330 -7590 17350
rect -7570 17330 -7560 17350
rect -7600 17190 -7560 17330
rect -7600 17170 -7590 17190
rect -7570 17170 -7560 17190
rect -7600 17160 -7560 17170
rect -7520 17350 -7480 17360
rect -7520 17330 -7510 17350
rect -7490 17330 -7480 17350
rect -7520 17190 -7480 17330
rect -7520 17170 -7510 17190
rect -7490 17170 -7480 17190
rect -7520 17160 -7480 17170
rect -7440 17350 -7400 17360
rect -7440 17330 -7430 17350
rect -7410 17330 -7400 17350
rect -7440 17190 -7400 17330
rect -7440 17170 -7430 17190
rect -7410 17170 -7400 17190
rect -7440 17160 -7400 17170
rect -7360 17350 -7320 17360
rect -7360 17330 -7350 17350
rect -7330 17330 -7320 17350
rect -7360 17190 -7320 17330
rect -7360 17170 -7350 17190
rect -7330 17170 -7320 17190
rect -7360 17160 -7320 17170
rect -7280 17350 -7240 17360
rect -7280 17330 -7270 17350
rect -7250 17330 -7240 17350
rect -7280 17190 -7240 17330
rect -7280 17170 -7270 17190
rect -7250 17170 -7240 17190
rect -7280 17160 -7240 17170
rect -7200 17350 -7160 17360
rect -7200 17330 -7190 17350
rect -7170 17330 -7160 17350
rect -7200 17190 -7160 17330
rect -7200 17170 -7190 17190
rect -7170 17170 -7160 17190
rect -7200 17160 -7160 17170
rect -7120 17350 -7080 17360
rect -7120 17330 -7110 17350
rect -7090 17330 -7080 17350
rect -7120 17190 -7080 17330
rect -7120 17170 -7110 17190
rect -7090 17170 -7080 17190
rect -7120 17160 -7080 17170
rect -7040 17350 -7000 17360
rect -7040 17330 -7030 17350
rect -7010 17330 -7000 17350
rect -7040 17190 -7000 17330
rect -7040 17170 -7030 17190
rect -7010 17170 -7000 17190
rect -7040 17160 -7000 17170
rect -6960 17350 -6920 17360
rect -6960 17330 -6950 17350
rect -6930 17330 -6920 17350
rect -6960 17190 -6920 17330
rect -6960 17170 -6950 17190
rect -6930 17170 -6920 17190
rect -6960 17160 -6920 17170
rect -6880 17350 -6840 17360
rect -6880 17330 -6870 17350
rect -6850 17330 -6840 17350
rect -6880 17190 -6840 17330
rect -6880 17170 -6870 17190
rect -6850 17170 -6840 17190
rect -6880 17160 -6840 17170
rect -6800 17350 -6760 17360
rect -6800 17330 -6790 17350
rect -6770 17330 -6760 17350
rect -6800 17190 -6760 17330
rect -6800 17170 -6790 17190
rect -6770 17170 -6760 17190
rect -6800 17160 -6760 17170
rect -6720 17350 -6680 17360
rect -6720 17330 -6710 17350
rect -6690 17330 -6680 17350
rect -6720 17190 -6680 17330
rect -6720 17170 -6710 17190
rect -6690 17170 -6680 17190
rect -6720 17160 -6680 17170
rect -6640 17350 -6600 17360
rect -6640 17330 -6630 17350
rect -6610 17330 -6600 17350
rect -6640 17190 -6600 17330
rect -6640 17170 -6630 17190
rect -6610 17170 -6600 17190
rect -6640 17160 -6600 17170
rect -6560 17350 -6520 17360
rect -6560 17330 -6550 17350
rect -6530 17330 -6520 17350
rect -6560 17190 -6520 17330
rect -6560 17170 -6550 17190
rect -6530 17170 -6520 17190
rect -6560 17160 -6520 17170
rect -6480 17350 -6440 17360
rect -6480 17330 -6470 17350
rect -6450 17330 -6440 17350
rect -6480 17190 -6440 17330
rect -6480 17170 -6470 17190
rect -6450 17170 -6440 17190
rect -6480 17160 -6440 17170
rect -6400 17350 -6360 17360
rect -6400 17330 -6390 17350
rect -6370 17330 -6360 17350
rect -6400 17190 -6360 17330
rect -6400 17170 -6390 17190
rect -6370 17170 -6360 17190
rect -6400 17160 -6360 17170
rect -6320 17350 -6280 17360
rect -6320 17330 -6310 17350
rect -6290 17330 -6280 17350
rect -6320 17190 -6280 17330
rect -6320 17170 -6310 17190
rect -6290 17170 -6280 17190
rect -6320 17160 -6280 17170
rect -6240 17350 -6200 17360
rect -6240 17330 -6230 17350
rect -6210 17330 -6200 17350
rect -6240 17190 -6200 17330
rect -6240 17170 -6230 17190
rect -6210 17170 -6200 17190
rect -6240 17160 -6200 17170
rect -6160 17350 -6120 17360
rect -6160 17330 -6150 17350
rect -6130 17330 -6120 17350
rect -6160 17190 -6120 17330
rect -6160 17170 -6150 17190
rect -6130 17170 -6120 17190
rect -6160 17160 -6120 17170
rect -6080 17350 -6040 17360
rect -6080 17330 -6070 17350
rect -6050 17330 -6040 17350
rect -6080 17190 -6040 17330
rect -6080 17170 -6070 17190
rect -6050 17170 -6040 17190
rect -6080 17160 -6040 17170
rect -6000 17350 -5960 17360
rect -6000 17330 -5990 17350
rect -5970 17330 -5960 17350
rect -6000 17190 -5960 17330
rect -6000 17170 -5990 17190
rect -5970 17170 -5960 17190
rect -6000 17160 -5960 17170
rect -5920 17350 -5880 17360
rect -5920 17330 -5910 17350
rect -5890 17330 -5880 17350
rect -5920 17190 -5880 17330
rect -5920 17170 -5910 17190
rect -5890 17170 -5880 17190
rect -5920 17160 -5880 17170
rect -5840 17350 -5800 17360
rect -5840 17330 -5830 17350
rect -5810 17330 -5800 17350
rect -5840 17190 -5800 17330
rect -5840 17170 -5830 17190
rect -5810 17170 -5800 17190
rect -5840 17160 -5800 17170
rect -5760 17350 -5720 17360
rect -5760 17330 -5750 17350
rect -5730 17330 -5720 17350
rect -5760 17190 -5720 17330
rect -5760 17170 -5750 17190
rect -5730 17170 -5720 17190
rect -5760 17160 -5720 17170
rect -5440 17350 -5400 17360
rect -5440 17330 -5430 17350
rect -5410 17330 -5400 17350
rect -5440 17190 -5400 17330
rect -5440 17170 -5430 17190
rect -5410 17170 -5400 17190
rect -5440 17160 -5400 17170
rect -5280 17350 -5240 17360
rect -5280 17330 -5270 17350
rect -5250 17330 -5240 17350
rect -5280 17190 -5240 17330
rect -5280 17170 -5270 17190
rect -5250 17170 -5240 17190
rect -5280 17160 -5240 17170
rect -14960 16470 -14920 16480
rect -14960 16450 -14950 16470
rect -14930 16450 -14920 16470
rect -14960 16310 -14920 16450
rect -14960 16290 -14950 16310
rect -14930 16290 -14920 16310
rect -14960 16150 -14920 16290
rect -14960 16130 -14950 16150
rect -14930 16130 -14920 16150
rect -14960 15990 -14920 16130
rect -14960 15970 -14950 15990
rect -14930 15970 -14920 15990
rect -14960 15960 -14920 15970
rect -14880 16470 -14840 16480
rect -14880 16450 -14870 16470
rect -14850 16450 -14840 16470
rect -14880 16310 -14840 16450
rect -14880 16290 -14870 16310
rect -14850 16290 -14840 16310
rect -14880 16150 -14840 16290
rect -14880 16130 -14870 16150
rect -14850 16130 -14840 16150
rect -14880 15990 -14840 16130
rect -14880 15970 -14870 15990
rect -14850 15970 -14840 15990
rect -14880 15960 -14840 15970
rect -14800 16470 -14760 16480
rect -14800 16450 -14790 16470
rect -14770 16450 -14760 16470
rect -14800 16310 -14760 16450
rect -14800 16290 -14790 16310
rect -14770 16290 -14760 16310
rect -14800 16150 -14760 16290
rect -14800 16130 -14790 16150
rect -14770 16130 -14760 16150
rect -14800 15990 -14760 16130
rect -14800 15970 -14790 15990
rect -14770 15970 -14760 15990
rect -14800 15960 -14760 15970
rect -14720 16470 -14680 16480
rect -14720 16450 -14710 16470
rect -14690 16450 -14680 16470
rect -14720 16310 -14680 16450
rect -14720 16290 -14710 16310
rect -14690 16290 -14680 16310
rect -14720 16150 -14680 16290
rect -14720 16130 -14710 16150
rect -14690 16130 -14680 16150
rect -14720 15990 -14680 16130
rect -14720 15970 -14710 15990
rect -14690 15970 -14680 15990
rect -14720 15960 -14680 15970
rect -14640 16470 -14600 16480
rect -14640 16450 -14630 16470
rect -14610 16450 -14600 16470
rect -14640 16310 -14600 16450
rect -14640 16290 -14630 16310
rect -14610 16290 -14600 16310
rect -14640 16150 -14600 16290
rect -14640 16130 -14630 16150
rect -14610 16130 -14600 16150
rect -14640 15990 -14600 16130
rect -14640 15970 -14630 15990
rect -14610 15970 -14600 15990
rect -14640 15960 -14600 15970
rect -14560 16470 -14520 16480
rect -14560 16450 -14550 16470
rect -14530 16450 -14520 16470
rect -14560 16310 -14520 16450
rect -14560 16290 -14550 16310
rect -14530 16290 -14520 16310
rect -14560 16150 -14520 16290
rect -14560 16130 -14550 16150
rect -14530 16130 -14520 16150
rect -14560 15990 -14520 16130
rect -14560 15970 -14550 15990
rect -14530 15970 -14520 15990
rect -14560 15960 -14520 15970
rect -14480 16470 -14440 16480
rect -14480 16450 -14470 16470
rect -14450 16450 -14440 16470
rect -14480 16310 -14440 16450
rect -14480 16290 -14470 16310
rect -14450 16290 -14440 16310
rect -14480 16150 -14440 16290
rect -14480 16130 -14470 16150
rect -14450 16130 -14440 16150
rect -14480 15990 -14440 16130
rect -14480 15970 -14470 15990
rect -14450 15970 -14440 15990
rect -14480 15960 -14440 15970
rect -14400 16470 -14360 16480
rect -14400 16450 -14390 16470
rect -14370 16450 -14360 16470
rect -14400 16310 -14360 16450
rect -14400 16290 -14390 16310
rect -14370 16290 -14360 16310
rect -14400 16150 -14360 16290
rect -14400 16130 -14390 16150
rect -14370 16130 -14360 16150
rect -14400 15990 -14360 16130
rect -14400 15970 -14390 15990
rect -14370 15970 -14360 15990
rect -14400 15960 -14360 15970
rect -14320 16470 -14280 16480
rect -14320 16450 -14310 16470
rect -14290 16450 -14280 16470
rect -14320 16310 -14280 16450
rect -14320 16290 -14310 16310
rect -14290 16290 -14280 16310
rect -14320 16150 -14280 16290
rect -14320 16130 -14310 16150
rect -14290 16130 -14280 16150
rect -14320 15990 -14280 16130
rect -14320 15970 -14310 15990
rect -14290 15970 -14280 15990
rect -14320 15960 -14280 15970
rect -14240 16470 -14200 16480
rect -14240 16450 -14230 16470
rect -14210 16450 -14200 16470
rect -14240 16310 -14200 16450
rect -14240 16290 -14230 16310
rect -14210 16290 -14200 16310
rect -14240 16150 -14200 16290
rect -14240 16130 -14230 16150
rect -14210 16130 -14200 16150
rect -14240 15990 -14200 16130
rect -14240 15970 -14230 15990
rect -14210 15970 -14200 15990
rect -14240 15960 -14200 15970
rect -14160 16470 -14120 16480
rect -14160 16450 -14150 16470
rect -14130 16450 -14120 16470
rect -14160 16310 -14120 16450
rect -14160 16290 -14150 16310
rect -14130 16290 -14120 16310
rect -14160 16150 -14120 16290
rect -14160 16130 -14150 16150
rect -14130 16130 -14120 16150
rect -14160 15990 -14120 16130
rect -14160 15970 -14150 15990
rect -14130 15970 -14120 15990
rect -14160 15960 -14120 15970
rect -14080 16470 -14040 16480
rect -14080 16450 -14070 16470
rect -14050 16450 -14040 16470
rect -14080 16310 -14040 16450
rect -14080 16290 -14070 16310
rect -14050 16290 -14040 16310
rect -14080 16150 -14040 16290
rect -14080 16130 -14070 16150
rect -14050 16130 -14040 16150
rect -14080 15990 -14040 16130
rect -14080 15970 -14070 15990
rect -14050 15970 -14040 15990
rect -14080 15960 -14040 15970
rect -14000 16470 -13960 16480
rect -14000 16450 -13990 16470
rect -13970 16450 -13960 16470
rect -14000 16310 -13960 16450
rect -14000 16290 -13990 16310
rect -13970 16290 -13960 16310
rect -14000 16150 -13960 16290
rect -14000 16130 -13990 16150
rect -13970 16130 -13960 16150
rect -14000 15990 -13960 16130
rect -14000 15970 -13990 15990
rect -13970 15970 -13960 15990
rect -14000 15960 -13960 15970
rect -13920 16470 -13880 16480
rect -13920 16450 -13910 16470
rect -13890 16450 -13880 16470
rect -13920 16310 -13880 16450
rect -13920 16290 -13910 16310
rect -13890 16290 -13880 16310
rect -13920 16150 -13880 16290
rect -13920 16130 -13910 16150
rect -13890 16130 -13880 16150
rect -13920 15990 -13880 16130
rect -13920 15970 -13910 15990
rect -13890 15970 -13880 15990
rect -13920 15960 -13880 15970
rect -13840 16470 -13800 16480
rect -13840 16450 -13830 16470
rect -13810 16450 -13800 16470
rect -13840 16310 -13800 16450
rect -13840 16290 -13830 16310
rect -13810 16290 -13800 16310
rect -13840 16150 -13800 16290
rect -13840 16130 -13830 16150
rect -13810 16130 -13800 16150
rect -13840 15990 -13800 16130
rect -13840 15970 -13830 15990
rect -13810 15970 -13800 15990
rect -13840 15960 -13800 15970
rect -13760 16470 -13720 16480
rect -13760 16450 -13750 16470
rect -13730 16450 -13720 16470
rect -13760 16310 -13720 16450
rect -13760 16290 -13750 16310
rect -13730 16290 -13720 16310
rect -13760 16150 -13720 16290
rect -13760 16130 -13750 16150
rect -13730 16130 -13720 16150
rect -13760 15990 -13720 16130
rect -13760 15970 -13750 15990
rect -13730 15970 -13720 15990
rect -13760 15960 -13720 15970
rect -13680 16470 -13640 16480
rect -13680 16450 -13670 16470
rect -13650 16450 -13640 16470
rect -13680 16310 -13640 16450
rect -13680 16290 -13670 16310
rect -13650 16290 -13640 16310
rect -13680 16150 -13640 16290
rect -13680 16130 -13670 16150
rect -13650 16130 -13640 16150
rect -13680 15990 -13640 16130
rect -13680 15970 -13670 15990
rect -13650 15970 -13640 15990
rect -13680 15960 -13640 15970
rect -13600 16470 -13560 16480
rect -13600 16450 -13590 16470
rect -13570 16450 -13560 16470
rect -13600 16310 -13560 16450
rect -13600 16290 -13590 16310
rect -13570 16290 -13560 16310
rect -13600 16150 -13560 16290
rect -13600 16130 -13590 16150
rect -13570 16130 -13560 16150
rect -13600 15990 -13560 16130
rect -13600 15970 -13590 15990
rect -13570 15970 -13560 15990
rect -13600 15960 -13560 15970
rect -13520 16470 -13480 16480
rect -13520 16450 -13510 16470
rect -13490 16450 -13480 16470
rect -13520 16310 -13480 16450
rect -13520 16290 -13510 16310
rect -13490 16290 -13480 16310
rect -13520 16150 -13480 16290
rect -13520 16130 -13510 16150
rect -13490 16130 -13480 16150
rect -13520 15990 -13480 16130
rect -13520 15970 -13510 15990
rect -13490 15970 -13480 15990
rect -13520 15960 -13480 15970
rect -13440 16470 -13400 16480
rect -13440 16450 -13430 16470
rect -13410 16450 -13400 16470
rect -13440 16310 -13400 16450
rect -13440 16290 -13430 16310
rect -13410 16290 -13400 16310
rect -13440 16150 -13400 16290
rect -13440 16130 -13430 16150
rect -13410 16130 -13400 16150
rect -13440 15990 -13400 16130
rect -13440 15970 -13430 15990
rect -13410 15970 -13400 15990
rect -13440 15960 -13400 15970
rect -13360 16470 -13320 16480
rect -13360 16450 -13350 16470
rect -13330 16450 -13320 16470
rect -13360 16310 -13320 16450
rect -13360 16290 -13350 16310
rect -13330 16290 -13320 16310
rect -13360 16150 -13320 16290
rect -13360 16130 -13350 16150
rect -13330 16130 -13320 16150
rect -13360 15990 -13320 16130
rect -13360 15970 -13350 15990
rect -13330 15970 -13320 15990
rect -13360 15960 -13320 15970
rect -13280 16470 -13240 16480
rect -13280 16450 -13270 16470
rect -13250 16450 -13240 16470
rect -13280 16310 -13240 16450
rect -13280 16290 -13270 16310
rect -13250 16290 -13240 16310
rect -13280 16150 -13240 16290
rect -13280 16130 -13270 16150
rect -13250 16130 -13240 16150
rect -13280 15990 -13240 16130
rect -13280 15970 -13270 15990
rect -13250 15970 -13240 15990
rect -13280 15960 -13240 15970
rect -13200 16470 -13160 16480
rect -13200 16450 -13190 16470
rect -13170 16450 -13160 16470
rect -13200 16310 -13160 16450
rect -13200 16290 -13190 16310
rect -13170 16290 -13160 16310
rect -13200 16150 -13160 16290
rect -13200 16130 -13190 16150
rect -13170 16130 -13160 16150
rect -13200 15990 -13160 16130
rect -13200 15970 -13190 15990
rect -13170 15970 -13160 15990
rect -13200 15960 -13160 15970
rect -13120 16470 -13080 16480
rect -13120 16450 -13110 16470
rect -13090 16450 -13080 16470
rect -13120 16310 -13080 16450
rect -13120 16290 -13110 16310
rect -13090 16290 -13080 16310
rect -13120 16150 -13080 16290
rect -13120 16130 -13110 16150
rect -13090 16130 -13080 16150
rect -13120 15990 -13080 16130
rect -13120 15970 -13110 15990
rect -13090 15970 -13080 15990
rect -13120 15960 -13080 15970
rect -13040 16470 -13000 16480
rect -13040 16450 -13030 16470
rect -13010 16450 -13000 16470
rect -13040 16310 -13000 16450
rect -13040 16290 -13030 16310
rect -13010 16290 -13000 16310
rect -13040 16150 -13000 16290
rect -13040 16130 -13030 16150
rect -13010 16130 -13000 16150
rect -13040 15990 -13000 16130
rect -13040 15970 -13030 15990
rect -13010 15970 -13000 15990
rect -13040 15960 -13000 15970
rect -12960 16470 -12920 16480
rect -12960 16450 -12950 16470
rect -12930 16450 -12920 16470
rect -12960 16310 -12920 16450
rect -12960 16290 -12950 16310
rect -12930 16290 -12920 16310
rect -12960 16150 -12920 16290
rect -12960 16130 -12950 16150
rect -12930 16130 -12920 16150
rect -12960 15990 -12920 16130
rect -12960 15970 -12950 15990
rect -12930 15970 -12920 15990
rect -12960 15960 -12920 15970
rect -12880 16470 -12840 16480
rect -12880 16450 -12870 16470
rect -12850 16450 -12840 16470
rect -12880 16310 -12840 16450
rect -12880 16290 -12870 16310
rect -12850 16290 -12840 16310
rect -12880 16150 -12840 16290
rect -12880 16130 -12870 16150
rect -12850 16130 -12840 16150
rect -12880 15990 -12840 16130
rect -12880 15970 -12870 15990
rect -12850 15970 -12840 15990
rect -12880 15960 -12840 15970
rect -12800 16470 -12760 16480
rect -12800 16450 -12790 16470
rect -12770 16450 -12760 16470
rect -12800 16310 -12760 16450
rect -12800 16290 -12790 16310
rect -12770 16290 -12760 16310
rect -12800 16150 -12760 16290
rect -12800 16130 -12790 16150
rect -12770 16130 -12760 16150
rect -12800 15990 -12760 16130
rect -12800 15970 -12790 15990
rect -12770 15970 -12760 15990
rect -12800 15960 -12760 15970
rect -12720 16470 -12680 16480
rect -12720 16450 -12710 16470
rect -12690 16450 -12680 16470
rect -12720 16310 -12680 16450
rect -12720 16290 -12710 16310
rect -12690 16290 -12680 16310
rect -12720 16150 -12680 16290
rect -12720 16130 -12710 16150
rect -12690 16130 -12680 16150
rect -12720 15990 -12680 16130
rect -12720 15970 -12710 15990
rect -12690 15970 -12680 15990
rect -12720 15960 -12680 15970
rect -12640 16470 -12600 16480
rect -12640 16450 -12630 16470
rect -12610 16450 -12600 16470
rect -12640 16310 -12600 16450
rect -12640 16290 -12630 16310
rect -12610 16290 -12600 16310
rect -12640 16150 -12600 16290
rect -12640 16130 -12630 16150
rect -12610 16130 -12600 16150
rect -12640 15990 -12600 16130
rect -12640 15970 -12630 15990
rect -12610 15970 -12600 15990
rect -12640 15960 -12600 15970
rect -12560 16470 -12520 16480
rect -12560 16450 -12550 16470
rect -12530 16450 -12520 16470
rect -12560 16310 -12520 16450
rect -12560 16290 -12550 16310
rect -12530 16290 -12520 16310
rect -12560 16150 -12520 16290
rect -12560 16130 -12550 16150
rect -12530 16130 -12520 16150
rect -12560 15990 -12520 16130
rect -12560 15970 -12550 15990
rect -12530 15970 -12520 15990
rect -12560 15960 -12520 15970
rect -12480 16470 -12440 16480
rect -12480 16450 -12470 16470
rect -12450 16450 -12440 16470
rect -12480 16310 -12440 16450
rect -12480 16290 -12470 16310
rect -12450 16290 -12440 16310
rect -12480 16150 -12440 16290
rect -12480 16130 -12470 16150
rect -12450 16130 -12440 16150
rect -12480 15990 -12440 16130
rect -12480 15970 -12470 15990
rect -12450 15970 -12440 15990
rect -12480 15960 -12440 15970
rect -12400 16470 -12360 16480
rect -12400 16450 -12390 16470
rect -12370 16450 -12360 16470
rect -12400 16310 -12360 16450
rect -12400 16290 -12390 16310
rect -12370 16290 -12360 16310
rect -12400 16150 -12360 16290
rect -12400 16130 -12390 16150
rect -12370 16130 -12360 16150
rect -12400 15990 -12360 16130
rect -12400 15970 -12390 15990
rect -12370 15970 -12360 15990
rect -12400 15960 -12360 15970
rect -12320 16470 -12280 16480
rect -12320 16450 -12310 16470
rect -12290 16450 -12280 16470
rect -12320 16310 -12280 16450
rect -12320 16290 -12310 16310
rect -12290 16290 -12280 16310
rect -12320 16150 -12280 16290
rect -12320 16130 -12310 16150
rect -12290 16130 -12280 16150
rect -12320 15990 -12280 16130
rect -12320 15970 -12310 15990
rect -12290 15970 -12280 15990
rect -12320 15960 -12280 15970
rect -12240 16470 -12200 16480
rect -12240 16450 -12230 16470
rect -12210 16450 -12200 16470
rect -12240 16310 -12200 16450
rect -12240 16290 -12230 16310
rect -12210 16290 -12200 16310
rect -12240 16150 -12200 16290
rect -12240 16130 -12230 16150
rect -12210 16130 -12200 16150
rect -12240 15990 -12200 16130
rect -12240 15970 -12230 15990
rect -12210 15970 -12200 15990
rect -12240 15960 -12200 15970
rect -12160 16470 -12120 16480
rect -12160 16450 -12150 16470
rect -12130 16450 -12120 16470
rect -12160 16310 -12120 16450
rect -12160 16290 -12150 16310
rect -12130 16290 -12120 16310
rect -12160 16150 -12120 16290
rect -12160 16130 -12150 16150
rect -12130 16130 -12120 16150
rect -12160 15990 -12120 16130
rect -12160 15970 -12150 15990
rect -12130 15970 -12120 15990
rect -12160 15960 -12120 15970
rect -12080 16470 -12040 16480
rect -12080 16450 -12070 16470
rect -12050 16450 -12040 16470
rect -12080 16310 -12040 16450
rect -12080 16290 -12070 16310
rect -12050 16290 -12040 16310
rect -12080 16150 -12040 16290
rect -12080 16130 -12070 16150
rect -12050 16130 -12040 16150
rect -12080 15990 -12040 16130
rect -12080 15970 -12070 15990
rect -12050 15970 -12040 15990
rect -12080 15960 -12040 15970
rect -12000 16470 -11960 16480
rect -12000 16450 -11990 16470
rect -11970 16450 -11960 16470
rect -12000 16310 -11960 16450
rect -12000 16290 -11990 16310
rect -11970 16290 -11960 16310
rect -12000 16150 -11960 16290
rect -12000 16130 -11990 16150
rect -11970 16130 -11960 16150
rect -12000 15990 -11960 16130
rect -12000 15970 -11990 15990
rect -11970 15970 -11960 15990
rect -12000 15960 -11960 15970
rect -11920 16470 -11880 16480
rect -11920 16450 -11910 16470
rect -11890 16450 -11880 16470
rect -11920 16310 -11880 16450
rect -11920 16290 -11910 16310
rect -11890 16290 -11880 16310
rect -11920 16150 -11880 16290
rect -11920 16130 -11910 16150
rect -11890 16130 -11880 16150
rect -11920 15990 -11880 16130
rect -11920 15970 -11910 15990
rect -11890 15970 -11880 15990
rect -11920 15960 -11880 15970
rect -11840 16470 -11800 16480
rect -11840 16450 -11830 16470
rect -11810 16450 -11800 16470
rect -11840 16310 -11800 16450
rect -11840 16290 -11830 16310
rect -11810 16290 -11800 16310
rect -11840 16150 -11800 16290
rect -11840 16130 -11830 16150
rect -11810 16130 -11800 16150
rect -11840 15990 -11800 16130
rect -11840 15970 -11830 15990
rect -11810 15970 -11800 15990
rect -11840 15960 -11800 15970
rect -11760 16470 -11720 16480
rect -11760 16450 -11750 16470
rect -11730 16450 -11720 16470
rect -11760 16310 -11720 16450
rect -11760 16290 -11750 16310
rect -11730 16290 -11720 16310
rect -11760 16150 -11720 16290
rect -11760 16130 -11750 16150
rect -11730 16130 -11720 16150
rect -11760 15990 -11720 16130
rect -11760 15970 -11750 15990
rect -11730 15970 -11720 15990
rect -11760 15960 -11720 15970
rect -11680 16470 -11640 16480
rect -11680 16450 -11670 16470
rect -11650 16450 -11640 16470
rect -11680 16310 -11640 16450
rect -11680 16290 -11670 16310
rect -11650 16290 -11640 16310
rect -11680 16150 -11640 16290
rect -11680 16130 -11670 16150
rect -11650 16130 -11640 16150
rect -11680 15990 -11640 16130
rect -11680 15970 -11670 15990
rect -11650 15970 -11640 15990
rect -11680 15960 -11640 15970
rect -11600 16470 -11560 16480
rect -11600 16450 -11590 16470
rect -11570 16450 -11560 16470
rect -11600 16310 -11560 16450
rect -11600 16290 -11590 16310
rect -11570 16290 -11560 16310
rect -11600 16150 -11560 16290
rect -11600 16130 -11590 16150
rect -11570 16130 -11560 16150
rect -11600 15990 -11560 16130
rect -11600 15970 -11590 15990
rect -11570 15970 -11560 15990
rect -11600 15960 -11560 15970
rect -11520 16470 -11480 16480
rect -11520 16450 -11510 16470
rect -11490 16450 -11480 16470
rect -11520 16310 -11480 16450
rect -11520 16290 -11510 16310
rect -11490 16290 -11480 16310
rect -11520 16150 -11480 16290
rect -11520 16130 -11510 16150
rect -11490 16130 -11480 16150
rect -11520 15990 -11480 16130
rect -11520 15970 -11510 15990
rect -11490 15970 -11480 15990
rect -11520 15960 -11480 15970
rect -11440 16470 -11400 16480
rect -11440 16450 -11430 16470
rect -11410 16450 -11400 16470
rect -11440 16310 -11400 16450
rect -11440 16290 -11430 16310
rect -11410 16290 -11400 16310
rect -11440 16150 -11400 16290
rect -11440 16130 -11430 16150
rect -11410 16130 -11400 16150
rect -11440 15990 -11400 16130
rect -11440 15970 -11430 15990
rect -11410 15970 -11400 15990
rect -11440 15960 -11400 15970
rect -11360 16470 -11320 16480
rect -11360 16450 -11350 16470
rect -11330 16450 -11320 16470
rect -11360 16310 -11320 16450
rect -11360 16290 -11350 16310
rect -11330 16290 -11320 16310
rect -11360 16150 -11320 16290
rect -11360 16130 -11350 16150
rect -11330 16130 -11320 16150
rect -11360 15990 -11320 16130
rect -11360 15970 -11350 15990
rect -11330 15970 -11320 15990
rect -11360 15960 -11320 15970
rect -11280 16470 -11240 16480
rect -11280 16450 -11270 16470
rect -11250 16450 -11240 16470
rect -11280 16310 -11240 16450
rect -11280 16290 -11270 16310
rect -11250 16290 -11240 16310
rect -11280 16150 -11240 16290
rect -11280 16130 -11270 16150
rect -11250 16130 -11240 16150
rect -11280 15990 -11240 16130
rect -11280 15970 -11270 15990
rect -11250 15970 -11240 15990
rect -11280 15960 -11240 15970
rect -11200 16470 -11160 16480
rect -11200 16450 -11190 16470
rect -11170 16450 -11160 16470
rect -11200 16310 -11160 16450
rect -11200 16290 -11190 16310
rect -11170 16290 -11160 16310
rect -11200 16150 -11160 16290
rect -11200 16130 -11190 16150
rect -11170 16130 -11160 16150
rect -11200 15990 -11160 16130
rect -11200 15970 -11190 15990
rect -11170 15970 -11160 15990
rect -11200 15960 -11160 15970
rect -11120 16470 -11080 16480
rect -11120 16450 -11110 16470
rect -11090 16450 -11080 16470
rect -11120 16310 -11080 16450
rect -11120 16290 -11110 16310
rect -11090 16290 -11080 16310
rect -11120 16150 -11080 16290
rect -11120 16130 -11110 16150
rect -11090 16130 -11080 16150
rect -11120 15990 -11080 16130
rect -11120 15970 -11110 15990
rect -11090 15970 -11080 15990
rect -11120 15960 -11080 15970
rect -11040 16470 -11000 16480
rect -11040 16450 -11030 16470
rect -11010 16450 -11000 16470
rect -11040 16310 -11000 16450
rect -11040 16290 -11030 16310
rect -11010 16290 -11000 16310
rect -11040 16150 -11000 16290
rect -11040 16130 -11030 16150
rect -11010 16130 -11000 16150
rect -11040 15990 -11000 16130
rect -11040 15970 -11030 15990
rect -11010 15970 -11000 15990
rect -11040 15960 -11000 15970
rect -10960 16470 -10920 16480
rect -10960 16450 -10950 16470
rect -10930 16450 -10920 16470
rect -10960 16310 -10920 16450
rect -10960 16290 -10950 16310
rect -10930 16290 -10920 16310
rect -10960 16150 -10920 16290
rect -10960 16130 -10950 16150
rect -10930 16130 -10920 16150
rect -10960 15990 -10920 16130
rect -10960 15970 -10950 15990
rect -10930 15970 -10920 15990
rect -10960 15960 -10920 15970
rect -10880 16470 -10840 16480
rect -10880 16450 -10870 16470
rect -10850 16450 -10840 16470
rect -10880 16310 -10840 16450
rect -10880 16290 -10870 16310
rect -10850 16290 -10840 16310
rect -10880 16150 -10840 16290
rect -10880 16130 -10870 16150
rect -10850 16130 -10840 16150
rect -10880 15990 -10840 16130
rect -10880 15970 -10870 15990
rect -10850 15970 -10840 15990
rect -10880 15960 -10840 15970
rect -10800 16470 -10760 16480
rect -10800 16450 -10790 16470
rect -10770 16450 -10760 16470
rect -10800 16310 -10760 16450
rect -10800 16290 -10790 16310
rect -10770 16290 -10760 16310
rect -10800 16150 -10760 16290
rect -10800 16130 -10790 16150
rect -10770 16130 -10760 16150
rect -10800 15990 -10760 16130
rect -10800 15970 -10790 15990
rect -10770 15970 -10760 15990
rect -10800 15960 -10760 15970
rect -10720 16470 -10680 16480
rect -10720 16450 -10710 16470
rect -10690 16450 -10680 16470
rect -10720 16310 -10680 16450
rect -10720 16290 -10710 16310
rect -10690 16290 -10680 16310
rect -10720 16150 -10680 16290
rect -10720 16130 -10710 16150
rect -10690 16130 -10680 16150
rect -10720 15990 -10680 16130
rect -10720 15970 -10710 15990
rect -10690 15970 -10680 15990
rect -10720 15960 -10680 15970
rect -10640 16470 -10600 16480
rect -10640 16450 -10630 16470
rect -10610 16450 -10600 16470
rect -10640 16310 -10600 16450
rect -10640 16290 -10630 16310
rect -10610 16290 -10600 16310
rect -10640 16150 -10600 16290
rect -10640 16130 -10630 16150
rect -10610 16130 -10600 16150
rect -10640 15990 -10600 16130
rect -10640 15970 -10630 15990
rect -10610 15970 -10600 15990
rect -10640 15960 -10600 15970
rect -10560 16470 -10520 16480
rect -10560 16450 -10550 16470
rect -10530 16450 -10520 16470
rect -10560 16310 -10520 16450
rect -10560 16290 -10550 16310
rect -10530 16290 -10520 16310
rect -10560 16150 -10520 16290
rect -10560 16130 -10550 16150
rect -10530 16130 -10520 16150
rect -10560 15990 -10520 16130
rect -10560 15970 -10550 15990
rect -10530 15970 -10520 15990
rect -10560 15960 -10520 15970
rect -10480 16470 -10440 16480
rect -10480 16450 -10470 16470
rect -10450 16450 -10440 16470
rect -10480 16310 -10440 16450
rect -10480 16290 -10470 16310
rect -10450 16290 -10440 16310
rect -10480 16150 -10440 16290
rect -10480 16130 -10470 16150
rect -10450 16130 -10440 16150
rect -10480 15990 -10440 16130
rect -10480 15970 -10470 15990
rect -10450 15970 -10440 15990
rect -10480 15960 -10440 15970
rect -10400 16470 -10360 16480
rect -10400 16450 -10390 16470
rect -10370 16450 -10360 16470
rect -10400 16310 -10360 16450
rect -10400 16290 -10390 16310
rect -10370 16290 -10360 16310
rect -10400 16150 -10360 16290
rect -10400 16130 -10390 16150
rect -10370 16130 -10360 16150
rect -10400 15990 -10360 16130
rect -10400 15970 -10390 15990
rect -10370 15970 -10360 15990
rect -10400 15960 -10360 15970
rect -10320 16470 -10280 16480
rect -10320 16450 -10310 16470
rect -10290 16450 -10280 16470
rect -10320 16310 -10280 16450
rect -10320 16290 -10310 16310
rect -10290 16290 -10280 16310
rect -10320 16150 -10280 16290
rect -10320 16130 -10310 16150
rect -10290 16130 -10280 16150
rect -10320 15990 -10280 16130
rect -10320 15970 -10310 15990
rect -10290 15970 -10280 15990
rect -10320 15960 -10280 15970
rect -10240 16470 -10200 16480
rect -10240 16450 -10230 16470
rect -10210 16450 -10200 16470
rect -10240 16310 -10200 16450
rect -10240 16290 -10230 16310
rect -10210 16290 -10200 16310
rect -10240 16150 -10200 16290
rect -10240 16130 -10230 16150
rect -10210 16130 -10200 16150
rect -10240 15990 -10200 16130
rect -10240 15970 -10230 15990
rect -10210 15970 -10200 15990
rect -10240 15960 -10200 15970
rect -10160 16470 -10120 16480
rect -10160 16450 -10150 16470
rect -10130 16450 -10120 16470
rect -10160 16310 -10120 16450
rect -10160 16290 -10150 16310
rect -10130 16290 -10120 16310
rect -10160 16150 -10120 16290
rect -10160 16130 -10150 16150
rect -10130 16130 -10120 16150
rect -10160 15990 -10120 16130
rect -10160 15970 -10150 15990
rect -10130 15970 -10120 15990
rect -10160 15960 -10120 15970
rect -10080 16470 -10040 16480
rect -10080 16450 -10070 16470
rect -10050 16450 -10040 16470
rect -10080 16310 -10040 16450
rect -10080 16290 -10070 16310
rect -10050 16290 -10040 16310
rect -10080 16150 -10040 16290
rect -10080 16130 -10070 16150
rect -10050 16130 -10040 16150
rect -10080 15990 -10040 16130
rect -10080 15970 -10070 15990
rect -10050 15970 -10040 15990
rect -10080 15960 -10040 15970
rect -10000 16470 -9960 16480
rect -10000 16450 -9990 16470
rect -9970 16450 -9960 16470
rect -10000 16310 -9960 16450
rect -10000 16290 -9990 16310
rect -9970 16290 -9960 16310
rect -10000 16150 -9960 16290
rect -10000 16130 -9990 16150
rect -9970 16130 -9960 16150
rect -10000 15990 -9960 16130
rect -10000 15970 -9990 15990
rect -9970 15970 -9960 15990
rect -10000 15960 -9960 15970
rect -9920 16470 -9880 16480
rect -9920 16450 -9910 16470
rect -9890 16450 -9880 16470
rect -9920 16310 -9880 16450
rect -9920 16290 -9910 16310
rect -9890 16290 -9880 16310
rect -9920 16150 -9880 16290
rect -9920 16130 -9910 16150
rect -9890 16130 -9880 16150
rect -9920 15990 -9880 16130
rect -9920 15970 -9910 15990
rect -9890 15970 -9880 15990
rect -9920 15960 -9880 15970
rect -9840 16470 -9800 16480
rect -9840 16450 -9830 16470
rect -9810 16450 -9800 16470
rect -9840 16310 -9800 16450
rect -9840 16290 -9830 16310
rect -9810 16290 -9800 16310
rect -9840 16150 -9800 16290
rect -9840 16130 -9830 16150
rect -9810 16130 -9800 16150
rect -9840 15990 -9800 16130
rect -9840 15970 -9830 15990
rect -9810 15970 -9800 15990
rect -9840 15960 -9800 15970
rect -9760 16470 -9720 16480
rect -9760 16450 -9750 16470
rect -9730 16450 -9720 16470
rect -9760 16310 -9720 16450
rect -9760 16290 -9750 16310
rect -9730 16290 -9720 16310
rect -9760 16150 -9720 16290
rect -9760 16130 -9750 16150
rect -9730 16130 -9720 16150
rect -9760 15990 -9720 16130
rect -9760 15970 -9750 15990
rect -9730 15970 -9720 15990
rect -9760 15960 -9720 15970
rect -9680 16470 -9640 16480
rect -9680 16450 -9670 16470
rect -9650 16450 -9640 16470
rect -9680 16310 -9640 16450
rect -9680 16290 -9670 16310
rect -9650 16290 -9640 16310
rect -9680 16150 -9640 16290
rect -9680 16130 -9670 16150
rect -9650 16130 -9640 16150
rect -9680 15990 -9640 16130
rect -9680 15970 -9670 15990
rect -9650 15970 -9640 15990
rect -9680 15960 -9640 15970
rect -9600 16470 -9560 16480
rect -9600 16450 -9590 16470
rect -9570 16450 -9560 16470
rect -9600 16310 -9560 16450
rect -9600 16290 -9590 16310
rect -9570 16290 -9560 16310
rect -9600 16150 -9560 16290
rect -9600 16130 -9590 16150
rect -9570 16130 -9560 16150
rect -9600 15990 -9560 16130
rect -9600 15970 -9590 15990
rect -9570 15970 -9560 15990
rect -9600 15960 -9560 15970
rect -9520 16470 -9480 16480
rect -9520 16450 -9510 16470
rect -9490 16450 -9480 16470
rect -9520 16310 -9480 16450
rect -9520 16290 -9510 16310
rect -9490 16290 -9480 16310
rect -9520 16150 -9480 16290
rect -9520 16130 -9510 16150
rect -9490 16130 -9480 16150
rect -9520 15990 -9480 16130
rect -9520 15970 -9510 15990
rect -9490 15970 -9480 15990
rect -9520 15960 -9480 15970
rect -9440 16470 -9400 16480
rect -9440 16450 -9430 16470
rect -9410 16450 -9400 16470
rect -9440 16310 -9400 16450
rect -9440 16290 -9430 16310
rect -9410 16290 -9400 16310
rect -9440 16150 -9400 16290
rect -9440 16130 -9430 16150
rect -9410 16130 -9400 16150
rect -9440 15990 -9400 16130
rect -9440 15970 -9430 15990
rect -9410 15970 -9400 15990
rect -9440 15960 -9400 15970
rect -9360 16470 -9320 16480
rect -9360 16450 -9350 16470
rect -9330 16450 -9320 16470
rect -9360 16310 -9320 16450
rect -9360 16290 -9350 16310
rect -9330 16290 -9320 16310
rect -9360 16150 -9320 16290
rect -9360 16130 -9350 16150
rect -9330 16130 -9320 16150
rect -9360 15990 -9320 16130
rect -9360 15970 -9350 15990
rect -9330 15970 -9320 15990
rect -9360 15960 -9320 15970
rect -9280 16470 -9240 16480
rect -9280 16450 -9270 16470
rect -9250 16450 -9240 16470
rect -9280 16310 -9240 16450
rect -9280 16290 -9270 16310
rect -9250 16290 -9240 16310
rect -9280 16150 -9240 16290
rect -9280 16130 -9270 16150
rect -9250 16130 -9240 16150
rect -9280 15990 -9240 16130
rect -9280 15970 -9270 15990
rect -9250 15970 -9240 15990
rect -9280 15960 -9240 15970
rect -9200 16470 -9160 16480
rect -9200 16450 -9190 16470
rect -9170 16450 -9160 16470
rect -9200 16310 -9160 16450
rect -9200 16290 -9190 16310
rect -9170 16290 -9160 16310
rect -9200 16150 -9160 16290
rect -9200 16130 -9190 16150
rect -9170 16130 -9160 16150
rect -9200 15990 -9160 16130
rect -9200 15970 -9190 15990
rect -9170 15970 -9160 15990
rect -9200 15960 -9160 15970
rect -9120 16470 -9080 16480
rect -9120 16450 -9110 16470
rect -9090 16450 -9080 16470
rect -9120 16310 -9080 16450
rect -9120 16290 -9110 16310
rect -9090 16290 -9080 16310
rect -9120 16150 -9080 16290
rect -9120 16130 -9110 16150
rect -9090 16130 -9080 16150
rect -9120 15990 -9080 16130
rect -9120 15970 -9110 15990
rect -9090 15970 -9080 15990
rect -9120 15960 -9080 15970
rect -9040 16470 -9000 16480
rect -9040 16450 -9030 16470
rect -9010 16450 -9000 16470
rect -9040 16310 -9000 16450
rect -9040 16290 -9030 16310
rect -9010 16290 -9000 16310
rect -9040 16150 -9000 16290
rect -9040 16130 -9030 16150
rect -9010 16130 -9000 16150
rect -9040 15990 -9000 16130
rect -9040 15970 -9030 15990
rect -9010 15970 -9000 15990
rect -9040 15960 -9000 15970
rect -8960 16470 -8920 16480
rect -8960 16450 -8950 16470
rect -8930 16450 -8920 16470
rect -8960 16310 -8920 16450
rect -8960 16290 -8950 16310
rect -8930 16290 -8920 16310
rect -8960 16150 -8920 16290
rect -8960 16130 -8950 16150
rect -8930 16130 -8920 16150
rect -8960 15990 -8920 16130
rect -8960 15970 -8950 15990
rect -8930 15970 -8920 15990
rect -8960 15960 -8920 15970
rect -8880 16470 -8840 16480
rect -8880 16450 -8870 16470
rect -8850 16450 -8840 16470
rect -8880 16310 -8840 16450
rect -8880 16290 -8870 16310
rect -8850 16290 -8840 16310
rect -8880 16150 -8840 16290
rect -8880 16130 -8870 16150
rect -8850 16130 -8840 16150
rect -8880 15990 -8840 16130
rect -8880 15970 -8870 15990
rect -8850 15970 -8840 15990
rect -8880 15960 -8840 15970
rect -8800 16470 -8760 16480
rect -8800 16450 -8790 16470
rect -8770 16450 -8760 16470
rect -8800 16310 -8760 16450
rect -8800 16290 -8790 16310
rect -8770 16290 -8760 16310
rect -8800 16150 -8760 16290
rect -8800 16130 -8790 16150
rect -8770 16130 -8760 16150
rect -8800 15990 -8760 16130
rect -8800 15970 -8790 15990
rect -8770 15970 -8760 15990
rect -8800 15960 -8760 15970
rect -8720 16470 -8680 16480
rect -8720 16450 -8710 16470
rect -8690 16450 -8680 16470
rect -8720 16310 -8680 16450
rect -8720 16290 -8710 16310
rect -8690 16290 -8680 16310
rect -8720 16150 -8680 16290
rect -8720 16130 -8710 16150
rect -8690 16130 -8680 16150
rect -8720 15990 -8680 16130
rect -8720 15970 -8710 15990
rect -8690 15970 -8680 15990
rect -8720 15960 -8680 15970
rect -8640 16470 -8600 16480
rect -8640 16450 -8630 16470
rect -8610 16450 -8600 16470
rect -8640 16310 -8600 16450
rect -8640 16290 -8630 16310
rect -8610 16290 -8600 16310
rect -8640 16150 -8600 16290
rect -8640 16130 -8630 16150
rect -8610 16130 -8600 16150
rect -8640 15990 -8600 16130
rect -8640 15970 -8630 15990
rect -8610 15970 -8600 15990
rect -8640 15960 -8600 15970
rect -8560 16470 -8520 16480
rect -8560 16450 -8550 16470
rect -8530 16450 -8520 16470
rect -8560 16310 -8520 16450
rect -8560 16290 -8550 16310
rect -8530 16290 -8520 16310
rect -8560 16150 -8520 16290
rect -8560 16130 -8550 16150
rect -8530 16130 -8520 16150
rect -8560 15990 -8520 16130
rect -8560 15970 -8550 15990
rect -8530 15970 -8520 15990
rect -8560 15960 -8520 15970
rect -8480 16470 -8440 16480
rect -8480 16450 -8470 16470
rect -8450 16450 -8440 16470
rect -8480 16310 -8440 16450
rect -8480 16290 -8470 16310
rect -8450 16290 -8440 16310
rect -8480 16150 -8440 16290
rect -8480 16130 -8470 16150
rect -8450 16130 -8440 16150
rect -8480 15990 -8440 16130
rect -8480 15970 -8470 15990
rect -8450 15970 -8440 15990
rect -8480 15960 -8440 15970
rect -8400 16470 -8360 16480
rect -8400 16450 -8390 16470
rect -8370 16450 -8360 16470
rect -8400 16310 -8360 16450
rect -8400 16290 -8390 16310
rect -8370 16290 -8360 16310
rect -8400 16150 -8360 16290
rect -8400 16130 -8390 16150
rect -8370 16130 -8360 16150
rect -8400 15990 -8360 16130
rect -8400 15970 -8390 15990
rect -8370 15970 -8360 15990
rect -8400 15960 -8360 15970
rect -8320 16470 -8280 16480
rect -8320 16450 -8310 16470
rect -8290 16450 -8280 16470
rect -8320 16310 -8280 16450
rect -8320 16290 -8310 16310
rect -8290 16290 -8280 16310
rect -8320 16150 -8280 16290
rect -8320 16130 -8310 16150
rect -8290 16130 -8280 16150
rect -8320 15990 -8280 16130
rect -8320 15970 -8310 15990
rect -8290 15970 -8280 15990
rect -8320 15960 -8280 15970
rect -8240 16470 -8200 16480
rect -8240 16450 -8230 16470
rect -8210 16450 -8200 16470
rect -8240 16310 -8200 16450
rect -8240 16290 -8230 16310
rect -8210 16290 -8200 16310
rect -8240 16150 -8200 16290
rect -8240 16130 -8230 16150
rect -8210 16130 -8200 16150
rect -8240 15990 -8200 16130
rect -8240 15970 -8230 15990
rect -8210 15970 -8200 15990
rect -8240 15960 -8200 15970
rect -8160 16470 -8120 16480
rect -8160 16450 -8150 16470
rect -8130 16450 -8120 16470
rect -8160 16310 -8120 16450
rect -8160 16290 -8150 16310
rect -8130 16290 -8120 16310
rect -8160 16150 -8120 16290
rect -8160 16130 -8150 16150
rect -8130 16130 -8120 16150
rect -8160 15990 -8120 16130
rect -8160 15970 -8150 15990
rect -8130 15970 -8120 15990
rect -8160 15960 -8120 15970
rect -8080 16470 -8040 16480
rect -8080 16450 -8070 16470
rect -8050 16450 -8040 16470
rect -8080 16310 -8040 16450
rect -8080 16290 -8070 16310
rect -8050 16290 -8040 16310
rect -8080 16150 -8040 16290
rect -8080 16130 -8070 16150
rect -8050 16130 -8040 16150
rect -8080 15990 -8040 16130
rect -8080 15970 -8070 15990
rect -8050 15970 -8040 15990
rect -8080 15960 -8040 15970
rect -8000 16470 -7960 16480
rect -8000 16450 -7990 16470
rect -7970 16450 -7960 16470
rect -8000 16310 -7960 16450
rect -8000 16290 -7990 16310
rect -7970 16290 -7960 16310
rect -8000 16150 -7960 16290
rect -8000 16130 -7990 16150
rect -7970 16130 -7960 16150
rect -8000 15990 -7960 16130
rect -8000 15970 -7990 15990
rect -7970 15970 -7960 15990
rect -8000 15960 -7960 15970
rect -7920 16470 -7880 16480
rect -7920 16450 -7910 16470
rect -7890 16450 -7880 16470
rect -7920 16310 -7880 16450
rect -7920 16290 -7910 16310
rect -7890 16290 -7880 16310
rect -7920 16150 -7880 16290
rect -7920 16130 -7910 16150
rect -7890 16130 -7880 16150
rect -7920 15990 -7880 16130
rect -7920 15970 -7910 15990
rect -7890 15970 -7880 15990
rect -7920 15960 -7880 15970
rect -7840 16470 -7800 16480
rect -7840 16450 -7830 16470
rect -7810 16450 -7800 16470
rect -7840 16310 -7800 16450
rect -7840 16290 -7830 16310
rect -7810 16290 -7800 16310
rect -7840 16150 -7800 16290
rect -7840 16130 -7830 16150
rect -7810 16130 -7800 16150
rect -7840 15990 -7800 16130
rect -7840 15970 -7830 15990
rect -7810 15970 -7800 15990
rect -7840 15960 -7800 15970
rect -7760 16470 -7720 16480
rect -7760 16450 -7750 16470
rect -7730 16450 -7720 16470
rect -7760 16310 -7720 16450
rect -7760 16290 -7750 16310
rect -7730 16290 -7720 16310
rect -7760 16150 -7720 16290
rect -7760 16130 -7750 16150
rect -7730 16130 -7720 16150
rect -7760 15990 -7720 16130
rect -7760 15970 -7750 15990
rect -7730 15970 -7720 15990
rect -7760 15960 -7720 15970
rect -7680 16470 -7640 16480
rect -7680 16450 -7670 16470
rect -7650 16450 -7640 16470
rect -7680 16310 -7640 16450
rect -7680 16290 -7670 16310
rect -7650 16290 -7640 16310
rect -7680 16150 -7640 16290
rect -7680 16130 -7670 16150
rect -7650 16130 -7640 16150
rect -7680 15990 -7640 16130
rect -7680 15970 -7670 15990
rect -7650 15970 -7640 15990
rect -7680 15960 -7640 15970
rect -7600 16470 -7560 16480
rect -7600 16450 -7590 16470
rect -7570 16450 -7560 16470
rect -7600 16310 -7560 16450
rect -7600 16290 -7590 16310
rect -7570 16290 -7560 16310
rect -7600 16150 -7560 16290
rect -7600 16130 -7590 16150
rect -7570 16130 -7560 16150
rect -7600 15990 -7560 16130
rect -7600 15970 -7590 15990
rect -7570 15970 -7560 15990
rect -7600 15960 -7560 15970
rect -7520 16470 -7480 16480
rect -7520 16450 -7510 16470
rect -7490 16450 -7480 16470
rect -7520 16310 -7480 16450
rect -7520 16290 -7510 16310
rect -7490 16290 -7480 16310
rect -7520 16150 -7480 16290
rect -7520 16130 -7510 16150
rect -7490 16130 -7480 16150
rect -7520 15990 -7480 16130
rect -7520 15970 -7510 15990
rect -7490 15970 -7480 15990
rect -7520 15960 -7480 15970
rect -7440 16470 -7400 16480
rect -7440 16450 -7430 16470
rect -7410 16450 -7400 16470
rect -7440 16310 -7400 16450
rect -7440 16290 -7430 16310
rect -7410 16290 -7400 16310
rect -7440 16150 -7400 16290
rect -7440 16130 -7430 16150
rect -7410 16130 -7400 16150
rect -7440 15990 -7400 16130
rect -7440 15970 -7430 15990
rect -7410 15970 -7400 15990
rect -7440 15960 -7400 15970
rect -7360 16470 -7320 16480
rect -7360 16450 -7350 16470
rect -7330 16450 -7320 16470
rect -7360 16310 -7320 16450
rect -7360 16290 -7350 16310
rect -7330 16290 -7320 16310
rect -7360 16150 -7320 16290
rect -7360 16130 -7350 16150
rect -7330 16130 -7320 16150
rect -7360 15990 -7320 16130
rect -7360 15970 -7350 15990
rect -7330 15970 -7320 15990
rect -7360 15960 -7320 15970
rect -7280 16470 -7240 16480
rect -7280 16450 -7270 16470
rect -7250 16450 -7240 16470
rect -7280 16310 -7240 16450
rect -7280 16290 -7270 16310
rect -7250 16290 -7240 16310
rect -7280 16150 -7240 16290
rect -7280 16130 -7270 16150
rect -7250 16130 -7240 16150
rect -7280 15990 -7240 16130
rect -7280 15970 -7270 15990
rect -7250 15970 -7240 15990
rect -7280 15960 -7240 15970
rect -7200 16470 -7160 16480
rect -7200 16450 -7190 16470
rect -7170 16450 -7160 16470
rect -7200 16310 -7160 16450
rect -7200 16290 -7190 16310
rect -7170 16290 -7160 16310
rect -7200 16150 -7160 16290
rect -7200 16130 -7190 16150
rect -7170 16130 -7160 16150
rect -7200 15990 -7160 16130
rect -7200 15970 -7190 15990
rect -7170 15970 -7160 15990
rect -7200 15960 -7160 15970
rect -7120 16470 -7080 16480
rect -7120 16450 -7110 16470
rect -7090 16450 -7080 16470
rect -7120 16310 -7080 16450
rect -7120 16290 -7110 16310
rect -7090 16290 -7080 16310
rect -7120 16150 -7080 16290
rect -7120 16130 -7110 16150
rect -7090 16130 -7080 16150
rect -7120 15990 -7080 16130
rect -7120 15970 -7110 15990
rect -7090 15970 -7080 15990
rect -7120 15960 -7080 15970
rect -7040 16470 -7000 16480
rect -7040 16450 -7030 16470
rect -7010 16450 -7000 16470
rect -7040 16310 -7000 16450
rect -7040 16290 -7030 16310
rect -7010 16290 -7000 16310
rect -7040 16150 -7000 16290
rect -7040 16130 -7030 16150
rect -7010 16130 -7000 16150
rect -7040 15990 -7000 16130
rect -7040 15970 -7030 15990
rect -7010 15970 -7000 15990
rect -7040 15960 -7000 15970
rect -6960 16470 -6920 16480
rect -6960 16450 -6950 16470
rect -6930 16450 -6920 16470
rect -6960 16310 -6920 16450
rect -6960 16290 -6950 16310
rect -6930 16290 -6920 16310
rect -6960 16150 -6920 16290
rect -6960 16130 -6950 16150
rect -6930 16130 -6920 16150
rect -6960 15990 -6920 16130
rect -6960 15970 -6950 15990
rect -6930 15970 -6920 15990
rect -6960 15960 -6920 15970
rect -6880 16470 -6840 16480
rect -6880 16450 -6870 16470
rect -6850 16450 -6840 16470
rect -6880 16310 -6840 16450
rect -6880 16290 -6870 16310
rect -6850 16290 -6840 16310
rect -6880 16150 -6840 16290
rect -6880 16130 -6870 16150
rect -6850 16130 -6840 16150
rect -6880 15990 -6840 16130
rect -6880 15970 -6870 15990
rect -6850 15970 -6840 15990
rect -6880 15960 -6840 15970
rect -6800 16470 -6760 16480
rect -6800 16450 -6790 16470
rect -6770 16450 -6760 16470
rect -6800 16310 -6760 16450
rect -6800 16290 -6790 16310
rect -6770 16290 -6760 16310
rect -6800 16150 -6760 16290
rect -6800 16130 -6790 16150
rect -6770 16130 -6760 16150
rect -6800 15990 -6760 16130
rect -6800 15970 -6790 15990
rect -6770 15970 -6760 15990
rect -6800 15960 -6760 15970
rect -6720 16470 -6680 16480
rect -6720 16450 -6710 16470
rect -6690 16450 -6680 16470
rect -6720 16310 -6680 16450
rect -6720 16290 -6710 16310
rect -6690 16290 -6680 16310
rect -6720 16150 -6680 16290
rect -6720 16130 -6710 16150
rect -6690 16130 -6680 16150
rect -6720 15990 -6680 16130
rect -6720 15970 -6710 15990
rect -6690 15970 -6680 15990
rect -6720 15960 -6680 15970
rect -6640 16470 -6600 16480
rect -6640 16450 -6630 16470
rect -6610 16450 -6600 16470
rect -6640 16310 -6600 16450
rect -6640 16290 -6630 16310
rect -6610 16290 -6600 16310
rect -6640 16150 -6600 16290
rect -6640 16130 -6630 16150
rect -6610 16130 -6600 16150
rect -6640 15990 -6600 16130
rect -6640 15970 -6630 15990
rect -6610 15970 -6600 15990
rect -6640 15960 -6600 15970
rect -6560 16470 -6520 16480
rect -6560 16450 -6550 16470
rect -6530 16450 -6520 16470
rect -6560 16310 -6520 16450
rect -6560 16290 -6550 16310
rect -6530 16290 -6520 16310
rect -6560 16150 -6520 16290
rect -6560 16130 -6550 16150
rect -6530 16130 -6520 16150
rect -6560 15990 -6520 16130
rect -6560 15970 -6550 15990
rect -6530 15970 -6520 15990
rect -6560 15960 -6520 15970
rect -6480 16470 -6440 16480
rect -6480 16450 -6470 16470
rect -6450 16450 -6440 16470
rect -6480 16310 -6440 16450
rect -6480 16290 -6470 16310
rect -6450 16290 -6440 16310
rect -6480 16150 -6440 16290
rect -6480 16130 -6470 16150
rect -6450 16130 -6440 16150
rect -6480 15990 -6440 16130
rect -6480 15970 -6470 15990
rect -6450 15970 -6440 15990
rect -6480 15960 -6440 15970
rect -6400 16470 -6360 16480
rect -6400 16450 -6390 16470
rect -6370 16450 -6360 16470
rect -6400 16310 -6360 16450
rect -6400 16290 -6390 16310
rect -6370 16290 -6360 16310
rect -6400 16150 -6360 16290
rect -6400 16130 -6390 16150
rect -6370 16130 -6360 16150
rect -6400 15990 -6360 16130
rect -6400 15970 -6390 15990
rect -6370 15970 -6360 15990
rect -6400 15960 -6360 15970
rect -6320 16470 -6280 16480
rect -6320 16450 -6310 16470
rect -6290 16450 -6280 16470
rect -6320 16310 -6280 16450
rect -6320 16290 -6310 16310
rect -6290 16290 -6280 16310
rect -6320 16150 -6280 16290
rect -6320 16130 -6310 16150
rect -6290 16130 -6280 16150
rect -6320 15990 -6280 16130
rect -6320 15970 -6310 15990
rect -6290 15970 -6280 15990
rect -6320 15960 -6280 15970
rect -6240 16470 -6200 16480
rect -6240 16450 -6230 16470
rect -6210 16450 -6200 16470
rect -6240 16310 -6200 16450
rect -6240 16290 -6230 16310
rect -6210 16290 -6200 16310
rect -6240 16150 -6200 16290
rect -6240 16130 -6230 16150
rect -6210 16130 -6200 16150
rect -6240 15990 -6200 16130
rect -6240 15970 -6230 15990
rect -6210 15970 -6200 15990
rect -6240 15960 -6200 15970
rect -6160 16470 -6120 16480
rect -6160 16450 -6150 16470
rect -6130 16450 -6120 16470
rect -6160 16310 -6120 16450
rect -6160 16290 -6150 16310
rect -6130 16290 -6120 16310
rect -6160 16150 -6120 16290
rect -6160 16130 -6150 16150
rect -6130 16130 -6120 16150
rect -6160 15990 -6120 16130
rect -6160 15970 -6150 15990
rect -6130 15970 -6120 15990
rect -6160 15960 -6120 15970
rect -6080 16470 -6040 16480
rect -6080 16450 -6070 16470
rect -6050 16450 -6040 16470
rect -6080 16310 -6040 16450
rect -6080 16290 -6070 16310
rect -6050 16290 -6040 16310
rect -6080 16150 -6040 16290
rect -6080 16130 -6070 16150
rect -6050 16130 -6040 16150
rect -6080 15990 -6040 16130
rect -6080 15970 -6070 15990
rect -6050 15970 -6040 15990
rect -6080 15960 -6040 15970
rect -6000 16470 -5960 16480
rect -6000 16450 -5990 16470
rect -5970 16450 -5960 16470
rect -6000 16310 -5960 16450
rect -6000 16290 -5990 16310
rect -5970 16290 -5960 16310
rect -6000 16150 -5960 16290
rect -6000 16130 -5990 16150
rect -5970 16130 -5960 16150
rect -6000 15990 -5960 16130
rect -6000 15970 -5990 15990
rect -5970 15970 -5960 15990
rect -6000 15960 -5960 15970
rect -5920 16470 -5880 16480
rect -5920 16450 -5910 16470
rect -5890 16450 -5880 16470
rect -5920 16310 -5880 16450
rect -5920 16290 -5910 16310
rect -5890 16290 -5880 16310
rect -5920 16150 -5880 16290
rect -5920 16130 -5910 16150
rect -5890 16130 -5880 16150
rect -5920 15990 -5880 16130
rect -5920 15970 -5910 15990
rect -5890 15970 -5880 15990
rect -5920 15960 -5880 15970
rect -5840 16470 -5800 16480
rect -5840 16450 -5830 16470
rect -5810 16450 -5800 16470
rect -5840 16310 -5800 16450
rect -5840 16290 -5830 16310
rect -5810 16290 -5800 16310
rect -5840 16150 -5800 16290
rect -5840 16130 -5830 16150
rect -5810 16130 -5800 16150
rect -5840 15990 -5800 16130
rect -5840 15970 -5830 15990
rect -5810 15970 -5800 15990
rect -5840 15960 -5800 15970
rect -5760 16470 -5720 16480
rect -5760 16450 -5750 16470
rect -5730 16450 -5720 16470
rect -5760 16310 -5720 16450
rect -5760 16290 -5750 16310
rect -5730 16290 -5720 16310
rect -5760 16150 -5720 16290
rect -5600 16470 -5560 16480
rect -5600 16450 -5590 16470
rect -5570 16450 -5560 16470
rect -5600 16310 -5560 16450
rect -5600 16290 -5590 16310
rect -5570 16290 -5560 16310
rect -5760 16130 -5750 16150
rect -5730 16130 -5720 16150
rect -5760 15990 -5720 16130
rect -5760 15970 -5750 15990
rect -5730 15970 -5720 15990
rect -5760 15960 -5720 15970
rect -5680 16150 -5640 16160
rect -5680 16130 -5670 16150
rect -5650 16130 -5640 16150
rect -5680 15990 -5640 16130
rect -5680 15970 -5670 15990
rect -5650 15970 -5640 15990
rect -5680 15960 -5640 15970
rect -5600 16150 -5560 16290
rect -5600 16130 -5590 16150
rect -5570 16130 -5560 16150
rect -5600 15990 -5560 16130
rect -5600 15970 -5590 15990
rect -5570 15970 -5560 15990
rect -5600 15960 -5560 15970
rect -5440 16470 -5400 16480
rect -5440 16450 -5430 16470
rect -5410 16450 -5400 16470
rect -5440 16310 -5400 16450
rect -5440 16290 -5430 16310
rect -5410 16290 -5400 16310
rect -5440 16150 -5400 16290
rect -5440 16130 -5430 16150
rect -5410 16130 -5400 16150
rect -5440 15990 -5400 16130
rect -5440 15970 -5430 15990
rect -5410 15970 -5400 15990
rect -5440 15960 -5400 15970
rect -5360 16470 -5320 16480
rect -5360 16450 -5350 16470
rect -5330 16450 -5320 16470
rect -5360 16310 -5320 16450
rect -5360 16290 -5350 16310
rect -5330 16290 -5320 16310
rect -5360 16150 -5320 16290
rect -5360 16130 -5350 16150
rect -5330 16130 -5320 16150
rect -5360 15990 -5320 16130
rect -5360 15970 -5350 15990
rect -5330 15970 -5320 15990
rect -5360 15960 -5320 15970
rect -5280 16470 -5240 16480
rect -5280 16450 -5270 16470
rect -5250 16450 -5240 16470
rect -5280 16310 -5240 16450
rect -5280 16290 -5270 16310
rect -5250 16290 -5240 16310
rect -5280 16150 -5240 16290
rect -5280 16130 -5270 16150
rect -5250 16130 -5240 16150
rect -5280 15990 -5240 16130
rect -5280 15970 -5270 15990
rect -5250 15970 -5240 15990
rect -5280 15960 -5240 15970
rect -5200 16470 -5160 16480
rect -5200 16450 -5190 16470
rect -5170 16450 -5160 16470
rect -5200 16310 -5160 16450
rect -5200 16290 -5190 16310
rect -5170 16290 -5160 16310
rect -5200 16150 -5160 16290
rect -5200 16130 -5190 16150
rect -5170 16130 -5160 16150
rect -5200 15990 -5160 16130
rect -5200 15970 -5190 15990
rect -5170 15970 -5160 15990
rect -5200 15960 -5160 15970
rect -5120 16470 -5080 16480
rect -5120 16450 -5110 16470
rect -5090 16450 -5080 16470
rect -5120 16310 -5080 16450
rect -5120 16290 -5110 16310
rect -5090 16290 -5080 16310
rect -5120 16150 -5080 16290
rect -5120 16130 -5110 16150
rect -5090 16130 -5080 16150
rect -5120 15990 -5080 16130
rect -5120 15970 -5110 15990
rect -5090 15970 -5080 15990
rect -5120 15960 -5080 15970
rect -5040 16470 -5000 16480
rect -5040 16450 -5030 16470
rect -5010 16450 -5000 16470
rect -5040 16310 -5000 16450
rect -5040 16290 -5030 16310
rect -5010 16290 -5000 16310
rect -5040 16150 -5000 16290
rect -5040 16130 -5030 16150
rect -5010 16130 -5000 16150
rect -5040 15990 -5000 16130
rect -5040 15970 -5030 15990
rect -5010 15970 -5000 15990
rect -5040 15960 -5000 15970
rect -4960 16470 -4920 16480
rect -4960 16450 -4950 16470
rect -4930 16450 -4920 16470
rect -4960 16310 -4920 16450
rect -4960 16290 -4950 16310
rect -4930 16290 -4920 16310
rect -4960 16150 -4920 16290
rect -4960 16130 -4950 16150
rect -4930 16130 -4920 16150
rect -4960 15990 -4920 16130
rect -4960 15970 -4950 15990
rect -4930 15970 -4920 15990
rect -4960 15960 -4920 15970
rect -4880 16470 -4840 16480
rect -4880 16450 -4870 16470
rect -4850 16450 -4840 16470
rect -4880 16310 -4840 16450
rect -4880 16290 -4870 16310
rect -4850 16290 -4840 16310
rect -4880 16150 -4840 16290
rect -4880 16130 -4870 16150
rect -4850 16130 -4840 16150
rect -4880 15990 -4840 16130
rect -4880 15970 -4870 15990
rect -4850 15970 -4840 15990
rect -4880 15960 -4840 15970
rect -4800 16470 -4760 16480
rect -4800 16450 -4790 16470
rect -4770 16450 -4760 16470
rect -4800 16310 -4760 16450
rect -4800 16290 -4790 16310
rect -4770 16290 -4760 16310
rect -4800 16150 -4760 16290
rect -4800 16130 -4790 16150
rect -4770 16130 -4760 16150
rect -4800 15990 -4760 16130
rect -4800 15970 -4790 15990
rect -4770 15970 -4760 15990
rect -4800 15960 -4760 15970
rect -4720 16470 -4680 16480
rect -4720 16450 -4710 16470
rect -4690 16450 -4680 16470
rect -4720 16310 -4680 16450
rect -4720 16290 -4710 16310
rect -4690 16290 -4680 16310
rect -4720 16150 -4680 16290
rect -4720 16130 -4710 16150
rect -4690 16130 -4680 16150
rect -4720 15990 -4680 16130
rect -4720 15970 -4710 15990
rect -4690 15970 -4680 15990
rect -4720 15960 -4680 15970
rect -4640 16470 -4600 16480
rect -4640 16450 -4630 16470
rect -4610 16450 -4600 16470
rect -4640 16310 -4600 16450
rect -4640 16290 -4630 16310
rect -4610 16290 -4600 16310
rect -4640 16150 -4600 16290
rect -4640 16130 -4630 16150
rect -4610 16130 -4600 16150
rect -4640 15990 -4600 16130
rect -4640 15970 -4630 15990
rect -4610 15970 -4600 15990
rect -4640 15960 -4600 15970
rect -4560 16470 -4520 16480
rect -4560 16450 -4550 16470
rect -4530 16450 -4520 16470
rect -4560 16310 -4520 16450
rect -4560 16290 -4550 16310
rect -4530 16290 -4520 16310
rect -4560 16150 -4520 16290
rect -4560 16130 -4550 16150
rect -4530 16130 -4520 16150
rect -4560 15990 -4520 16130
rect -4560 15970 -4550 15990
rect -4530 15970 -4520 15990
rect -4560 15960 -4520 15970
rect -4480 16470 -4440 16480
rect -4480 16450 -4470 16470
rect -4450 16450 -4440 16470
rect -4480 16310 -4440 16450
rect -4480 16290 -4470 16310
rect -4450 16290 -4440 16310
rect -4480 16150 -4440 16290
rect -4480 16130 -4470 16150
rect -4450 16130 -4440 16150
rect -4480 15990 -4440 16130
rect -4480 15970 -4470 15990
rect -4450 15970 -4440 15990
rect -4480 15960 -4440 15970
rect -4400 16470 -4360 16480
rect -4400 16450 -4390 16470
rect -4370 16450 -4360 16470
rect -4400 16310 -4360 16450
rect -4400 16290 -4390 16310
rect -4370 16290 -4360 16310
rect -4400 16150 -4360 16290
rect -4400 16130 -4390 16150
rect -4370 16130 -4360 16150
rect -4400 15990 -4360 16130
rect -4400 15970 -4390 15990
rect -4370 15970 -4360 15990
rect -4400 15960 -4360 15970
rect -4320 16470 -4280 16480
rect -4320 16450 -4310 16470
rect -4290 16450 -4280 16470
rect -4320 16310 -4280 16450
rect -4320 16290 -4310 16310
rect -4290 16290 -4280 16310
rect -4320 16150 -4280 16290
rect -4320 16130 -4310 16150
rect -4290 16130 -4280 16150
rect -4320 15990 -4280 16130
rect -4320 15970 -4310 15990
rect -4290 15970 -4280 15990
rect -4320 15960 -4280 15970
rect -4240 16470 -4200 16480
rect -4240 16450 -4230 16470
rect -4210 16450 -4200 16470
rect -4240 16310 -4200 16450
rect -4240 16290 -4230 16310
rect -4210 16290 -4200 16310
rect -4240 16150 -4200 16290
rect -4240 16130 -4230 16150
rect -4210 16130 -4200 16150
rect -4240 15990 -4200 16130
rect -4240 15970 -4230 15990
rect -4210 15970 -4200 15990
rect -4240 15960 -4200 15970
rect -4160 16470 -4120 16480
rect -4160 16450 -4150 16470
rect -4130 16450 -4120 16470
rect -4160 16310 -4120 16450
rect -4160 16290 -4150 16310
rect -4130 16290 -4120 16310
rect -4160 16150 -4120 16290
rect -4160 16130 -4150 16150
rect -4130 16130 -4120 16150
rect -4160 15990 -4120 16130
rect -4160 15970 -4150 15990
rect -4130 15970 -4120 15990
rect -4160 15960 -4120 15970
rect -4080 16470 -4040 16480
rect -4080 16450 -4070 16470
rect -4050 16450 -4040 16470
rect -4080 16310 -4040 16450
rect -4080 16290 -4070 16310
rect -4050 16290 -4040 16310
rect -4080 16150 -4040 16290
rect -4080 16130 -4070 16150
rect -4050 16130 -4040 16150
rect -4080 15990 -4040 16130
rect -4080 15970 -4070 15990
rect -4050 15970 -4040 15990
rect -4080 15960 -4040 15970
rect -4000 16470 -3960 16480
rect -4000 16450 -3990 16470
rect -3970 16450 -3960 16470
rect -4000 16310 -3960 16450
rect -4000 16290 -3990 16310
rect -3970 16290 -3960 16310
rect -4000 16150 -3960 16290
rect -4000 16130 -3990 16150
rect -3970 16130 -3960 16150
rect -4000 15990 -3960 16130
rect -4000 15970 -3990 15990
rect -3970 15970 -3960 15990
rect -4000 15960 -3960 15970
rect -3920 16470 -3880 16480
rect -3920 16450 -3910 16470
rect -3890 16450 -3880 16470
rect -3920 16310 -3880 16450
rect -3920 16290 -3910 16310
rect -3890 16290 -3880 16310
rect -3920 16150 -3880 16290
rect -3920 16130 -3910 16150
rect -3890 16130 -3880 16150
rect -3920 15990 -3880 16130
rect -3920 15970 -3910 15990
rect -3890 15970 -3880 15990
rect -3920 15960 -3880 15970
rect -3840 16470 -3800 16480
rect -3840 16450 -3830 16470
rect -3810 16450 -3800 16470
rect -3840 16310 -3800 16450
rect -3840 16290 -3830 16310
rect -3810 16290 -3800 16310
rect -3840 16150 -3800 16290
rect -3840 16130 -3830 16150
rect -3810 16130 -3800 16150
rect -3840 15990 -3800 16130
rect -3840 15970 -3830 15990
rect -3810 15970 -3800 15990
rect -3840 15960 -3800 15970
rect -3760 16470 -3720 16480
rect -3760 16450 -3750 16470
rect -3730 16450 -3720 16470
rect -3760 16310 -3720 16450
rect -3760 16290 -3750 16310
rect -3730 16290 -3720 16310
rect -3760 16150 -3720 16290
rect -3760 16130 -3750 16150
rect -3730 16130 -3720 16150
rect -3760 15990 -3720 16130
rect -3760 15970 -3750 15990
rect -3730 15970 -3720 15990
rect -3760 15960 -3720 15970
rect -3680 16470 -3640 16480
rect -3680 16450 -3670 16470
rect -3650 16450 -3640 16470
rect -3680 16310 -3640 16450
rect -3680 16290 -3670 16310
rect -3650 16290 -3640 16310
rect -3680 16150 -3640 16290
rect -3680 16130 -3670 16150
rect -3650 16130 -3640 16150
rect -3680 15990 -3640 16130
rect -3680 15970 -3670 15990
rect -3650 15970 -3640 15990
rect -3680 15960 -3640 15970
rect -3600 16470 -3560 16480
rect -3600 16450 -3590 16470
rect -3570 16450 -3560 16470
rect -3600 16310 -3560 16450
rect -3600 16290 -3590 16310
rect -3570 16290 -3560 16310
rect -3600 16150 -3560 16290
rect -3600 16130 -3590 16150
rect -3570 16130 -3560 16150
rect -3600 15990 -3560 16130
rect -3600 15970 -3590 15990
rect -3570 15970 -3560 15990
rect -3600 15960 -3560 15970
rect -3520 16470 -3480 16480
rect -3520 16450 -3510 16470
rect -3490 16450 -3480 16470
rect -3520 16310 -3480 16450
rect -3520 16290 -3510 16310
rect -3490 16290 -3480 16310
rect -3520 16150 -3480 16290
rect -3520 16130 -3510 16150
rect -3490 16130 -3480 16150
rect -3520 15990 -3480 16130
rect -3520 15970 -3510 15990
rect -3490 15970 -3480 15990
rect -3520 15960 -3480 15970
rect -3440 16470 -3400 16480
rect -3440 16450 -3430 16470
rect -3410 16450 -3400 16470
rect -3440 16310 -3400 16450
rect -3440 16290 -3430 16310
rect -3410 16290 -3400 16310
rect -3440 16150 -3400 16290
rect -3440 16130 -3430 16150
rect -3410 16130 -3400 16150
rect -3440 15990 -3400 16130
rect -3440 15970 -3430 15990
rect -3410 15970 -3400 15990
rect -3440 15960 -3400 15970
rect -3360 16470 -3320 16480
rect -3360 16450 -3350 16470
rect -3330 16450 -3320 16470
rect -3360 16310 -3320 16450
rect -3360 16290 -3350 16310
rect -3330 16290 -3320 16310
rect -3360 16150 -3320 16290
rect -3360 16130 -3350 16150
rect -3330 16130 -3320 16150
rect -3360 15990 -3320 16130
rect -3360 15970 -3350 15990
rect -3330 15970 -3320 15990
rect -3360 15960 -3320 15970
rect -3280 16470 -3240 16480
rect -3280 16450 -3270 16470
rect -3250 16450 -3240 16470
rect -3280 16310 -3240 16450
rect -3280 16290 -3270 16310
rect -3250 16290 -3240 16310
rect -3280 16150 -3240 16290
rect -3280 16130 -3270 16150
rect -3250 16130 -3240 16150
rect -3280 15990 -3240 16130
rect -3280 15970 -3270 15990
rect -3250 15970 -3240 15990
rect -3280 15960 -3240 15970
rect -3200 16470 -3160 16480
rect -3200 16450 -3190 16470
rect -3170 16450 -3160 16470
rect -3200 16310 -3160 16450
rect -3200 16290 -3190 16310
rect -3170 16290 -3160 16310
rect -3200 16150 -3160 16290
rect -3200 16130 -3190 16150
rect -3170 16130 -3160 16150
rect -3200 15990 -3160 16130
rect -3200 15970 -3190 15990
rect -3170 15970 -3160 15990
rect -3200 15960 -3160 15970
rect -3120 16470 -3080 16480
rect -3120 16450 -3110 16470
rect -3090 16450 -3080 16470
rect -3120 16310 -3080 16450
rect -3120 16290 -3110 16310
rect -3090 16290 -3080 16310
rect -3120 16150 -3080 16290
rect -3120 16130 -3110 16150
rect -3090 16130 -3080 16150
rect -3120 15990 -3080 16130
rect -3120 15970 -3110 15990
rect -3090 15970 -3080 15990
rect -3120 15960 -3080 15970
rect -3040 16470 -3000 16480
rect -3040 16450 -3030 16470
rect -3010 16450 -3000 16470
rect -3040 16310 -3000 16450
rect -3040 16290 -3030 16310
rect -3010 16290 -3000 16310
rect -3040 16150 -3000 16290
rect -3040 16130 -3030 16150
rect -3010 16130 -3000 16150
rect -3040 15990 -3000 16130
rect -3040 15970 -3030 15990
rect -3010 15970 -3000 15990
rect -3040 15960 -3000 15970
rect -2960 16470 -2920 16480
rect -2960 16450 -2950 16470
rect -2930 16450 -2920 16470
rect -2960 16310 -2920 16450
rect -2960 16290 -2950 16310
rect -2930 16290 -2920 16310
rect -2960 16150 -2920 16290
rect -2960 16130 -2950 16150
rect -2930 16130 -2920 16150
rect -2960 15990 -2920 16130
rect -2960 15970 -2950 15990
rect -2930 15970 -2920 15990
rect -2960 15960 -2920 15970
rect -2880 16470 -2840 16480
rect -2880 16450 -2870 16470
rect -2850 16450 -2840 16470
rect -2880 16310 -2840 16450
rect -2880 16290 -2870 16310
rect -2850 16290 -2840 16310
rect -2880 16150 -2840 16290
rect -2880 16130 -2870 16150
rect -2850 16130 -2840 16150
rect -2880 15990 -2840 16130
rect -2880 15970 -2870 15990
rect -2850 15970 -2840 15990
rect -2880 15960 -2840 15970
rect -2800 16470 -2760 16480
rect -2800 16450 -2790 16470
rect -2770 16450 -2760 16470
rect -2800 16310 -2760 16450
rect -2800 16290 -2790 16310
rect -2770 16290 -2760 16310
rect -2800 16150 -2760 16290
rect -2800 16130 -2790 16150
rect -2770 16130 -2760 16150
rect -2800 15990 -2760 16130
rect -2800 15970 -2790 15990
rect -2770 15970 -2760 15990
rect -2800 15960 -2760 15970
rect -2720 16470 -2680 16480
rect -2720 16450 -2710 16470
rect -2690 16450 -2680 16470
rect -2720 16310 -2680 16450
rect -2720 16290 -2710 16310
rect -2690 16290 -2680 16310
rect -2720 16150 -2680 16290
rect -2720 16130 -2710 16150
rect -2690 16130 -2680 16150
rect -2720 15990 -2680 16130
rect -2720 15970 -2710 15990
rect -2690 15970 -2680 15990
rect -2720 15960 -2680 15970
rect -2640 16470 -2600 16480
rect -2640 16450 -2630 16470
rect -2610 16450 -2600 16470
rect -2640 16310 -2600 16450
rect -2640 16290 -2630 16310
rect -2610 16290 -2600 16310
rect -2640 16150 -2600 16290
rect -2640 16130 -2630 16150
rect -2610 16130 -2600 16150
rect -2640 15990 -2600 16130
rect -2640 15970 -2630 15990
rect -2610 15970 -2600 15990
rect -2640 15960 -2600 15970
rect -2560 16470 -2520 16480
rect -2560 16450 -2550 16470
rect -2530 16450 -2520 16470
rect -2560 16310 -2520 16450
rect -2560 16290 -2550 16310
rect -2530 16290 -2520 16310
rect -2560 16150 -2520 16290
rect -2560 16130 -2550 16150
rect -2530 16130 -2520 16150
rect -2560 15990 -2520 16130
rect -2560 15970 -2550 15990
rect -2530 15970 -2520 15990
rect -2560 15960 -2520 15970
rect -2480 16470 -2440 16480
rect -2480 16450 -2470 16470
rect -2450 16450 -2440 16470
rect -2480 16310 -2440 16450
rect -2480 16290 -2470 16310
rect -2450 16290 -2440 16310
rect -2480 16150 -2440 16290
rect -2480 16130 -2470 16150
rect -2450 16130 -2440 16150
rect -2480 15990 -2440 16130
rect -2480 15970 -2470 15990
rect -2450 15970 -2440 15990
rect -2480 15960 -2440 15970
rect -2400 16470 -2360 16480
rect -2400 16450 -2390 16470
rect -2370 16450 -2360 16470
rect -2400 16310 -2360 16450
rect -2400 16290 -2390 16310
rect -2370 16290 -2360 16310
rect -2400 16150 -2360 16290
rect -2400 16130 -2390 16150
rect -2370 16130 -2360 16150
rect -2400 15990 -2360 16130
rect -2400 15970 -2390 15990
rect -2370 15970 -2360 15990
rect -2400 15960 -2360 15970
rect -2320 16470 -2280 16480
rect -2320 16450 -2310 16470
rect -2290 16450 -2280 16470
rect -2320 16310 -2280 16450
rect -2320 16290 -2310 16310
rect -2290 16290 -2280 16310
rect -2320 16150 -2280 16290
rect -2320 16130 -2310 16150
rect -2290 16130 -2280 16150
rect -2320 15990 -2280 16130
rect -2320 15970 -2310 15990
rect -2290 15970 -2280 15990
rect -2320 15960 -2280 15970
rect -2240 16470 -2200 16480
rect -2240 16450 -2230 16470
rect -2210 16450 -2200 16470
rect -2240 16310 -2200 16450
rect -2240 16290 -2230 16310
rect -2210 16290 -2200 16310
rect -2240 16150 -2200 16290
rect -2240 16130 -2230 16150
rect -2210 16130 -2200 16150
rect -2240 15990 -2200 16130
rect -2240 15970 -2230 15990
rect -2210 15970 -2200 15990
rect -2240 15960 -2200 15970
rect -2160 16470 -2120 16480
rect -2160 16450 -2150 16470
rect -2130 16450 -2120 16470
rect -2160 16310 -2120 16450
rect -2160 16290 -2150 16310
rect -2130 16290 -2120 16310
rect -2160 16150 -2120 16290
rect -2160 16130 -2150 16150
rect -2130 16130 -2120 16150
rect -2160 15990 -2120 16130
rect -2160 15970 -2150 15990
rect -2130 15970 -2120 15990
rect -2160 15960 -2120 15970
rect -2080 16470 -2040 16480
rect -2080 16450 -2070 16470
rect -2050 16450 -2040 16470
rect -2080 16310 -2040 16450
rect -2080 16290 -2070 16310
rect -2050 16290 -2040 16310
rect -2080 16150 -2040 16290
rect -2080 16130 -2070 16150
rect -2050 16130 -2040 16150
rect -2080 15990 -2040 16130
rect -2080 15970 -2070 15990
rect -2050 15970 -2040 15990
rect -2080 15960 -2040 15970
rect -2000 16470 -1960 16480
rect -2000 16450 -1990 16470
rect -1970 16450 -1960 16470
rect -2000 16310 -1960 16450
rect -2000 16290 -1990 16310
rect -1970 16290 -1960 16310
rect -2000 16150 -1960 16290
rect -2000 16130 -1990 16150
rect -1970 16130 -1960 16150
rect -2000 15990 -1960 16130
rect -2000 15970 -1990 15990
rect -1970 15970 -1960 15990
rect -2000 15960 -1960 15970
rect -1920 15920 -1880 17440
rect -1840 16470 -1800 16480
rect -1840 16450 -1830 16470
rect -1810 16450 -1800 16470
rect -1840 16310 -1800 16450
rect -1840 16290 -1830 16310
rect -1810 16290 -1800 16310
rect -1840 16150 -1800 16290
rect -1840 16130 -1830 16150
rect -1810 16130 -1800 16150
rect -1840 15990 -1800 16130
rect -1840 15970 -1830 15990
rect -1810 15970 -1800 15990
rect -1840 15960 -1800 15970
rect -1760 16470 -1720 16480
rect -1760 16450 -1750 16470
rect -1730 16450 -1720 16470
rect -1760 16310 -1720 16450
rect -1760 16290 -1750 16310
rect -1730 16290 -1720 16310
rect -1760 16150 -1720 16290
rect -1760 16130 -1750 16150
rect -1730 16130 -1720 16150
rect -1760 15990 -1720 16130
rect -1760 15970 -1750 15990
rect -1730 15970 -1720 15990
rect -1760 15960 -1720 15970
rect -1680 16470 -1640 16480
rect -1680 16450 -1670 16470
rect -1650 16450 -1640 16470
rect -1680 16310 -1640 16450
rect -1680 16290 -1670 16310
rect -1650 16290 -1640 16310
rect -1680 16150 -1640 16290
rect -1680 16130 -1670 16150
rect -1650 16130 -1640 16150
rect -1680 15990 -1640 16130
rect -1680 15970 -1670 15990
rect -1650 15970 -1640 15990
rect -1680 15960 -1640 15970
rect -1600 16470 -1560 16480
rect -1600 16450 -1590 16470
rect -1570 16450 -1560 16470
rect -1600 16310 -1560 16450
rect -1600 16290 -1590 16310
rect -1570 16290 -1560 16310
rect -1600 16150 -1560 16290
rect -1600 16130 -1590 16150
rect -1570 16130 -1560 16150
rect -1600 15990 -1560 16130
rect -1600 15970 -1590 15990
rect -1570 15970 -1560 15990
rect -1600 15960 -1560 15970
rect -1520 16470 -1480 16480
rect -1520 16450 -1510 16470
rect -1490 16450 -1480 16470
rect -1520 16310 -1480 16450
rect -1520 16290 -1510 16310
rect -1490 16290 -1480 16310
rect -1520 16150 -1480 16290
rect -1520 16130 -1510 16150
rect -1490 16130 -1480 16150
rect -1520 15990 -1480 16130
rect -1520 15970 -1510 15990
rect -1490 15970 -1480 15990
rect -1520 15960 -1480 15970
rect -1440 16470 -1400 16480
rect -1440 16450 -1430 16470
rect -1410 16450 -1400 16470
rect -1440 16310 -1400 16450
rect -1440 16290 -1430 16310
rect -1410 16290 -1400 16310
rect -1440 16150 -1400 16290
rect -1440 16130 -1430 16150
rect -1410 16130 -1400 16150
rect -1440 15990 -1400 16130
rect -1440 15970 -1430 15990
rect -1410 15970 -1400 15990
rect -1440 15960 -1400 15970
rect -1360 16470 -1320 16480
rect -1360 16450 -1350 16470
rect -1330 16450 -1320 16470
rect -1360 16310 -1320 16450
rect -1360 16290 -1350 16310
rect -1330 16290 -1320 16310
rect -1360 16150 -1320 16290
rect -1360 16130 -1350 16150
rect -1330 16130 -1320 16150
rect -1360 15990 -1320 16130
rect -1360 15970 -1350 15990
rect -1330 15970 -1320 15990
rect -1360 15960 -1320 15970
rect -1200 16470 -1160 16480
rect -1200 16450 -1190 16470
rect -1170 16450 -1160 16470
rect -1200 16310 -1160 16450
rect -1200 16290 -1190 16310
rect -1170 16290 -1160 16310
rect -1200 16150 -1160 16290
rect -1200 16130 -1190 16150
rect -1170 16130 -1160 16150
rect -1200 15990 -1160 16130
rect -1200 15970 -1190 15990
rect -1170 15970 -1160 15990
rect -1200 15960 -1160 15970
rect -1040 16470 -1000 16480
rect -1040 16450 -1030 16470
rect -1010 16450 -1000 16470
rect -1040 16310 -1000 16450
rect -1040 16290 -1030 16310
rect -1010 16290 -1000 16310
rect -1040 16150 -1000 16290
rect -1040 16130 -1030 16150
rect -1010 16130 -1000 16150
rect -1040 15990 -1000 16130
rect -1040 15970 -1030 15990
rect -1010 15970 -1000 15990
rect -1040 15960 -1000 15970
rect -880 16470 -840 16480
rect -880 16450 -870 16470
rect -850 16450 -840 16470
rect -880 16310 -840 16450
rect -880 16290 -870 16310
rect -850 16290 -840 16310
rect -880 16150 -840 16290
rect -880 16130 -870 16150
rect -850 16130 -840 16150
rect -880 15990 -840 16130
rect -880 15970 -870 15990
rect -850 15970 -840 15990
rect -880 15960 -840 15970
rect -720 16470 -680 16480
rect -720 16450 -710 16470
rect -690 16450 -680 16470
rect -720 16310 -680 16450
rect -720 16290 -710 16310
rect -690 16290 -680 16310
rect -720 16150 -680 16290
rect -720 16130 -710 16150
rect -690 16130 -680 16150
rect -720 15990 -680 16130
rect -720 15970 -710 15990
rect -690 15970 -680 15990
rect -720 15960 -680 15970
rect -560 16470 -520 16480
rect -560 16450 -550 16470
rect -530 16450 -520 16470
rect -560 16310 -520 16450
rect -560 16290 -550 16310
rect -530 16290 -520 16310
rect -560 16150 -520 16290
rect -560 16130 -550 16150
rect -530 16130 -520 16150
rect -560 15990 -520 16130
rect -560 15970 -550 15990
rect -530 15970 -520 15990
rect -560 15960 -520 15970
<< viali >>
rect -14950 21410 -14930 21430
rect -14950 21250 -14930 21270
rect -14950 21090 -14930 21110
rect -14950 20930 -14930 20950
rect -14870 21410 -14850 21430
rect -14870 21250 -14850 21270
rect -14870 21090 -14850 21110
rect -14870 20930 -14850 20950
rect -14790 21410 -14770 21430
rect -14790 21250 -14770 21270
rect -14790 21090 -14770 21110
rect -14790 20930 -14770 20950
rect -14710 21410 -14690 21430
rect -14710 21250 -14690 21270
rect -14710 21090 -14690 21110
rect -14710 20930 -14690 20950
rect -14630 21410 -14610 21430
rect -14630 21250 -14610 21270
rect -14630 21090 -14610 21110
rect -14630 20930 -14610 20950
rect -14550 21410 -14530 21430
rect -14550 21250 -14530 21270
rect -14550 21090 -14530 21110
rect -14550 20930 -14530 20950
rect -14470 21410 -14450 21430
rect -14470 21250 -14450 21270
rect -14470 21090 -14450 21110
rect -14470 20930 -14450 20950
rect -14390 21410 -14370 21430
rect -14390 21250 -14370 21270
rect -14390 21090 -14370 21110
rect -14390 20930 -14370 20950
rect -14310 21410 -14290 21430
rect -14310 21250 -14290 21270
rect -14310 21090 -14290 21110
rect -14310 20930 -14290 20950
rect -14230 21410 -14210 21430
rect -14230 21250 -14210 21270
rect -14230 21090 -14210 21110
rect -14230 20930 -14210 20950
rect -14150 21410 -14130 21430
rect -14150 21250 -14130 21270
rect -14150 21090 -14130 21110
rect -14150 20930 -14130 20950
rect -14070 21410 -14050 21430
rect -14070 21250 -14050 21270
rect -14070 21090 -14050 21110
rect -14070 20930 -14050 20950
rect -13990 21410 -13970 21430
rect -13990 21250 -13970 21270
rect -13990 21090 -13970 21110
rect -13990 20930 -13970 20950
rect -13910 21410 -13890 21430
rect -13910 21250 -13890 21270
rect -13910 21090 -13890 21110
rect -13910 20930 -13890 20950
rect -13830 21410 -13810 21430
rect -13830 21250 -13810 21270
rect -13830 21090 -13810 21110
rect -13830 20930 -13810 20950
rect -13750 21410 -13730 21430
rect -13750 21250 -13730 21270
rect -13750 21090 -13730 21110
rect -13750 20930 -13730 20950
rect -13670 21410 -13650 21430
rect -13670 21250 -13650 21270
rect -13670 21090 -13650 21110
rect -13670 20930 -13650 20950
rect -13590 21410 -13570 21430
rect -13590 21250 -13570 21270
rect -13590 21090 -13570 21110
rect -13590 20930 -13570 20950
rect -13510 21410 -13490 21430
rect -13510 21250 -13490 21270
rect -13510 21090 -13490 21110
rect -13510 20930 -13490 20950
rect -13430 21410 -13410 21430
rect -13430 21250 -13410 21270
rect -13430 21090 -13410 21110
rect -13430 20930 -13410 20950
rect -13350 21410 -13330 21430
rect -13350 21250 -13330 21270
rect -13350 21090 -13330 21110
rect -13350 20930 -13330 20950
rect -13270 21410 -13250 21430
rect -13270 21250 -13250 21270
rect -13270 21090 -13250 21110
rect -13270 20930 -13250 20950
rect -13190 21410 -13170 21430
rect -13190 21250 -13170 21270
rect -13190 21090 -13170 21110
rect -13190 20930 -13170 20950
rect -13110 21410 -13090 21430
rect -13110 21250 -13090 21270
rect -13110 21090 -13090 21110
rect -13110 20930 -13090 20950
rect -13030 21410 -13010 21430
rect -13030 21250 -13010 21270
rect -13030 21090 -13010 21110
rect -13030 20930 -13010 20950
rect -12950 21410 -12930 21430
rect -12950 21250 -12930 21270
rect -12950 21090 -12930 21110
rect -12950 20930 -12930 20950
rect -12870 21410 -12850 21430
rect -12870 21250 -12850 21270
rect -12870 21090 -12850 21110
rect -12870 20930 -12850 20950
rect -12790 21410 -12770 21430
rect -12790 21250 -12770 21270
rect -12790 21090 -12770 21110
rect -12790 20930 -12770 20950
rect -12710 21410 -12690 21430
rect -12710 21250 -12690 21270
rect -12710 21090 -12690 21110
rect -12710 20930 -12690 20950
rect -12630 21410 -12610 21430
rect -12630 21250 -12610 21270
rect -12630 21090 -12610 21110
rect -12630 20930 -12610 20950
rect -12550 21410 -12530 21430
rect -12550 21250 -12530 21270
rect -12550 21090 -12530 21110
rect -12550 20930 -12530 20950
rect -12470 21410 -12450 21430
rect -12470 21250 -12450 21270
rect -12470 21090 -12450 21110
rect -12470 20930 -12450 20950
rect -12390 21410 -12370 21430
rect -12390 21250 -12370 21270
rect -12390 21090 -12370 21110
rect -12390 20930 -12370 20950
rect -12310 21410 -12290 21430
rect -12310 21250 -12290 21270
rect -12310 21090 -12290 21110
rect -12310 20930 -12290 20950
rect -12230 21410 -12210 21430
rect -12230 21250 -12210 21270
rect -12230 21090 -12210 21110
rect -12230 20930 -12210 20950
rect -12150 21410 -12130 21430
rect -12150 21250 -12130 21270
rect -12150 21090 -12130 21110
rect -12150 20930 -12130 20950
rect -12070 21410 -12050 21430
rect -12070 21250 -12050 21270
rect -12070 21090 -12050 21110
rect -12070 20930 -12050 20950
rect -11990 21410 -11970 21430
rect -11990 21250 -11970 21270
rect -11990 21090 -11970 21110
rect -11990 20930 -11970 20950
rect -11910 21410 -11890 21430
rect -11910 21250 -11890 21270
rect -11910 21090 -11890 21110
rect -11910 20930 -11890 20950
rect -11830 21410 -11810 21430
rect -11830 21250 -11810 21270
rect -11830 21090 -11810 21110
rect -11830 20930 -11810 20950
rect -11750 21410 -11730 21430
rect -11750 21250 -11730 21270
rect -11750 21090 -11730 21110
rect -11750 20930 -11730 20950
rect -11670 21410 -11650 21430
rect -11670 21250 -11650 21270
rect -11670 21090 -11650 21110
rect -11670 20930 -11650 20950
rect -11590 21410 -11570 21430
rect -11590 21250 -11570 21270
rect -11590 21090 -11570 21110
rect -11590 20930 -11570 20950
rect -11510 21410 -11490 21430
rect -11510 21250 -11490 21270
rect -11510 21090 -11490 21110
rect -11510 20930 -11490 20950
rect -11430 21410 -11410 21430
rect -11430 21250 -11410 21270
rect -11430 21090 -11410 21110
rect -11430 20930 -11410 20950
rect -11350 21410 -11330 21430
rect -11350 21250 -11330 21270
rect -11350 21090 -11330 21110
rect -11350 20930 -11330 20950
rect -11270 21410 -11250 21430
rect -11270 21250 -11250 21270
rect -11270 21090 -11250 21110
rect -11270 20930 -11250 20950
rect -11190 21410 -11170 21430
rect -11190 21250 -11170 21270
rect -11190 21090 -11170 21110
rect -11190 20930 -11170 20950
rect -11110 21410 -11090 21430
rect -11110 21250 -11090 21270
rect -11110 21090 -11090 21110
rect -11110 20930 -11090 20950
rect -11030 21410 -11010 21430
rect -11030 21250 -11010 21270
rect -11030 21090 -11010 21110
rect -11030 20930 -11010 20950
rect -10950 21410 -10930 21430
rect -10950 21250 -10930 21270
rect -10950 21090 -10930 21110
rect -10950 20930 -10930 20950
rect -10870 21410 -10850 21430
rect -10870 21250 -10850 21270
rect -10870 21090 -10850 21110
rect -10870 20930 -10850 20950
rect -10790 21410 -10770 21430
rect -10790 21250 -10770 21270
rect -10790 21090 -10770 21110
rect -10790 20930 -10770 20950
rect -10710 21410 -10690 21430
rect -10710 21250 -10690 21270
rect -10710 21090 -10690 21110
rect -10710 20930 -10690 20950
rect -10630 21410 -10610 21430
rect -10630 21250 -10610 21270
rect -10630 21090 -10610 21110
rect -10630 20930 -10610 20950
rect -10550 21410 -10530 21430
rect -10550 21250 -10530 21270
rect -10550 21090 -10530 21110
rect -10550 20930 -10530 20950
rect -10470 21410 -10450 21430
rect -10470 21250 -10450 21270
rect -10470 21090 -10450 21110
rect -10470 20930 -10450 20950
rect -10390 21410 -10370 21430
rect -10390 21250 -10370 21270
rect -10390 21090 -10370 21110
rect -10390 20930 -10370 20950
rect -10310 21410 -10290 21430
rect -10310 21250 -10290 21270
rect -10310 21090 -10290 21110
rect -10310 20930 -10290 20950
rect -10230 21410 -10210 21430
rect -10230 21250 -10210 21270
rect -10230 21090 -10210 21110
rect -10230 20930 -10210 20950
rect -10150 21410 -10130 21430
rect -10150 21250 -10130 21270
rect -10150 21090 -10130 21110
rect -10150 20930 -10130 20950
rect -10070 21410 -10050 21430
rect -10070 21250 -10050 21270
rect -10070 21090 -10050 21110
rect -10070 20930 -10050 20950
rect -9990 21410 -9970 21430
rect -9990 21250 -9970 21270
rect -9990 21090 -9970 21110
rect -9990 20930 -9970 20950
rect -9910 21410 -9890 21430
rect -9910 21250 -9890 21270
rect -9910 21090 -9890 21110
rect -9910 20930 -9890 20950
rect -9830 21410 -9810 21430
rect -9830 21250 -9810 21270
rect -9830 21090 -9810 21110
rect -9830 20930 -9810 20950
rect -9750 21410 -9730 21430
rect -9750 21250 -9730 21270
rect -9750 21090 -9730 21110
rect -9750 20930 -9730 20950
rect -9670 21410 -9650 21430
rect -9670 21250 -9650 21270
rect -9670 21090 -9650 21110
rect -9670 20930 -9650 20950
rect -9590 21410 -9570 21430
rect -9590 21250 -9570 21270
rect -9590 21090 -9570 21110
rect -9590 20930 -9570 20950
rect -9510 21410 -9490 21430
rect -9510 21250 -9490 21270
rect -9510 21090 -9490 21110
rect -9510 20930 -9490 20950
rect -9430 21410 -9410 21430
rect -9430 21250 -9410 21270
rect -9430 21090 -9410 21110
rect -9430 20930 -9410 20950
rect -9350 21410 -9330 21430
rect -9350 21250 -9330 21270
rect -9350 21090 -9330 21110
rect -9350 20930 -9330 20950
rect -9270 21410 -9250 21430
rect -9270 21250 -9250 21270
rect -9270 21090 -9250 21110
rect -9270 20930 -9250 20950
rect -9190 21410 -9170 21430
rect -9190 21250 -9170 21270
rect -9190 21090 -9170 21110
rect -9190 20930 -9170 20950
rect -9110 21410 -9090 21430
rect -9110 21250 -9090 21270
rect -9110 21090 -9090 21110
rect -9110 20930 -9090 20950
rect -9030 21410 -9010 21430
rect -9030 21250 -9010 21270
rect -9030 21090 -9010 21110
rect -9030 20930 -9010 20950
rect -8950 21410 -8930 21430
rect -8950 21250 -8930 21270
rect -8950 21090 -8930 21110
rect -8950 20930 -8930 20950
rect -8870 21410 -8850 21430
rect -8870 21250 -8850 21270
rect -8870 21090 -8850 21110
rect -8870 20930 -8850 20950
rect -8790 21410 -8770 21430
rect -8790 21250 -8770 21270
rect -8790 21090 -8770 21110
rect -8790 20930 -8770 20950
rect -8710 21410 -8690 21430
rect -8710 21250 -8690 21270
rect -8710 21090 -8690 21110
rect -8710 20930 -8690 20950
rect -8630 21410 -8610 21430
rect -8630 21250 -8610 21270
rect -8630 21090 -8610 21110
rect -8630 20930 -8610 20950
rect -8550 21410 -8530 21430
rect -8550 21250 -8530 21270
rect -8550 21090 -8530 21110
rect -8550 20930 -8530 20950
rect -8470 21410 -8450 21430
rect -8470 21250 -8450 21270
rect -8470 21090 -8450 21110
rect -8470 20930 -8450 20950
rect -8390 21410 -8370 21430
rect -8390 21250 -8370 21270
rect -8390 21090 -8370 21110
rect -8390 20930 -8370 20950
rect -8310 21410 -8290 21430
rect -8310 21250 -8290 21270
rect -8310 21090 -8290 21110
rect -8310 20930 -8290 20950
rect -8230 21410 -8210 21430
rect -8230 21250 -8210 21270
rect -8230 21090 -8210 21110
rect -8230 20930 -8210 20950
rect -8150 21410 -8130 21430
rect -8150 21250 -8130 21270
rect -8150 21090 -8130 21110
rect -8150 20930 -8130 20950
rect -8070 21410 -8050 21430
rect -8070 21250 -8050 21270
rect -8070 21090 -8050 21110
rect -8070 20930 -8050 20950
rect -7990 21410 -7970 21430
rect -7990 21250 -7970 21270
rect -7990 21090 -7970 21110
rect -7990 20930 -7970 20950
rect -7910 21410 -7890 21430
rect -7910 21250 -7890 21270
rect -7910 21090 -7890 21110
rect -7910 20930 -7890 20950
rect -7830 21410 -7810 21430
rect -7830 21250 -7810 21270
rect -7830 21090 -7810 21110
rect -7830 20930 -7810 20950
rect -7750 21410 -7730 21430
rect -7750 21250 -7730 21270
rect -7750 21090 -7730 21110
rect -7750 20930 -7730 20950
rect -7670 21410 -7650 21430
rect -7670 21250 -7650 21270
rect -7670 21090 -7650 21110
rect -7670 20930 -7650 20950
rect -7590 21410 -7570 21430
rect -7590 21250 -7570 21270
rect -7590 21090 -7570 21110
rect -7590 20930 -7570 20950
rect -7510 21410 -7490 21430
rect -7510 21250 -7490 21270
rect -7510 21090 -7490 21110
rect -7510 20930 -7490 20950
rect -7430 21410 -7410 21430
rect -7430 21250 -7410 21270
rect -7430 21090 -7410 21110
rect -7430 20930 -7410 20950
rect -7350 21410 -7330 21430
rect -7350 21250 -7330 21270
rect -7350 21090 -7330 21110
rect -7350 20930 -7330 20950
rect -7270 21410 -7250 21430
rect -7270 21250 -7250 21270
rect -7270 21090 -7250 21110
rect -7270 20930 -7250 20950
rect -7190 21410 -7170 21430
rect -7190 21250 -7170 21270
rect -7190 21090 -7170 21110
rect -7190 20930 -7170 20950
rect -7110 21410 -7090 21430
rect -7110 21250 -7090 21270
rect -7110 21090 -7090 21110
rect -7110 20930 -7090 20950
rect -7030 21410 -7010 21430
rect -7030 21250 -7010 21270
rect -7030 21090 -7010 21110
rect -7030 20930 -7010 20950
rect -6950 21410 -6930 21430
rect -6950 21250 -6930 21270
rect -6950 21090 -6930 21110
rect -6950 20930 -6930 20950
rect -6870 21410 -6850 21430
rect -6870 21250 -6850 21270
rect -6870 21090 -6850 21110
rect -6870 20930 -6850 20950
rect -6790 21410 -6770 21430
rect -6790 21250 -6770 21270
rect -6790 21090 -6770 21110
rect -6790 20930 -6770 20950
rect -6710 21410 -6690 21430
rect -6710 21250 -6690 21270
rect -6710 21090 -6690 21110
rect -6710 20930 -6690 20950
rect -6630 21410 -6610 21430
rect -6630 21250 -6610 21270
rect -6630 21090 -6610 21110
rect -6630 20930 -6610 20950
rect -6550 21410 -6530 21430
rect -6550 21250 -6530 21270
rect -6550 21090 -6530 21110
rect -6550 20930 -6530 20950
rect -6470 21410 -6450 21430
rect -6470 21250 -6450 21270
rect -6470 21090 -6450 21110
rect -6470 20930 -6450 20950
rect -6390 21410 -6370 21430
rect -6390 21250 -6370 21270
rect -6390 21090 -6370 21110
rect -6390 20930 -6370 20950
rect -6310 21410 -6290 21430
rect -6310 21250 -6290 21270
rect -6310 21090 -6290 21110
rect -6310 20930 -6290 20950
rect -6230 21410 -6210 21430
rect -6230 21250 -6210 21270
rect -6230 21090 -6210 21110
rect -6230 20930 -6210 20950
rect -6150 21410 -6130 21430
rect -6150 21250 -6130 21270
rect -6150 21090 -6130 21110
rect -6150 20930 -6130 20950
rect -5670 21410 -5650 21430
rect -5670 21250 -5650 21270
rect -5670 21090 -5650 21110
rect -5670 20930 -5650 20950
rect -5590 21410 -5570 21430
rect -5590 21250 -5570 21270
rect -5590 21090 -5570 21110
rect -5590 20930 -5570 20950
rect -5510 21410 -5490 21430
rect -5510 21250 -5490 21270
rect -5510 21090 -5490 21110
rect -5510 20930 -5490 20950
rect -5430 21410 -5410 21430
rect -5430 21250 -5410 21270
rect -5430 21090 -5410 21110
rect -5430 20930 -5410 20950
rect -5350 21410 -5330 21430
rect -5350 21250 -5330 21270
rect -5350 21090 -5330 21110
rect -5350 20930 -5330 20950
rect -5270 21410 -5250 21430
rect -5270 21250 -5250 21270
rect -5270 21090 -5250 21110
rect -5270 20930 -5250 20950
rect -5190 21410 -5170 21430
rect -5190 21250 -5170 21270
rect -5190 21090 -5170 21110
rect -5190 20930 -5170 20950
rect -5110 21410 -5090 21430
rect -5110 21250 -5090 21270
rect -5110 21090 -5090 21110
rect -5110 20930 -5090 20950
rect -5030 21410 -5010 21430
rect -5030 21250 -5010 21270
rect -5030 21090 -5010 21110
rect -5030 20930 -5010 20950
rect -4950 21410 -4930 21430
rect -4950 21250 -4930 21270
rect -4950 21090 -4930 21110
rect -4950 20930 -4930 20950
rect -4870 21410 -4850 21430
rect -4870 21250 -4850 21270
rect -4870 21090 -4850 21110
rect -4870 20930 -4850 20950
rect -4790 21410 -4770 21430
rect -4790 21250 -4770 21270
rect -4790 21090 -4770 21110
rect -4790 20930 -4770 20950
rect -4710 21410 -4690 21430
rect -4710 21250 -4690 21270
rect -4710 21090 -4690 21110
rect -4710 20930 -4690 20950
rect -4630 21410 -4610 21430
rect -4630 21250 -4610 21270
rect -4630 21090 -4610 21110
rect -4630 20930 -4610 20950
rect -4550 21410 -4530 21430
rect -4550 21250 -4530 21270
rect -4550 21090 -4530 21110
rect -4550 20930 -4530 20950
rect -4470 21410 -4450 21430
rect -4470 21250 -4450 21270
rect -4470 21090 -4450 21110
rect -4470 20930 -4450 20950
rect -4390 21410 -4370 21430
rect -4390 21250 -4370 21270
rect -4390 21090 -4370 21110
rect -4390 20930 -4370 20950
rect -4310 21410 -4290 21430
rect -4310 21250 -4290 21270
rect -4310 21090 -4290 21110
rect -4310 20930 -4290 20950
rect -4230 21410 -4210 21430
rect -4230 21250 -4210 21270
rect -4230 21090 -4210 21110
rect -4230 20930 -4210 20950
rect -4150 21410 -4130 21430
rect -4150 21250 -4130 21270
rect -4150 21090 -4130 21110
rect -4150 20930 -4130 20950
rect -4070 21410 -4050 21430
rect -4070 21250 -4050 21270
rect -4070 21090 -4050 21110
rect -4070 20930 -4050 20950
rect -3990 21410 -3970 21430
rect -3990 21250 -3970 21270
rect -3990 21090 -3970 21110
rect -3990 20930 -3970 20950
rect -3910 21410 -3890 21430
rect -3910 21250 -3890 21270
rect -3910 21090 -3890 21110
rect -3910 20930 -3890 20950
rect -3830 21410 -3810 21430
rect -3830 21250 -3810 21270
rect -3830 21090 -3810 21110
rect -3830 20930 -3810 20950
rect -3750 21410 -3730 21430
rect -3750 21250 -3730 21270
rect -3750 21090 -3730 21110
rect -3750 20930 -3730 20950
rect -3670 21410 -3650 21430
rect -3670 21250 -3650 21270
rect -3670 21090 -3650 21110
rect -3670 20930 -3650 20950
rect -3590 21410 -3570 21430
rect -3590 21250 -3570 21270
rect -3590 21090 -3570 21110
rect -3590 20930 -3570 20950
rect -3510 21410 -3490 21430
rect -3510 21250 -3490 21270
rect -3510 21090 -3490 21110
rect -3510 20930 -3490 20950
rect -3430 21410 -3410 21430
rect -3430 21250 -3410 21270
rect -3430 21090 -3410 21110
rect -3430 20930 -3410 20950
rect -3350 21410 -3330 21430
rect -3350 21250 -3330 21270
rect -3350 21090 -3330 21110
rect -3350 20930 -3330 20950
rect -3270 21410 -3250 21430
rect -3270 21250 -3250 21270
rect -3270 21090 -3250 21110
rect -3270 20930 -3250 20950
rect -3190 21410 -3170 21430
rect -3190 21250 -3170 21270
rect -3190 21090 -3170 21110
rect -3190 20930 -3170 20950
rect -3110 21410 -3090 21430
rect -3110 21250 -3090 21270
rect -3110 21090 -3090 21110
rect -3110 20930 -3090 20950
rect -3030 21410 -3010 21430
rect -3030 21250 -3010 21270
rect -3030 21090 -3010 21110
rect -3030 20930 -3010 20950
rect -2950 21410 -2930 21430
rect -2950 21250 -2930 21270
rect -2950 21090 -2930 21110
rect -2950 20930 -2930 20950
rect -2870 21410 -2850 21430
rect -2870 21250 -2850 21270
rect -2870 21090 -2850 21110
rect -2870 20930 -2850 20950
rect -2790 21410 -2770 21430
rect -2790 21250 -2770 21270
rect -2790 21090 -2770 21110
rect -2790 20930 -2770 20950
rect -2710 21410 -2690 21430
rect -2710 21250 -2690 21270
rect -2710 21090 -2690 21110
rect -2710 20930 -2690 20950
rect -2630 21410 -2610 21430
rect -2630 21250 -2610 21270
rect -2630 21090 -2610 21110
rect -2630 20930 -2610 20950
rect -2550 21410 -2530 21430
rect -2550 21250 -2530 21270
rect -2550 21090 -2530 21110
rect -2550 20930 -2530 20950
rect -2470 21410 -2450 21430
rect -2470 21250 -2450 21270
rect -2470 21090 -2450 21110
rect -2470 20930 -2450 20950
rect -2390 21410 -2370 21430
rect -2390 21250 -2370 21270
rect -2390 21090 -2370 21110
rect -2390 20930 -2370 20950
rect -2310 21410 -2290 21430
rect -2310 21250 -2290 21270
rect -2310 21090 -2290 21110
rect -2310 20930 -2290 20950
rect -2230 21410 -2210 21430
rect -2230 21250 -2210 21270
rect -2230 21090 -2210 21110
rect -2230 20930 -2210 20950
rect -2150 21410 -2130 21430
rect -2150 21250 -2130 21270
rect -2150 21090 -2130 21110
rect -2150 20930 -2130 20950
rect -2070 21410 -2050 21430
rect -2070 21250 -2050 21270
rect -2070 21090 -2050 21110
rect -2070 20930 -2050 20950
rect -1990 21410 -1970 21430
rect -1990 21250 -1970 21270
rect -1990 21090 -1970 21110
rect -1990 20930 -1970 20950
rect -16550 20650 -16530 20670
rect -16550 20490 -16530 20510
rect -16470 20650 -16450 20670
rect -16470 20490 -16450 20510
rect -16390 20650 -16370 20670
rect -16390 20490 -16370 20510
rect -16310 20650 -16290 20670
rect -16310 20490 -16290 20510
rect -16230 20650 -16210 20670
rect -16230 20490 -16210 20510
rect -16150 20650 -16130 20670
rect -16150 20490 -16130 20510
rect -16070 20650 -16050 20670
rect -16070 20490 -16050 20510
rect -15990 20650 -15970 20670
rect -15990 20490 -15970 20510
rect -15910 20650 -15890 20670
rect -15910 20490 -15890 20510
rect -15830 20650 -15810 20670
rect -15830 20490 -15810 20510
rect -15750 20650 -15730 20670
rect -15750 20490 -15730 20510
rect -15670 20650 -15650 20670
rect -15670 20490 -15650 20510
rect -15590 20650 -15570 20670
rect -15590 20490 -15570 20510
rect -14950 20650 -14930 20670
rect -14950 20490 -14930 20510
rect -14870 20650 -14850 20670
rect -14870 20490 -14850 20510
rect -14790 20650 -14770 20670
rect -14790 20490 -14770 20510
rect -14710 20650 -14690 20670
rect -14710 20490 -14690 20510
rect -14630 20650 -14610 20670
rect -14630 20490 -14610 20510
rect -14550 20650 -14530 20670
rect -14550 20490 -14530 20510
rect -14470 20650 -14450 20670
rect -14470 20490 -14450 20510
rect -14390 20650 -14370 20670
rect -14390 20490 -14370 20510
rect -14310 20650 -14290 20670
rect -14310 20490 -14290 20510
rect -14230 20650 -14210 20670
rect -14230 20490 -14210 20510
rect -14150 20650 -14130 20670
rect -14150 20490 -14130 20510
rect -14070 20650 -14050 20670
rect -14070 20490 -14050 20510
rect -13990 20650 -13970 20670
rect -13990 20490 -13970 20510
rect -13910 20650 -13890 20670
rect -13910 20490 -13890 20510
rect -13830 20650 -13810 20670
rect -13830 20490 -13810 20510
rect -13750 20650 -13730 20670
rect -13750 20490 -13730 20510
rect -13670 20650 -13650 20670
rect -13670 20490 -13650 20510
rect -13590 20650 -13570 20670
rect -13590 20490 -13570 20510
rect -13510 20650 -13490 20670
rect -13510 20490 -13490 20510
rect -13430 20650 -13410 20670
rect -13430 20490 -13410 20510
rect -13350 20650 -13330 20670
rect -13350 20490 -13330 20510
rect -13270 20650 -13250 20670
rect -13270 20490 -13250 20510
rect -13190 20650 -13170 20670
rect -13190 20490 -13170 20510
rect -13110 20650 -13090 20670
rect -13110 20490 -13090 20510
rect -13030 20650 -13010 20670
rect -13030 20490 -13010 20510
rect -12950 20650 -12930 20670
rect -12950 20490 -12930 20510
rect -12870 20650 -12850 20670
rect -12870 20490 -12850 20510
rect -12790 20650 -12770 20670
rect -12790 20490 -12770 20510
rect -12710 20650 -12690 20670
rect -12710 20490 -12690 20510
rect -12630 20650 -12610 20670
rect -12630 20490 -12610 20510
rect -12550 20650 -12530 20670
rect -12550 20490 -12530 20510
rect -12470 20650 -12450 20670
rect -12470 20490 -12450 20510
rect -12390 20650 -12370 20670
rect -12390 20490 -12370 20510
rect -12310 20650 -12290 20670
rect -12310 20490 -12290 20510
rect -12230 20650 -12210 20670
rect -12230 20490 -12210 20510
rect -12150 20650 -12130 20670
rect -12150 20490 -12130 20510
rect -12070 20650 -12050 20670
rect -12070 20490 -12050 20510
rect -11990 20650 -11970 20670
rect -11990 20490 -11970 20510
rect -11910 20650 -11890 20670
rect -11910 20490 -11890 20510
rect -11830 20650 -11810 20670
rect -11830 20490 -11810 20510
rect -11750 20650 -11730 20670
rect -11750 20490 -11730 20510
rect -11670 20650 -11650 20670
rect -11670 20490 -11650 20510
rect -11590 20650 -11570 20670
rect -11590 20490 -11570 20510
rect -11510 20650 -11490 20670
rect -11510 20490 -11490 20510
rect -11430 20650 -11410 20670
rect -11430 20490 -11410 20510
rect -11350 20650 -11330 20670
rect -11350 20490 -11330 20510
rect -11270 20650 -11250 20670
rect -11270 20490 -11250 20510
rect -11190 20650 -11170 20670
rect -11190 20490 -11170 20510
rect -11110 20650 -11090 20670
rect -11110 20490 -11090 20510
rect -11030 20650 -11010 20670
rect -11030 20490 -11010 20510
rect -10950 20650 -10930 20670
rect -10950 20490 -10930 20510
rect -10870 20650 -10850 20670
rect -10870 20490 -10850 20510
rect -10790 20650 -10770 20670
rect -10790 20490 -10770 20510
rect -10710 20650 -10690 20670
rect -10710 20490 -10690 20510
rect -10630 20650 -10610 20670
rect -10630 20490 -10610 20510
rect -10550 20650 -10530 20670
rect -10550 20490 -10530 20510
rect -10470 20650 -10450 20670
rect -10470 20490 -10450 20510
rect -10390 20650 -10370 20670
rect -10390 20490 -10370 20510
rect -10310 20650 -10290 20670
rect -10310 20490 -10290 20510
rect -10230 20650 -10210 20670
rect -10230 20490 -10210 20510
rect -10150 20650 -10130 20670
rect -10150 20490 -10130 20510
rect -10070 20650 -10050 20670
rect -10070 20490 -10050 20510
rect -9990 20650 -9970 20670
rect -9990 20490 -9970 20510
rect -9910 20650 -9890 20670
rect -9910 20490 -9890 20510
rect -9830 20650 -9810 20670
rect -9830 20490 -9810 20510
rect -9750 20650 -9730 20670
rect -9750 20490 -9730 20510
rect -9670 20650 -9650 20670
rect -9670 20490 -9650 20510
rect -9590 20650 -9570 20670
rect -9590 20490 -9570 20510
rect -9510 20650 -9490 20670
rect -9510 20490 -9490 20510
rect -9430 20650 -9410 20670
rect -9430 20490 -9410 20510
rect -9350 20650 -9330 20670
rect -9350 20490 -9330 20510
rect -9270 20650 -9250 20670
rect -9270 20490 -9250 20510
rect -9190 20650 -9170 20670
rect -9190 20490 -9170 20510
rect -9110 20650 -9090 20670
rect -9110 20490 -9090 20510
rect -9030 20650 -9010 20670
rect -9030 20490 -9010 20510
rect -8950 20650 -8930 20670
rect -8950 20490 -8930 20510
rect -8870 20650 -8850 20670
rect -8870 20490 -8850 20510
rect -8790 20650 -8770 20670
rect -8790 20490 -8770 20510
rect -8710 20650 -8690 20670
rect -8710 20490 -8690 20510
rect -8630 20650 -8610 20670
rect -8630 20490 -8610 20510
rect -8550 20650 -8530 20670
rect -8550 20490 -8530 20510
rect -8470 20650 -8450 20670
rect -8470 20490 -8450 20510
rect -8390 20650 -8370 20670
rect -8390 20490 -8370 20510
rect -8310 20650 -8290 20670
rect -8310 20490 -8290 20510
rect -8230 20650 -8210 20670
rect -8230 20490 -8210 20510
rect -8150 20650 -8130 20670
rect -8150 20490 -8130 20510
rect -8070 20650 -8050 20670
rect -8070 20490 -8050 20510
rect -7990 20650 -7970 20670
rect -7990 20490 -7970 20510
rect -7910 20650 -7890 20670
rect -7910 20490 -7890 20510
rect -7830 20650 -7810 20670
rect -7830 20490 -7810 20510
rect -7750 20650 -7730 20670
rect -7750 20490 -7730 20510
rect -7670 20650 -7650 20670
rect -7670 20490 -7650 20510
rect -7590 20650 -7570 20670
rect -7590 20490 -7570 20510
rect -7510 20650 -7490 20670
rect -7510 20490 -7490 20510
rect -7430 20650 -7410 20670
rect -7430 20490 -7410 20510
rect -7350 20650 -7330 20670
rect -7350 20490 -7330 20510
rect -7270 20650 -7250 20670
rect -7270 20490 -7250 20510
rect -7190 20650 -7170 20670
rect -7190 20490 -7170 20510
rect -7110 20650 -7090 20670
rect -7110 20490 -7090 20510
rect -7030 20650 -7010 20670
rect -7030 20490 -7010 20510
rect -6950 20650 -6930 20670
rect -6950 20490 -6930 20510
rect -6870 20650 -6850 20670
rect -6870 20490 -6850 20510
rect -6790 20650 -6770 20670
rect -6790 20490 -6770 20510
rect -6710 20650 -6690 20670
rect -6710 20490 -6690 20510
rect -6630 20650 -6610 20670
rect -6630 20490 -6610 20510
rect -6550 20650 -6530 20670
rect -6550 20490 -6530 20510
rect -6470 20650 -6450 20670
rect -6470 20490 -6450 20510
rect -6390 20650 -6370 20670
rect -6390 20490 -6370 20510
rect -6310 20650 -6290 20670
rect -6310 20490 -6290 20510
rect -6230 20650 -6210 20670
rect -6230 20490 -6210 20510
rect -6150 20650 -6130 20670
rect -6150 20490 -6130 20510
rect -5670 20650 -5650 20670
rect -5670 20490 -5650 20510
rect -5590 20650 -5570 20670
rect -5590 20490 -5570 20510
rect -5510 20650 -5490 20670
rect -5510 20490 -5490 20510
rect -5430 20650 -5410 20670
rect -5430 20490 -5410 20510
rect -5350 20650 -5330 20670
rect -5350 20490 -5330 20510
rect -5270 20650 -5250 20670
rect -5270 20490 -5250 20510
rect -5190 20650 -5170 20670
rect -5190 20490 -5170 20510
rect -5110 20650 -5090 20670
rect -5110 20490 -5090 20510
rect -5030 20650 -5010 20670
rect -5030 20490 -5010 20510
rect -4950 20650 -4930 20670
rect -4950 20490 -4930 20510
rect -4870 20650 -4850 20670
rect -4870 20490 -4850 20510
rect -4790 20650 -4770 20670
rect -4790 20490 -4770 20510
rect -4710 20650 -4690 20670
rect -4710 20490 -4690 20510
rect -4630 20650 -4610 20670
rect -4630 20490 -4610 20510
rect -4550 20650 -4530 20670
rect -4550 20490 -4530 20510
rect -4470 20650 -4450 20670
rect -4470 20490 -4450 20510
rect -4390 20650 -4370 20670
rect -4390 20490 -4370 20510
rect -4310 20650 -4290 20670
rect -4310 20490 -4290 20510
rect -4230 20650 -4210 20670
rect -4230 20490 -4210 20510
rect -4150 20650 -4130 20670
rect -4150 20490 -4130 20510
rect -4070 20650 -4050 20670
rect -4070 20490 -4050 20510
rect -3990 20650 -3970 20670
rect -3990 20490 -3970 20510
rect -3910 20650 -3890 20670
rect -3910 20490 -3890 20510
rect -3830 20650 -3810 20670
rect -3830 20490 -3810 20510
rect -3750 20650 -3730 20670
rect -3750 20490 -3730 20510
rect -3670 20650 -3650 20670
rect -3670 20490 -3650 20510
rect -3590 20650 -3570 20670
rect -3590 20490 -3570 20510
rect -3510 20650 -3490 20670
rect -3510 20490 -3490 20510
rect -3430 20650 -3410 20670
rect -3430 20490 -3410 20510
rect -3350 20650 -3330 20670
rect -3350 20490 -3330 20510
rect -3270 20650 -3250 20670
rect -3270 20490 -3250 20510
rect -3190 20650 -3170 20670
rect -3190 20490 -3170 20510
rect -3110 20650 -3090 20670
rect -3110 20490 -3090 20510
rect -3030 20650 -3010 20670
rect -3030 20490 -3010 20510
rect -2950 20650 -2930 20670
rect -2950 20490 -2930 20510
rect -2870 20650 -2850 20670
rect -2870 20490 -2850 20510
rect -2790 20650 -2770 20670
rect -2790 20490 -2770 20510
rect -2710 20650 -2690 20670
rect -2710 20490 -2690 20510
rect -2630 20650 -2610 20670
rect -2630 20490 -2610 20510
rect -2550 20650 -2530 20670
rect -2550 20490 -2530 20510
rect -2470 20650 -2450 20670
rect -2470 20490 -2450 20510
rect -2390 20650 -2370 20670
rect -2390 20490 -2370 20510
rect -2310 20650 -2290 20670
rect -2310 20490 -2290 20510
rect -2230 20650 -2210 20670
rect -2230 20490 -2210 20510
rect -2150 20650 -2130 20670
rect -2150 20490 -2130 20510
rect -2070 20650 -2050 20670
rect -2070 20490 -2050 20510
rect -1990 20650 -1970 20670
rect -1990 20490 -1970 20510
rect -1830 21410 -1810 21430
rect -1830 21250 -1810 21270
rect -1830 21090 -1810 21110
rect -1830 20930 -1810 20950
rect -1750 21410 -1730 21430
rect -1750 21250 -1730 21270
rect -1750 21090 -1730 21110
rect -1750 20930 -1730 20950
rect -1670 21410 -1650 21430
rect -1670 21250 -1650 21270
rect -1670 21090 -1650 21110
rect -1670 20930 -1650 20950
rect -1510 21410 -1490 21430
rect -1510 21250 -1490 21270
rect -1510 21090 -1490 21110
rect -1510 20930 -1490 20950
rect -1350 21410 -1330 21430
rect -1350 21250 -1330 21270
rect -1350 21090 -1330 21110
rect -1350 20930 -1330 20950
rect -1270 21410 -1250 21430
rect -1270 21250 -1250 21270
rect -1270 21090 -1250 21110
rect -1270 20930 -1250 20950
rect -1190 21410 -1170 21430
rect -1190 21250 -1170 21270
rect -1190 21090 -1170 21110
rect -1190 20930 -1170 20950
rect -1110 21410 -1090 21430
rect -1110 21250 -1090 21270
rect -1110 21090 -1090 21110
rect -1110 20930 -1090 20950
rect -1030 21410 -1010 21430
rect -1030 21250 -1010 21270
rect -1030 21090 -1010 21110
rect -1030 20930 -1010 20950
rect -870 21410 -850 21430
rect -870 21250 -850 21270
rect -870 21090 -850 21110
rect -870 20930 -850 20950
rect -710 21410 -690 21430
rect -710 21250 -690 21270
rect -710 21090 -690 21110
rect -710 20930 -690 20950
rect -550 21410 -530 21430
rect -550 21250 -530 21270
rect -550 21090 -530 21110
rect -550 20930 -530 20950
rect -1910 20650 -1890 20670
rect -1910 20490 -1890 20510
rect -5270 20330 -5250 20350
rect -5270 20170 -5250 20190
rect -5110 20330 -5090 20350
rect -5110 20170 -5090 20190
rect -5030 20330 -5010 20350
rect -5030 20170 -5010 20190
rect -4950 20330 -4930 20350
rect -4950 20170 -4930 20190
rect -4870 20330 -4850 20350
rect -4870 20170 -4850 20190
rect -4790 20330 -4770 20350
rect -4790 20170 -4770 20190
rect -4710 20330 -4690 20350
rect -4710 20170 -4690 20190
rect -4630 20330 -4610 20350
rect -4630 20170 -4610 20190
rect -4550 20330 -4530 20350
rect -4550 20170 -4530 20190
rect -4470 20330 -4450 20350
rect -4470 20170 -4450 20190
rect -4390 20330 -4370 20350
rect -4390 20170 -4370 20190
rect -4310 20330 -4290 20350
rect -4310 20170 -4290 20190
rect -4230 20330 -4210 20350
rect -4230 20170 -4210 20190
rect -4150 20330 -4130 20350
rect -4150 20170 -4130 20190
rect -4070 20330 -4050 20350
rect -4070 20170 -4050 20190
rect -3990 20330 -3970 20350
rect -3990 20170 -3970 20190
rect -3910 20330 -3890 20350
rect -3910 20170 -3890 20190
rect -3830 20330 -3810 20350
rect -3830 20170 -3810 20190
rect -3750 20330 -3730 20350
rect -3750 20170 -3730 20190
rect -3670 20330 -3650 20350
rect -3670 20170 -3650 20190
rect -3590 20330 -3570 20350
rect -3590 20170 -3570 20190
rect -3510 20330 -3490 20350
rect -3510 20170 -3490 20190
rect -3430 20330 -3410 20350
rect -3430 20170 -3410 20190
rect -3350 20330 -3330 20350
rect -3350 20170 -3330 20190
rect -3270 20330 -3250 20350
rect -3270 20170 -3250 20190
rect -3190 20330 -3170 20350
rect -3190 20170 -3170 20190
rect -3110 20330 -3090 20350
rect -3110 20170 -3090 20190
rect -3030 20330 -3010 20350
rect -3030 20170 -3010 20190
rect -2950 20330 -2930 20350
rect -2950 20170 -2930 20190
rect -2870 20330 -2850 20350
rect -2870 20170 -2850 20190
rect -2790 20330 -2770 20350
rect -2790 20170 -2770 20190
rect -2710 20330 -2690 20350
rect -2710 20170 -2690 20190
rect -2630 20330 -2610 20350
rect -2630 20170 -2610 20190
rect -2550 20330 -2530 20350
rect -2550 20170 -2530 20190
rect -2470 20330 -2450 20350
rect -2470 20170 -2450 20190
rect -2390 20330 -2370 20350
rect -2390 20170 -2370 20190
rect -2310 20330 -2290 20350
rect -2310 20170 -2290 20190
rect -2230 20330 -2210 20350
rect -2230 20170 -2210 20190
rect -2150 20330 -2130 20350
rect -2150 20170 -2130 20190
rect -2070 20330 -2050 20350
rect -2070 20170 -2050 20190
rect -1990 20330 -1970 20350
rect -1990 20170 -1970 20190
rect -1830 20650 -1810 20670
rect -1830 20490 -1810 20510
rect -1750 20650 -1730 20670
rect -1750 20490 -1730 20510
rect 20530 20650 20550 20670
rect 20530 20490 20550 20510
rect 20610 20650 20630 20670
rect 20610 20490 20630 20510
rect 20690 20650 20710 20670
rect 20690 20490 20710 20510
rect 20770 20650 20790 20670
rect 20770 20490 20790 20510
rect 20850 20650 20870 20670
rect 20850 20490 20870 20510
rect 20930 20650 20950 20670
rect 20930 20490 20950 20510
rect 21010 20650 21030 20670
rect 21010 20490 21030 20510
rect 21090 20650 21110 20670
rect 21090 20490 21110 20510
rect 21170 20650 21190 20670
rect 21170 20490 21190 20510
rect 21250 20650 21270 20670
rect 21250 20490 21270 20510
rect 21330 20650 21350 20670
rect 21330 20490 21350 20510
rect 21410 20650 21430 20670
rect 21410 20490 21430 20510
rect 21490 20650 21510 20670
rect 21490 20490 21510 20510
rect 21570 20650 21590 20670
rect 21570 20490 21590 20510
rect -1830 20330 -1810 20350
rect -1830 20170 -1810 20190
rect -1750 20330 -1730 20350
rect -1750 20170 -1730 20190
rect 20530 20010 20550 20030
rect 20530 19850 20550 19870
rect 20610 20010 20630 20030
rect 20610 19850 20630 19870
rect 20690 20010 20710 20030
rect 20690 19850 20710 19870
rect 20770 20010 20790 20030
rect 20770 19850 20790 19870
rect 20850 20010 20870 20030
rect 20850 19850 20870 19870
rect 20930 20010 20950 20030
rect 20930 19850 20950 19870
rect 21010 20010 21030 20030
rect 21010 19850 21030 19870
rect 21090 20010 21110 20030
rect 21090 19850 21110 19870
rect 21170 20010 21190 20030
rect 21170 19850 21190 19870
rect 21250 20010 21270 20030
rect 21250 19850 21270 19870
rect 21330 20010 21350 20030
rect 21330 19850 21350 19870
rect 21410 20010 21430 20030
rect 21410 19850 21430 19870
rect 21490 20010 21510 20030
rect 21490 19850 21510 19870
rect 21570 20010 21590 20030
rect 21570 19850 21590 19870
rect -16550 18850 -16530 18870
rect -16550 18690 -16530 18710
rect -16550 18530 -16530 18550
rect -16470 18850 -16450 18870
rect -16470 18690 -16450 18710
rect -16470 18530 -16450 18550
rect -16390 18850 -16370 18870
rect -16390 18690 -16370 18710
rect -16390 18530 -16370 18550
rect -16310 18850 -16290 18870
rect -16310 18690 -16290 18710
rect -16310 18530 -16290 18550
rect -16230 18850 -16210 18870
rect -16230 18690 -16210 18710
rect -16230 18530 -16210 18550
rect -16150 18850 -16130 18870
rect -16150 18690 -16130 18710
rect -16150 18530 -16130 18550
rect -16070 18850 -16050 18870
rect -16070 18690 -16050 18710
rect -16070 18530 -16050 18550
rect -15990 18850 -15970 18870
rect -15990 18690 -15970 18710
rect -15990 18530 -15970 18550
rect -15910 18850 -15890 18870
rect -15910 18690 -15890 18710
rect -15910 18530 -15890 18550
rect -15830 18850 -15810 18870
rect -15830 18690 -15810 18710
rect -15830 18530 -15810 18550
rect -15750 18850 -15730 18870
rect -15750 18690 -15730 18710
rect -15750 18530 -15730 18550
rect -15670 18850 -15650 18870
rect -15670 18690 -15650 18710
rect -15670 18530 -15650 18550
rect -15590 18850 -15570 18870
rect -15590 18690 -15570 18710
rect -15590 18530 -15570 18550
rect 20530 18010 20550 18030
rect 20530 17850 20550 17870
rect 20610 18010 20630 18030
rect 20610 17850 20630 17870
rect 20690 18010 20710 18030
rect 20690 17850 20710 17870
rect 20770 18010 20790 18030
rect 20770 17850 20790 17870
rect 20850 18010 20870 18030
rect 20850 17850 20870 17870
rect 20930 18010 20950 18030
rect 20930 17850 20950 17870
rect 21010 18010 21030 18030
rect 21010 17850 21030 17870
rect 21090 18010 21110 18030
rect 21090 17850 21110 17870
rect 21170 18010 21190 18030
rect 21170 17850 21190 17870
rect 21250 18010 21270 18030
rect 21250 17850 21270 17870
rect 21330 18010 21350 18030
rect 21330 17850 21350 17870
rect 21410 18010 21430 18030
rect 21410 17850 21430 17870
rect 21490 18010 21510 18030
rect 21490 17850 21510 17870
rect 21570 18010 21590 18030
rect 21570 17850 21590 17870
rect -16550 17330 -16530 17350
rect -16550 17170 -16530 17190
rect -16470 17330 -16450 17350
rect -16470 17170 -16450 17190
rect -16390 17330 -16370 17350
rect -16390 17170 -16370 17190
rect -16310 17330 -16290 17350
rect -16310 17170 -16290 17190
rect -16230 17330 -16210 17350
rect -16230 17170 -16210 17190
rect -16150 17330 -16130 17350
rect -16150 17170 -16130 17190
rect -16070 17330 -16050 17350
rect -16070 17170 -16050 17190
rect -15990 17330 -15970 17350
rect -15990 17170 -15970 17190
rect -15910 17330 -15890 17350
rect -15910 17170 -15890 17190
rect -15830 17330 -15810 17350
rect -15830 17170 -15810 17190
rect -15750 17330 -15730 17350
rect -15750 17170 -15730 17190
rect -15670 17330 -15650 17350
rect -15670 17170 -15650 17190
rect -15590 17330 -15570 17350
rect -15590 17170 -15570 17190
rect -14950 17330 -14930 17350
rect -14950 17170 -14930 17190
rect -14870 17330 -14850 17350
rect -14870 17170 -14850 17190
rect -14790 17330 -14770 17350
rect -14790 17170 -14770 17190
rect -14710 17330 -14690 17350
rect -14710 17170 -14690 17190
rect -14630 17330 -14610 17350
rect -14630 17170 -14610 17190
rect -14550 17330 -14530 17350
rect -14550 17170 -14530 17190
rect -14470 17330 -14450 17350
rect -14470 17170 -14450 17190
rect -14390 17330 -14370 17350
rect -14390 17170 -14370 17190
rect -14310 17330 -14290 17350
rect -14310 17170 -14290 17190
rect -14230 17330 -14210 17350
rect -14230 17170 -14210 17190
rect -14150 17330 -14130 17350
rect -14150 17170 -14130 17190
rect -14070 17330 -14050 17350
rect -14070 17170 -14050 17190
rect -13990 17330 -13970 17350
rect -13990 17170 -13970 17190
rect -13910 17330 -13890 17350
rect -13910 17170 -13890 17190
rect -13830 17330 -13810 17350
rect -13830 17170 -13810 17190
rect -13750 17330 -13730 17350
rect -13750 17170 -13730 17190
rect -13670 17330 -13650 17350
rect -13670 17170 -13650 17190
rect -13590 17330 -13570 17350
rect -13590 17170 -13570 17190
rect -13510 17330 -13490 17350
rect -13510 17170 -13490 17190
rect -13430 17330 -13410 17350
rect -13430 17170 -13410 17190
rect -13350 17330 -13330 17350
rect -13350 17170 -13330 17190
rect -13270 17330 -13250 17350
rect -13270 17170 -13250 17190
rect -13190 17330 -13170 17350
rect -13190 17170 -13170 17190
rect -13110 17330 -13090 17350
rect -13110 17170 -13090 17190
rect -13030 17330 -13010 17350
rect -13030 17170 -13010 17190
rect -12950 17330 -12930 17350
rect -12950 17170 -12930 17190
rect -12870 17330 -12850 17350
rect -12870 17170 -12850 17190
rect -12790 17330 -12770 17350
rect -12790 17170 -12770 17190
rect -12710 17330 -12690 17350
rect -12710 17170 -12690 17190
rect -12630 17330 -12610 17350
rect -12630 17170 -12610 17190
rect -12550 17330 -12530 17350
rect -12550 17170 -12530 17190
rect -12470 17330 -12450 17350
rect -12470 17170 -12450 17190
rect -12390 17330 -12370 17350
rect -12390 17170 -12370 17190
rect -12310 17330 -12290 17350
rect -12310 17170 -12290 17190
rect -12230 17330 -12210 17350
rect -12230 17170 -12210 17190
rect -12150 17330 -12130 17350
rect -12150 17170 -12130 17190
rect -12070 17330 -12050 17350
rect -12070 17170 -12050 17190
rect -11990 17330 -11970 17350
rect -11990 17170 -11970 17190
rect -11910 17330 -11890 17350
rect -11910 17170 -11890 17190
rect -11830 17330 -11810 17350
rect -11830 17170 -11810 17190
rect -11750 17330 -11730 17350
rect -11750 17170 -11730 17190
rect -11670 17330 -11650 17350
rect -11670 17170 -11650 17190
rect -11590 17330 -11570 17350
rect -11590 17170 -11570 17190
rect -11510 17330 -11490 17350
rect -11510 17170 -11490 17190
rect -11430 17330 -11410 17350
rect -11430 17170 -11410 17190
rect -11350 17330 -11330 17350
rect -11350 17170 -11330 17190
rect -11270 17330 -11250 17350
rect -11270 17170 -11250 17190
rect -11190 17330 -11170 17350
rect -11190 17170 -11170 17190
rect -11110 17330 -11090 17350
rect -11110 17170 -11090 17190
rect -11030 17330 -11010 17350
rect -11030 17170 -11010 17190
rect -10950 17330 -10930 17350
rect -10950 17170 -10930 17190
rect -10870 17330 -10850 17350
rect -10870 17170 -10850 17190
rect -10790 17330 -10770 17350
rect -10790 17170 -10770 17190
rect -10710 17330 -10690 17350
rect -10710 17170 -10690 17190
rect -10630 17330 -10610 17350
rect -10630 17170 -10610 17190
rect -10550 17330 -10530 17350
rect -10550 17170 -10530 17190
rect -10470 17330 -10450 17350
rect -10470 17170 -10450 17190
rect -10390 17330 -10370 17350
rect -10390 17170 -10370 17190
rect -10310 17330 -10290 17350
rect -10310 17170 -10290 17190
rect -10230 17330 -10210 17350
rect -10230 17170 -10210 17190
rect -10150 17330 -10130 17350
rect -10150 17170 -10130 17190
rect -10070 17330 -10050 17350
rect -10070 17170 -10050 17190
rect -9990 17330 -9970 17350
rect -9990 17170 -9970 17190
rect -9910 17330 -9890 17350
rect -9910 17170 -9890 17190
rect -9830 17330 -9810 17350
rect -9830 17170 -9810 17190
rect -9750 17330 -9730 17350
rect -9750 17170 -9730 17190
rect -9670 17330 -9650 17350
rect -9670 17170 -9650 17190
rect -9590 17330 -9570 17350
rect -9590 17170 -9570 17190
rect -9510 17330 -9490 17350
rect -9510 17170 -9490 17190
rect -9430 17330 -9410 17350
rect -9430 17170 -9410 17190
rect -9350 17330 -9330 17350
rect -9350 17170 -9330 17190
rect -9270 17330 -9250 17350
rect -9270 17170 -9250 17190
rect -9190 17330 -9170 17350
rect -9190 17170 -9170 17190
rect -9110 17330 -9090 17350
rect -9110 17170 -9090 17190
rect -9030 17330 -9010 17350
rect -9030 17170 -9010 17190
rect -8950 17330 -8930 17350
rect -8950 17170 -8930 17190
rect -8870 17330 -8850 17350
rect -8870 17170 -8850 17190
rect -8790 17330 -8770 17350
rect -8790 17170 -8770 17190
rect -8710 17330 -8690 17350
rect -8710 17170 -8690 17190
rect -8630 17330 -8610 17350
rect -8630 17170 -8610 17190
rect -8550 17330 -8530 17350
rect -8550 17170 -8530 17190
rect -8470 17330 -8450 17350
rect -8470 17170 -8450 17190
rect -8390 17330 -8370 17350
rect -8390 17170 -8370 17190
rect -8310 17330 -8290 17350
rect -8310 17170 -8290 17190
rect -8230 17330 -8210 17350
rect -8230 17170 -8210 17190
rect -8150 17330 -8130 17350
rect -8150 17170 -8130 17190
rect -8070 17330 -8050 17350
rect -8070 17170 -8050 17190
rect -7990 17330 -7970 17350
rect -7990 17170 -7970 17190
rect -7910 17330 -7890 17350
rect -7910 17170 -7890 17190
rect -7830 17330 -7810 17350
rect -7830 17170 -7810 17190
rect -7750 17330 -7730 17350
rect -7750 17170 -7730 17190
rect -7670 17330 -7650 17350
rect -7670 17170 -7650 17190
rect -7590 17330 -7570 17350
rect -7590 17170 -7570 17190
rect -7510 17330 -7490 17350
rect -7510 17170 -7490 17190
rect -7430 17330 -7410 17350
rect -7430 17170 -7410 17190
rect -7350 17330 -7330 17350
rect -7350 17170 -7330 17190
rect -7270 17330 -7250 17350
rect -7270 17170 -7250 17190
rect -7190 17330 -7170 17350
rect -7190 17170 -7170 17190
rect -7110 17330 -7090 17350
rect -7110 17170 -7090 17190
rect -7030 17330 -7010 17350
rect -7030 17170 -7010 17190
rect -6950 17330 -6930 17350
rect -6950 17170 -6930 17190
rect -6870 17330 -6850 17350
rect -6870 17170 -6850 17190
rect -6790 17330 -6770 17350
rect -6790 17170 -6770 17190
rect -6710 17330 -6690 17350
rect -6710 17170 -6690 17190
rect -6630 17330 -6610 17350
rect -6630 17170 -6610 17190
rect -6550 17330 -6530 17350
rect -6550 17170 -6530 17190
rect -6470 17330 -6450 17350
rect -6470 17170 -6450 17190
rect -6390 17330 -6370 17350
rect -6390 17170 -6370 17190
rect -6310 17330 -6290 17350
rect -6310 17170 -6290 17190
rect -6230 17330 -6210 17350
rect -6230 17170 -6210 17190
rect -6150 17330 -6130 17350
rect -6150 17170 -6130 17190
rect -6070 17330 -6050 17350
rect -6070 17170 -6050 17190
rect -5990 17330 -5970 17350
rect -5990 17170 -5970 17190
rect -5910 17330 -5890 17350
rect -5910 17170 -5890 17190
rect -5830 17330 -5810 17350
rect -5830 17170 -5810 17190
rect -5750 17330 -5730 17350
rect -5750 17170 -5730 17190
rect -5430 17330 -5410 17350
rect -5430 17170 -5410 17190
rect -5270 17330 -5250 17350
rect -5270 17170 -5250 17190
rect -14950 16450 -14930 16470
rect -14950 16290 -14930 16310
rect -14950 16130 -14930 16150
rect -14950 15970 -14930 15990
rect -14870 16450 -14850 16470
rect -14870 16290 -14850 16310
rect -14870 16130 -14850 16150
rect -14870 15970 -14850 15990
rect -14790 16450 -14770 16470
rect -14790 16290 -14770 16310
rect -14790 16130 -14770 16150
rect -14790 15970 -14770 15990
rect -14710 16450 -14690 16470
rect -14710 16290 -14690 16310
rect -14710 16130 -14690 16150
rect -14710 15970 -14690 15990
rect -14630 16450 -14610 16470
rect -14630 16290 -14610 16310
rect -14630 16130 -14610 16150
rect -14630 15970 -14610 15990
rect -14550 16450 -14530 16470
rect -14550 16290 -14530 16310
rect -14550 16130 -14530 16150
rect -14550 15970 -14530 15990
rect -14470 16450 -14450 16470
rect -14470 16290 -14450 16310
rect -14470 16130 -14450 16150
rect -14470 15970 -14450 15990
rect -14390 16450 -14370 16470
rect -14390 16290 -14370 16310
rect -14390 16130 -14370 16150
rect -14390 15970 -14370 15990
rect -14310 16450 -14290 16470
rect -14310 16290 -14290 16310
rect -14310 16130 -14290 16150
rect -14310 15970 -14290 15990
rect -14230 16450 -14210 16470
rect -14230 16290 -14210 16310
rect -14230 16130 -14210 16150
rect -14230 15970 -14210 15990
rect -14150 16450 -14130 16470
rect -14150 16290 -14130 16310
rect -14150 16130 -14130 16150
rect -14150 15970 -14130 15990
rect -14070 16450 -14050 16470
rect -14070 16290 -14050 16310
rect -14070 16130 -14050 16150
rect -14070 15970 -14050 15990
rect -13990 16450 -13970 16470
rect -13990 16290 -13970 16310
rect -13990 16130 -13970 16150
rect -13990 15970 -13970 15990
rect -13910 16450 -13890 16470
rect -13910 16290 -13890 16310
rect -13910 16130 -13890 16150
rect -13910 15970 -13890 15990
rect -13830 16450 -13810 16470
rect -13830 16290 -13810 16310
rect -13830 16130 -13810 16150
rect -13830 15970 -13810 15990
rect -13750 16450 -13730 16470
rect -13750 16290 -13730 16310
rect -13750 16130 -13730 16150
rect -13750 15970 -13730 15990
rect -13670 16450 -13650 16470
rect -13670 16290 -13650 16310
rect -13670 16130 -13650 16150
rect -13670 15970 -13650 15990
rect -13590 16450 -13570 16470
rect -13590 16290 -13570 16310
rect -13590 16130 -13570 16150
rect -13590 15970 -13570 15990
rect -13510 16450 -13490 16470
rect -13510 16290 -13490 16310
rect -13510 16130 -13490 16150
rect -13510 15970 -13490 15990
rect -13430 16450 -13410 16470
rect -13430 16290 -13410 16310
rect -13430 16130 -13410 16150
rect -13430 15970 -13410 15990
rect -13350 16450 -13330 16470
rect -13350 16290 -13330 16310
rect -13350 16130 -13330 16150
rect -13350 15970 -13330 15990
rect -13270 16450 -13250 16470
rect -13270 16290 -13250 16310
rect -13270 16130 -13250 16150
rect -13270 15970 -13250 15990
rect -13190 16450 -13170 16470
rect -13190 16290 -13170 16310
rect -13190 16130 -13170 16150
rect -13190 15970 -13170 15990
rect -13110 16450 -13090 16470
rect -13110 16290 -13090 16310
rect -13110 16130 -13090 16150
rect -13110 15970 -13090 15990
rect -13030 16450 -13010 16470
rect -13030 16290 -13010 16310
rect -13030 16130 -13010 16150
rect -13030 15970 -13010 15990
rect -12950 16450 -12930 16470
rect -12950 16290 -12930 16310
rect -12950 16130 -12930 16150
rect -12950 15970 -12930 15990
rect -12870 16450 -12850 16470
rect -12870 16290 -12850 16310
rect -12870 16130 -12850 16150
rect -12870 15970 -12850 15990
rect -12790 16450 -12770 16470
rect -12790 16290 -12770 16310
rect -12790 16130 -12770 16150
rect -12790 15970 -12770 15990
rect -12710 16450 -12690 16470
rect -12710 16290 -12690 16310
rect -12710 16130 -12690 16150
rect -12710 15970 -12690 15990
rect -12630 16450 -12610 16470
rect -12630 16290 -12610 16310
rect -12630 16130 -12610 16150
rect -12630 15970 -12610 15990
rect -12550 16450 -12530 16470
rect -12550 16290 -12530 16310
rect -12550 16130 -12530 16150
rect -12550 15970 -12530 15990
rect -12470 16450 -12450 16470
rect -12470 16290 -12450 16310
rect -12470 16130 -12450 16150
rect -12470 15970 -12450 15990
rect -12390 16450 -12370 16470
rect -12390 16290 -12370 16310
rect -12390 16130 -12370 16150
rect -12390 15970 -12370 15990
rect -12310 16450 -12290 16470
rect -12310 16290 -12290 16310
rect -12310 16130 -12290 16150
rect -12310 15970 -12290 15990
rect -12230 16450 -12210 16470
rect -12230 16290 -12210 16310
rect -12230 16130 -12210 16150
rect -12230 15970 -12210 15990
rect -12150 16450 -12130 16470
rect -12150 16290 -12130 16310
rect -12150 16130 -12130 16150
rect -12150 15970 -12130 15990
rect -12070 16450 -12050 16470
rect -12070 16290 -12050 16310
rect -12070 16130 -12050 16150
rect -12070 15970 -12050 15990
rect -11990 16450 -11970 16470
rect -11990 16290 -11970 16310
rect -11990 16130 -11970 16150
rect -11990 15970 -11970 15990
rect -11910 16450 -11890 16470
rect -11910 16290 -11890 16310
rect -11910 16130 -11890 16150
rect -11910 15970 -11890 15990
rect -11830 16450 -11810 16470
rect -11830 16290 -11810 16310
rect -11830 16130 -11810 16150
rect -11830 15970 -11810 15990
rect -11750 16450 -11730 16470
rect -11750 16290 -11730 16310
rect -11750 16130 -11730 16150
rect -11750 15970 -11730 15990
rect -11670 16450 -11650 16470
rect -11670 16290 -11650 16310
rect -11670 16130 -11650 16150
rect -11670 15970 -11650 15990
rect -11590 16450 -11570 16470
rect -11590 16290 -11570 16310
rect -11590 16130 -11570 16150
rect -11590 15970 -11570 15990
rect -11510 16450 -11490 16470
rect -11510 16290 -11490 16310
rect -11510 16130 -11490 16150
rect -11510 15970 -11490 15990
rect -11430 16450 -11410 16470
rect -11430 16290 -11410 16310
rect -11430 16130 -11410 16150
rect -11430 15970 -11410 15990
rect -11350 16450 -11330 16470
rect -11350 16290 -11330 16310
rect -11350 16130 -11330 16150
rect -11350 15970 -11330 15990
rect -11270 16450 -11250 16470
rect -11270 16290 -11250 16310
rect -11270 16130 -11250 16150
rect -11270 15970 -11250 15990
rect -11190 16450 -11170 16470
rect -11190 16290 -11170 16310
rect -11190 16130 -11170 16150
rect -11190 15970 -11170 15990
rect -11110 16450 -11090 16470
rect -11110 16290 -11090 16310
rect -11110 16130 -11090 16150
rect -11110 15970 -11090 15990
rect -11030 16450 -11010 16470
rect -11030 16290 -11010 16310
rect -11030 16130 -11010 16150
rect -11030 15970 -11010 15990
rect -10950 16450 -10930 16470
rect -10950 16290 -10930 16310
rect -10950 16130 -10930 16150
rect -10950 15970 -10930 15990
rect -10870 16450 -10850 16470
rect -10870 16290 -10850 16310
rect -10870 16130 -10850 16150
rect -10870 15970 -10850 15990
rect -10790 16450 -10770 16470
rect -10790 16290 -10770 16310
rect -10790 16130 -10770 16150
rect -10790 15970 -10770 15990
rect -10710 16450 -10690 16470
rect -10710 16290 -10690 16310
rect -10710 16130 -10690 16150
rect -10710 15970 -10690 15990
rect -10630 16450 -10610 16470
rect -10630 16290 -10610 16310
rect -10630 16130 -10610 16150
rect -10630 15970 -10610 15990
rect -10550 16450 -10530 16470
rect -10550 16290 -10530 16310
rect -10550 16130 -10530 16150
rect -10550 15970 -10530 15990
rect -10470 16450 -10450 16470
rect -10470 16290 -10450 16310
rect -10470 16130 -10450 16150
rect -10470 15970 -10450 15990
rect -10390 16450 -10370 16470
rect -10390 16290 -10370 16310
rect -10390 16130 -10370 16150
rect -10390 15970 -10370 15990
rect -10310 16450 -10290 16470
rect -10310 16290 -10290 16310
rect -10310 16130 -10290 16150
rect -10310 15970 -10290 15990
rect -10230 16450 -10210 16470
rect -10230 16290 -10210 16310
rect -10230 16130 -10210 16150
rect -10230 15970 -10210 15990
rect -10150 16450 -10130 16470
rect -10150 16290 -10130 16310
rect -10150 16130 -10130 16150
rect -10150 15970 -10130 15990
rect -10070 16450 -10050 16470
rect -10070 16290 -10050 16310
rect -10070 16130 -10050 16150
rect -10070 15970 -10050 15990
rect -9990 16450 -9970 16470
rect -9990 16290 -9970 16310
rect -9990 16130 -9970 16150
rect -9990 15970 -9970 15990
rect -9910 16450 -9890 16470
rect -9910 16290 -9890 16310
rect -9910 16130 -9890 16150
rect -9910 15970 -9890 15990
rect -9830 16450 -9810 16470
rect -9830 16290 -9810 16310
rect -9830 16130 -9810 16150
rect -9830 15970 -9810 15990
rect -9750 16450 -9730 16470
rect -9750 16290 -9730 16310
rect -9750 16130 -9730 16150
rect -9750 15970 -9730 15990
rect -9670 16450 -9650 16470
rect -9670 16290 -9650 16310
rect -9670 16130 -9650 16150
rect -9670 15970 -9650 15990
rect -9590 16450 -9570 16470
rect -9590 16290 -9570 16310
rect -9590 16130 -9570 16150
rect -9590 15970 -9570 15990
rect -9510 16450 -9490 16470
rect -9510 16290 -9490 16310
rect -9510 16130 -9490 16150
rect -9510 15970 -9490 15990
rect -9430 16450 -9410 16470
rect -9430 16290 -9410 16310
rect -9430 16130 -9410 16150
rect -9430 15970 -9410 15990
rect -9350 16450 -9330 16470
rect -9350 16290 -9330 16310
rect -9350 16130 -9330 16150
rect -9350 15970 -9330 15990
rect -9270 16450 -9250 16470
rect -9270 16290 -9250 16310
rect -9270 16130 -9250 16150
rect -9270 15970 -9250 15990
rect -9190 16450 -9170 16470
rect -9190 16290 -9170 16310
rect -9190 16130 -9170 16150
rect -9190 15970 -9170 15990
rect -9110 16450 -9090 16470
rect -9110 16290 -9090 16310
rect -9110 16130 -9090 16150
rect -9110 15970 -9090 15990
rect -9030 16450 -9010 16470
rect -9030 16290 -9010 16310
rect -9030 16130 -9010 16150
rect -9030 15970 -9010 15990
rect -8950 16450 -8930 16470
rect -8950 16290 -8930 16310
rect -8950 16130 -8930 16150
rect -8950 15970 -8930 15990
rect -8870 16450 -8850 16470
rect -8870 16290 -8850 16310
rect -8870 16130 -8850 16150
rect -8870 15970 -8850 15990
rect -8790 16450 -8770 16470
rect -8790 16290 -8770 16310
rect -8790 16130 -8770 16150
rect -8790 15970 -8770 15990
rect -8710 16450 -8690 16470
rect -8710 16290 -8690 16310
rect -8710 16130 -8690 16150
rect -8710 15970 -8690 15990
rect -8630 16450 -8610 16470
rect -8630 16290 -8610 16310
rect -8630 16130 -8610 16150
rect -8630 15970 -8610 15990
rect -8550 16450 -8530 16470
rect -8550 16290 -8530 16310
rect -8550 16130 -8530 16150
rect -8550 15970 -8530 15990
rect -8470 16450 -8450 16470
rect -8470 16290 -8450 16310
rect -8470 16130 -8450 16150
rect -8470 15970 -8450 15990
rect -8390 16450 -8370 16470
rect -8390 16290 -8370 16310
rect -8390 16130 -8370 16150
rect -8390 15970 -8370 15990
rect -8310 16450 -8290 16470
rect -8310 16290 -8290 16310
rect -8310 16130 -8290 16150
rect -8310 15970 -8290 15990
rect -8230 16450 -8210 16470
rect -8230 16290 -8210 16310
rect -8230 16130 -8210 16150
rect -8230 15970 -8210 15990
rect -8150 16450 -8130 16470
rect -8150 16290 -8130 16310
rect -8150 16130 -8130 16150
rect -8150 15970 -8130 15990
rect -8070 16450 -8050 16470
rect -8070 16290 -8050 16310
rect -8070 16130 -8050 16150
rect -8070 15970 -8050 15990
rect -7990 16450 -7970 16470
rect -7990 16290 -7970 16310
rect -7990 16130 -7970 16150
rect -7990 15970 -7970 15990
rect -7910 16450 -7890 16470
rect -7910 16290 -7890 16310
rect -7910 16130 -7890 16150
rect -7910 15970 -7890 15990
rect -7830 16450 -7810 16470
rect -7830 16290 -7810 16310
rect -7830 16130 -7810 16150
rect -7830 15970 -7810 15990
rect -7750 16450 -7730 16470
rect -7750 16290 -7730 16310
rect -7750 16130 -7730 16150
rect -7750 15970 -7730 15990
rect -7670 16450 -7650 16470
rect -7670 16290 -7650 16310
rect -7670 16130 -7650 16150
rect -7670 15970 -7650 15990
rect -7590 16450 -7570 16470
rect -7590 16290 -7570 16310
rect -7590 16130 -7570 16150
rect -7590 15970 -7570 15990
rect -7510 16450 -7490 16470
rect -7510 16290 -7490 16310
rect -7510 16130 -7490 16150
rect -7510 15970 -7490 15990
rect -7430 16450 -7410 16470
rect -7430 16290 -7410 16310
rect -7430 16130 -7410 16150
rect -7430 15970 -7410 15990
rect -7350 16450 -7330 16470
rect -7350 16290 -7330 16310
rect -7350 16130 -7330 16150
rect -7350 15970 -7330 15990
rect -7270 16450 -7250 16470
rect -7270 16290 -7250 16310
rect -7270 16130 -7250 16150
rect -7270 15970 -7250 15990
rect -7190 16450 -7170 16470
rect -7190 16290 -7170 16310
rect -7190 16130 -7170 16150
rect -7190 15970 -7170 15990
rect -7110 16450 -7090 16470
rect -7110 16290 -7090 16310
rect -7110 16130 -7090 16150
rect -7110 15970 -7090 15990
rect -7030 16450 -7010 16470
rect -7030 16290 -7010 16310
rect -7030 16130 -7010 16150
rect -7030 15970 -7010 15990
rect -6950 16450 -6930 16470
rect -6950 16290 -6930 16310
rect -6950 16130 -6930 16150
rect -6950 15970 -6930 15990
rect -6870 16450 -6850 16470
rect -6870 16290 -6850 16310
rect -6870 16130 -6850 16150
rect -6870 15970 -6850 15990
rect -6790 16450 -6770 16470
rect -6790 16290 -6770 16310
rect -6790 16130 -6770 16150
rect -6790 15970 -6770 15990
rect -6710 16450 -6690 16470
rect -6710 16290 -6690 16310
rect -6710 16130 -6690 16150
rect -6710 15970 -6690 15990
rect -6630 16450 -6610 16470
rect -6630 16290 -6610 16310
rect -6630 16130 -6610 16150
rect -6630 15970 -6610 15990
rect -6550 16450 -6530 16470
rect -6550 16290 -6530 16310
rect -6550 16130 -6530 16150
rect -6550 15970 -6530 15990
rect -6470 16450 -6450 16470
rect -6470 16290 -6450 16310
rect -6470 16130 -6450 16150
rect -6470 15970 -6450 15990
rect -6390 16450 -6370 16470
rect -6390 16290 -6370 16310
rect -6390 16130 -6370 16150
rect -6390 15970 -6370 15990
rect -6310 16450 -6290 16470
rect -6310 16290 -6290 16310
rect -6310 16130 -6290 16150
rect -6310 15970 -6290 15990
rect -6230 16450 -6210 16470
rect -6230 16290 -6210 16310
rect -6230 16130 -6210 16150
rect -6230 15970 -6210 15990
rect -6150 16450 -6130 16470
rect -6150 16290 -6130 16310
rect -6150 16130 -6130 16150
rect -6150 15970 -6130 15990
rect -6070 16450 -6050 16470
rect -6070 16290 -6050 16310
rect -6070 16130 -6050 16150
rect -6070 15970 -6050 15990
rect -5990 16450 -5970 16470
rect -5990 16290 -5970 16310
rect -5990 16130 -5970 16150
rect -5990 15970 -5970 15990
rect -5910 16450 -5890 16470
rect -5910 16290 -5890 16310
rect -5910 16130 -5890 16150
rect -5910 15970 -5890 15990
rect -5830 16450 -5810 16470
rect -5830 16290 -5810 16310
rect -5830 16130 -5810 16150
rect -5830 15970 -5810 15990
rect -5750 16450 -5730 16470
rect -5750 16290 -5730 16310
rect -5590 16450 -5570 16470
rect -5590 16290 -5570 16310
rect -5750 16130 -5730 16150
rect -5750 15970 -5730 15990
rect -5670 16130 -5650 16150
rect -5670 15970 -5650 15990
rect -5590 16130 -5570 16150
rect -5590 15970 -5570 15990
rect -5430 16450 -5410 16470
rect -5430 16290 -5410 16310
rect -5430 16130 -5410 16150
rect -5430 15970 -5410 15990
rect -5350 16450 -5330 16470
rect -5350 16290 -5330 16310
rect -5350 16130 -5330 16150
rect -5350 15970 -5330 15990
rect -5270 16450 -5250 16470
rect -5270 16290 -5250 16310
rect -5270 16130 -5250 16150
rect -5270 15970 -5250 15990
rect -5190 16450 -5170 16470
rect -5190 16290 -5170 16310
rect -5190 16130 -5170 16150
rect -5190 15970 -5170 15990
rect -5110 16450 -5090 16470
rect -5110 16290 -5090 16310
rect -5110 16130 -5090 16150
rect -5110 15970 -5090 15990
rect -5030 16450 -5010 16470
rect -5030 16290 -5010 16310
rect -5030 16130 -5010 16150
rect -5030 15970 -5010 15990
rect -4950 16450 -4930 16470
rect -4950 16290 -4930 16310
rect -4950 16130 -4930 16150
rect -4950 15970 -4930 15990
rect -4870 16450 -4850 16470
rect -4870 16290 -4850 16310
rect -4870 16130 -4850 16150
rect -4870 15970 -4850 15990
rect -4790 16450 -4770 16470
rect -4790 16290 -4770 16310
rect -4790 16130 -4770 16150
rect -4790 15970 -4770 15990
rect -4710 16450 -4690 16470
rect -4710 16290 -4690 16310
rect -4710 16130 -4690 16150
rect -4710 15970 -4690 15990
rect -4630 16450 -4610 16470
rect -4630 16290 -4610 16310
rect -4630 16130 -4610 16150
rect -4630 15970 -4610 15990
rect -4550 16450 -4530 16470
rect -4550 16290 -4530 16310
rect -4550 16130 -4530 16150
rect -4550 15970 -4530 15990
rect -4470 16450 -4450 16470
rect -4470 16290 -4450 16310
rect -4470 16130 -4450 16150
rect -4470 15970 -4450 15990
rect -4390 16450 -4370 16470
rect -4390 16290 -4370 16310
rect -4390 16130 -4370 16150
rect -4390 15970 -4370 15990
rect -4310 16450 -4290 16470
rect -4310 16290 -4290 16310
rect -4310 16130 -4290 16150
rect -4310 15970 -4290 15990
rect -4230 16450 -4210 16470
rect -4230 16290 -4210 16310
rect -4230 16130 -4210 16150
rect -4230 15970 -4210 15990
rect -4150 16450 -4130 16470
rect -4150 16290 -4130 16310
rect -4150 16130 -4130 16150
rect -4150 15970 -4130 15990
rect -4070 16450 -4050 16470
rect -4070 16290 -4050 16310
rect -4070 16130 -4050 16150
rect -4070 15970 -4050 15990
rect -3990 16450 -3970 16470
rect -3990 16290 -3970 16310
rect -3990 16130 -3970 16150
rect -3990 15970 -3970 15990
rect -3910 16450 -3890 16470
rect -3910 16290 -3890 16310
rect -3910 16130 -3890 16150
rect -3910 15970 -3890 15990
rect -3830 16450 -3810 16470
rect -3830 16290 -3810 16310
rect -3830 16130 -3810 16150
rect -3830 15970 -3810 15990
rect -3750 16450 -3730 16470
rect -3750 16290 -3730 16310
rect -3750 16130 -3730 16150
rect -3750 15970 -3730 15990
rect -3670 16450 -3650 16470
rect -3670 16290 -3650 16310
rect -3670 16130 -3650 16150
rect -3670 15970 -3650 15990
rect -3590 16450 -3570 16470
rect -3590 16290 -3570 16310
rect -3590 16130 -3570 16150
rect -3590 15970 -3570 15990
rect -3510 16450 -3490 16470
rect -3510 16290 -3490 16310
rect -3510 16130 -3490 16150
rect -3510 15970 -3490 15990
rect -3430 16450 -3410 16470
rect -3430 16290 -3410 16310
rect -3430 16130 -3410 16150
rect -3430 15970 -3410 15990
rect -3350 16450 -3330 16470
rect -3350 16290 -3330 16310
rect -3350 16130 -3330 16150
rect -3350 15970 -3330 15990
rect -3270 16450 -3250 16470
rect -3270 16290 -3250 16310
rect -3270 16130 -3250 16150
rect -3270 15970 -3250 15990
rect -3190 16450 -3170 16470
rect -3190 16290 -3170 16310
rect -3190 16130 -3170 16150
rect -3190 15970 -3170 15990
rect -3110 16450 -3090 16470
rect -3110 16290 -3090 16310
rect -3110 16130 -3090 16150
rect -3110 15970 -3090 15990
rect -3030 16450 -3010 16470
rect -3030 16290 -3010 16310
rect -3030 16130 -3010 16150
rect -3030 15970 -3010 15990
rect -2950 16450 -2930 16470
rect -2950 16290 -2930 16310
rect -2950 16130 -2930 16150
rect -2950 15970 -2930 15990
rect -2870 16450 -2850 16470
rect -2870 16290 -2850 16310
rect -2870 16130 -2850 16150
rect -2870 15970 -2850 15990
rect -2790 16450 -2770 16470
rect -2790 16290 -2770 16310
rect -2790 16130 -2770 16150
rect -2790 15970 -2770 15990
rect -2710 16450 -2690 16470
rect -2710 16290 -2690 16310
rect -2710 16130 -2690 16150
rect -2710 15970 -2690 15990
rect -2630 16450 -2610 16470
rect -2630 16290 -2610 16310
rect -2630 16130 -2610 16150
rect -2630 15970 -2610 15990
rect -2550 16450 -2530 16470
rect -2550 16290 -2530 16310
rect -2550 16130 -2530 16150
rect -2550 15970 -2530 15990
rect -2470 16450 -2450 16470
rect -2470 16290 -2450 16310
rect -2470 16130 -2450 16150
rect -2470 15970 -2450 15990
rect -2390 16450 -2370 16470
rect -2390 16290 -2370 16310
rect -2390 16130 -2370 16150
rect -2390 15970 -2370 15990
rect -2310 16450 -2290 16470
rect -2310 16290 -2290 16310
rect -2310 16130 -2290 16150
rect -2310 15970 -2290 15990
rect -2230 16450 -2210 16470
rect -2230 16290 -2210 16310
rect -2230 16130 -2210 16150
rect -2230 15970 -2210 15990
rect -2150 16450 -2130 16470
rect -2150 16290 -2130 16310
rect -2150 16130 -2130 16150
rect -2150 15970 -2130 15990
rect -2070 16450 -2050 16470
rect -2070 16290 -2050 16310
rect -2070 16130 -2050 16150
rect -2070 15970 -2050 15990
rect -1990 16450 -1970 16470
rect -1990 16290 -1970 16310
rect -1990 16130 -1970 16150
rect -1990 15970 -1970 15990
rect -1830 16450 -1810 16470
rect -1830 16290 -1810 16310
rect -1830 16130 -1810 16150
rect -1830 15970 -1810 15990
rect -1750 16450 -1730 16470
rect -1750 16290 -1730 16310
rect -1750 16130 -1730 16150
rect -1750 15970 -1730 15990
rect -1670 16450 -1650 16470
rect -1670 16290 -1650 16310
rect -1670 16130 -1650 16150
rect -1670 15970 -1650 15990
rect -1590 16450 -1570 16470
rect -1590 16290 -1570 16310
rect -1590 16130 -1570 16150
rect -1590 15970 -1570 15990
rect -1510 16450 -1490 16470
rect -1510 16290 -1490 16310
rect -1510 16130 -1490 16150
rect -1510 15970 -1490 15990
rect -1430 16450 -1410 16470
rect -1430 16290 -1410 16310
rect -1430 16130 -1410 16150
rect -1430 15970 -1410 15990
rect -1350 16450 -1330 16470
rect -1350 16290 -1330 16310
rect -1350 16130 -1330 16150
rect -1350 15970 -1330 15990
rect -1190 16450 -1170 16470
rect -1190 16290 -1170 16310
rect -1190 16130 -1170 16150
rect -1190 15970 -1170 15990
rect -1030 16450 -1010 16470
rect -1030 16290 -1010 16310
rect -1030 16130 -1010 16150
rect -1030 15970 -1010 15990
rect -870 16450 -850 16470
rect -870 16290 -850 16310
rect -870 16130 -850 16150
rect -870 15970 -850 15990
rect -710 16450 -690 16470
rect -710 16290 -690 16310
rect -710 16130 -690 16150
rect -710 15970 -690 15990
rect -550 16450 -530 16470
rect -550 16290 -530 16310
rect -550 16130 -530 16150
rect -550 15970 -530 15990
<< metal1 >>
rect -14960 21435 -14920 21440
rect -14960 21405 -14955 21435
rect -14925 21405 -14920 21435
rect -14960 21400 -14920 21405
rect -14880 21435 -14840 21440
rect -14880 21405 -14875 21435
rect -14845 21405 -14840 21435
rect -14880 21400 -14840 21405
rect -14800 21435 -14760 21440
rect -14800 21405 -14795 21435
rect -14765 21405 -14760 21435
rect -14800 21400 -14760 21405
rect -14720 21435 -14680 21440
rect -14720 21405 -14715 21435
rect -14685 21405 -14680 21435
rect -14720 21400 -14680 21405
rect -14640 21435 -14600 21440
rect -14640 21405 -14635 21435
rect -14605 21405 -14600 21435
rect -14640 21400 -14600 21405
rect -14560 21435 -14520 21440
rect -14560 21405 -14555 21435
rect -14525 21405 -14520 21435
rect -14560 21400 -14520 21405
rect -14480 21435 -14440 21440
rect -14480 21405 -14475 21435
rect -14445 21405 -14440 21435
rect -14480 21400 -14440 21405
rect -14400 21435 -14360 21440
rect -14400 21405 -14395 21435
rect -14365 21405 -14360 21435
rect -14400 21400 -14360 21405
rect -14320 21435 -14280 21440
rect -14320 21405 -14315 21435
rect -14285 21405 -14280 21435
rect -14320 21400 -14280 21405
rect -14240 21435 -14200 21440
rect -14240 21405 -14235 21435
rect -14205 21405 -14200 21435
rect -14240 21400 -14200 21405
rect -14160 21435 -14120 21440
rect -14160 21405 -14155 21435
rect -14125 21405 -14120 21435
rect -14160 21400 -14120 21405
rect -14080 21435 -14040 21440
rect -14080 21405 -14075 21435
rect -14045 21405 -14040 21435
rect -14080 21400 -14040 21405
rect -14000 21435 -13960 21440
rect -14000 21405 -13995 21435
rect -13965 21405 -13960 21435
rect -14000 21400 -13960 21405
rect -13920 21435 -13880 21440
rect -13920 21405 -13915 21435
rect -13885 21405 -13880 21435
rect -13920 21400 -13880 21405
rect -13840 21435 -13800 21440
rect -13840 21405 -13835 21435
rect -13805 21405 -13800 21435
rect -13840 21400 -13800 21405
rect -13760 21435 -13720 21440
rect -13760 21405 -13755 21435
rect -13725 21405 -13720 21435
rect -13760 21400 -13720 21405
rect -13680 21435 -13640 21440
rect -13680 21405 -13675 21435
rect -13645 21405 -13640 21435
rect -13680 21400 -13640 21405
rect -13600 21435 -13560 21440
rect -13600 21405 -13595 21435
rect -13565 21405 -13560 21435
rect -13600 21400 -13560 21405
rect -13520 21435 -13480 21440
rect -13520 21405 -13515 21435
rect -13485 21405 -13480 21435
rect -13520 21400 -13480 21405
rect -13440 21435 -13400 21440
rect -13440 21405 -13435 21435
rect -13405 21405 -13400 21435
rect -13440 21400 -13400 21405
rect -13360 21435 -13320 21440
rect -13360 21405 -13355 21435
rect -13325 21405 -13320 21435
rect -13360 21400 -13320 21405
rect -13280 21435 -13240 21440
rect -13280 21405 -13275 21435
rect -13245 21405 -13240 21435
rect -13280 21400 -13240 21405
rect -13200 21435 -13160 21440
rect -13200 21405 -13195 21435
rect -13165 21405 -13160 21435
rect -13200 21400 -13160 21405
rect -13120 21435 -13080 21440
rect -13120 21405 -13115 21435
rect -13085 21405 -13080 21435
rect -13120 21400 -13080 21405
rect -13040 21435 -13000 21440
rect -13040 21405 -13035 21435
rect -13005 21405 -13000 21435
rect -13040 21400 -13000 21405
rect -12960 21435 -12920 21440
rect -12960 21405 -12955 21435
rect -12925 21405 -12920 21435
rect -12960 21400 -12920 21405
rect -12880 21435 -12840 21440
rect -12880 21405 -12875 21435
rect -12845 21405 -12840 21435
rect -12880 21400 -12840 21405
rect -12800 21435 -12760 21440
rect -12800 21405 -12795 21435
rect -12765 21405 -12760 21435
rect -12800 21400 -12760 21405
rect -12720 21435 -12680 21440
rect -12720 21405 -12715 21435
rect -12685 21405 -12680 21435
rect -12720 21400 -12680 21405
rect -12640 21435 -12600 21440
rect -12640 21405 -12635 21435
rect -12605 21405 -12600 21435
rect -12640 21400 -12600 21405
rect -12560 21435 -12520 21440
rect -12560 21405 -12555 21435
rect -12525 21405 -12520 21435
rect -12560 21400 -12520 21405
rect -12480 21435 -12440 21440
rect -12480 21405 -12475 21435
rect -12445 21405 -12440 21435
rect -12480 21400 -12440 21405
rect -12400 21435 -12360 21440
rect -12400 21405 -12395 21435
rect -12365 21405 -12360 21435
rect -12400 21400 -12360 21405
rect -12320 21435 -12280 21440
rect -12320 21405 -12315 21435
rect -12285 21405 -12280 21435
rect -12320 21400 -12280 21405
rect -12240 21435 -12200 21440
rect -12240 21405 -12235 21435
rect -12205 21405 -12200 21435
rect -12240 21400 -12200 21405
rect -12160 21435 -12120 21440
rect -12160 21405 -12155 21435
rect -12125 21405 -12120 21435
rect -12160 21400 -12120 21405
rect -12080 21435 -12040 21440
rect -12080 21405 -12075 21435
rect -12045 21405 -12040 21435
rect -12080 21400 -12040 21405
rect -12000 21435 -11960 21440
rect -12000 21405 -11995 21435
rect -11965 21405 -11960 21435
rect -12000 21400 -11960 21405
rect -11920 21435 -11880 21440
rect -11920 21405 -11915 21435
rect -11885 21405 -11880 21435
rect -11920 21400 -11880 21405
rect -11840 21435 -11800 21440
rect -11840 21405 -11835 21435
rect -11805 21405 -11800 21435
rect -11840 21400 -11800 21405
rect -11760 21435 -11720 21440
rect -11760 21405 -11755 21435
rect -11725 21405 -11720 21435
rect -11760 21400 -11720 21405
rect -11680 21435 -11640 21440
rect -11680 21405 -11675 21435
rect -11645 21405 -11640 21435
rect -11680 21400 -11640 21405
rect -11600 21435 -11560 21440
rect -11600 21405 -11595 21435
rect -11565 21405 -11560 21435
rect -11600 21400 -11560 21405
rect -11520 21435 -11480 21440
rect -11520 21405 -11515 21435
rect -11485 21405 -11480 21435
rect -11520 21400 -11480 21405
rect -11440 21435 -11400 21440
rect -11440 21405 -11435 21435
rect -11405 21405 -11400 21435
rect -11440 21400 -11400 21405
rect -11360 21435 -11320 21440
rect -11360 21405 -11355 21435
rect -11325 21405 -11320 21435
rect -11360 21400 -11320 21405
rect -11280 21435 -11240 21440
rect -11280 21405 -11275 21435
rect -11245 21405 -11240 21435
rect -11280 21400 -11240 21405
rect -11200 21435 -11160 21440
rect -11200 21405 -11195 21435
rect -11165 21405 -11160 21435
rect -11200 21400 -11160 21405
rect -11120 21435 -11080 21440
rect -11120 21405 -11115 21435
rect -11085 21405 -11080 21435
rect -11120 21400 -11080 21405
rect -11040 21435 -11000 21440
rect -11040 21405 -11035 21435
rect -11005 21405 -11000 21435
rect -11040 21400 -11000 21405
rect -10960 21435 -10920 21440
rect -10960 21405 -10955 21435
rect -10925 21405 -10920 21435
rect -10960 21400 -10920 21405
rect -10880 21435 -10840 21440
rect -10880 21405 -10875 21435
rect -10845 21405 -10840 21435
rect -10880 21400 -10840 21405
rect -10800 21435 -10760 21440
rect -10800 21405 -10795 21435
rect -10765 21405 -10760 21435
rect -10800 21400 -10760 21405
rect -10720 21435 -10680 21440
rect -10720 21405 -10715 21435
rect -10685 21405 -10680 21435
rect -10720 21400 -10680 21405
rect -10640 21435 -10600 21440
rect -10640 21405 -10635 21435
rect -10605 21405 -10600 21435
rect -10640 21400 -10600 21405
rect -10560 21435 -10520 21440
rect -10560 21405 -10555 21435
rect -10525 21405 -10520 21435
rect -10560 21400 -10520 21405
rect -10480 21435 -10440 21440
rect -10480 21405 -10475 21435
rect -10445 21405 -10440 21435
rect -10480 21400 -10440 21405
rect -10400 21435 -10360 21440
rect -10400 21405 -10395 21435
rect -10365 21405 -10360 21435
rect -10400 21400 -10360 21405
rect -10320 21435 -10280 21440
rect -10320 21405 -10315 21435
rect -10285 21405 -10280 21435
rect -10320 21400 -10280 21405
rect -10240 21435 -10200 21440
rect -10240 21405 -10235 21435
rect -10205 21405 -10200 21435
rect -10240 21400 -10200 21405
rect -10160 21435 -10120 21440
rect -10160 21405 -10155 21435
rect -10125 21405 -10120 21435
rect -10160 21400 -10120 21405
rect -10080 21435 -10040 21440
rect -10080 21405 -10075 21435
rect -10045 21405 -10040 21435
rect -10080 21400 -10040 21405
rect -10000 21435 -9960 21440
rect -10000 21405 -9995 21435
rect -9965 21405 -9960 21435
rect -10000 21400 -9960 21405
rect -9920 21435 -9880 21440
rect -9920 21405 -9915 21435
rect -9885 21405 -9880 21435
rect -9920 21400 -9880 21405
rect -9840 21435 -9800 21440
rect -9840 21405 -9835 21435
rect -9805 21405 -9800 21435
rect -9840 21400 -9800 21405
rect -9760 21435 -9720 21440
rect -9760 21405 -9755 21435
rect -9725 21405 -9720 21435
rect -9760 21400 -9720 21405
rect -9680 21435 -9640 21440
rect -9680 21405 -9675 21435
rect -9645 21405 -9640 21435
rect -9680 21400 -9640 21405
rect -9600 21435 -9560 21440
rect -9600 21405 -9595 21435
rect -9565 21405 -9560 21435
rect -9600 21400 -9560 21405
rect -9520 21435 -9480 21440
rect -9520 21405 -9515 21435
rect -9485 21405 -9480 21435
rect -9520 21400 -9480 21405
rect -9440 21435 -9400 21440
rect -9440 21405 -9435 21435
rect -9405 21405 -9400 21435
rect -9440 21400 -9400 21405
rect -9360 21435 -9320 21440
rect -9360 21405 -9355 21435
rect -9325 21405 -9320 21435
rect -9360 21400 -9320 21405
rect -9280 21435 -9240 21440
rect -9280 21405 -9275 21435
rect -9245 21405 -9240 21435
rect -9280 21400 -9240 21405
rect -9200 21435 -9160 21440
rect -9200 21405 -9195 21435
rect -9165 21405 -9160 21435
rect -9200 21400 -9160 21405
rect -9120 21435 -9080 21440
rect -9120 21405 -9115 21435
rect -9085 21405 -9080 21435
rect -9120 21400 -9080 21405
rect -9040 21435 -9000 21440
rect -9040 21405 -9035 21435
rect -9005 21405 -9000 21435
rect -9040 21400 -9000 21405
rect -8960 21435 -8920 21440
rect -8960 21405 -8955 21435
rect -8925 21405 -8920 21435
rect -8960 21400 -8920 21405
rect -8880 21435 -8840 21440
rect -8880 21405 -8875 21435
rect -8845 21405 -8840 21435
rect -8880 21400 -8840 21405
rect -8800 21435 -8760 21440
rect -8800 21405 -8795 21435
rect -8765 21405 -8760 21435
rect -8800 21400 -8760 21405
rect -8720 21435 -8680 21440
rect -8720 21405 -8715 21435
rect -8685 21405 -8680 21435
rect -8720 21400 -8680 21405
rect -8640 21435 -8600 21440
rect -8640 21405 -8635 21435
rect -8605 21405 -8600 21435
rect -8640 21400 -8600 21405
rect -8560 21435 -8520 21440
rect -8560 21405 -8555 21435
rect -8525 21405 -8520 21435
rect -8560 21400 -8520 21405
rect -8480 21435 -8440 21440
rect -8480 21405 -8475 21435
rect -8445 21405 -8440 21435
rect -8480 21400 -8440 21405
rect -8400 21435 -8360 21440
rect -8400 21405 -8395 21435
rect -8365 21405 -8360 21435
rect -8400 21400 -8360 21405
rect -8320 21435 -8280 21440
rect -8320 21405 -8315 21435
rect -8285 21405 -8280 21435
rect -8320 21400 -8280 21405
rect -8240 21435 -8200 21440
rect -8240 21405 -8235 21435
rect -8205 21405 -8200 21435
rect -8240 21400 -8200 21405
rect -8160 21435 -8120 21440
rect -8160 21405 -8155 21435
rect -8125 21405 -8120 21435
rect -8160 21400 -8120 21405
rect -8080 21435 -8040 21440
rect -8080 21405 -8075 21435
rect -8045 21405 -8040 21435
rect -8080 21400 -8040 21405
rect -8000 21435 -7960 21440
rect -8000 21405 -7995 21435
rect -7965 21405 -7960 21435
rect -8000 21400 -7960 21405
rect -7920 21435 -7880 21440
rect -7920 21405 -7915 21435
rect -7885 21405 -7880 21435
rect -7920 21400 -7880 21405
rect -7840 21435 -7800 21440
rect -7840 21405 -7835 21435
rect -7805 21405 -7800 21435
rect -7840 21400 -7800 21405
rect -7760 21435 -7720 21440
rect -7760 21405 -7755 21435
rect -7725 21405 -7720 21435
rect -7760 21400 -7720 21405
rect -7680 21435 -7640 21440
rect -7680 21405 -7675 21435
rect -7645 21405 -7640 21435
rect -7680 21400 -7640 21405
rect -7600 21435 -7560 21440
rect -7600 21405 -7595 21435
rect -7565 21405 -7560 21435
rect -7600 21400 -7560 21405
rect -7520 21435 -7480 21440
rect -7520 21405 -7515 21435
rect -7485 21405 -7480 21435
rect -7520 21400 -7480 21405
rect -7440 21435 -7400 21440
rect -7440 21405 -7435 21435
rect -7405 21405 -7400 21435
rect -7440 21400 -7400 21405
rect -7360 21435 -7320 21440
rect -7360 21405 -7355 21435
rect -7325 21405 -7320 21435
rect -7360 21400 -7320 21405
rect -7280 21435 -7240 21440
rect -7280 21405 -7275 21435
rect -7245 21405 -7240 21435
rect -7280 21400 -7240 21405
rect -7200 21435 -7160 21440
rect -7200 21405 -7195 21435
rect -7165 21405 -7160 21435
rect -7200 21400 -7160 21405
rect -7120 21435 -7080 21440
rect -7120 21405 -7115 21435
rect -7085 21405 -7080 21435
rect -7120 21400 -7080 21405
rect -7040 21435 -7000 21440
rect -7040 21405 -7035 21435
rect -7005 21405 -7000 21435
rect -7040 21400 -7000 21405
rect -6960 21435 -6920 21440
rect -6960 21405 -6955 21435
rect -6925 21405 -6920 21435
rect -6960 21400 -6920 21405
rect -6880 21435 -6840 21440
rect -6880 21405 -6875 21435
rect -6845 21405 -6840 21435
rect -6880 21400 -6840 21405
rect -6800 21435 -6760 21440
rect -6800 21405 -6795 21435
rect -6765 21405 -6760 21435
rect -6800 21400 -6760 21405
rect -6720 21435 -6680 21440
rect -6720 21405 -6715 21435
rect -6685 21405 -6680 21435
rect -6720 21400 -6680 21405
rect -6640 21435 -6600 21440
rect -6640 21405 -6635 21435
rect -6605 21405 -6600 21435
rect -6640 21400 -6600 21405
rect -6560 21435 -6520 21440
rect -6560 21405 -6555 21435
rect -6525 21405 -6520 21435
rect -6560 21400 -6520 21405
rect -6480 21435 -6440 21440
rect -6480 21405 -6475 21435
rect -6445 21405 -6440 21435
rect -6480 21400 -6440 21405
rect -6400 21435 -6360 21440
rect -6400 21405 -6395 21435
rect -6365 21405 -6360 21435
rect -6400 21400 -6360 21405
rect -6320 21435 -6280 21440
rect -6320 21405 -6315 21435
rect -6285 21405 -6280 21435
rect -6320 21400 -6280 21405
rect -6240 21435 -6200 21440
rect -6240 21405 -6235 21435
rect -6205 21405 -6200 21435
rect -6240 21400 -6200 21405
rect -6160 21435 -6120 21440
rect -6160 21405 -6155 21435
rect -6125 21405 -6120 21435
rect -6160 21400 -6120 21405
rect -5680 21435 -5640 21440
rect -5680 21405 -5675 21435
rect -5645 21405 -5640 21435
rect -5680 21400 -5640 21405
rect -5600 21435 -5560 21440
rect -5600 21405 -5595 21435
rect -5565 21405 -5560 21435
rect -5600 21400 -5560 21405
rect -5520 21435 -5480 21440
rect -5520 21405 -5515 21435
rect -5485 21405 -5480 21435
rect -5520 21400 -5480 21405
rect -5440 21435 -5400 21440
rect -5440 21405 -5435 21435
rect -5405 21405 -5400 21435
rect -5440 21400 -5400 21405
rect -5360 21435 -5320 21440
rect -5360 21405 -5355 21435
rect -5325 21405 -5320 21435
rect -5360 21400 -5320 21405
rect -5280 21435 -5240 21440
rect -5280 21405 -5275 21435
rect -5245 21405 -5240 21435
rect -5280 21400 -5240 21405
rect -5200 21435 -5160 21440
rect -5200 21405 -5195 21435
rect -5165 21405 -5160 21435
rect -5200 21400 -5160 21405
rect -5120 21435 -5080 21440
rect -5120 21405 -5115 21435
rect -5085 21405 -5080 21435
rect -5120 21400 -5080 21405
rect -5040 21435 -5000 21440
rect -5040 21405 -5035 21435
rect -5005 21405 -5000 21435
rect -5040 21400 -5000 21405
rect -4960 21435 -4920 21440
rect -4960 21405 -4955 21435
rect -4925 21405 -4920 21435
rect -4960 21400 -4920 21405
rect -4880 21435 -4840 21440
rect -4880 21405 -4875 21435
rect -4845 21405 -4840 21435
rect -4880 21400 -4840 21405
rect -4800 21435 -4760 21440
rect -4800 21405 -4795 21435
rect -4765 21405 -4760 21435
rect -4800 21400 -4760 21405
rect -4720 21435 -4680 21440
rect -4720 21405 -4715 21435
rect -4685 21405 -4680 21435
rect -4720 21400 -4680 21405
rect -4640 21435 -4600 21440
rect -4640 21405 -4635 21435
rect -4605 21405 -4600 21435
rect -4640 21400 -4600 21405
rect -4560 21435 -4520 21440
rect -4560 21405 -4555 21435
rect -4525 21405 -4520 21435
rect -4560 21400 -4520 21405
rect -4480 21435 -4440 21440
rect -4480 21405 -4475 21435
rect -4445 21405 -4440 21435
rect -4480 21400 -4440 21405
rect -4400 21435 -4360 21440
rect -4400 21405 -4395 21435
rect -4365 21405 -4360 21435
rect -4400 21400 -4360 21405
rect -4320 21435 -4280 21440
rect -4320 21405 -4315 21435
rect -4285 21405 -4280 21435
rect -4320 21400 -4280 21405
rect -4240 21435 -4200 21440
rect -4240 21405 -4235 21435
rect -4205 21405 -4200 21435
rect -4240 21400 -4200 21405
rect -4160 21435 -4120 21440
rect -4160 21405 -4155 21435
rect -4125 21405 -4120 21435
rect -4160 21400 -4120 21405
rect -4080 21435 -4040 21440
rect -4080 21405 -4075 21435
rect -4045 21405 -4040 21435
rect -4080 21400 -4040 21405
rect -4000 21435 -3960 21440
rect -4000 21405 -3995 21435
rect -3965 21405 -3960 21435
rect -4000 21400 -3960 21405
rect -3920 21435 -3880 21440
rect -3920 21405 -3915 21435
rect -3885 21405 -3880 21435
rect -3920 21400 -3880 21405
rect -3840 21435 -3800 21440
rect -3840 21405 -3835 21435
rect -3805 21405 -3800 21435
rect -3840 21400 -3800 21405
rect -3760 21435 -3720 21440
rect -3760 21405 -3755 21435
rect -3725 21405 -3720 21435
rect -3760 21400 -3720 21405
rect -3680 21435 -3640 21440
rect -3680 21405 -3675 21435
rect -3645 21405 -3640 21435
rect -3680 21400 -3640 21405
rect -3600 21435 -3560 21440
rect -3600 21405 -3595 21435
rect -3565 21405 -3560 21435
rect -3600 21400 -3560 21405
rect -3520 21435 -3480 21440
rect -3520 21405 -3515 21435
rect -3485 21405 -3480 21435
rect -3520 21400 -3480 21405
rect -3440 21435 -3400 21440
rect -3440 21405 -3435 21435
rect -3405 21405 -3400 21435
rect -3440 21400 -3400 21405
rect -3360 21435 -3320 21440
rect -3360 21405 -3355 21435
rect -3325 21405 -3320 21435
rect -3360 21400 -3320 21405
rect -3280 21435 -3240 21440
rect -3280 21405 -3275 21435
rect -3245 21405 -3240 21435
rect -3280 21400 -3240 21405
rect -3200 21435 -3160 21440
rect -3200 21405 -3195 21435
rect -3165 21405 -3160 21435
rect -3200 21400 -3160 21405
rect -3120 21435 -3080 21440
rect -3120 21405 -3115 21435
rect -3085 21405 -3080 21435
rect -3120 21400 -3080 21405
rect -3040 21435 -3000 21440
rect -3040 21405 -3035 21435
rect -3005 21405 -3000 21435
rect -3040 21400 -3000 21405
rect -2960 21435 -2920 21440
rect -2960 21405 -2955 21435
rect -2925 21405 -2920 21435
rect -2960 21400 -2920 21405
rect -2880 21435 -2840 21440
rect -2880 21405 -2875 21435
rect -2845 21405 -2840 21435
rect -2880 21400 -2840 21405
rect -2800 21435 -2760 21440
rect -2800 21405 -2795 21435
rect -2765 21405 -2760 21435
rect -2800 21400 -2760 21405
rect -2720 21435 -2680 21440
rect -2720 21405 -2715 21435
rect -2685 21405 -2680 21435
rect -2720 21400 -2680 21405
rect -2640 21435 -2600 21440
rect -2640 21405 -2635 21435
rect -2605 21405 -2600 21435
rect -2640 21400 -2600 21405
rect -2560 21435 -2520 21440
rect -2560 21405 -2555 21435
rect -2525 21405 -2520 21435
rect -2560 21400 -2520 21405
rect -2480 21435 -2440 21440
rect -2480 21405 -2475 21435
rect -2445 21405 -2440 21435
rect -2480 21400 -2440 21405
rect -2400 21435 -2360 21440
rect -2400 21405 -2395 21435
rect -2365 21405 -2360 21435
rect -2400 21400 -2360 21405
rect -2320 21435 -2280 21440
rect -2320 21405 -2315 21435
rect -2285 21405 -2280 21435
rect -2320 21400 -2280 21405
rect -2240 21435 -2200 21440
rect -2240 21405 -2235 21435
rect -2205 21405 -2200 21435
rect -2240 21400 -2200 21405
rect -2160 21435 -2120 21440
rect -2160 21405 -2155 21435
rect -2125 21405 -2120 21435
rect -2160 21400 -2120 21405
rect -2080 21435 -2040 21440
rect -2080 21405 -2075 21435
rect -2045 21405 -2040 21435
rect -2080 21400 -2040 21405
rect -2000 21435 -1960 21440
rect -2000 21405 -1995 21435
rect -1965 21405 -1960 21435
rect -2000 21400 -1960 21405
rect -1840 21435 -1800 21440
rect -1840 21405 -1835 21435
rect -1805 21405 -1800 21435
rect -1840 21400 -1800 21405
rect -1760 21435 -1720 21440
rect -1760 21405 -1755 21435
rect -1725 21405 -1720 21435
rect -1760 21400 -1720 21405
rect -1680 21435 -1640 21440
rect -1680 21405 -1675 21435
rect -1645 21405 -1640 21435
rect -1680 21400 -1640 21405
rect -1520 21435 -1480 21440
rect -1520 21405 -1515 21435
rect -1485 21405 -1480 21435
rect -1520 21400 -1480 21405
rect -1360 21435 -1320 21440
rect -1360 21405 -1355 21435
rect -1325 21405 -1320 21435
rect -1360 21400 -1320 21405
rect -1280 21435 -1240 21440
rect -1280 21405 -1275 21435
rect -1245 21405 -1240 21435
rect -1280 21400 -1240 21405
rect -1200 21435 -1160 21440
rect -1200 21405 -1195 21435
rect -1165 21405 -1160 21435
rect -1200 21400 -1160 21405
rect -1120 21435 -1080 21440
rect -1120 21405 -1115 21435
rect -1085 21405 -1080 21435
rect -1120 21400 -1080 21405
rect -1040 21435 -1000 21440
rect -1040 21405 -1035 21435
rect -1005 21405 -1000 21435
rect -1040 21400 -1000 21405
rect -880 21435 -840 21440
rect -880 21405 -875 21435
rect -845 21405 -840 21435
rect -880 21400 -840 21405
rect -720 21435 -680 21440
rect -720 21405 -715 21435
rect -685 21405 -680 21435
rect -720 21400 -680 21405
rect -560 21435 -520 21440
rect -560 21405 -555 21435
rect -525 21405 -520 21435
rect -560 21400 -520 21405
rect -14960 21275 -14920 21280
rect -14960 21245 -14955 21275
rect -14925 21245 -14920 21275
rect -14960 21240 -14920 21245
rect -14880 21275 -14840 21280
rect -14880 21245 -14875 21275
rect -14845 21245 -14840 21275
rect -14880 21240 -14840 21245
rect -14800 21275 -14760 21280
rect -14800 21245 -14795 21275
rect -14765 21245 -14760 21275
rect -14800 21240 -14760 21245
rect -14720 21275 -14680 21280
rect -14720 21245 -14715 21275
rect -14685 21245 -14680 21275
rect -14720 21240 -14680 21245
rect -14640 21275 -14600 21280
rect -14640 21245 -14635 21275
rect -14605 21245 -14600 21275
rect -14640 21240 -14600 21245
rect -14560 21275 -14520 21280
rect -14560 21245 -14555 21275
rect -14525 21245 -14520 21275
rect -14560 21240 -14520 21245
rect -14480 21275 -14440 21280
rect -14480 21245 -14475 21275
rect -14445 21245 -14440 21275
rect -14480 21240 -14440 21245
rect -14400 21275 -14360 21280
rect -14400 21245 -14395 21275
rect -14365 21245 -14360 21275
rect -14400 21240 -14360 21245
rect -14320 21275 -14280 21280
rect -14320 21245 -14315 21275
rect -14285 21245 -14280 21275
rect -14320 21240 -14280 21245
rect -14240 21275 -14200 21280
rect -14240 21245 -14235 21275
rect -14205 21245 -14200 21275
rect -14240 21240 -14200 21245
rect -14160 21275 -14120 21280
rect -14160 21245 -14155 21275
rect -14125 21245 -14120 21275
rect -14160 21240 -14120 21245
rect -14080 21275 -14040 21280
rect -14080 21245 -14075 21275
rect -14045 21245 -14040 21275
rect -14080 21240 -14040 21245
rect -14000 21275 -13960 21280
rect -14000 21245 -13995 21275
rect -13965 21245 -13960 21275
rect -14000 21240 -13960 21245
rect -13920 21275 -13880 21280
rect -13920 21245 -13915 21275
rect -13885 21245 -13880 21275
rect -13920 21240 -13880 21245
rect -13840 21275 -13800 21280
rect -13840 21245 -13835 21275
rect -13805 21245 -13800 21275
rect -13840 21240 -13800 21245
rect -13760 21275 -13720 21280
rect -13760 21245 -13755 21275
rect -13725 21245 -13720 21275
rect -13760 21240 -13720 21245
rect -13680 21275 -13640 21280
rect -13680 21245 -13675 21275
rect -13645 21245 -13640 21275
rect -13680 21240 -13640 21245
rect -13600 21275 -13560 21280
rect -13600 21245 -13595 21275
rect -13565 21245 -13560 21275
rect -13600 21240 -13560 21245
rect -13520 21275 -13480 21280
rect -13520 21245 -13515 21275
rect -13485 21245 -13480 21275
rect -13520 21240 -13480 21245
rect -13440 21275 -13400 21280
rect -13440 21245 -13435 21275
rect -13405 21245 -13400 21275
rect -13440 21240 -13400 21245
rect -13360 21275 -13320 21280
rect -13360 21245 -13355 21275
rect -13325 21245 -13320 21275
rect -13360 21240 -13320 21245
rect -13280 21275 -13240 21280
rect -13280 21245 -13275 21275
rect -13245 21245 -13240 21275
rect -13280 21240 -13240 21245
rect -13200 21275 -13160 21280
rect -13200 21245 -13195 21275
rect -13165 21245 -13160 21275
rect -13200 21240 -13160 21245
rect -13120 21275 -13080 21280
rect -13120 21245 -13115 21275
rect -13085 21245 -13080 21275
rect -13120 21240 -13080 21245
rect -13040 21275 -13000 21280
rect -13040 21245 -13035 21275
rect -13005 21245 -13000 21275
rect -13040 21240 -13000 21245
rect -12960 21275 -12920 21280
rect -12960 21245 -12955 21275
rect -12925 21245 -12920 21275
rect -12960 21240 -12920 21245
rect -12880 21275 -12840 21280
rect -12880 21245 -12875 21275
rect -12845 21245 -12840 21275
rect -12880 21240 -12840 21245
rect -12800 21275 -12760 21280
rect -12800 21245 -12795 21275
rect -12765 21245 -12760 21275
rect -12800 21240 -12760 21245
rect -12720 21275 -12680 21280
rect -12720 21245 -12715 21275
rect -12685 21245 -12680 21275
rect -12720 21240 -12680 21245
rect -12640 21275 -12600 21280
rect -12640 21245 -12635 21275
rect -12605 21245 -12600 21275
rect -12640 21240 -12600 21245
rect -12560 21275 -12520 21280
rect -12560 21245 -12555 21275
rect -12525 21245 -12520 21275
rect -12560 21240 -12520 21245
rect -12480 21275 -12440 21280
rect -12480 21245 -12475 21275
rect -12445 21245 -12440 21275
rect -12480 21240 -12440 21245
rect -12400 21275 -12360 21280
rect -12400 21245 -12395 21275
rect -12365 21245 -12360 21275
rect -12400 21240 -12360 21245
rect -12320 21275 -12280 21280
rect -12320 21245 -12315 21275
rect -12285 21245 -12280 21275
rect -12320 21240 -12280 21245
rect -12240 21275 -12200 21280
rect -12240 21245 -12235 21275
rect -12205 21245 -12200 21275
rect -12240 21240 -12200 21245
rect -12160 21275 -12120 21280
rect -12160 21245 -12155 21275
rect -12125 21245 -12120 21275
rect -12160 21240 -12120 21245
rect -12080 21275 -12040 21280
rect -12080 21245 -12075 21275
rect -12045 21245 -12040 21275
rect -12080 21240 -12040 21245
rect -12000 21275 -11960 21280
rect -12000 21245 -11995 21275
rect -11965 21245 -11960 21275
rect -12000 21240 -11960 21245
rect -11920 21275 -11880 21280
rect -11920 21245 -11915 21275
rect -11885 21245 -11880 21275
rect -11920 21240 -11880 21245
rect -11840 21275 -11800 21280
rect -11840 21245 -11835 21275
rect -11805 21245 -11800 21275
rect -11840 21240 -11800 21245
rect -11760 21275 -11720 21280
rect -11760 21245 -11755 21275
rect -11725 21245 -11720 21275
rect -11760 21240 -11720 21245
rect -11680 21275 -11640 21280
rect -11680 21245 -11675 21275
rect -11645 21245 -11640 21275
rect -11680 21240 -11640 21245
rect -11600 21275 -11560 21280
rect -11600 21245 -11595 21275
rect -11565 21245 -11560 21275
rect -11600 21240 -11560 21245
rect -11520 21275 -11480 21280
rect -11520 21245 -11515 21275
rect -11485 21245 -11480 21275
rect -11520 21240 -11480 21245
rect -11440 21275 -11400 21280
rect -11440 21245 -11435 21275
rect -11405 21245 -11400 21275
rect -11440 21240 -11400 21245
rect -11360 21275 -11320 21280
rect -11360 21245 -11355 21275
rect -11325 21245 -11320 21275
rect -11360 21240 -11320 21245
rect -11280 21275 -11240 21280
rect -11280 21245 -11275 21275
rect -11245 21245 -11240 21275
rect -11280 21240 -11240 21245
rect -11200 21275 -11160 21280
rect -11200 21245 -11195 21275
rect -11165 21245 -11160 21275
rect -11200 21240 -11160 21245
rect -11120 21275 -11080 21280
rect -11120 21245 -11115 21275
rect -11085 21245 -11080 21275
rect -11120 21240 -11080 21245
rect -11040 21275 -11000 21280
rect -11040 21245 -11035 21275
rect -11005 21245 -11000 21275
rect -11040 21240 -11000 21245
rect -10960 21275 -10920 21280
rect -10960 21245 -10955 21275
rect -10925 21245 -10920 21275
rect -10960 21240 -10920 21245
rect -10880 21275 -10840 21280
rect -10880 21245 -10875 21275
rect -10845 21245 -10840 21275
rect -10880 21240 -10840 21245
rect -10800 21275 -10760 21280
rect -10800 21245 -10795 21275
rect -10765 21245 -10760 21275
rect -10800 21240 -10760 21245
rect -10720 21275 -10680 21280
rect -10720 21245 -10715 21275
rect -10685 21245 -10680 21275
rect -10720 21240 -10680 21245
rect -10640 21275 -10600 21280
rect -10640 21245 -10635 21275
rect -10605 21245 -10600 21275
rect -10640 21240 -10600 21245
rect -10560 21275 -10520 21280
rect -10560 21245 -10555 21275
rect -10525 21245 -10520 21275
rect -10560 21240 -10520 21245
rect -10480 21275 -10440 21280
rect -10480 21245 -10475 21275
rect -10445 21245 -10440 21275
rect -10480 21240 -10440 21245
rect -10400 21275 -10360 21280
rect -10400 21245 -10395 21275
rect -10365 21245 -10360 21275
rect -10400 21240 -10360 21245
rect -10320 21275 -10280 21280
rect -10320 21245 -10315 21275
rect -10285 21245 -10280 21275
rect -10320 21240 -10280 21245
rect -10240 21275 -10200 21280
rect -10240 21245 -10235 21275
rect -10205 21245 -10200 21275
rect -10240 21240 -10200 21245
rect -10160 21275 -10120 21280
rect -10160 21245 -10155 21275
rect -10125 21245 -10120 21275
rect -10160 21240 -10120 21245
rect -10080 21275 -10040 21280
rect -10080 21245 -10075 21275
rect -10045 21245 -10040 21275
rect -10080 21240 -10040 21245
rect -10000 21275 -9960 21280
rect -10000 21245 -9995 21275
rect -9965 21245 -9960 21275
rect -10000 21240 -9960 21245
rect -9920 21275 -9880 21280
rect -9920 21245 -9915 21275
rect -9885 21245 -9880 21275
rect -9920 21240 -9880 21245
rect -9840 21275 -9800 21280
rect -9840 21245 -9835 21275
rect -9805 21245 -9800 21275
rect -9840 21240 -9800 21245
rect -9760 21275 -9720 21280
rect -9760 21245 -9755 21275
rect -9725 21245 -9720 21275
rect -9760 21240 -9720 21245
rect -9680 21275 -9640 21280
rect -9680 21245 -9675 21275
rect -9645 21245 -9640 21275
rect -9680 21240 -9640 21245
rect -9600 21275 -9560 21280
rect -9600 21245 -9595 21275
rect -9565 21245 -9560 21275
rect -9600 21240 -9560 21245
rect -9520 21275 -9480 21280
rect -9520 21245 -9515 21275
rect -9485 21245 -9480 21275
rect -9520 21240 -9480 21245
rect -9440 21275 -9400 21280
rect -9440 21245 -9435 21275
rect -9405 21245 -9400 21275
rect -9440 21240 -9400 21245
rect -9360 21275 -9320 21280
rect -9360 21245 -9355 21275
rect -9325 21245 -9320 21275
rect -9360 21240 -9320 21245
rect -9280 21275 -9240 21280
rect -9280 21245 -9275 21275
rect -9245 21245 -9240 21275
rect -9280 21240 -9240 21245
rect -9200 21275 -9160 21280
rect -9200 21245 -9195 21275
rect -9165 21245 -9160 21275
rect -9200 21240 -9160 21245
rect -9120 21275 -9080 21280
rect -9120 21245 -9115 21275
rect -9085 21245 -9080 21275
rect -9120 21240 -9080 21245
rect -9040 21275 -9000 21280
rect -9040 21245 -9035 21275
rect -9005 21245 -9000 21275
rect -9040 21240 -9000 21245
rect -8960 21275 -8920 21280
rect -8960 21245 -8955 21275
rect -8925 21245 -8920 21275
rect -8960 21240 -8920 21245
rect -8880 21275 -8840 21280
rect -8880 21245 -8875 21275
rect -8845 21245 -8840 21275
rect -8880 21240 -8840 21245
rect -8800 21275 -8760 21280
rect -8800 21245 -8795 21275
rect -8765 21245 -8760 21275
rect -8800 21240 -8760 21245
rect -8720 21275 -8680 21280
rect -8720 21245 -8715 21275
rect -8685 21245 -8680 21275
rect -8720 21240 -8680 21245
rect -8640 21275 -8600 21280
rect -8640 21245 -8635 21275
rect -8605 21245 -8600 21275
rect -8640 21240 -8600 21245
rect -8560 21275 -8520 21280
rect -8560 21245 -8555 21275
rect -8525 21245 -8520 21275
rect -8560 21240 -8520 21245
rect -8480 21275 -8440 21280
rect -8480 21245 -8475 21275
rect -8445 21245 -8440 21275
rect -8480 21240 -8440 21245
rect -8400 21275 -8360 21280
rect -8400 21245 -8395 21275
rect -8365 21245 -8360 21275
rect -8400 21240 -8360 21245
rect -8320 21275 -8280 21280
rect -8320 21245 -8315 21275
rect -8285 21245 -8280 21275
rect -8320 21240 -8280 21245
rect -8240 21275 -8200 21280
rect -8240 21245 -8235 21275
rect -8205 21245 -8200 21275
rect -8240 21240 -8200 21245
rect -8160 21275 -8120 21280
rect -8160 21245 -8155 21275
rect -8125 21245 -8120 21275
rect -8160 21240 -8120 21245
rect -8080 21275 -8040 21280
rect -8080 21245 -8075 21275
rect -8045 21245 -8040 21275
rect -8080 21240 -8040 21245
rect -8000 21275 -7960 21280
rect -8000 21245 -7995 21275
rect -7965 21245 -7960 21275
rect -8000 21240 -7960 21245
rect -7920 21275 -7880 21280
rect -7920 21245 -7915 21275
rect -7885 21245 -7880 21275
rect -7920 21240 -7880 21245
rect -7840 21275 -7800 21280
rect -7840 21245 -7835 21275
rect -7805 21245 -7800 21275
rect -7840 21240 -7800 21245
rect -7760 21275 -7720 21280
rect -7760 21245 -7755 21275
rect -7725 21245 -7720 21275
rect -7760 21240 -7720 21245
rect -7680 21275 -7640 21280
rect -7680 21245 -7675 21275
rect -7645 21245 -7640 21275
rect -7680 21240 -7640 21245
rect -7600 21275 -7560 21280
rect -7600 21245 -7595 21275
rect -7565 21245 -7560 21275
rect -7600 21240 -7560 21245
rect -7520 21275 -7480 21280
rect -7520 21245 -7515 21275
rect -7485 21245 -7480 21275
rect -7520 21240 -7480 21245
rect -7440 21275 -7400 21280
rect -7440 21245 -7435 21275
rect -7405 21245 -7400 21275
rect -7440 21240 -7400 21245
rect -7360 21275 -7320 21280
rect -7360 21245 -7355 21275
rect -7325 21245 -7320 21275
rect -7360 21240 -7320 21245
rect -7280 21275 -7240 21280
rect -7280 21245 -7275 21275
rect -7245 21245 -7240 21275
rect -7280 21240 -7240 21245
rect -7200 21275 -7160 21280
rect -7200 21245 -7195 21275
rect -7165 21245 -7160 21275
rect -7200 21240 -7160 21245
rect -7120 21275 -7080 21280
rect -7120 21245 -7115 21275
rect -7085 21245 -7080 21275
rect -7120 21240 -7080 21245
rect -7040 21275 -7000 21280
rect -7040 21245 -7035 21275
rect -7005 21245 -7000 21275
rect -7040 21240 -7000 21245
rect -6960 21275 -6920 21280
rect -6960 21245 -6955 21275
rect -6925 21245 -6920 21275
rect -6960 21240 -6920 21245
rect -6880 21275 -6840 21280
rect -6880 21245 -6875 21275
rect -6845 21245 -6840 21275
rect -6880 21240 -6840 21245
rect -6800 21275 -6760 21280
rect -6800 21245 -6795 21275
rect -6765 21245 -6760 21275
rect -6800 21240 -6760 21245
rect -6720 21275 -6680 21280
rect -6720 21245 -6715 21275
rect -6685 21245 -6680 21275
rect -6720 21240 -6680 21245
rect -6640 21275 -6600 21280
rect -6640 21245 -6635 21275
rect -6605 21245 -6600 21275
rect -6640 21240 -6600 21245
rect -6560 21275 -6520 21280
rect -6560 21245 -6555 21275
rect -6525 21245 -6520 21275
rect -6560 21240 -6520 21245
rect -6480 21275 -6440 21280
rect -6480 21245 -6475 21275
rect -6445 21245 -6440 21275
rect -6480 21240 -6440 21245
rect -6400 21275 -6360 21280
rect -6400 21245 -6395 21275
rect -6365 21245 -6360 21275
rect -6400 21240 -6360 21245
rect -6320 21275 -6280 21280
rect -6320 21245 -6315 21275
rect -6285 21245 -6280 21275
rect -6320 21240 -6280 21245
rect -6240 21275 -6200 21280
rect -6240 21245 -6235 21275
rect -6205 21245 -6200 21275
rect -6240 21240 -6200 21245
rect -6160 21275 -6120 21280
rect -6160 21245 -6155 21275
rect -6125 21245 -6120 21275
rect -6160 21240 -6120 21245
rect -5680 21275 -5640 21280
rect -5680 21245 -5675 21275
rect -5645 21245 -5640 21275
rect -5680 21240 -5640 21245
rect -5600 21275 -5560 21280
rect -5600 21245 -5595 21275
rect -5565 21245 -5560 21275
rect -5600 21240 -5560 21245
rect -5520 21275 -5480 21280
rect -5520 21245 -5515 21275
rect -5485 21245 -5480 21275
rect -5520 21240 -5480 21245
rect -5440 21275 -5400 21280
rect -5440 21245 -5435 21275
rect -5405 21245 -5400 21275
rect -5440 21240 -5400 21245
rect -5360 21275 -5320 21280
rect -5360 21245 -5355 21275
rect -5325 21245 -5320 21275
rect -5360 21240 -5320 21245
rect -5280 21275 -5240 21280
rect -5280 21245 -5275 21275
rect -5245 21245 -5240 21275
rect -5280 21240 -5240 21245
rect -5200 21275 -5160 21280
rect -5200 21245 -5195 21275
rect -5165 21245 -5160 21275
rect -5200 21240 -5160 21245
rect -5120 21275 -5080 21280
rect -5120 21245 -5115 21275
rect -5085 21245 -5080 21275
rect -5120 21240 -5080 21245
rect -5040 21275 -5000 21280
rect -5040 21245 -5035 21275
rect -5005 21245 -5000 21275
rect -5040 21240 -5000 21245
rect -4960 21275 -4920 21280
rect -4960 21245 -4955 21275
rect -4925 21245 -4920 21275
rect -4960 21240 -4920 21245
rect -4880 21275 -4840 21280
rect -4880 21245 -4875 21275
rect -4845 21245 -4840 21275
rect -4880 21240 -4840 21245
rect -4800 21275 -4760 21280
rect -4800 21245 -4795 21275
rect -4765 21245 -4760 21275
rect -4800 21240 -4760 21245
rect -4720 21275 -4680 21280
rect -4720 21245 -4715 21275
rect -4685 21245 -4680 21275
rect -4720 21240 -4680 21245
rect -4640 21275 -4600 21280
rect -4640 21245 -4635 21275
rect -4605 21245 -4600 21275
rect -4640 21240 -4600 21245
rect -4560 21275 -4520 21280
rect -4560 21245 -4555 21275
rect -4525 21245 -4520 21275
rect -4560 21240 -4520 21245
rect -4480 21275 -4440 21280
rect -4480 21245 -4475 21275
rect -4445 21245 -4440 21275
rect -4480 21240 -4440 21245
rect -4400 21275 -4360 21280
rect -4400 21245 -4395 21275
rect -4365 21245 -4360 21275
rect -4400 21240 -4360 21245
rect -4320 21275 -4280 21280
rect -4320 21245 -4315 21275
rect -4285 21245 -4280 21275
rect -4320 21240 -4280 21245
rect -4240 21275 -4200 21280
rect -4240 21245 -4235 21275
rect -4205 21245 -4200 21275
rect -4240 21240 -4200 21245
rect -4160 21275 -4120 21280
rect -4160 21245 -4155 21275
rect -4125 21245 -4120 21275
rect -4160 21240 -4120 21245
rect -4080 21275 -4040 21280
rect -4080 21245 -4075 21275
rect -4045 21245 -4040 21275
rect -4080 21240 -4040 21245
rect -4000 21275 -3960 21280
rect -4000 21245 -3995 21275
rect -3965 21245 -3960 21275
rect -4000 21240 -3960 21245
rect -3920 21275 -3880 21280
rect -3920 21245 -3915 21275
rect -3885 21245 -3880 21275
rect -3920 21240 -3880 21245
rect -3840 21275 -3800 21280
rect -3840 21245 -3835 21275
rect -3805 21245 -3800 21275
rect -3840 21240 -3800 21245
rect -3760 21275 -3720 21280
rect -3760 21245 -3755 21275
rect -3725 21245 -3720 21275
rect -3760 21240 -3720 21245
rect -3680 21275 -3640 21280
rect -3680 21245 -3675 21275
rect -3645 21245 -3640 21275
rect -3680 21240 -3640 21245
rect -3600 21275 -3560 21280
rect -3600 21245 -3595 21275
rect -3565 21245 -3560 21275
rect -3600 21240 -3560 21245
rect -3520 21275 -3480 21280
rect -3520 21245 -3515 21275
rect -3485 21245 -3480 21275
rect -3520 21240 -3480 21245
rect -3440 21275 -3400 21280
rect -3440 21245 -3435 21275
rect -3405 21245 -3400 21275
rect -3440 21240 -3400 21245
rect -3360 21275 -3320 21280
rect -3360 21245 -3355 21275
rect -3325 21245 -3320 21275
rect -3360 21240 -3320 21245
rect -3280 21275 -3240 21280
rect -3280 21245 -3275 21275
rect -3245 21245 -3240 21275
rect -3280 21240 -3240 21245
rect -3200 21275 -3160 21280
rect -3200 21245 -3195 21275
rect -3165 21245 -3160 21275
rect -3200 21240 -3160 21245
rect -3120 21275 -3080 21280
rect -3120 21245 -3115 21275
rect -3085 21245 -3080 21275
rect -3120 21240 -3080 21245
rect -3040 21275 -3000 21280
rect -3040 21245 -3035 21275
rect -3005 21245 -3000 21275
rect -3040 21240 -3000 21245
rect -2960 21275 -2920 21280
rect -2960 21245 -2955 21275
rect -2925 21245 -2920 21275
rect -2960 21240 -2920 21245
rect -2880 21275 -2840 21280
rect -2880 21245 -2875 21275
rect -2845 21245 -2840 21275
rect -2880 21240 -2840 21245
rect -2800 21275 -2760 21280
rect -2800 21245 -2795 21275
rect -2765 21245 -2760 21275
rect -2800 21240 -2760 21245
rect -2720 21275 -2680 21280
rect -2720 21245 -2715 21275
rect -2685 21245 -2680 21275
rect -2720 21240 -2680 21245
rect -2640 21275 -2600 21280
rect -2640 21245 -2635 21275
rect -2605 21245 -2600 21275
rect -2640 21240 -2600 21245
rect -2560 21275 -2520 21280
rect -2560 21245 -2555 21275
rect -2525 21245 -2520 21275
rect -2560 21240 -2520 21245
rect -2480 21275 -2440 21280
rect -2480 21245 -2475 21275
rect -2445 21245 -2440 21275
rect -2480 21240 -2440 21245
rect -2400 21275 -2360 21280
rect -2400 21245 -2395 21275
rect -2365 21245 -2360 21275
rect -2400 21240 -2360 21245
rect -2320 21275 -2280 21280
rect -2320 21245 -2315 21275
rect -2285 21245 -2280 21275
rect -2320 21240 -2280 21245
rect -2240 21275 -2200 21280
rect -2240 21245 -2235 21275
rect -2205 21245 -2200 21275
rect -2240 21240 -2200 21245
rect -2160 21275 -2120 21280
rect -2160 21245 -2155 21275
rect -2125 21245 -2120 21275
rect -2160 21240 -2120 21245
rect -2080 21275 -2040 21280
rect -2080 21245 -2075 21275
rect -2045 21245 -2040 21275
rect -2080 21240 -2040 21245
rect -2000 21275 -1960 21280
rect -2000 21245 -1995 21275
rect -1965 21245 -1960 21275
rect -2000 21240 -1960 21245
rect -1840 21275 -1800 21280
rect -1840 21245 -1835 21275
rect -1805 21245 -1800 21275
rect -1840 21240 -1800 21245
rect -1760 21275 -1720 21280
rect -1760 21245 -1755 21275
rect -1725 21245 -1720 21275
rect -1760 21240 -1720 21245
rect -1680 21275 -1640 21280
rect -1680 21245 -1675 21275
rect -1645 21245 -1640 21275
rect -1680 21240 -1640 21245
rect -1520 21275 -1480 21280
rect -1520 21245 -1515 21275
rect -1485 21245 -1480 21275
rect -1520 21240 -1480 21245
rect -1360 21275 -1320 21280
rect -1360 21245 -1355 21275
rect -1325 21245 -1320 21275
rect -1360 21240 -1320 21245
rect -1280 21275 -1240 21280
rect -1280 21245 -1275 21275
rect -1245 21245 -1240 21275
rect -1280 21240 -1240 21245
rect -1200 21275 -1160 21280
rect -1200 21245 -1195 21275
rect -1165 21245 -1160 21275
rect -1200 21240 -1160 21245
rect -1120 21275 -1080 21280
rect -1120 21245 -1115 21275
rect -1085 21245 -1080 21275
rect -1120 21240 -1080 21245
rect -1040 21275 -1000 21280
rect -1040 21245 -1035 21275
rect -1005 21245 -1000 21275
rect -1040 21240 -1000 21245
rect -880 21275 -840 21280
rect -880 21245 -875 21275
rect -845 21245 -840 21275
rect -880 21240 -840 21245
rect -720 21275 -680 21280
rect -720 21245 -715 21275
rect -685 21245 -680 21275
rect -720 21240 -680 21245
rect -560 21275 -520 21280
rect -560 21245 -555 21275
rect -525 21245 -520 21275
rect -560 21240 -520 21245
rect -14960 21115 -14920 21120
rect -14960 21085 -14955 21115
rect -14925 21085 -14920 21115
rect -14960 21080 -14920 21085
rect -14880 21115 -14840 21120
rect -14880 21085 -14875 21115
rect -14845 21085 -14840 21115
rect -14880 21080 -14840 21085
rect -14800 21115 -14760 21120
rect -14800 21085 -14795 21115
rect -14765 21085 -14760 21115
rect -14800 21080 -14760 21085
rect -14720 21115 -14680 21120
rect -14720 21085 -14715 21115
rect -14685 21085 -14680 21115
rect -14720 21080 -14680 21085
rect -14640 21115 -14600 21120
rect -14640 21085 -14635 21115
rect -14605 21085 -14600 21115
rect -14640 21080 -14600 21085
rect -14560 21115 -14520 21120
rect -14560 21085 -14555 21115
rect -14525 21085 -14520 21115
rect -14560 21080 -14520 21085
rect -14480 21115 -14440 21120
rect -14480 21085 -14475 21115
rect -14445 21085 -14440 21115
rect -14480 21080 -14440 21085
rect -14400 21115 -14360 21120
rect -14400 21085 -14395 21115
rect -14365 21085 -14360 21115
rect -14400 21080 -14360 21085
rect -14320 21115 -14280 21120
rect -14320 21085 -14315 21115
rect -14285 21085 -14280 21115
rect -14320 21080 -14280 21085
rect -14240 21115 -14200 21120
rect -14240 21085 -14235 21115
rect -14205 21085 -14200 21115
rect -14240 21080 -14200 21085
rect -14160 21115 -14120 21120
rect -14160 21085 -14155 21115
rect -14125 21085 -14120 21115
rect -14160 21080 -14120 21085
rect -14080 21115 -14040 21120
rect -14080 21085 -14075 21115
rect -14045 21085 -14040 21115
rect -14080 21080 -14040 21085
rect -14000 21115 -13960 21120
rect -14000 21085 -13995 21115
rect -13965 21085 -13960 21115
rect -14000 21080 -13960 21085
rect -13920 21115 -13880 21120
rect -13920 21085 -13915 21115
rect -13885 21085 -13880 21115
rect -13920 21080 -13880 21085
rect -13840 21115 -13800 21120
rect -13840 21085 -13835 21115
rect -13805 21085 -13800 21115
rect -13840 21080 -13800 21085
rect -13760 21115 -13720 21120
rect -13760 21085 -13755 21115
rect -13725 21085 -13720 21115
rect -13760 21080 -13720 21085
rect -13680 21115 -13640 21120
rect -13680 21085 -13675 21115
rect -13645 21085 -13640 21115
rect -13680 21080 -13640 21085
rect -13600 21115 -13560 21120
rect -13600 21085 -13595 21115
rect -13565 21085 -13560 21115
rect -13600 21080 -13560 21085
rect -13520 21115 -13480 21120
rect -13520 21085 -13515 21115
rect -13485 21085 -13480 21115
rect -13520 21080 -13480 21085
rect -13440 21115 -13400 21120
rect -13440 21085 -13435 21115
rect -13405 21085 -13400 21115
rect -13440 21080 -13400 21085
rect -13360 21115 -13320 21120
rect -13360 21085 -13355 21115
rect -13325 21085 -13320 21115
rect -13360 21080 -13320 21085
rect -13280 21115 -13240 21120
rect -13280 21085 -13275 21115
rect -13245 21085 -13240 21115
rect -13280 21080 -13240 21085
rect -13200 21115 -13160 21120
rect -13200 21085 -13195 21115
rect -13165 21085 -13160 21115
rect -13200 21080 -13160 21085
rect -13120 21115 -13080 21120
rect -13120 21085 -13115 21115
rect -13085 21085 -13080 21115
rect -13120 21080 -13080 21085
rect -13040 21115 -13000 21120
rect -13040 21085 -13035 21115
rect -13005 21085 -13000 21115
rect -13040 21080 -13000 21085
rect -12960 21115 -12920 21120
rect -12960 21085 -12955 21115
rect -12925 21085 -12920 21115
rect -12960 21080 -12920 21085
rect -12880 21115 -12840 21120
rect -12880 21085 -12875 21115
rect -12845 21085 -12840 21115
rect -12880 21080 -12840 21085
rect -12800 21115 -12760 21120
rect -12800 21085 -12795 21115
rect -12765 21085 -12760 21115
rect -12800 21080 -12760 21085
rect -12720 21115 -12680 21120
rect -12720 21085 -12715 21115
rect -12685 21085 -12680 21115
rect -12720 21080 -12680 21085
rect -12640 21115 -12600 21120
rect -12640 21085 -12635 21115
rect -12605 21085 -12600 21115
rect -12640 21080 -12600 21085
rect -12560 21115 -12520 21120
rect -12560 21085 -12555 21115
rect -12525 21085 -12520 21115
rect -12560 21080 -12520 21085
rect -12480 21115 -12440 21120
rect -12480 21085 -12475 21115
rect -12445 21085 -12440 21115
rect -12480 21080 -12440 21085
rect -12400 21115 -12360 21120
rect -12400 21085 -12395 21115
rect -12365 21085 -12360 21115
rect -12400 21080 -12360 21085
rect -12320 21115 -12280 21120
rect -12320 21085 -12315 21115
rect -12285 21085 -12280 21115
rect -12320 21080 -12280 21085
rect -12240 21115 -12200 21120
rect -12240 21085 -12235 21115
rect -12205 21085 -12200 21115
rect -12240 21080 -12200 21085
rect -12160 21115 -12120 21120
rect -12160 21085 -12155 21115
rect -12125 21085 -12120 21115
rect -12160 21080 -12120 21085
rect -12080 21115 -12040 21120
rect -12080 21085 -12075 21115
rect -12045 21085 -12040 21115
rect -12080 21080 -12040 21085
rect -12000 21115 -11960 21120
rect -12000 21085 -11995 21115
rect -11965 21085 -11960 21115
rect -12000 21080 -11960 21085
rect -11920 21115 -11880 21120
rect -11920 21085 -11915 21115
rect -11885 21085 -11880 21115
rect -11920 21080 -11880 21085
rect -11840 21115 -11800 21120
rect -11840 21085 -11835 21115
rect -11805 21085 -11800 21115
rect -11840 21080 -11800 21085
rect -11760 21115 -11720 21120
rect -11760 21085 -11755 21115
rect -11725 21085 -11720 21115
rect -11760 21080 -11720 21085
rect -11680 21115 -11640 21120
rect -11680 21085 -11675 21115
rect -11645 21085 -11640 21115
rect -11680 21080 -11640 21085
rect -11600 21115 -11560 21120
rect -11600 21085 -11595 21115
rect -11565 21085 -11560 21115
rect -11600 21080 -11560 21085
rect -11520 21115 -11480 21120
rect -11520 21085 -11515 21115
rect -11485 21085 -11480 21115
rect -11520 21080 -11480 21085
rect -11440 21115 -11400 21120
rect -11440 21085 -11435 21115
rect -11405 21085 -11400 21115
rect -11440 21080 -11400 21085
rect -11360 21115 -11320 21120
rect -11360 21085 -11355 21115
rect -11325 21085 -11320 21115
rect -11360 21080 -11320 21085
rect -11280 21115 -11240 21120
rect -11280 21085 -11275 21115
rect -11245 21085 -11240 21115
rect -11280 21080 -11240 21085
rect -11200 21115 -11160 21120
rect -11200 21085 -11195 21115
rect -11165 21085 -11160 21115
rect -11200 21080 -11160 21085
rect -11120 21115 -11080 21120
rect -11120 21085 -11115 21115
rect -11085 21085 -11080 21115
rect -11120 21080 -11080 21085
rect -11040 21115 -11000 21120
rect -11040 21085 -11035 21115
rect -11005 21085 -11000 21115
rect -11040 21080 -11000 21085
rect -10960 21115 -10920 21120
rect -10960 21085 -10955 21115
rect -10925 21085 -10920 21115
rect -10960 21080 -10920 21085
rect -10880 21115 -10840 21120
rect -10880 21085 -10875 21115
rect -10845 21085 -10840 21115
rect -10880 21080 -10840 21085
rect -10800 21115 -10760 21120
rect -10800 21085 -10795 21115
rect -10765 21085 -10760 21115
rect -10800 21080 -10760 21085
rect -10720 21115 -10680 21120
rect -10720 21085 -10715 21115
rect -10685 21085 -10680 21115
rect -10720 21080 -10680 21085
rect -10640 21115 -10600 21120
rect -10640 21085 -10635 21115
rect -10605 21085 -10600 21115
rect -10640 21080 -10600 21085
rect -10560 21115 -10520 21120
rect -10560 21085 -10555 21115
rect -10525 21085 -10520 21115
rect -10560 21080 -10520 21085
rect -10480 21115 -10440 21120
rect -10480 21085 -10475 21115
rect -10445 21085 -10440 21115
rect -10480 21080 -10440 21085
rect -10400 21115 -10360 21120
rect -10400 21085 -10395 21115
rect -10365 21085 -10360 21115
rect -10400 21080 -10360 21085
rect -10320 21115 -10280 21120
rect -10320 21085 -10315 21115
rect -10285 21085 -10280 21115
rect -10320 21080 -10280 21085
rect -10240 21115 -10200 21120
rect -10240 21085 -10235 21115
rect -10205 21085 -10200 21115
rect -10240 21080 -10200 21085
rect -10160 21115 -10120 21120
rect -10160 21085 -10155 21115
rect -10125 21085 -10120 21115
rect -10160 21080 -10120 21085
rect -10080 21115 -10040 21120
rect -10080 21085 -10075 21115
rect -10045 21085 -10040 21115
rect -10080 21080 -10040 21085
rect -10000 21115 -9960 21120
rect -10000 21085 -9995 21115
rect -9965 21085 -9960 21115
rect -10000 21080 -9960 21085
rect -9920 21115 -9880 21120
rect -9920 21085 -9915 21115
rect -9885 21085 -9880 21115
rect -9920 21080 -9880 21085
rect -9840 21115 -9800 21120
rect -9840 21085 -9835 21115
rect -9805 21085 -9800 21115
rect -9840 21080 -9800 21085
rect -9760 21115 -9720 21120
rect -9760 21085 -9755 21115
rect -9725 21085 -9720 21115
rect -9760 21080 -9720 21085
rect -9680 21115 -9640 21120
rect -9680 21085 -9675 21115
rect -9645 21085 -9640 21115
rect -9680 21080 -9640 21085
rect -9600 21115 -9560 21120
rect -9600 21085 -9595 21115
rect -9565 21085 -9560 21115
rect -9600 21080 -9560 21085
rect -9520 21115 -9480 21120
rect -9520 21085 -9515 21115
rect -9485 21085 -9480 21115
rect -9520 21080 -9480 21085
rect -9440 21115 -9400 21120
rect -9440 21085 -9435 21115
rect -9405 21085 -9400 21115
rect -9440 21080 -9400 21085
rect -9360 21115 -9320 21120
rect -9360 21085 -9355 21115
rect -9325 21085 -9320 21115
rect -9360 21080 -9320 21085
rect -9280 21115 -9240 21120
rect -9280 21085 -9275 21115
rect -9245 21085 -9240 21115
rect -9280 21080 -9240 21085
rect -9200 21115 -9160 21120
rect -9200 21085 -9195 21115
rect -9165 21085 -9160 21115
rect -9200 21080 -9160 21085
rect -9120 21115 -9080 21120
rect -9120 21085 -9115 21115
rect -9085 21085 -9080 21115
rect -9120 21080 -9080 21085
rect -9040 21115 -9000 21120
rect -9040 21085 -9035 21115
rect -9005 21085 -9000 21115
rect -9040 21080 -9000 21085
rect -8960 21115 -8920 21120
rect -8960 21085 -8955 21115
rect -8925 21085 -8920 21115
rect -8960 21080 -8920 21085
rect -8880 21115 -8840 21120
rect -8880 21085 -8875 21115
rect -8845 21085 -8840 21115
rect -8880 21080 -8840 21085
rect -8800 21115 -8760 21120
rect -8800 21085 -8795 21115
rect -8765 21085 -8760 21115
rect -8800 21080 -8760 21085
rect -8720 21115 -8680 21120
rect -8720 21085 -8715 21115
rect -8685 21085 -8680 21115
rect -8720 21080 -8680 21085
rect -8640 21115 -8600 21120
rect -8640 21085 -8635 21115
rect -8605 21085 -8600 21115
rect -8640 21080 -8600 21085
rect -8560 21115 -8520 21120
rect -8560 21085 -8555 21115
rect -8525 21085 -8520 21115
rect -8560 21080 -8520 21085
rect -8480 21115 -8440 21120
rect -8480 21085 -8475 21115
rect -8445 21085 -8440 21115
rect -8480 21080 -8440 21085
rect -8400 21115 -8360 21120
rect -8400 21085 -8395 21115
rect -8365 21085 -8360 21115
rect -8400 21080 -8360 21085
rect -8320 21115 -8280 21120
rect -8320 21085 -8315 21115
rect -8285 21085 -8280 21115
rect -8320 21080 -8280 21085
rect -8240 21115 -8200 21120
rect -8240 21085 -8235 21115
rect -8205 21085 -8200 21115
rect -8240 21080 -8200 21085
rect -8160 21115 -8120 21120
rect -8160 21085 -8155 21115
rect -8125 21085 -8120 21115
rect -8160 21080 -8120 21085
rect -8080 21115 -8040 21120
rect -8080 21085 -8075 21115
rect -8045 21085 -8040 21115
rect -8080 21080 -8040 21085
rect -8000 21115 -7960 21120
rect -8000 21085 -7995 21115
rect -7965 21085 -7960 21115
rect -8000 21080 -7960 21085
rect -7920 21115 -7880 21120
rect -7920 21085 -7915 21115
rect -7885 21085 -7880 21115
rect -7920 21080 -7880 21085
rect -7840 21115 -7800 21120
rect -7840 21085 -7835 21115
rect -7805 21085 -7800 21115
rect -7840 21080 -7800 21085
rect -7760 21115 -7720 21120
rect -7760 21085 -7755 21115
rect -7725 21085 -7720 21115
rect -7760 21080 -7720 21085
rect -7680 21115 -7640 21120
rect -7680 21085 -7675 21115
rect -7645 21085 -7640 21115
rect -7680 21080 -7640 21085
rect -7600 21115 -7560 21120
rect -7600 21085 -7595 21115
rect -7565 21085 -7560 21115
rect -7600 21080 -7560 21085
rect -7520 21115 -7480 21120
rect -7520 21085 -7515 21115
rect -7485 21085 -7480 21115
rect -7520 21080 -7480 21085
rect -7440 21115 -7400 21120
rect -7440 21085 -7435 21115
rect -7405 21085 -7400 21115
rect -7440 21080 -7400 21085
rect -7360 21115 -7320 21120
rect -7360 21085 -7355 21115
rect -7325 21085 -7320 21115
rect -7360 21080 -7320 21085
rect -7280 21115 -7240 21120
rect -7280 21085 -7275 21115
rect -7245 21085 -7240 21115
rect -7280 21080 -7240 21085
rect -7200 21115 -7160 21120
rect -7200 21085 -7195 21115
rect -7165 21085 -7160 21115
rect -7200 21080 -7160 21085
rect -7120 21115 -7080 21120
rect -7120 21085 -7115 21115
rect -7085 21085 -7080 21115
rect -7120 21080 -7080 21085
rect -7040 21115 -7000 21120
rect -7040 21085 -7035 21115
rect -7005 21085 -7000 21115
rect -7040 21080 -7000 21085
rect -6960 21115 -6920 21120
rect -6960 21085 -6955 21115
rect -6925 21085 -6920 21115
rect -6960 21080 -6920 21085
rect -6880 21115 -6840 21120
rect -6880 21085 -6875 21115
rect -6845 21085 -6840 21115
rect -6880 21080 -6840 21085
rect -6800 21115 -6760 21120
rect -6800 21085 -6795 21115
rect -6765 21085 -6760 21115
rect -6800 21080 -6760 21085
rect -6720 21115 -6680 21120
rect -6720 21085 -6715 21115
rect -6685 21085 -6680 21115
rect -6720 21080 -6680 21085
rect -6640 21115 -6600 21120
rect -6640 21085 -6635 21115
rect -6605 21085 -6600 21115
rect -6640 21080 -6600 21085
rect -6560 21115 -6520 21120
rect -6560 21085 -6555 21115
rect -6525 21085 -6520 21115
rect -6560 21080 -6520 21085
rect -6480 21115 -6440 21120
rect -6480 21085 -6475 21115
rect -6445 21085 -6440 21115
rect -6480 21080 -6440 21085
rect -6400 21115 -6360 21120
rect -6400 21085 -6395 21115
rect -6365 21085 -6360 21115
rect -6400 21080 -6360 21085
rect -6320 21115 -6280 21120
rect -6320 21085 -6315 21115
rect -6285 21085 -6280 21115
rect -6320 21080 -6280 21085
rect -6240 21115 -6200 21120
rect -6240 21085 -6235 21115
rect -6205 21085 -6200 21115
rect -6240 21080 -6200 21085
rect -6160 21115 -6120 21120
rect -6160 21085 -6155 21115
rect -6125 21085 -6120 21115
rect -6160 21080 -6120 21085
rect -5680 21115 -5640 21120
rect -5680 21085 -5675 21115
rect -5645 21085 -5640 21115
rect -5680 21080 -5640 21085
rect -5600 21115 -5560 21120
rect -5600 21085 -5595 21115
rect -5565 21085 -5560 21115
rect -5600 21080 -5560 21085
rect -5520 21115 -5480 21120
rect -5520 21085 -5515 21115
rect -5485 21085 -5480 21115
rect -5520 21080 -5480 21085
rect -5440 21115 -5400 21120
rect -5440 21085 -5435 21115
rect -5405 21085 -5400 21115
rect -5440 21080 -5400 21085
rect -5360 21115 -5320 21120
rect -5360 21085 -5355 21115
rect -5325 21085 -5320 21115
rect -5360 21080 -5320 21085
rect -5280 21115 -5240 21120
rect -5280 21085 -5275 21115
rect -5245 21085 -5240 21115
rect -5280 21080 -5240 21085
rect -5200 21115 -5160 21120
rect -5200 21085 -5195 21115
rect -5165 21085 -5160 21115
rect -5200 21080 -5160 21085
rect -5120 21115 -5080 21120
rect -5120 21085 -5115 21115
rect -5085 21085 -5080 21115
rect -5120 21080 -5080 21085
rect -5040 21115 -5000 21120
rect -5040 21085 -5035 21115
rect -5005 21085 -5000 21115
rect -5040 21080 -5000 21085
rect -4960 21115 -4920 21120
rect -4960 21085 -4955 21115
rect -4925 21085 -4920 21115
rect -4960 21080 -4920 21085
rect -4880 21115 -4840 21120
rect -4880 21085 -4875 21115
rect -4845 21085 -4840 21115
rect -4880 21080 -4840 21085
rect -4800 21115 -4760 21120
rect -4800 21085 -4795 21115
rect -4765 21085 -4760 21115
rect -4800 21080 -4760 21085
rect -4720 21115 -4680 21120
rect -4720 21085 -4715 21115
rect -4685 21085 -4680 21115
rect -4720 21080 -4680 21085
rect -4640 21115 -4600 21120
rect -4640 21085 -4635 21115
rect -4605 21085 -4600 21115
rect -4640 21080 -4600 21085
rect -4560 21115 -4520 21120
rect -4560 21085 -4555 21115
rect -4525 21085 -4520 21115
rect -4560 21080 -4520 21085
rect -4480 21115 -4440 21120
rect -4480 21085 -4475 21115
rect -4445 21085 -4440 21115
rect -4480 21080 -4440 21085
rect -4400 21115 -4360 21120
rect -4400 21085 -4395 21115
rect -4365 21085 -4360 21115
rect -4400 21080 -4360 21085
rect -4320 21115 -4280 21120
rect -4320 21085 -4315 21115
rect -4285 21085 -4280 21115
rect -4320 21080 -4280 21085
rect -4240 21115 -4200 21120
rect -4240 21085 -4235 21115
rect -4205 21085 -4200 21115
rect -4240 21080 -4200 21085
rect -4160 21115 -4120 21120
rect -4160 21085 -4155 21115
rect -4125 21085 -4120 21115
rect -4160 21080 -4120 21085
rect -4080 21115 -4040 21120
rect -4080 21085 -4075 21115
rect -4045 21085 -4040 21115
rect -4080 21080 -4040 21085
rect -4000 21115 -3960 21120
rect -4000 21085 -3995 21115
rect -3965 21085 -3960 21115
rect -4000 21080 -3960 21085
rect -3920 21115 -3880 21120
rect -3920 21085 -3915 21115
rect -3885 21085 -3880 21115
rect -3920 21080 -3880 21085
rect -3840 21115 -3800 21120
rect -3840 21085 -3835 21115
rect -3805 21085 -3800 21115
rect -3840 21080 -3800 21085
rect -3760 21115 -3720 21120
rect -3760 21085 -3755 21115
rect -3725 21085 -3720 21115
rect -3760 21080 -3720 21085
rect -3680 21115 -3640 21120
rect -3680 21085 -3675 21115
rect -3645 21085 -3640 21115
rect -3680 21080 -3640 21085
rect -3600 21115 -3560 21120
rect -3600 21085 -3595 21115
rect -3565 21085 -3560 21115
rect -3600 21080 -3560 21085
rect -3520 21115 -3480 21120
rect -3520 21085 -3515 21115
rect -3485 21085 -3480 21115
rect -3520 21080 -3480 21085
rect -3440 21115 -3400 21120
rect -3440 21085 -3435 21115
rect -3405 21085 -3400 21115
rect -3440 21080 -3400 21085
rect -3360 21115 -3320 21120
rect -3360 21085 -3355 21115
rect -3325 21085 -3320 21115
rect -3360 21080 -3320 21085
rect -3280 21115 -3240 21120
rect -3280 21085 -3275 21115
rect -3245 21085 -3240 21115
rect -3280 21080 -3240 21085
rect -3200 21115 -3160 21120
rect -3200 21085 -3195 21115
rect -3165 21085 -3160 21115
rect -3200 21080 -3160 21085
rect -3120 21115 -3080 21120
rect -3120 21085 -3115 21115
rect -3085 21085 -3080 21115
rect -3120 21080 -3080 21085
rect -3040 21115 -3000 21120
rect -3040 21085 -3035 21115
rect -3005 21085 -3000 21115
rect -3040 21080 -3000 21085
rect -2960 21115 -2920 21120
rect -2960 21085 -2955 21115
rect -2925 21085 -2920 21115
rect -2960 21080 -2920 21085
rect -2880 21115 -2840 21120
rect -2880 21085 -2875 21115
rect -2845 21085 -2840 21115
rect -2880 21080 -2840 21085
rect -2800 21115 -2760 21120
rect -2800 21085 -2795 21115
rect -2765 21085 -2760 21115
rect -2800 21080 -2760 21085
rect -2720 21115 -2680 21120
rect -2720 21085 -2715 21115
rect -2685 21085 -2680 21115
rect -2720 21080 -2680 21085
rect -2640 21115 -2600 21120
rect -2640 21085 -2635 21115
rect -2605 21085 -2600 21115
rect -2640 21080 -2600 21085
rect -2560 21115 -2520 21120
rect -2560 21085 -2555 21115
rect -2525 21085 -2520 21115
rect -2560 21080 -2520 21085
rect -2480 21115 -2440 21120
rect -2480 21085 -2475 21115
rect -2445 21085 -2440 21115
rect -2480 21080 -2440 21085
rect -2400 21115 -2360 21120
rect -2400 21085 -2395 21115
rect -2365 21085 -2360 21115
rect -2400 21080 -2360 21085
rect -2320 21115 -2280 21120
rect -2320 21085 -2315 21115
rect -2285 21085 -2280 21115
rect -2320 21080 -2280 21085
rect -2240 21115 -2200 21120
rect -2240 21085 -2235 21115
rect -2205 21085 -2200 21115
rect -2240 21080 -2200 21085
rect -2160 21115 -2120 21120
rect -2160 21085 -2155 21115
rect -2125 21085 -2120 21115
rect -2160 21080 -2120 21085
rect -2080 21115 -2040 21120
rect -2080 21085 -2075 21115
rect -2045 21085 -2040 21115
rect -2080 21080 -2040 21085
rect -2000 21115 -1960 21120
rect -2000 21085 -1995 21115
rect -1965 21085 -1960 21115
rect -2000 21080 -1960 21085
rect -1840 21115 -1800 21120
rect -1840 21085 -1835 21115
rect -1805 21085 -1800 21115
rect -1840 21080 -1800 21085
rect -1760 21115 -1720 21120
rect -1760 21085 -1755 21115
rect -1725 21085 -1720 21115
rect -1760 21080 -1720 21085
rect -1680 21115 -1640 21120
rect -1680 21085 -1675 21115
rect -1645 21085 -1640 21115
rect -1680 21080 -1640 21085
rect -1520 21115 -1480 21120
rect -1520 21085 -1515 21115
rect -1485 21085 -1480 21115
rect -1520 21080 -1480 21085
rect -1360 21115 -1320 21120
rect -1360 21085 -1355 21115
rect -1325 21085 -1320 21115
rect -1360 21080 -1320 21085
rect -1280 21115 -1240 21120
rect -1280 21085 -1275 21115
rect -1245 21085 -1240 21115
rect -1280 21080 -1240 21085
rect -1200 21115 -1160 21120
rect -1200 21085 -1195 21115
rect -1165 21085 -1160 21115
rect -1200 21080 -1160 21085
rect -1120 21115 -1080 21120
rect -1120 21085 -1115 21115
rect -1085 21085 -1080 21115
rect -1120 21080 -1080 21085
rect -1040 21115 -1000 21120
rect -1040 21085 -1035 21115
rect -1005 21085 -1000 21115
rect -1040 21080 -1000 21085
rect -880 21115 -840 21120
rect -880 21085 -875 21115
rect -845 21085 -840 21115
rect -880 21080 -840 21085
rect -720 21115 -680 21120
rect -720 21085 -715 21115
rect -685 21085 -680 21115
rect -720 21080 -680 21085
rect -560 21115 -520 21120
rect -560 21085 -555 21115
rect -525 21085 -520 21115
rect -560 21080 -520 21085
rect -14960 20955 -14920 20960
rect -14960 20925 -14955 20955
rect -14925 20925 -14920 20955
rect -14960 20920 -14920 20925
rect -14880 20955 -14840 20960
rect -14880 20925 -14875 20955
rect -14845 20925 -14840 20955
rect -14880 20920 -14840 20925
rect -14800 20955 -14760 20960
rect -14800 20925 -14795 20955
rect -14765 20925 -14760 20955
rect -14800 20920 -14760 20925
rect -14720 20955 -14680 20960
rect -14720 20925 -14715 20955
rect -14685 20925 -14680 20955
rect -14720 20920 -14680 20925
rect -14640 20955 -14600 20960
rect -14640 20925 -14635 20955
rect -14605 20925 -14600 20955
rect -14640 20920 -14600 20925
rect -14560 20955 -14520 20960
rect -14560 20925 -14555 20955
rect -14525 20925 -14520 20955
rect -14560 20920 -14520 20925
rect -14480 20955 -14440 20960
rect -14480 20925 -14475 20955
rect -14445 20925 -14440 20955
rect -14480 20920 -14440 20925
rect -14400 20955 -14360 20960
rect -14400 20925 -14395 20955
rect -14365 20925 -14360 20955
rect -14400 20920 -14360 20925
rect -14320 20955 -14280 20960
rect -14320 20925 -14315 20955
rect -14285 20925 -14280 20955
rect -14320 20920 -14280 20925
rect -14240 20955 -14200 20960
rect -14240 20925 -14235 20955
rect -14205 20925 -14200 20955
rect -14240 20920 -14200 20925
rect -14160 20955 -14120 20960
rect -14160 20925 -14155 20955
rect -14125 20925 -14120 20955
rect -14160 20920 -14120 20925
rect -14080 20955 -14040 20960
rect -14080 20925 -14075 20955
rect -14045 20925 -14040 20955
rect -14080 20920 -14040 20925
rect -14000 20955 -13960 20960
rect -14000 20925 -13995 20955
rect -13965 20925 -13960 20955
rect -14000 20920 -13960 20925
rect -13920 20955 -13880 20960
rect -13920 20925 -13915 20955
rect -13885 20925 -13880 20955
rect -13920 20920 -13880 20925
rect -13840 20955 -13800 20960
rect -13840 20925 -13835 20955
rect -13805 20925 -13800 20955
rect -13840 20920 -13800 20925
rect -13760 20955 -13720 20960
rect -13760 20925 -13755 20955
rect -13725 20925 -13720 20955
rect -13760 20920 -13720 20925
rect -13680 20955 -13640 20960
rect -13680 20925 -13675 20955
rect -13645 20925 -13640 20955
rect -13680 20920 -13640 20925
rect -13600 20955 -13560 20960
rect -13600 20925 -13595 20955
rect -13565 20925 -13560 20955
rect -13600 20920 -13560 20925
rect -13520 20955 -13480 20960
rect -13520 20925 -13515 20955
rect -13485 20925 -13480 20955
rect -13520 20920 -13480 20925
rect -13440 20955 -13400 20960
rect -13440 20925 -13435 20955
rect -13405 20925 -13400 20955
rect -13440 20920 -13400 20925
rect -13360 20955 -13320 20960
rect -13360 20925 -13355 20955
rect -13325 20925 -13320 20955
rect -13360 20920 -13320 20925
rect -13280 20955 -13240 20960
rect -13280 20925 -13275 20955
rect -13245 20925 -13240 20955
rect -13280 20920 -13240 20925
rect -13200 20955 -13160 20960
rect -13200 20925 -13195 20955
rect -13165 20925 -13160 20955
rect -13200 20920 -13160 20925
rect -13120 20955 -13080 20960
rect -13120 20925 -13115 20955
rect -13085 20925 -13080 20955
rect -13120 20920 -13080 20925
rect -13040 20955 -13000 20960
rect -13040 20925 -13035 20955
rect -13005 20925 -13000 20955
rect -13040 20920 -13000 20925
rect -12960 20955 -12920 20960
rect -12960 20925 -12955 20955
rect -12925 20925 -12920 20955
rect -12960 20920 -12920 20925
rect -12880 20955 -12840 20960
rect -12880 20925 -12875 20955
rect -12845 20925 -12840 20955
rect -12880 20920 -12840 20925
rect -12800 20955 -12760 20960
rect -12800 20925 -12795 20955
rect -12765 20925 -12760 20955
rect -12800 20920 -12760 20925
rect -12720 20955 -12680 20960
rect -12720 20925 -12715 20955
rect -12685 20925 -12680 20955
rect -12720 20920 -12680 20925
rect -12640 20955 -12600 20960
rect -12640 20925 -12635 20955
rect -12605 20925 -12600 20955
rect -12640 20920 -12600 20925
rect -12560 20955 -12520 20960
rect -12560 20925 -12555 20955
rect -12525 20925 -12520 20955
rect -12560 20920 -12520 20925
rect -12480 20955 -12440 20960
rect -12480 20925 -12475 20955
rect -12445 20925 -12440 20955
rect -12480 20920 -12440 20925
rect -12400 20955 -12360 20960
rect -12400 20925 -12395 20955
rect -12365 20925 -12360 20955
rect -12400 20920 -12360 20925
rect -12320 20955 -12280 20960
rect -12320 20925 -12315 20955
rect -12285 20925 -12280 20955
rect -12320 20920 -12280 20925
rect -12240 20955 -12200 20960
rect -12240 20925 -12235 20955
rect -12205 20925 -12200 20955
rect -12240 20920 -12200 20925
rect -12160 20955 -12120 20960
rect -12160 20925 -12155 20955
rect -12125 20925 -12120 20955
rect -12160 20920 -12120 20925
rect -12080 20955 -12040 20960
rect -12080 20925 -12075 20955
rect -12045 20925 -12040 20955
rect -12080 20920 -12040 20925
rect -12000 20955 -11960 20960
rect -12000 20925 -11995 20955
rect -11965 20925 -11960 20955
rect -12000 20920 -11960 20925
rect -11920 20955 -11880 20960
rect -11920 20925 -11915 20955
rect -11885 20925 -11880 20955
rect -11920 20920 -11880 20925
rect -11840 20955 -11800 20960
rect -11840 20925 -11835 20955
rect -11805 20925 -11800 20955
rect -11840 20920 -11800 20925
rect -11760 20955 -11720 20960
rect -11760 20925 -11755 20955
rect -11725 20925 -11720 20955
rect -11760 20920 -11720 20925
rect -11680 20955 -11640 20960
rect -11680 20925 -11675 20955
rect -11645 20925 -11640 20955
rect -11680 20920 -11640 20925
rect -11600 20955 -11560 20960
rect -11600 20925 -11595 20955
rect -11565 20925 -11560 20955
rect -11600 20920 -11560 20925
rect -11520 20955 -11480 20960
rect -11520 20925 -11515 20955
rect -11485 20925 -11480 20955
rect -11520 20920 -11480 20925
rect -11440 20955 -11400 20960
rect -11440 20925 -11435 20955
rect -11405 20925 -11400 20955
rect -11440 20920 -11400 20925
rect -11360 20955 -11320 20960
rect -11360 20925 -11355 20955
rect -11325 20925 -11320 20955
rect -11360 20920 -11320 20925
rect -11280 20955 -11240 20960
rect -11280 20925 -11275 20955
rect -11245 20925 -11240 20955
rect -11280 20920 -11240 20925
rect -11200 20955 -11160 20960
rect -11200 20925 -11195 20955
rect -11165 20925 -11160 20955
rect -11200 20920 -11160 20925
rect -11120 20955 -11080 20960
rect -11120 20925 -11115 20955
rect -11085 20925 -11080 20955
rect -11120 20920 -11080 20925
rect -11040 20955 -11000 20960
rect -11040 20925 -11035 20955
rect -11005 20925 -11000 20955
rect -11040 20920 -11000 20925
rect -10960 20955 -10920 20960
rect -10960 20925 -10955 20955
rect -10925 20925 -10920 20955
rect -10960 20920 -10920 20925
rect -10880 20955 -10840 20960
rect -10880 20925 -10875 20955
rect -10845 20925 -10840 20955
rect -10880 20920 -10840 20925
rect -10800 20955 -10760 20960
rect -10800 20925 -10795 20955
rect -10765 20925 -10760 20955
rect -10800 20920 -10760 20925
rect -10720 20955 -10680 20960
rect -10720 20925 -10715 20955
rect -10685 20925 -10680 20955
rect -10720 20920 -10680 20925
rect -10640 20955 -10600 20960
rect -10640 20925 -10635 20955
rect -10605 20925 -10600 20955
rect -10640 20920 -10600 20925
rect -10560 20955 -10520 20960
rect -10560 20925 -10555 20955
rect -10525 20925 -10520 20955
rect -10560 20920 -10520 20925
rect -10480 20955 -10440 20960
rect -10480 20925 -10475 20955
rect -10445 20925 -10440 20955
rect -10480 20920 -10440 20925
rect -10400 20955 -10360 20960
rect -10400 20925 -10395 20955
rect -10365 20925 -10360 20955
rect -10400 20920 -10360 20925
rect -10320 20955 -10280 20960
rect -10320 20925 -10315 20955
rect -10285 20925 -10280 20955
rect -10320 20920 -10280 20925
rect -10240 20955 -10200 20960
rect -10240 20925 -10235 20955
rect -10205 20925 -10200 20955
rect -10240 20920 -10200 20925
rect -10160 20955 -10120 20960
rect -10160 20925 -10155 20955
rect -10125 20925 -10120 20955
rect -10160 20920 -10120 20925
rect -10080 20955 -10040 20960
rect -10080 20925 -10075 20955
rect -10045 20925 -10040 20955
rect -10080 20920 -10040 20925
rect -10000 20955 -9960 20960
rect -10000 20925 -9995 20955
rect -9965 20925 -9960 20955
rect -10000 20920 -9960 20925
rect -9920 20955 -9880 20960
rect -9920 20925 -9915 20955
rect -9885 20925 -9880 20955
rect -9920 20920 -9880 20925
rect -9840 20955 -9800 20960
rect -9840 20925 -9835 20955
rect -9805 20925 -9800 20955
rect -9840 20920 -9800 20925
rect -9760 20955 -9720 20960
rect -9760 20925 -9755 20955
rect -9725 20925 -9720 20955
rect -9760 20920 -9720 20925
rect -9680 20955 -9640 20960
rect -9680 20925 -9675 20955
rect -9645 20925 -9640 20955
rect -9680 20920 -9640 20925
rect -9600 20955 -9560 20960
rect -9600 20925 -9595 20955
rect -9565 20925 -9560 20955
rect -9600 20920 -9560 20925
rect -9520 20955 -9480 20960
rect -9520 20925 -9515 20955
rect -9485 20925 -9480 20955
rect -9520 20920 -9480 20925
rect -9440 20955 -9400 20960
rect -9440 20925 -9435 20955
rect -9405 20925 -9400 20955
rect -9440 20920 -9400 20925
rect -9360 20955 -9320 20960
rect -9360 20925 -9355 20955
rect -9325 20925 -9320 20955
rect -9360 20920 -9320 20925
rect -9280 20955 -9240 20960
rect -9280 20925 -9275 20955
rect -9245 20925 -9240 20955
rect -9280 20920 -9240 20925
rect -9200 20955 -9160 20960
rect -9200 20925 -9195 20955
rect -9165 20925 -9160 20955
rect -9200 20920 -9160 20925
rect -9120 20955 -9080 20960
rect -9120 20925 -9115 20955
rect -9085 20925 -9080 20955
rect -9120 20920 -9080 20925
rect -9040 20955 -9000 20960
rect -9040 20925 -9035 20955
rect -9005 20925 -9000 20955
rect -9040 20920 -9000 20925
rect -8960 20955 -8920 20960
rect -8960 20925 -8955 20955
rect -8925 20925 -8920 20955
rect -8960 20920 -8920 20925
rect -8880 20955 -8840 20960
rect -8880 20925 -8875 20955
rect -8845 20925 -8840 20955
rect -8880 20920 -8840 20925
rect -8800 20955 -8760 20960
rect -8800 20925 -8795 20955
rect -8765 20925 -8760 20955
rect -8800 20920 -8760 20925
rect -8720 20955 -8680 20960
rect -8720 20925 -8715 20955
rect -8685 20925 -8680 20955
rect -8720 20920 -8680 20925
rect -8640 20955 -8600 20960
rect -8640 20925 -8635 20955
rect -8605 20925 -8600 20955
rect -8640 20920 -8600 20925
rect -8560 20955 -8520 20960
rect -8560 20925 -8555 20955
rect -8525 20925 -8520 20955
rect -8560 20920 -8520 20925
rect -8480 20955 -8440 20960
rect -8480 20925 -8475 20955
rect -8445 20925 -8440 20955
rect -8480 20920 -8440 20925
rect -8400 20955 -8360 20960
rect -8400 20925 -8395 20955
rect -8365 20925 -8360 20955
rect -8400 20920 -8360 20925
rect -8320 20955 -8280 20960
rect -8320 20925 -8315 20955
rect -8285 20925 -8280 20955
rect -8320 20920 -8280 20925
rect -8240 20955 -8200 20960
rect -8240 20925 -8235 20955
rect -8205 20925 -8200 20955
rect -8240 20920 -8200 20925
rect -8160 20955 -8120 20960
rect -8160 20925 -8155 20955
rect -8125 20925 -8120 20955
rect -8160 20920 -8120 20925
rect -8080 20955 -8040 20960
rect -8080 20925 -8075 20955
rect -8045 20925 -8040 20955
rect -8080 20920 -8040 20925
rect -8000 20955 -7960 20960
rect -8000 20925 -7995 20955
rect -7965 20925 -7960 20955
rect -8000 20920 -7960 20925
rect -7920 20955 -7880 20960
rect -7920 20925 -7915 20955
rect -7885 20925 -7880 20955
rect -7920 20920 -7880 20925
rect -7840 20955 -7800 20960
rect -7840 20925 -7835 20955
rect -7805 20925 -7800 20955
rect -7840 20920 -7800 20925
rect -7760 20955 -7720 20960
rect -7760 20925 -7755 20955
rect -7725 20925 -7720 20955
rect -7760 20920 -7720 20925
rect -7680 20955 -7640 20960
rect -7680 20925 -7675 20955
rect -7645 20925 -7640 20955
rect -7680 20920 -7640 20925
rect -7600 20955 -7560 20960
rect -7600 20925 -7595 20955
rect -7565 20925 -7560 20955
rect -7600 20920 -7560 20925
rect -7520 20955 -7480 20960
rect -7520 20925 -7515 20955
rect -7485 20925 -7480 20955
rect -7520 20920 -7480 20925
rect -7440 20955 -7400 20960
rect -7440 20925 -7435 20955
rect -7405 20925 -7400 20955
rect -7440 20920 -7400 20925
rect -7360 20955 -7320 20960
rect -7360 20925 -7355 20955
rect -7325 20925 -7320 20955
rect -7360 20920 -7320 20925
rect -7280 20955 -7240 20960
rect -7280 20925 -7275 20955
rect -7245 20925 -7240 20955
rect -7280 20920 -7240 20925
rect -7200 20955 -7160 20960
rect -7200 20925 -7195 20955
rect -7165 20925 -7160 20955
rect -7200 20920 -7160 20925
rect -7120 20955 -7080 20960
rect -7120 20925 -7115 20955
rect -7085 20925 -7080 20955
rect -7120 20920 -7080 20925
rect -7040 20955 -7000 20960
rect -7040 20925 -7035 20955
rect -7005 20925 -7000 20955
rect -7040 20920 -7000 20925
rect -6960 20955 -6920 20960
rect -6960 20925 -6955 20955
rect -6925 20925 -6920 20955
rect -6960 20920 -6920 20925
rect -6880 20955 -6840 20960
rect -6880 20925 -6875 20955
rect -6845 20925 -6840 20955
rect -6880 20920 -6840 20925
rect -6800 20955 -6760 20960
rect -6800 20925 -6795 20955
rect -6765 20925 -6760 20955
rect -6800 20920 -6760 20925
rect -6720 20955 -6680 20960
rect -6720 20925 -6715 20955
rect -6685 20925 -6680 20955
rect -6720 20920 -6680 20925
rect -6640 20955 -6600 20960
rect -6640 20925 -6635 20955
rect -6605 20925 -6600 20955
rect -6640 20920 -6600 20925
rect -6560 20955 -6520 20960
rect -6560 20925 -6555 20955
rect -6525 20925 -6520 20955
rect -6560 20920 -6520 20925
rect -6480 20955 -6440 20960
rect -6480 20925 -6475 20955
rect -6445 20925 -6440 20955
rect -6480 20920 -6440 20925
rect -6400 20955 -6360 20960
rect -6400 20925 -6395 20955
rect -6365 20925 -6360 20955
rect -6400 20920 -6360 20925
rect -6320 20955 -6280 20960
rect -6320 20925 -6315 20955
rect -6285 20925 -6280 20955
rect -6320 20920 -6280 20925
rect -6240 20955 -6200 20960
rect -6240 20925 -6235 20955
rect -6205 20925 -6200 20955
rect -6240 20920 -6200 20925
rect -6160 20955 -6120 20960
rect -6160 20925 -6155 20955
rect -6125 20925 -6120 20955
rect -6160 20920 -6120 20925
rect -5680 20955 -5640 20960
rect -5680 20925 -5675 20955
rect -5645 20925 -5640 20955
rect -5680 20920 -5640 20925
rect -5600 20955 -5560 20960
rect -5600 20925 -5595 20955
rect -5565 20925 -5560 20955
rect -5600 20920 -5560 20925
rect -5520 20955 -5480 20960
rect -5520 20925 -5515 20955
rect -5485 20925 -5480 20955
rect -5520 20920 -5480 20925
rect -5440 20955 -5400 20960
rect -5440 20925 -5435 20955
rect -5405 20925 -5400 20955
rect -5440 20920 -5400 20925
rect -5360 20955 -5320 20960
rect -5360 20925 -5355 20955
rect -5325 20925 -5320 20955
rect -5360 20920 -5320 20925
rect -5280 20955 -5240 20960
rect -5280 20925 -5275 20955
rect -5245 20925 -5240 20955
rect -5280 20920 -5240 20925
rect -5200 20955 -5160 20960
rect -5200 20925 -5195 20955
rect -5165 20925 -5160 20955
rect -5200 20920 -5160 20925
rect -5120 20955 -5080 20960
rect -5120 20925 -5115 20955
rect -5085 20925 -5080 20955
rect -5120 20920 -5080 20925
rect -5040 20955 -5000 20960
rect -5040 20925 -5035 20955
rect -5005 20925 -5000 20955
rect -5040 20920 -5000 20925
rect -4960 20955 -4920 20960
rect -4960 20925 -4955 20955
rect -4925 20925 -4920 20955
rect -4960 20920 -4920 20925
rect -4880 20955 -4840 20960
rect -4880 20925 -4875 20955
rect -4845 20925 -4840 20955
rect -4880 20920 -4840 20925
rect -4800 20955 -4760 20960
rect -4800 20925 -4795 20955
rect -4765 20925 -4760 20955
rect -4800 20920 -4760 20925
rect -4720 20955 -4680 20960
rect -4720 20925 -4715 20955
rect -4685 20925 -4680 20955
rect -4720 20920 -4680 20925
rect -4640 20955 -4600 20960
rect -4640 20925 -4635 20955
rect -4605 20925 -4600 20955
rect -4640 20920 -4600 20925
rect -4560 20955 -4520 20960
rect -4560 20925 -4555 20955
rect -4525 20925 -4520 20955
rect -4560 20920 -4520 20925
rect -4480 20955 -4440 20960
rect -4480 20925 -4475 20955
rect -4445 20925 -4440 20955
rect -4480 20920 -4440 20925
rect -4400 20955 -4360 20960
rect -4400 20925 -4395 20955
rect -4365 20925 -4360 20955
rect -4400 20920 -4360 20925
rect -4320 20955 -4280 20960
rect -4320 20925 -4315 20955
rect -4285 20925 -4280 20955
rect -4320 20920 -4280 20925
rect -4240 20955 -4200 20960
rect -4240 20925 -4235 20955
rect -4205 20925 -4200 20955
rect -4240 20920 -4200 20925
rect -4160 20955 -4120 20960
rect -4160 20925 -4155 20955
rect -4125 20925 -4120 20955
rect -4160 20920 -4120 20925
rect -4080 20955 -4040 20960
rect -4080 20925 -4075 20955
rect -4045 20925 -4040 20955
rect -4080 20920 -4040 20925
rect -4000 20955 -3960 20960
rect -4000 20925 -3995 20955
rect -3965 20925 -3960 20955
rect -4000 20920 -3960 20925
rect -3920 20955 -3880 20960
rect -3920 20925 -3915 20955
rect -3885 20925 -3880 20955
rect -3920 20920 -3880 20925
rect -3840 20955 -3800 20960
rect -3840 20925 -3835 20955
rect -3805 20925 -3800 20955
rect -3840 20920 -3800 20925
rect -3760 20955 -3720 20960
rect -3760 20925 -3755 20955
rect -3725 20925 -3720 20955
rect -3760 20920 -3720 20925
rect -3680 20955 -3640 20960
rect -3680 20925 -3675 20955
rect -3645 20925 -3640 20955
rect -3680 20920 -3640 20925
rect -3600 20955 -3560 20960
rect -3600 20925 -3595 20955
rect -3565 20925 -3560 20955
rect -3600 20920 -3560 20925
rect -3520 20955 -3480 20960
rect -3520 20925 -3515 20955
rect -3485 20925 -3480 20955
rect -3520 20920 -3480 20925
rect -3440 20955 -3400 20960
rect -3440 20925 -3435 20955
rect -3405 20925 -3400 20955
rect -3440 20920 -3400 20925
rect -3360 20955 -3320 20960
rect -3360 20925 -3355 20955
rect -3325 20925 -3320 20955
rect -3360 20920 -3320 20925
rect -3280 20955 -3240 20960
rect -3280 20925 -3275 20955
rect -3245 20925 -3240 20955
rect -3280 20920 -3240 20925
rect -3200 20955 -3160 20960
rect -3200 20925 -3195 20955
rect -3165 20925 -3160 20955
rect -3200 20920 -3160 20925
rect -3120 20955 -3080 20960
rect -3120 20925 -3115 20955
rect -3085 20925 -3080 20955
rect -3120 20920 -3080 20925
rect -3040 20955 -3000 20960
rect -3040 20925 -3035 20955
rect -3005 20925 -3000 20955
rect -3040 20920 -3000 20925
rect -2960 20955 -2920 20960
rect -2960 20925 -2955 20955
rect -2925 20925 -2920 20955
rect -2960 20920 -2920 20925
rect -2880 20955 -2840 20960
rect -2880 20925 -2875 20955
rect -2845 20925 -2840 20955
rect -2880 20920 -2840 20925
rect -2800 20955 -2760 20960
rect -2800 20925 -2795 20955
rect -2765 20925 -2760 20955
rect -2800 20920 -2760 20925
rect -2720 20955 -2680 20960
rect -2720 20925 -2715 20955
rect -2685 20925 -2680 20955
rect -2720 20920 -2680 20925
rect -2640 20955 -2600 20960
rect -2640 20925 -2635 20955
rect -2605 20925 -2600 20955
rect -2640 20920 -2600 20925
rect -2560 20955 -2520 20960
rect -2560 20925 -2555 20955
rect -2525 20925 -2520 20955
rect -2560 20920 -2520 20925
rect -2480 20955 -2440 20960
rect -2480 20925 -2475 20955
rect -2445 20925 -2440 20955
rect -2480 20920 -2440 20925
rect -2400 20955 -2360 20960
rect -2400 20925 -2395 20955
rect -2365 20925 -2360 20955
rect -2400 20920 -2360 20925
rect -2320 20955 -2280 20960
rect -2320 20925 -2315 20955
rect -2285 20925 -2280 20955
rect -2320 20920 -2280 20925
rect -2240 20955 -2200 20960
rect -2240 20925 -2235 20955
rect -2205 20925 -2200 20955
rect -2240 20920 -2200 20925
rect -2160 20955 -2120 20960
rect -2160 20925 -2155 20955
rect -2125 20925 -2120 20955
rect -2160 20920 -2120 20925
rect -2080 20955 -2040 20960
rect -2080 20925 -2075 20955
rect -2045 20925 -2040 20955
rect -2080 20920 -2040 20925
rect -2000 20955 -1960 20960
rect -2000 20925 -1995 20955
rect -1965 20925 -1960 20955
rect -2000 20920 -1960 20925
rect -1840 20955 -1800 20960
rect -1840 20925 -1835 20955
rect -1805 20925 -1800 20955
rect -1840 20920 -1800 20925
rect -1760 20955 -1720 20960
rect -1760 20925 -1755 20955
rect -1725 20925 -1720 20955
rect -1760 20920 -1720 20925
rect -1680 20955 -1640 20960
rect -1680 20925 -1675 20955
rect -1645 20925 -1640 20955
rect -1680 20920 -1640 20925
rect -1520 20955 -1480 20960
rect -1520 20925 -1515 20955
rect -1485 20925 -1480 20955
rect -1520 20920 -1480 20925
rect -1360 20955 -1320 20960
rect -1360 20925 -1355 20955
rect -1325 20925 -1320 20955
rect -1360 20920 -1320 20925
rect -1280 20955 -1240 20960
rect -1280 20925 -1275 20955
rect -1245 20925 -1240 20955
rect -1280 20920 -1240 20925
rect -1200 20955 -1160 20960
rect -1200 20925 -1195 20955
rect -1165 20925 -1160 20955
rect -1200 20920 -1160 20925
rect -1120 20955 -1080 20960
rect -1120 20925 -1115 20955
rect -1085 20925 -1080 20955
rect -1120 20920 -1080 20925
rect -1040 20955 -1000 20960
rect -1040 20925 -1035 20955
rect -1005 20925 -1000 20955
rect -1040 20920 -1000 20925
rect -880 20955 -840 20960
rect -880 20925 -875 20955
rect -845 20925 -840 20955
rect -880 20920 -840 20925
rect -720 20955 -680 20960
rect -720 20925 -715 20955
rect -685 20925 -680 20955
rect -720 20920 -680 20925
rect -560 20955 -520 20960
rect -560 20925 -555 20955
rect -525 20925 -520 20955
rect -560 20920 -520 20925
rect -16560 20675 -16520 20680
rect -16560 20645 -16555 20675
rect -16525 20645 -16520 20675
rect -16560 20640 -16520 20645
rect -16480 20675 -16440 20680
rect -16480 20645 -16475 20675
rect -16445 20645 -16440 20675
rect -16480 20640 -16440 20645
rect -16400 20675 -16360 20680
rect -16400 20645 -16395 20675
rect -16365 20645 -16360 20675
rect -16400 20640 -16360 20645
rect -16320 20675 -16280 20680
rect -16320 20645 -16315 20675
rect -16285 20645 -16280 20675
rect -16320 20640 -16280 20645
rect -16240 20675 -16200 20680
rect -16240 20645 -16235 20675
rect -16205 20645 -16200 20675
rect -16240 20640 -16200 20645
rect -16160 20675 -16120 20680
rect -16160 20645 -16155 20675
rect -16125 20645 -16120 20675
rect -16160 20640 -16120 20645
rect -16080 20675 -16040 20680
rect -16080 20645 -16075 20675
rect -16045 20645 -16040 20675
rect -16080 20640 -16040 20645
rect -16000 20675 -15960 20680
rect -16000 20645 -15995 20675
rect -15965 20645 -15960 20675
rect -16000 20640 -15960 20645
rect -15920 20675 -15880 20680
rect -15920 20645 -15915 20675
rect -15885 20645 -15880 20675
rect -15920 20640 -15880 20645
rect -15840 20675 -15800 20680
rect -15840 20645 -15835 20675
rect -15805 20645 -15800 20675
rect -15840 20640 -15800 20645
rect -15760 20675 -15720 20680
rect -15760 20645 -15755 20675
rect -15725 20645 -15720 20675
rect -15760 20640 -15720 20645
rect -15680 20675 -15640 20680
rect -15680 20645 -15675 20675
rect -15645 20645 -15640 20675
rect -15680 20640 -15640 20645
rect -15600 20675 -15560 20680
rect -15600 20645 -15595 20675
rect -15565 20645 -15560 20675
rect -15600 20640 -15560 20645
rect -14960 20675 -14920 20680
rect -14960 20645 -14955 20675
rect -14925 20645 -14920 20675
rect -14960 20640 -14920 20645
rect -14880 20675 -14840 20680
rect -14880 20645 -14875 20675
rect -14845 20645 -14840 20675
rect -14880 20640 -14840 20645
rect -14800 20675 -14760 20680
rect -14800 20645 -14795 20675
rect -14765 20645 -14760 20675
rect -14800 20640 -14760 20645
rect -14720 20675 -14680 20680
rect -14720 20645 -14715 20675
rect -14685 20645 -14680 20675
rect -14720 20640 -14680 20645
rect -14640 20675 -14600 20680
rect -14640 20645 -14635 20675
rect -14605 20645 -14600 20675
rect -14640 20640 -14600 20645
rect -14560 20675 -14520 20680
rect -14560 20645 -14555 20675
rect -14525 20645 -14520 20675
rect -14560 20640 -14520 20645
rect -14480 20675 -14440 20680
rect -14480 20645 -14475 20675
rect -14445 20645 -14440 20675
rect -14480 20640 -14440 20645
rect -14400 20675 -14360 20680
rect -14400 20645 -14395 20675
rect -14365 20645 -14360 20675
rect -14400 20640 -14360 20645
rect -14320 20675 -14280 20680
rect -14320 20645 -14315 20675
rect -14285 20645 -14280 20675
rect -14320 20640 -14280 20645
rect -14240 20675 -14200 20680
rect -14240 20645 -14235 20675
rect -14205 20645 -14200 20675
rect -14240 20640 -14200 20645
rect -14160 20675 -14120 20680
rect -14160 20645 -14155 20675
rect -14125 20645 -14120 20675
rect -14160 20640 -14120 20645
rect -14080 20675 -14040 20680
rect -14080 20645 -14075 20675
rect -14045 20645 -14040 20675
rect -14080 20640 -14040 20645
rect -14000 20675 -13960 20680
rect -14000 20645 -13995 20675
rect -13965 20645 -13960 20675
rect -14000 20640 -13960 20645
rect -13920 20675 -13880 20680
rect -13920 20645 -13915 20675
rect -13885 20645 -13880 20675
rect -13920 20640 -13880 20645
rect -13840 20675 -13800 20680
rect -13840 20645 -13835 20675
rect -13805 20645 -13800 20675
rect -13840 20640 -13800 20645
rect -13760 20675 -13720 20680
rect -13760 20645 -13755 20675
rect -13725 20645 -13720 20675
rect -13760 20640 -13720 20645
rect -13680 20675 -13640 20680
rect -13680 20645 -13675 20675
rect -13645 20645 -13640 20675
rect -13680 20640 -13640 20645
rect -13600 20675 -13560 20680
rect -13600 20645 -13595 20675
rect -13565 20645 -13560 20675
rect -13600 20640 -13560 20645
rect -13520 20675 -13480 20680
rect -13520 20645 -13515 20675
rect -13485 20645 -13480 20675
rect -13520 20640 -13480 20645
rect -13440 20675 -13400 20680
rect -13440 20645 -13435 20675
rect -13405 20645 -13400 20675
rect -13440 20640 -13400 20645
rect -13360 20675 -13320 20680
rect -13360 20645 -13355 20675
rect -13325 20645 -13320 20675
rect -13360 20640 -13320 20645
rect -13280 20675 -13240 20680
rect -13280 20645 -13275 20675
rect -13245 20645 -13240 20675
rect -13280 20640 -13240 20645
rect -13200 20675 -13160 20680
rect -13200 20645 -13195 20675
rect -13165 20645 -13160 20675
rect -13200 20640 -13160 20645
rect -13120 20675 -13080 20680
rect -13120 20645 -13115 20675
rect -13085 20645 -13080 20675
rect -13120 20640 -13080 20645
rect -13040 20675 -13000 20680
rect -13040 20645 -13035 20675
rect -13005 20645 -13000 20675
rect -13040 20640 -13000 20645
rect -12960 20675 -12920 20680
rect -12960 20645 -12955 20675
rect -12925 20645 -12920 20675
rect -12960 20640 -12920 20645
rect -12880 20675 -12840 20680
rect -12880 20645 -12875 20675
rect -12845 20645 -12840 20675
rect -12880 20640 -12840 20645
rect -12800 20675 -12760 20680
rect -12800 20645 -12795 20675
rect -12765 20645 -12760 20675
rect -12800 20640 -12760 20645
rect -12720 20675 -12680 20680
rect -12720 20645 -12715 20675
rect -12685 20645 -12680 20675
rect -12720 20640 -12680 20645
rect -12640 20675 -12600 20680
rect -12640 20645 -12635 20675
rect -12605 20645 -12600 20675
rect -12640 20640 -12600 20645
rect -12560 20675 -12520 20680
rect -12560 20645 -12555 20675
rect -12525 20645 -12520 20675
rect -12560 20640 -12520 20645
rect -12480 20675 -12440 20680
rect -12480 20645 -12475 20675
rect -12445 20645 -12440 20675
rect -12480 20640 -12440 20645
rect -12400 20675 -12360 20680
rect -12400 20645 -12395 20675
rect -12365 20645 -12360 20675
rect -12400 20640 -12360 20645
rect -12320 20675 -12280 20680
rect -12320 20645 -12315 20675
rect -12285 20645 -12280 20675
rect -12320 20640 -12280 20645
rect -12240 20675 -12200 20680
rect -12240 20645 -12235 20675
rect -12205 20645 -12200 20675
rect -12240 20640 -12200 20645
rect -12160 20675 -12120 20680
rect -12160 20645 -12155 20675
rect -12125 20645 -12120 20675
rect -12160 20640 -12120 20645
rect -12080 20675 -12040 20680
rect -12080 20645 -12075 20675
rect -12045 20645 -12040 20675
rect -12080 20640 -12040 20645
rect -12000 20675 -11960 20680
rect -12000 20645 -11995 20675
rect -11965 20645 -11960 20675
rect -12000 20640 -11960 20645
rect -11920 20675 -11880 20680
rect -11920 20645 -11915 20675
rect -11885 20645 -11880 20675
rect -11920 20640 -11880 20645
rect -11840 20675 -11800 20680
rect -11840 20645 -11835 20675
rect -11805 20645 -11800 20675
rect -11840 20640 -11800 20645
rect -11760 20675 -11720 20680
rect -11760 20645 -11755 20675
rect -11725 20645 -11720 20675
rect -11760 20640 -11720 20645
rect -11680 20675 -11640 20680
rect -11680 20645 -11675 20675
rect -11645 20645 -11640 20675
rect -11680 20640 -11640 20645
rect -11600 20675 -11560 20680
rect -11600 20645 -11595 20675
rect -11565 20645 -11560 20675
rect -11600 20640 -11560 20645
rect -11520 20675 -11480 20680
rect -11520 20645 -11515 20675
rect -11485 20645 -11480 20675
rect -11520 20640 -11480 20645
rect -11440 20675 -11400 20680
rect -11440 20645 -11435 20675
rect -11405 20645 -11400 20675
rect -11440 20640 -11400 20645
rect -11360 20675 -11320 20680
rect -11360 20645 -11355 20675
rect -11325 20645 -11320 20675
rect -11360 20640 -11320 20645
rect -11280 20675 -11240 20680
rect -11280 20645 -11275 20675
rect -11245 20645 -11240 20675
rect -11280 20640 -11240 20645
rect -11200 20675 -11160 20680
rect -11200 20645 -11195 20675
rect -11165 20645 -11160 20675
rect -11200 20640 -11160 20645
rect -11120 20675 -11080 20680
rect -11120 20645 -11115 20675
rect -11085 20645 -11080 20675
rect -11120 20640 -11080 20645
rect -11040 20675 -11000 20680
rect -11040 20645 -11035 20675
rect -11005 20645 -11000 20675
rect -11040 20640 -11000 20645
rect -10960 20675 -10920 20680
rect -10960 20645 -10955 20675
rect -10925 20645 -10920 20675
rect -10960 20640 -10920 20645
rect -10880 20675 -10840 20680
rect -10880 20645 -10875 20675
rect -10845 20645 -10840 20675
rect -10880 20640 -10840 20645
rect -10800 20675 -10760 20680
rect -10800 20645 -10795 20675
rect -10765 20645 -10760 20675
rect -10800 20640 -10760 20645
rect -10720 20675 -10680 20680
rect -10720 20645 -10715 20675
rect -10685 20645 -10680 20675
rect -10720 20640 -10680 20645
rect -10640 20675 -10600 20680
rect -10640 20645 -10635 20675
rect -10605 20645 -10600 20675
rect -10640 20640 -10600 20645
rect -10560 20675 -10520 20680
rect -10560 20645 -10555 20675
rect -10525 20645 -10520 20675
rect -10560 20640 -10520 20645
rect -10480 20675 -10440 20680
rect -10480 20645 -10475 20675
rect -10445 20645 -10440 20675
rect -10480 20640 -10440 20645
rect -10400 20675 -10360 20680
rect -10400 20645 -10395 20675
rect -10365 20645 -10360 20675
rect -10400 20640 -10360 20645
rect -10320 20675 -10280 20680
rect -10320 20645 -10315 20675
rect -10285 20645 -10280 20675
rect -10320 20640 -10280 20645
rect -10240 20675 -10200 20680
rect -10240 20645 -10235 20675
rect -10205 20645 -10200 20675
rect -10240 20640 -10200 20645
rect -10160 20675 -10120 20680
rect -10160 20645 -10155 20675
rect -10125 20645 -10120 20675
rect -10160 20640 -10120 20645
rect -10080 20675 -10040 20680
rect -10080 20645 -10075 20675
rect -10045 20645 -10040 20675
rect -10080 20640 -10040 20645
rect -10000 20675 -9960 20680
rect -10000 20645 -9995 20675
rect -9965 20645 -9960 20675
rect -10000 20640 -9960 20645
rect -9920 20675 -9880 20680
rect -9920 20645 -9915 20675
rect -9885 20645 -9880 20675
rect -9920 20640 -9880 20645
rect -9840 20675 -9800 20680
rect -9840 20645 -9835 20675
rect -9805 20645 -9800 20675
rect -9840 20640 -9800 20645
rect -9760 20675 -9720 20680
rect -9760 20645 -9755 20675
rect -9725 20645 -9720 20675
rect -9760 20640 -9720 20645
rect -9680 20675 -9640 20680
rect -9680 20645 -9675 20675
rect -9645 20645 -9640 20675
rect -9680 20640 -9640 20645
rect -9600 20675 -9560 20680
rect -9600 20645 -9595 20675
rect -9565 20645 -9560 20675
rect -9600 20640 -9560 20645
rect -9520 20675 -9480 20680
rect -9520 20645 -9515 20675
rect -9485 20645 -9480 20675
rect -9520 20640 -9480 20645
rect -9440 20675 -9400 20680
rect -9440 20645 -9435 20675
rect -9405 20645 -9400 20675
rect -9440 20640 -9400 20645
rect -9360 20675 -9320 20680
rect -9360 20645 -9355 20675
rect -9325 20645 -9320 20675
rect -9360 20640 -9320 20645
rect -9280 20675 -9240 20680
rect -9280 20645 -9275 20675
rect -9245 20645 -9240 20675
rect -9280 20640 -9240 20645
rect -9200 20675 -9160 20680
rect -9200 20645 -9195 20675
rect -9165 20645 -9160 20675
rect -9200 20640 -9160 20645
rect -9120 20675 -9080 20680
rect -9120 20645 -9115 20675
rect -9085 20645 -9080 20675
rect -9120 20640 -9080 20645
rect -9040 20675 -9000 20680
rect -9040 20645 -9035 20675
rect -9005 20645 -9000 20675
rect -9040 20640 -9000 20645
rect -8960 20675 -8920 20680
rect -8960 20645 -8955 20675
rect -8925 20645 -8920 20675
rect -8960 20640 -8920 20645
rect -8880 20675 -8840 20680
rect -8880 20645 -8875 20675
rect -8845 20645 -8840 20675
rect -8880 20640 -8840 20645
rect -8800 20675 -8760 20680
rect -8800 20645 -8795 20675
rect -8765 20645 -8760 20675
rect -8800 20640 -8760 20645
rect -8720 20675 -8680 20680
rect -8720 20645 -8715 20675
rect -8685 20645 -8680 20675
rect -8720 20640 -8680 20645
rect -8640 20675 -8600 20680
rect -8640 20645 -8635 20675
rect -8605 20645 -8600 20675
rect -8640 20640 -8600 20645
rect -8560 20675 -8520 20680
rect -8560 20645 -8555 20675
rect -8525 20645 -8520 20675
rect -8560 20640 -8520 20645
rect -8480 20675 -8440 20680
rect -8480 20645 -8475 20675
rect -8445 20645 -8440 20675
rect -8480 20640 -8440 20645
rect -8400 20675 -8360 20680
rect -8400 20645 -8395 20675
rect -8365 20645 -8360 20675
rect -8400 20640 -8360 20645
rect -8320 20675 -8280 20680
rect -8320 20645 -8315 20675
rect -8285 20645 -8280 20675
rect -8320 20640 -8280 20645
rect -8240 20675 -8200 20680
rect -8240 20645 -8235 20675
rect -8205 20645 -8200 20675
rect -8240 20640 -8200 20645
rect -8160 20675 -8120 20680
rect -8160 20645 -8155 20675
rect -8125 20645 -8120 20675
rect -8160 20640 -8120 20645
rect -8080 20675 -8040 20680
rect -8080 20645 -8075 20675
rect -8045 20645 -8040 20675
rect -8080 20640 -8040 20645
rect -8000 20675 -7960 20680
rect -8000 20645 -7995 20675
rect -7965 20645 -7960 20675
rect -8000 20640 -7960 20645
rect -7920 20675 -7880 20680
rect -7920 20645 -7915 20675
rect -7885 20645 -7880 20675
rect -7920 20640 -7880 20645
rect -7840 20675 -7800 20680
rect -7840 20645 -7835 20675
rect -7805 20645 -7800 20675
rect -7840 20640 -7800 20645
rect -7760 20675 -7720 20680
rect -7760 20645 -7755 20675
rect -7725 20645 -7720 20675
rect -7760 20640 -7720 20645
rect -7680 20675 -7640 20680
rect -7680 20645 -7675 20675
rect -7645 20645 -7640 20675
rect -7680 20640 -7640 20645
rect -7600 20675 -7560 20680
rect -7600 20645 -7595 20675
rect -7565 20645 -7560 20675
rect -7600 20640 -7560 20645
rect -7520 20675 -7480 20680
rect -7520 20645 -7515 20675
rect -7485 20645 -7480 20675
rect -7520 20640 -7480 20645
rect -7440 20675 -7400 20680
rect -7440 20645 -7435 20675
rect -7405 20645 -7400 20675
rect -7440 20640 -7400 20645
rect -7360 20675 -7320 20680
rect -7360 20645 -7355 20675
rect -7325 20645 -7320 20675
rect -7360 20640 -7320 20645
rect -7280 20675 -7240 20680
rect -7280 20645 -7275 20675
rect -7245 20645 -7240 20675
rect -7280 20640 -7240 20645
rect -7200 20675 -7160 20680
rect -7200 20645 -7195 20675
rect -7165 20645 -7160 20675
rect -7200 20640 -7160 20645
rect -7120 20675 -7080 20680
rect -7120 20645 -7115 20675
rect -7085 20645 -7080 20675
rect -7120 20640 -7080 20645
rect -7040 20675 -7000 20680
rect -7040 20645 -7035 20675
rect -7005 20645 -7000 20675
rect -7040 20640 -7000 20645
rect -6960 20675 -6920 20680
rect -6960 20645 -6955 20675
rect -6925 20645 -6920 20675
rect -6960 20640 -6920 20645
rect -6880 20675 -6840 20680
rect -6880 20645 -6875 20675
rect -6845 20645 -6840 20675
rect -6880 20640 -6840 20645
rect -6800 20675 -6760 20680
rect -6800 20645 -6795 20675
rect -6765 20645 -6760 20675
rect -6800 20640 -6760 20645
rect -6720 20675 -6680 20680
rect -6720 20645 -6715 20675
rect -6685 20645 -6680 20675
rect -6720 20640 -6680 20645
rect -6640 20675 -6600 20680
rect -6640 20645 -6635 20675
rect -6605 20645 -6600 20675
rect -6640 20640 -6600 20645
rect -6560 20675 -6520 20680
rect -6560 20645 -6555 20675
rect -6525 20645 -6520 20675
rect -6560 20640 -6520 20645
rect -6480 20675 -6440 20680
rect -6480 20645 -6475 20675
rect -6445 20645 -6440 20675
rect -6480 20640 -6440 20645
rect -6400 20675 -6360 20680
rect -6400 20645 -6395 20675
rect -6365 20645 -6360 20675
rect -6400 20640 -6360 20645
rect -6320 20675 -6280 20680
rect -6320 20645 -6315 20675
rect -6285 20645 -6280 20675
rect -6320 20640 -6280 20645
rect -6240 20675 -6200 20680
rect -6240 20645 -6235 20675
rect -6205 20645 -6200 20675
rect -6240 20640 -6200 20645
rect -6160 20675 -6120 20680
rect -6160 20645 -6155 20675
rect -6125 20645 -6120 20675
rect -6160 20640 -6120 20645
rect -5680 20675 -5640 20680
rect -5680 20645 -5675 20675
rect -5645 20645 -5640 20675
rect -5680 20640 -5640 20645
rect -5600 20675 -5560 20680
rect -5600 20645 -5595 20675
rect -5565 20645 -5560 20675
rect -5600 20640 -5560 20645
rect -5520 20675 -5480 20680
rect -5520 20645 -5515 20675
rect -5485 20645 -5480 20675
rect -5520 20640 -5480 20645
rect -5440 20675 -5400 20680
rect -5440 20645 -5435 20675
rect -5405 20645 -5400 20675
rect -5440 20640 -5400 20645
rect -5360 20675 -5320 20680
rect -5360 20645 -5355 20675
rect -5325 20645 -5320 20675
rect -5360 20640 -5320 20645
rect -5280 20675 -5240 20680
rect -5280 20645 -5275 20675
rect -5245 20645 -5240 20675
rect -5280 20640 -5240 20645
rect -5200 20675 -5160 20680
rect -5200 20645 -5195 20675
rect -5165 20645 -5160 20675
rect -5200 20640 -5160 20645
rect -5120 20675 -5080 20680
rect -5120 20645 -5115 20675
rect -5085 20645 -5080 20675
rect -5120 20640 -5080 20645
rect -5040 20675 -5000 20680
rect -5040 20645 -5035 20675
rect -5005 20645 -5000 20675
rect -5040 20640 -5000 20645
rect -4960 20675 -4920 20680
rect -4960 20645 -4955 20675
rect -4925 20645 -4920 20675
rect -4960 20640 -4920 20645
rect -4880 20675 -4840 20680
rect -4880 20645 -4875 20675
rect -4845 20645 -4840 20675
rect -4880 20640 -4840 20645
rect -4800 20675 -4760 20680
rect -4800 20645 -4795 20675
rect -4765 20645 -4760 20675
rect -4800 20640 -4760 20645
rect -4720 20675 -4680 20680
rect -4720 20645 -4715 20675
rect -4685 20645 -4680 20675
rect -4720 20640 -4680 20645
rect -4640 20675 -4600 20680
rect -4640 20645 -4635 20675
rect -4605 20645 -4600 20675
rect -4640 20640 -4600 20645
rect -4560 20675 -4520 20680
rect -4560 20645 -4555 20675
rect -4525 20645 -4520 20675
rect -4560 20640 -4520 20645
rect -4480 20675 -4440 20680
rect -4480 20645 -4475 20675
rect -4445 20645 -4440 20675
rect -4480 20640 -4440 20645
rect -4400 20675 -4360 20680
rect -4400 20645 -4395 20675
rect -4365 20645 -4360 20675
rect -4400 20640 -4360 20645
rect -4320 20675 -4280 20680
rect -4320 20645 -4315 20675
rect -4285 20645 -4280 20675
rect -4320 20640 -4280 20645
rect -4240 20675 -4200 20680
rect -4240 20645 -4235 20675
rect -4205 20645 -4200 20675
rect -4240 20640 -4200 20645
rect -4160 20675 -4120 20680
rect -4160 20645 -4155 20675
rect -4125 20645 -4120 20675
rect -4160 20640 -4120 20645
rect -4080 20675 -4040 20680
rect -4080 20645 -4075 20675
rect -4045 20645 -4040 20675
rect -4080 20640 -4040 20645
rect -4000 20675 -3960 20680
rect -4000 20645 -3995 20675
rect -3965 20645 -3960 20675
rect -4000 20640 -3960 20645
rect -3920 20675 -3880 20680
rect -3920 20645 -3915 20675
rect -3885 20645 -3880 20675
rect -3920 20640 -3880 20645
rect -3840 20675 -3800 20680
rect -3840 20645 -3835 20675
rect -3805 20645 -3800 20675
rect -3840 20640 -3800 20645
rect -3760 20675 -3720 20680
rect -3760 20645 -3755 20675
rect -3725 20645 -3720 20675
rect -3760 20640 -3720 20645
rect -3680 20675 -3640 20680
rect -3680 20645 -3675 20675
rect -3645 20645 -3640 20675
rect -3680 20640 -3640 20645
rect -3600 20675 -3560 20680
rect -3600 20645 -3595 20675
rect -3565 20645 -3560 20675
rect -3600 20640 -3560 20645
rect -3520 20675 -3480 20680
rect -3520 20645 -3515 20675
rect -3485 20645 -3480 20675
rect -3520 20640 -3480 20645
rect -3440 20675 -3400 20680
rect -3440 20645 -3435 20675
rect -3405 20645 -3400 20675
rect -3440 20640 -3400 20645
rect -3360 20675 -3320 20680
rect -3360 20645 -3355 20675
rect -3325 20645 -3320 20675
rect -3360 20640 -3320 20645
rect -3280 20675 -3240 20680
rect -3280 20645 -3275 20675
rect -3245 20645 -3240 20675
rect -3280 20640 -3240 20645
rect -3200 20675 -3160 20680
rect -3200 20645 -3195 20675
rect -3165 20645 -3160 20675
rect -3200 20640 -3160 20645
rect -3120 20675 -3080 20680
rect -3120 20645 -3115 20675
rect -3085 20645 -3080 20675
rect -3120 20640 -3080 20645
rect -3040 20675 -3000 20680
rect -3040 20645 -3035 20675
rect -3005 20645 -3000 20675
rect -3040 20640 -3000 20645
rect -2960 20675 -2920 20680
rect -2960 20645 -2955 20675
rect -2925 20645 -2920 20675
rect -2960 20640 -2920 20645
rect -2880 20675 -2840 20680
rect -2880 20645 -2875 20675
rect -2845 20645 -2840 20675
rect -2880 20640 -2840 20645
rect -2800 20675 -2760 20680
rect -2800 20645 -2795 20675
rect -2765 20645 -2760 20675
rect -2800 20640 -2760 20645
rect -2720 20675 -2680 20680
rect -2720 20645 -2715 20675
rect -2685 20645 -2680 20675
rect -2720 20640 -2680 20645
rect -2640 20675 -2600 20680
rect -2640 20645 -2635 20675
rect -2605 20645 -2600 20675
rect -2640 20640 -2600 20645
rect -2560 20675 -2520 20680
rect -2560 20645 -2555 20675
rect -2525 20645 -2520 20675
rect -2560 20640 -2520 20645
rect -2480 20675 -2440 20680
rect -2480 20645 -2475 20675
rect -2445 20645 -2440 20675
rect -2480 20640 -2440 20645
rect -2400 20675 -2360 20680
rect -2400 20645 -2395 20675
rect -2365 20645 -2360 20675
rect -2400 20640 -2360 20645
rect -2320 20675 -2280 20680
rect -2320 20645 -2315 20675
rect -2285 20645 -2280 20675
rect -2320 20640 -2280 20645
rect -2240 20675 -2200 20680
rect -2240 20645 -2235 20675
rect -2205 20645 -2200 20675
rect -2240 20640 -2200 20645
rect -2160 20675 -2120 20680
rect -2160 20645 -2155 20675
rect -2125 20645 -2120 20675
rect -2160 20640 -2120 20645
rect -2080 20675 -2040 20680
rect -2080 20645 -2075 20675
rect -2045 20645 -2040 20675
rect -2080 20640 -2040 20645
rect -2000 20675 -1960 20680
rect -2000 20645 -1995 20675
rect -1965 20645 -1960 20675
rect -2000 20640 -1960 20645
rect -1920 20670 -1880 20680
rect -1920 20650 -1910 20670
rect -1890 20650 -1880 20670
rect -1920 20640 -1880 20650
rect -1840 20675 -1800 20680
rect -1840 20645 -1835 20675
rect -1805 20645 -1800 20675
rect -1840 20640 -1800 20645
rect -1760 20675 -1720 20680
rect -1760 20645 -1755 20675
rect -1725 20645 -1720 20675
rect -1760 20640 -1720 20645
rect 20520 20675 20560 20680
rect 20520 20645 20525 20675
rect 20555 20645 20560 20675
rect 20520 20640 20560 20645
rect 20600 20675 20640 20680
rect 20600 20645 20605 20675
rect 20635 20645 20640 20675
rect 20600 20640 20640 20645
rect 20680 20675 20720 20680
rect 20680 20645 20685 20675
rect 20715 20645 20720 20675
rect 20680 20640 20720 20645
rect 20760 20675 20800 20680
rect 20760 20645 20765 20675
rect 20795 20645 20800 20675
rect 20760 20640 20800 20645
rect 20840 20675 20880 20680
rect 20840 20645 20845 20675
rect 20875 20645 20880 20675
rect 20840 20640 20880 20645
rect 20920 20675 20960 20680
rect 20920 20645 20925 20675
rect 20955 20645 20960 20675
rect 20920 20640 20960 20645
rect 21000 20675 21040 20680
rect 21000 20645 21005 20675
rect 21035 20645 21040 20675
rect 21000 20640 21040 20645
rect 21080 20675 21120 20680
rect 21080 20645 21085 20675
rect 21115 20645 21120 20675
rect 21080 20640 21120 20645
rect 21160 20675 21200 20680
rect 21160 20645 21165 20675
rect 21195 20645 21200 20675
rect 21160 20640 21200 20645
rect 21240 20675 21280 20680
rect 21240 20645 21245 20675
rect 21275 20645 21280 20675
rect 21240 20640 21280 20645
rect 21320 20675 21360 20680
rect 21320 20645 21325 20675
rect 21355 20645 21360 20675
rect 21320 20640 21360 20645
rect 21400 20675 21440 20680
rect 21400 20645 21405 20675
rect 21435 20645 21440 20675
rect 21400 20640 21440 20645
rect 21480 20675 21520 20680
rect 21480 20645 21485 20675
rect 21515 20645 21520 20675
rect 21480 20640 21520 20645
rect 21560 20675 21600 20680
rect 21560 20645 21565 20675
rect 21595 20645 21600 20675
rect 21560 20640 21600 20645
rect -16560 20515 -16520 20520
rect -16560 20485 -16555 20515
rect -16525 20485 -16520 20515
rect -16560 20480 -16520 20485
rect -16480 20515 -16440 20520
rect -16480 20485 -16475 20515
rect -16445 20485 -16440 20515
rect -16480 20480 -16440 20485
rect -16400 20515 -16360 20520
rect -16400 20485 -16395 20515
rect -16365 20485 -16360 20515
rect -16400 20480 -16360 20485
rect -16320 20515 -16280 20520
rect -16320 20485 -16315 20515
rect -16285 20485 -16280 20515
rect -16320 20480 -16280 20485
rect -16240 20515 -16200 20520
rect -16240 20485 -16235 20515
rect -16205 20485 -16200 20515
rect -16240 20480 -16200 20485
rect -16160 20515 -16120 20520
rect -16160 20485 -16155 20515
rect -16125 20485 -16120 20515
rect -16160 20480 -16120 20485
rect -16080 20515 -16040 20520
rect -16080 20485 -16075 20515
rect -16045 20485 -16040 20515
rect -16080 20480 -16040 20485
rect -16000 20515 -15960 20520
rect -16000 20485 -15995 20515
rect -15965 20485 -15960 20515
rect -16000 20480 -15960 20485
rect -15920 20515 -15880 20520
rect -15920 20485 -15915 20515
rect -15885 20485 -15880 20515
rect -15920 20480 -15880 20485
rect -15840 20515 -15800 20520
rect -15840 20485 -15835 20515
rect -15805 20485 -15800 20515
rect -15840 20480 -15800 20485
rect -15760 20515 -15720 20520
rect -15760 20485 -15755 20515
rect -15725 20485 -15720 20515
rect -15760 20480 -15720 20485
rect -15680 20515 -15640 20520
rect -15680 20485 -15675 20515
rect -15645 20485 -15640 20515
rect -15680 20480 -15640 20485
rect -15600 20515 -15560 20520
rect -15600 20485 -15595 20515
rect -15565 20485 -15560 20515
rect -15600 20480 -15560 20485
rect -14960 20515 -14920 20520
rect -14960 20485 -14955 20515
rect -14925 20485 -14920 20515
rect -14960 20480 -14920 20485
rect -14880 20515 -14840 20520
rect -14880 20485 -14875 20515
rect -14845 20485 -14840 20515
rect -14880 20480 -14840 20485
rect -14800 20515 -14760 20520
rect -14800 20485 -14795 20515
rect -14765 20485 -14760 20515
rect -14800 20480 -14760 20485
rect -14720 20515 -14680 20520
rect -14720 20485 -14715 20515
rect -14685 20485 -14680 20515
rect -14720 20480 -14680 20485
rect -14640 20515 -14600 20520
rect -14640 20485 -14635 20515
rect -14605 20485 -14600 20515
rect -14640 20480 -14600 20485
rect -14560 20515 -14520 20520
rect -14560 20485 -14555 20515
rect -14525 20485 -14520 20515
rect -14560 20480 -14520 20485
rect -14480 20515 -14440 20520
rect -14480 20485 -14475 20515
rect -14445 20485 -14440 20515
rect -14480 20480 -14440 20485
rect -14400 20515 -14360 20520
rect -14400 20485 -14395 20515
rect -14365 20485 -14360 20515
rect -14400 20480 -14360 20485
rect -14320 20515 -14280 20520
rect -14320 20485 -14315 20515
rect -14285 20485 -14280 20515
rect -14320 20480 -14280 20485
rect -14240 20515 -14200 20520
rect -14240 20485 -14235 20515
rect -14205 20485 -14200 20515
rect -14240 20480 -14200 20485
rect -14160 20515 -14120 20520
rect -14160 20485 -14155 20515
rect -14125 20485 -14120 20515
rect -14160 20480 -14120 20485
rect -14080 20515 -14040 20520
rect -14080 20485 -14075 20515
rect -14045 20485 -14040 20515
rect -14080 20480 -14040 20485
rect -14000 20515 -13960 20520
rect -14000 20485 -13995 20515
rect -13965 20485 -13960 20515
rect -14000 20480 -13960 20485
rect -13920 20515 -13880 20520
rect -13920 20485 -13915 20515
rect -13885 20485 -13880 20515
rect -13920 20480 -13880 20485
rect -13840 20515 -13800 20520
rect -13840 20485 -13835 20515
rect -13805 20485 -13800 20515
rect -13840 20480 -13800 20485
rect -13760 20515 -13720 20520
rect -13760 20485 -13755 20515
rect -13725 20485 -13720 20515
rect -13760 20480 -13720 20485
rect -13680 20515 -13640 20520
rect -13680 20485 -13675 20515
rect -13645 20485 -13640 20515
rect -13680 20480 -13640 20485
rect -13600 20515 -13560 20520
rect -13600 20485 -13595 20515
rect -13565 20485 -13560 20515
rect -13600 20480 -13560 20485
rect -13520 20515 -13480 20520
rect -13520 20485 -13515 20515
rect -13485 20485 -13480 20515
rect -13520 20480 -13480 20485
rect -13440 20515 -13400 20520
rect -13440 20485 -13435 20515
rect -13405 20485 -13400 20515
rect -13440 20480 -13400 20485
rect -13360 20515 -13320 20520
rect -13360 20485 -13355 20515
rect -13325 20485 -13320 20515
rect -13360 20480 -13320 20485
rect -13280 20515 -13240 20520
rect -13280 20485 -13275 20515
rect -13245 20485 -13240 20515
rect -13280 20480 -13240 20485
rect -13200 20515 -13160 20520
rect -13200 20485 -13195 20515
rect -13165 20485 -13160 20515
rect -13200 20480 -13160 20485
rect -13120 20515 -13080 20520
rect -13120 20485 -13115 20515
rect -13085 20485 -13080 20515
rect -13120 20480 -13080 20485
rect -13040 20515 -13000 20520
rect -13040 20485 -13035 20515
rect -13005 20485 -13000 20515
rect -13040 20480 -13000 20485
rect -12960 20515 -12920 20520
rect -12960 20485 -12955 20515
rect -12925 20485 -12920 20515
rect -12960 20480 -12920 20485
rect -12880 20515 -12840 20520
rect -12880 20485 -12875 20515
rect -12845 20485 -12840 20515
rect -12880 20480 -12840 20485
rect -12800 20515 -12760 20520
rect -12800 20485 -12795 20515
rect -12765 20485 -12760 20515
rect -12800 20480 -12760 20485
rect -12720 20515 -12680 20520
rect -12720 20485 -12715 20515
rect -12685 20485 -12680 20515
rect -12720 20480 -12680 20485
rect -12640 20515 -12600 20520
rect -12640 20485 -12635 20515
rect -12605 20485 -12600 20515
rect -12640 20480 -12600 20485
rect -12560 20515 -12520 20520
rect -12560 20485 -12555 20515
rect -12525 20485 -12520 20515
rect -12560 20480 -12520 20485
rect -12480 20515 -12440 20520
rect -12480 20485 -12475 20515
rect -12445 20485 -12440 20515
rect -12480 20480 -12440 20485
rect -12400 20515 -12360 20520
rect -12400 20485 -12395 20515
rect -12365 20485 -12360 20515
rect -12400 20480 -12360 20485
rect -12320 20515 -12280 20520
rect -12320 20485 -12315 20515
rect -12285 20485 -12280 20515
rect -12320 20480 -12280 20485
rect -12240 20515 -12200 20520
rect -12240 20485 -12235 20515
rect -12205 20485 -12200 20515
rect -12240 20480 -12200 20485
rect -12160 20515 -12120 20520
rect -12160 20485 -12155 20515
rect -12125 20485 -12120 20515
rect -12160 20480 -12120 20485
rect -12080 20515 -12040 20520
rect -12080 20485 -12075 20515
rect -12045 20485 -12040 20515
rect -12080 20480 -12040 20485
rect -12000 20515 -11960 20520
rect -12000 20485 -11995 20515
rect -11965 20485 -11960 20515
rect -12000 20480 -11960 20485
rect -11920 20515 -11880 20520
rect -11920 20485 -11915 20515
rect -11885 20485 -11880 20515
rect -11920 20480 -11880 20485
rect -11840 20515 -11800 20520
rect -11840 20485 -11835 20515
rect -11805 20485 -11800 20515
rect -11840 20480 -11800 20485
rect -11760 20515 -11720 20520
rect -11760 20485 -11755 20515
rect -11725 20485 -11720 20515
rect -11760 20480 -11720 20485
rect -11680 20515 -11640 20520
rect -11680 20485 -11675 20515
rect -11645 20485 -11640 20515
rect -11680 20480 -11640 20485
rect -11600 20515 -11560 20520
rect -11600 20485 -11595 20515
rect -11565 20485 -11560 20515
rect -11600 20480 -11560 20485
rect -11520 20515 -11480 20520
rect -11520 20485 -11515 20515
rect -11485 20485 -11480 20515
rect -11520 20480 -11480 20485
rect -11440 20515 -11400 20520
rect -11440 20485 -11435 20515
rect -11405 20485 -11400 20515
rect -11440 20480 -11400 20485
rect -11360 20515 -11320 20520
rect -11360 20485 -11355 20515
rect -11325 20485 -11320 20515
rect -11360 20480 -11320 20485
rect -11280 20515 -11240 20520
rect -11280 20485 -11275 20515
rect -11245 20485 -11240 20515
rect -11280 20480 -11240 20485
rect -11200 20515 -11160 20520
rect -11200 20485 -11195 20515
rect -11165 20485 -11160 20515
rect -11200 20480 -11160 20485
rect -11120 20515 -11080 20520
rect -11120 20485 -11115 20515
rect -11085 20485 -11080 20515
rect -11120 20480 -11080 20485
rect -11040 20515 -11000 20520
rect -11040 20485 -11035 20515
rect -11005 20485 -11000 20515
rect -11040 20480 -11000 20485
rect -10960 20515 -10920 20520
rect -10960 20485 -10955 20515
rect -10925 20485 -10920 20515
rect -10960 20480 -10920 20485
rect -10880 20515 -10840 20520
rect -10880 20485 -10875 20515
rect -10845 20485 -10840 20515
rect -10880 20480 -10840 20485
rect -10800 20515 -10760 20520
rect -10800 20485 -10795 20515
rect -10765 20485 -10760 20515
rect -10800 20480 -10760 20485
rect -10720 20515 -10680 20520
rect -10720 20485 -10715 20515
rect -10685 20485 -10680 20515
rect -10720 20480 -10680 20485
rect -10640 20515 -10600 20520
rect -10640 20485 -10635 20515
rect -10605 20485 -10600 20515
rect -10640 20480 -10600 20485
rect -10560 20515 -10520 20520
rect -10560 20485 -10555 20515
rect -10525 20485 -10520 20515
rect -10560 20480 -10520 20485
rect -10480 20515 -10440 20520
rect -10480 20485 -10475 20515
rect -10445 20485 -10440 20515
rect -10480 20480 -10440 20485
rect -10400 20515 -10360 20520
rect -10400 20485 -10395 20515
rect -10365 20485 -10360 20515
rect -10400 20480 -10360 20485
rect -10320 20515 -10280 20520
rect -10320 20485 -10315 20515
rect -10285 20485 -10280 20515
rect -10320 20480 -10280 20485
rect -10240 20515 -10200 20520
rect -10240 20485 -10235 20515
rect -10205 20485 -10200 20515
rect -10240 20480 -10200 20485
rect -10160 20515 -10120 20520
rect -10160 20485 -10155 20515
rect -10125 20485 -10120 20515
rect -10160 20480 -10120 20485
rect -10080 20515 -10040 20520
rect -10080 20485 -10075 20515
rect -10045 20485 -10040 20515
rect -10080 20480 -10040 20485
rect -10000 20515 -9960 20520
rect -10000 20485 -9995 20515
rect -9965 20485 -9960 20515
rect -10000 20480 -9960 20485
rect -9920 20515 -9880 20520
rect -9920 20485 -9915 20515
rect -9885 20485 -9880 20515
rect -9920 20480 -9880 20485
rect -9840 20515 -9800 20520
rect -9840 20485 -9835 20515
rect -9805 20485 -9800 20515
rect -9840 20480 -9800 20485
rect -9760 20515 -9720 20520
rect -9760 20485 -9755 20515
rect -9725 20485 -9720 20515
rect -9760 20480 -9720 20485
rect -9680 20515 -9640 20520
rect -9680 20485 -9675 20515
rect -9645 20485 -9640 20515
rect -9680 20480 -9640 20485
rect -9600 20515 -9560 20520
rect -9600 20485 -9595 20515
rect -9565 20485 -9560 20515
rect -9600 20480 -9560 20485
rect -9520 20515 -9480 20520
rect -9520 20485 -9515 20515
rect -9485 20485 -9480 20515
rect -9520 20480 -9480 20485
rect -9440 20515 -9400 20520
rect -9440 20485 -9435 20515
rect -9405 20485 -9400 20515
rect -9440 20480 -9400 20485
rect -9360 20515 -9320 20520
rect -9360 20485 -9355 20515
rect -9325 20485 -9320 20515
rect -9360 20480 -9320 20485
rect -9280 20515 -9240 20520
rect -9280 20485 -9275 20515
rect -9245 20485 -9240 20515
rect -9280 20480 -9240 20485
rect -9200 20515 -9160 20520
rect -9200 20485 -9195 20515
rect -9165 20485 -9160 20515
rect -9200 20480 -9160 20485
rect -9120 20515 -9080 20520
rect -9120 20485 -9115 20515
rect -9085 20485 -9080 20515
rect -9120 20480 -9080 20485
rect -9040 20515 -9000 20520
rect -9040 20485 -9035 20515
rect -9005 20485 -9000 20515
rect -9040 20480 -9000 20485
rect -8960 20515 -8920 20520
rect -8960 20485 -8955 20515
rect -8925 20485 -8920 20515
rect -8960 20480 -8920 20485
rect -8880 20515 -8840 20520
rect -8880 20485 -8875 20515
rect -8845 20485 -8840 20515
rect -8880 20480 -8840 20485
rect -8800 20515 -8760 20520
rect -8800 20485 -8795 20515
rect -8765 20485 -8760 20515
rect -8800 20480 -8760 20485
rect -8720 20515 -8680 20520
rect -8720 20485 -8715 20515
rect -8685 20485 -8680 20515
rect -8720 20480 -8680 20485
rect -8640 20515 -8600 20520
rect -8640 20485 -8635 20515
rect -8605 20485 -8600 20515
rect -8640 20480 -8600 20485
rect -8560 20515 -8520 20520
rect -8560 20485 -8555 20515
rect -8525 20485 -8520 20515
rect -8560 20480 -8520 20485
rect -8480 20515 -8440 20520
rect -8480 20485 -8475 20515
rect -8445 20485 -8440 20515
rect -8480 20480 -8440 20485
rect -8400 20515 -8360 20520
rect -8400 20485 -8395 20515
rect -8365 20485 -8360 20515
rect -8400 20480 -8360 20485
rect -8320 20515 -8280 20520
rect -8320 20485 -8315 20515
rect -8285 20485 -8280 20515
rect -8320 20480 -8280 20485
rect -8240 20515 -8200 20520
rect -8240 20485 -8235 20515
rect -8205 20485 -8200 20515
rect -8240 20480 -8200 20485
rect -8160 20515 -8120 20520
rect -8160 20485 -8155 20515
rect -8125 20485 -8120 20515
rect -8160 20480 -8120 20485
rect -8080 20515 -8040 20520
rect -8080 20485 -8075 20515
rect -8045 20485 -8040 20515
rect -8080 20480 -8040 20485
rect -8000 20515 -7960 20520
rect -8000 20485 -7995 20515
rect -7965 20485 -7960 20515
rect -8000 20480 -7960 20485
rect -7920 20515 -7880 20520
rect -7920 20485 -7915 20515
rect -7885 20485 -7880 20515
rect -7920 20480 -7880 20485
rect -7840 20515 -7800 20520
rect -7840 20485 -7835 20515
rect -7805 20485 -7800 20515
rect -7840 20480 -7800 20485
rect -7760 20515 -7720 20520
rect -7760 20485 -7755 20515
rect -7725 20485 -7720 20515
rect -7760 20480 -7720 20485
rect -7680 20515 -7640 20520
rect -7680 20485 -7675 20515
rect -7645 20485 -7640 20515
rect -7680 20480 -7640 20485
rect -7600 20515 -7560 20520
rect -7600 20485 -7595 20515
rect -7565 20485 -7560 20515
rect -7600 20480 -7560 20485
rect -7520 20515 -7480 20520
rect -7520 20485 -7515 20515
rect -7485 20485 -7480 20515
rect -7520 20480 -7480 20485
rect -7440 20515 -7400 20520
rect -7440 20485 -7435 20515
rect -7405 20485 -7400 20515
rect -7440 20480 -7400 20485
rect -7360 20515 -7320 20520
rect -7360 20485 -7355 20515
rect -7325 20485 -7320 20515
rect -7360 20480 -7320 20485
rect -7280 20515 -7240 20520
rect -7280 20485 -7275 20515
rect -7245 20485 -7240 20515
rect -7280 20480 -7240 20485
rect -7200 20515 -7160 20520
rect -7200 20485 -7195 20515
rect -7165 20485 -7160 20515
rect -7200 20480 -7160 20485
rect -7120 20515 -7080 20520
rect -7120 20485 -7115 20515
rect -7085 20485 -7080 20515
rect -7120 20480 -7080 20485
rect -7040 20515 -7000 20520
rect -7040 20485 -7035 20515
rect -7005 20485 -7000 20515
rect -7040 20480 -7000 20485
rect -6960 20515 -6920 20520
rect -6960 20485 -6955 20515
rect -6925 20485 -6920 20515
rect -6960 20480 -6920 20485
rect -6880 20515 -6840 20520
rect -6880 20485 -6875 20515
rect -6845 20485 -6840 20515
rect -6880 20480 -6840 20485
rect -6800 20515 -6760 20520
rect -6800 20485 -6795 20515
rect -6765 20485 -6760 20515
rect -6800 20480 -6760 20485
rect -6720 20515 -6680 20520
rect -6720 20485 -6715 20515
rect -6685 20485 -6680 20515
rect -6720 20480 -6680 20485
rect -6640 20515 -6600 20520
rect -6640 20485 -6635 20515
rect -6605 20485 -6600 20515
rect -6640 20480 -6600 20485
rect -6560 20515 -6520 20520
rect -6560 20485 -6555 20515
rect -6525 20485 -6520 20515
rect -6560 20480 -6520 20485
rect -6480 20515 -6440 20520
rect -6480 20485 -6475 20515
rect -6445 20485 -6440 20515
rect -6480 20480 -6440 20485
rect -6400 20515 -6360 20520
rect -6400 20485 -6395 20515
rect -6365 20485 -6360 20515
rect -6400 20480 -6360 20485
rect -6320 20515 -6280 20520
rect -6320 20485 -6315 20515
rect -6285 20485 -6280 20515
rect -6320 20480 -6280 20485
rect -6240 20515 -6200 20520
rect -6240 20485 -6235 20515
rect -6205 20485 -6200 20515
rect -6240 20480 -6200 20485
rect -6160 20515 -6120 20520
rect -6160 20485 -6155 20515
rect -6125 20485 -6120 20515
rect -6160 20480 -6120 20485
rect -5680 20515 -5640 20520
rect -5680 20485 -5675 20515
rect -5645 20485 -5640 20515
rect -5680 20480 -5640 20485
rect -5600 20515 -5560 20520
rect -5600 20485 -5595 20515
rect -5565 20485 -5560 20515
rect -5600 20480 -5560 20485
rect -5520 20515 -5480 20520
rect -5520 20485 -5515 20515
rect -5485 20485 -5480 20515
rect -5520 20480 -5480 20485
rect -5440 20515 -5400 20520
rect -5440 20485 -5435 20515
rect -5405 20485 -5400 20515
rect -5440 20480 -5400 20485
rect -5360 20515 -5320 20520
rect -5360 20485 -5355 20515
rect -5325 20485 -5320 20515
rect -5360 20480 -5320 20485
rect -5280 20515 -5240 20520
rect -5280 20485 -5275 20515
rect -5245 20485 -5240 20515
rect -5280 20480 -5240 20485
rect -5200 20515 -5160 20520
rect -5200 20485 -5195 20515
rect -5165 20485 -5160 20515
rect -5200 20480 -5160 20485
rect -5120 20515 -5080 20520
rect -5120 20485 -5115 20515
rect -5085 20485 -5080 20515
rect -5120 20480 -5080 20485
rect -5040 20515 -5000 20520
rect -5040 20485 -5035 20515
rect -5005 20485 -5000 20515
rect -5040 20480 -5000 20485
rect -4960 20515 -4920 20520
rect -4960 20485 -4955 20515
rect -4925 20485 -4920 20515
rect -4960 20480 -4920 20485
rect -4880 20515 -4840 20520
rect -4880 20485 -4875 20515
rect -4845 20485 -4840 20515
rect -4880 20480 -4840 20485
rect -4800 20515 -4760 20520
rect -4800 20485 -4795 20515
rect -4765 20485 -4760 20515
rect -4800 20480 -4760 20485
rect -4720 20515 -4680 20520
rect -4720 20485 -4715 20515
rect -4685 20485 -4680 20515
rect -4720 20480 -4680 20485
rect -4640 20515 -4600 20520
rect -4640 20485 -4635 20515
rect -4605 20485 -4600 20515
rect -4640 20480 -4600 20485
rect -4560 20515 -4520 20520
rect -4560 20485 -4555 20515
rect -4525 20485 -4520 20515
rect -4560 20480 -4520 20485
rect -4480 20515 -4440 20520
rect -4480 20485 -4475 20515
rect -4445 20485 -4440 20515
rect -4480 20480 -4440 20485
rect -4400 20515 -4360 20520
rect -4400 20485 -4395 20515
rect -4365 20485 -4360 20515
rect -4400 20480 -4360 20485
rect -4320 20515 -4280 20520
rect -4320 20485 -4315 20515
rect -4285 20485 -4280 20515
rect -4320 20480 -4280 20485
rect -4240 20515 -4200 20520
rect -4240 20485 -4235 20515
rect -4205 20485 -4200 20515
rect -4240 20480 -4200 20485
rect -4160 20515 -4120 20520
rect -4160 20485 -4155 20515
rect -4125 20485 -4120 20515
rect -4160 20480 -4120 20485
rect -4080 20515 -4040 20520
rect -4080 20485 -4075 20515
rect -4045 20485 -4040 20515
rect -4080 20480 -4040 20485
rect -4000 20515 -3960 20520
rect -4000 20485 -3995 20515
rect -3965 20485 -3960 20515
rect -4000 20480 -3960 20485
rect -3920 20515 -3880 20520
rect -3920 20485 -3915 20515
rect -3885 20485 -3880 20515
rect -3920 20480 -3880 20485
rect -3840 20515 -3800 20520
rect -3840 20485 -3835 20515
rect -3805 20485 -3800 20515
rect -3840 20480 -3800 20485
rect -3760 20515 -3720 20520
rect -3760 20485 -3755 20515
rect -3725 20485 -3720 20515
rect -3760 20480 -3720 20485
rect -3680 20515 -3640 20520
rect -3680 20485 -3675 20515
rect -3645 20485 -3640 20515
rect -3680 20480 -3640 20485
rect -3600 20515 -3560 20520
rect -3600 20485 -3595 20515
rect -3565 20485 -3560 20515
rect -3600 20480 -3560 20485
rect -3520 20515 -3480 20520
rect -3520 20485 -3515 20515
rect -3485 20485 -3480 20515
rect -3520 20480 -3480 20485
rect -3440 20515 -3400 20520
rect -3440 20485 -3435 20515
rect -3405 20485 -3400 20515
rect -3440 20480 -3400 20485
rect -3360 20515 -3320 20520
rect -3360 20485 -3355 20515
rect -3325 20485 -3320 20515
rect -3360 20480 -3320 20485
rect -3280 20515 -3240 20520
rect -3280 20485 -3275 20515
rect -3245 20485 -3240 20515
rect -3280 20480 -3240 20485
rect -3200 20515 -3160 20520
rect -3200 20485 -3195 20515
rect -3165 20485 -3160 20515
rect -3200 20480 -3160 20485
rect -3120 20515 -3080 20520
rect -3120 20485 -3115 20515
rect -3085 20485 -3080 20515
rect -3120 20480 -3080 20485
rect -3040 20515 -3000 20520
rect -3040 20485 -3035 20515
rect -3005 20485 -3000 20515
rect -3040 20480 -3000 20485
rect -2960 20515 -2920 20520
rect -2960 20485 -2955 20515
rect -2925 20485 -2920 20515
rect -2960 20480 -2920 20485
rect -2880 20515 -2840 20520
rect -2880 20485 -2875 20515
rect -2845 20485 -2840 20515
rect -2880 20480 -2840 20485
rect -2800 20515 -2760 20520
rect -2800 20485 -2795 20515
rect -2765 20485 -2760 20515
rect -2800 20480 -2760 20485
rect -2720 20515 -2680 20520
rect -2720 20485 -2715 20515
rect -2685 20485 -2680 20515
rect -2720 20480 -2680 20485
rect -2640 20515 -2600 20520
rect -2640 20485 -2635 20515
rect -2605 20485 -2600 20515
rect -2640 20480 -2600 20485
rect -2560 20515 -2520 20520
rect -2560 20485 -2555 20515
rect -2525 20485 -2520 20515
rect -2560 20480 -2520 20485
rect -2480 20515 -2440 20520
rect -2480 20485 -2475 20515
rect -2445 20485 -2440 20515
rect -2480 20480 -2440 20485
rect -2400 20515 -2360 20520
rect -2400 20485 -2395 20515
rect -2365 20485 -2360 20515
rect -2400 20480 -2360 20485
rect -2320 20515 -2280 20520
rect -2320 20485 -2315 20515
rect -2285 20485 -2280 20515
rect -2320 20480 -2280 20485
rect -2240 20515 -2200 20520
rect -2240 20485 -2235 20515
rect -2205 20485 -2200 20515
rect -2240 20480 -2200 20485
rect -2160 20515 -2120 20520
rect -2160 20485 -2155 20515
rect -2125 20485 -2120 20515
rect -2160 20480 -2120 20485
rect -2080 20515 -2040 20520
rect -2080 20485 -2075 20515
rect -2045 20485 -2040 20515
rect -2080 20480 -2040 20485
rect -2000 20515 -1960 20520
rect -2000 20485 -1995 20515
rect -1965 20485 -1960 20515
rect -2000 20480 -1960 20485
rect -1920 20510 -1880 20520
rect -1920 20490 -1910 20510
rect -1890 20490 -1880 20510
rect -1920 20480 -1880 20490
rect -1840 20515 -1800 20520
rect -1840 20485 -1835 20515
rect -1805 20485 -1800 20515
rect -1840 20480 -1800 20485
rect -1760 20515 -1720 20520
rect -1760 20485 -1755 20515
rect -1725 20485 -1720 20515
rect -1760 20480 -1720 20485
rect 20520 20515 20560 20520
rect 20520 20485 20525 20515
rect 20555 20485 20560 20515
rect 20520 20480 20560 20485
rect 20600 20515 20640 20520
rect 20600 20485 20605 20515
rect 20635 20485 20640 20515
rect 20600 20480 20640 20485
rect 20680 20515 20720 20520
rect 20680 20485 20685 20515
rect 20715 20485 20720 20515
rect 20680 20480 20720 20485
rect 20760 20515 20800 20520
rect 20760 20485 20765 20515
rect 20795 20485 20800 20515
rect 20760 20480 20800 20485
rect 20840 20515 20880 20520
rect 20840 20485 20845 20515
rect 20875 20485 20880 20515
rect 20840 20480 20880 20485
rect 20920 20515 20960 20520
rect 20920 20485 20925 20515
rect 20955 20485 20960 20515
rect 20920 20480 20960 20485
rect 21000 20515 21040 20520
rect 21000 20485 21005 20515
rect 21035 20485 21040 20515
rect 21000 20480 21040 20485
rect 21080 20515 21120 20520
rect 21080 20485 21085 20515
rect 21115 20485 21120 20515
rect 21080 20480 21120 20485
rect 21160 20515 21200 20520
rect 21160 20485 21165 20515
rect 21195 20485 21200 20515
rect 21160 20480 21200 20485
rect 21240 20515 21280 20520
rect 21240 20485 21245 20515
rect 21275 20485 21280 20515
rect 21240 20480 21280 20485
rect 21320 20515 21360 20520
rect 21320 20485 21325 20515
rect 21355 20485 21360 20515
rect 21320 20480 21360 20485
rect 21400 20515 21440 20520
rect 21400 20485 21405 20515
rect 21435 20485 21440 20515
rect 21400 20480 21440 20485
rect 21480 20515 21520 20520
rect 21480 20485 21485 20515
rect 21515 20485 21520 20515
rect 21480 20480 21520 20485
rect 21560 20515 21600 20520
rect 21560 20485 21565 20515
rect 21595 20485 21600 20515
rect 21560 20480 21600 20485
rect -5280 20355 -5240 20360
rect -5280 20325 -5275 20355
rect -5245 20325 -5240 20355
rect -5280 20320 -5240 20325
rect -5120 20355 -5080 20360
rect -5120 20325 -5115 20355
rect -5085 20325 -5080 20355
rect -5120 20320 -5080 20325
rect -5040 20355 -5000 20360
rect -5040 20325 -5035 20355
rect -5005 20325 -5000 20355
rect -5040 20320 -5000 20325
rect -4960 20355 -4920 20360
rect -4960 20325 -4955 20355
rect -4925 20325 -4920 20355
rect -4960 20320 -4920 20325
rect -4880 20355 -4840 20360
rect -4880 20325 -4875 20355
rect -4845 20325 -4840 20355
rect -4880 20320 -4840 20325
rect -4800 20355 -4760 20360
rect -4800 20325 -4795 20355
rect -4765 20325 -4760 20355
rect -4800 20320 -4760 20325
rect -4720 20355 -4680 20360
rect -4720 20325 -4715 20355
rect -4685 20325 -4680 20355
rect -4720 20320 -4680 20325
rect -4640 20355 -4600 20360
rect -4640 20325 -4635 20355
rect -4605 20325 -4600 20355
rect -4640 20320 -4600 20325
rect -4560 20355 -4520 20360
rect -4560 20325 -4555 20355
rect -4525 20325 -4520 20355
rect -4560 20320 -4520 20325
rect -4480 20355 -4440 20360
rect -4480 20325 -4475 20355
rect -4445 20325 -4440 20355
rect -4480 20320 -4440 20325
rect -4400 20355 -4360 20360
rect -4400 20325 -4395 20355
rect -4365 20325 -4360 20355
rect -4400 20320 -4360 20325
rect -4320 20355 -4280 20360
rect -4320 20325 -4315 20355
rect -4285 20325 -4280 20355
rect -4320 20320 -4280 20325
rect -4240 20355 -4200 20360
rect -4240 20325 -4235 20355
rect -4205 20325 -4200 20355
rect -4240 20320 -4200 20325
rect -4160 20355 -4120 20360
rect -4160 20325 -4155 20355
rect -4125 20325 -4120 20355
rect -4160 20320 -4120 20325
rect -4080 20355 -4040 20360
rect -4080 20325 -4075 20355
rect -4045 20325 -4040 20355
rect -4080 20320 -4040 20325
rect -4000 20355 -3960 20360
rect -4000 20325 -3995 20355
rect -3965 20325 -3960 20355
rect -4000 20320 -3960 20325
rect -3920 20355 -3880 20360
rect -3920 20325 -3915 20355
rect -3885 20325 -3880 20355
rect -3920 20320 -3880 20325
rect -3840 20355 -3800 20360
rect -3840 20325 -3835 20355
rect -3805 20325 -3800 20355
rect -3840 20320 -3800 20325
rect -3760 20355 -3720 20360
rect -3760 20325 -3755 20355
rect -3725 20325 -3720 20355
rect -3760 20320 -3720 20325
rect -3680 20355 -3640 20360
rect -3680 20325 -3675 20355
rect -3645 20325 -3640 20355
rect -3680 20320 -3640 20325
rect -3600 20355 -3560 20360
rect -3600 20325 -3595 20355
rect -3565 20325 -3560 20355
rect -3600 20320 -3560 20325
rect -3520 20355 -3480 20360
rect -3520 20325 -3515 20355
rect -3485 20325 -3480 20355
rect -3520 20320 -3480 20325
rect -3440 20355 -3400 20360
rect -3440 20325 -3435 20355
rect -3405 20325 -3400 20355
rect -3440 20320 -3400 20325
rect -3360 20355 -3320 20360
rect -3360 20325 -3355 20355
rect -3325 20325 -3320 20355
rect -3360 20320 -3320 20325
rect -3280 20355 -3240 20360
rect -3280 20325 -3275 20355
rect -3245 20325 -3240 20355
rect -3280 20320 -3240 20325
rect -3200 20355 -3160 20360
rect -3200 20325 -3195 20355
rect -3165 20325 -3160 20355
rect -3200 20320 -3160 20325
rect -3120 20355 -3080 20360
rect -3120 20325 -3115 20355
rect -3085 20325 -3080 20355
rect -3120 20320 -3080 20325
rect -3040 20355 -3000 20360
rect -3040 20325 -3035 20355
rect -3005 20325 -3000 20355
rect -3040 20320 -3000 20325
rect -2960 20355 -2920 20360
rect -2960 20325 -2955 20355
rect -2925 20325 -2920 20355
rect -2960 20320 -2920 20325
rect -2880 20355 -2840 20360
rect -2880 20325 -2875 20355
rect -2845 20325 -2840 20355
rect -2880 20320 -2840 20325
rect -2800 20355 -2760 20360
rect -2800 20325 -2795 20355
rect -2765 20325 -2760 20355
rect -2800 20320 -2760 20325
rect -2720 20355 -2680 20360
rect -2720 20325 -2715 20355
rect -2685 20325 -2680 20355
rect -2720 20320 -2680 20325
rect -2640 20355 -2600 20360
rect -2640 20325 -2635 20355
rect -2605 20325 -2600 20355
rect -2640 20320 -2600 20325
rect -2560 20355 -2520 20360
rect -2560 20325 -2555 20355
rect -2525 20325 -2520 20355
rect -2560 20320 -2520 20325
rect -2480 20355 -2440 20360
rect -2480 20325 -2475 20355
rect -2445 20325 -2440 20355
rect -2480 20320 -2440 20325
rect -2400 20355 -2360 20360
rect -2400 20325 -2395 20355
rect -2365 20325 -2360 20355
rect -2400 20320 -2360 20325
rect -2320 20355 -2280 20360
rect -2320 20325 -2315 20355
rect -2285 20325 -2280 20355
rect -2320 20320 -2280 20325
rect -2240 20355 -2200 20360
rect -2240 20325 -2235 20355
rect -2205 20325 -2200 20355
rect -2240 20320 -2200 20325
rect -2160 20355 -2120 20360
rect -2160 20325 -2155 20355
rect -2125 20325 -2120 20355
rect -2160 20320 -2120 20325
rect -2080 20355 -2040 20360
rect -2080 20325 -2075 20355
rect -2045 20325 -2040 20355
rect -2080 20320 -2040 20325
rect -2000 20355 -1960 20360
rect -2000 20325 -1995 20355
rect -1965 20325 -1960 20355
rect -2000 20320 -1960 20325
rect -1840 20355 -1800 20360
rect -1840 20325 -1835 20355
rect -1805 20325 -1800 20355
rect -1840 20320 -1800 20325
rect -1760 20355 -1720 20360
rect -1760 20325 -1755 20355
rect -1725 20325 -1720 20355
rect -1760 20320 -1720 20325
rect -5280 20195 -5240 20200
rect -5280 20165 -5275 20195
rect -5245 20165 -5240 20195
rect -5280 20160 -5240 20165
rect -5120 20195 -5080 20200
rect -5120 20165 -5115 20195
rect -5085 20165 -5080 20195
rect -5120 20160 -5080 20165
rect -5040 20195 -5000 20200
rect -5040 20165 -5035 20195
rect -5005 20165 -5000 20195
rect -5040 20160 -5000 20165
rect -4960 20195 -4920 20200
rect -4960 20165 -4955 20195
rect -4925 20165 -4920 20195
rect -4960 20160 -4920 20165
rect -4880 20195 -4840 20200
rect -4880 20165 -4875 20195
rect -4845 20165 -4840 20195
rect -4880 20160 -4840 20165
rect -4800 20195 -4760 20200
rect -4800 20165 -4795 20195
rect -4765 20165 -4760 20195
rect -4800 20160 -4760 20165
rect -4720 20195 -4680 20200
rect -4720 20165 -4715 20195
rect -4685 20165 -4680 20195
rect -4720 20160 -4680 20165
rect -4640 20195 -4600 20200
rect -4640 20165 -4635 20195
rect -4605 20165 -4600 20195
rect -4640 20160 -4600 20165
rect -4560 20195 -4520 20200
rect -4560 20165 -4555 20195
rect -4525 20165 -4520 20195
rect -4560 20160 -4520 20165
rect -4480 20195 -4440 20200
rect -4480 20165 -4475 20195
rect -4445 20165 -4440 20195
rect -4480 20160 -4440 20165
rect -4400 20195 -4360 20200
rect -4400 20165 -4395 20195
rect -4365 20165 -4360 20195
rect -4400 20160 -4360 20165
rect -4320 20195 -4280 20200
rect -4320 20165 -4315 20195
rect -4285 20165 -4280 20195
rect -4320 20160 -4280 20165
rect -4240 20195 -4200 20200
rect -4240 20165 -4235 20195
rect -4205 20165 -4200 20195
rect -4240 20160 -4200 20165
rect -4160 20195 -4120 20200
rect -4160 20165 -4155 20195
rect -4125 20165 -4120 20195
rect -4160 20160 -4120 20165
rect -4080 20195 -4040 20200
rect -4080 20165 -4075 20195
rect -4045 20165 -4040 20195
rect -4080 20160 -4040 20165
rect -4000 20195 -3960 20200
rect -4000 20165 -3995 20195
rect -3965 20165 -3960 20195
rect -4000 20160 -3960 20165
rect -3920 20195 -3880 20200
rect -3920 20165 -3915 20195
rect -3885 20165 -3880 20195
rect -3920 20160 -3880 20165
rect -3840 20195 -3800 20200
rect -3840 20165 -3835 20195
rect -3805 20165 -3800 20195
rect -3840 20160 -3800 20165
rect -3760 20195 -3720 20200
rect -3760 20165 -3755 20195
rect -3725 20165 -3720 20195
rect -3760 20160 -3720 20165
rect -3680 20195 -3640 20200
rect -3680 20165 -3675 20195
rect -3645 20165 -3640 20195
rect -3680 20160 -3640 20165
rect -3600 20195 -3560 20200
rect -3600 20165 -3595 20195
rect -3565 20165 -3560 20195
rect -3600 20160 -3560 20165
rect -3520 20195 -3480 20200
rect -3520 20165 -3515 20195
rect -3485 20165 -3480 20195
rect -3520 20160 -3480 20165
rect -3440 20195 -3400 20200
rect -3440 20165 -3435 20195
rect -3405 20165 -3400 20195
rect -3440 20160 -3400 20165
rect -3360 20195 -3320 20200
rect -3360 20165 -3355 20195
rect -3325 20165 -3320 20195
rect -3360 20160 -3320 20165
rect -3280 20195 -3240 20200
rect -3280 20165 -3275 20195
rect -3245 20165 -3240 20195
rect -3280 20160 -3240 20165
rect -3200 20195 -3160 20200
rect -3200 20165 -3195 20195
rect -3165 20165 -3160 20195
rect -3200 20160 -3160 20165
rect -3120 20195 -3080 20200
rect -3120 20165 -3115 20195
rect -3085 20165 -3080 20195
rect -3120 20160 -3080 20165
rect -3040 20195 -3000 20200
rect -3040 20165 -3035 20195
rect -3005 20165 -3000 20195
rect -3040 20160 -3000 20165
rect -2960 20195 -2920 20200
rect -2960 20165 -2955 20195
rect -2925 20165 -2920 20195
rect -2960 20160 -2920 20165
rect -2880 20195 -2840 20200
rect -2880 20165 -2875 20195
rect -2845 20165 -2840 20195
rect -2880 20160 -2840 20165
rect -2800 20195 -2760 20200
rect -2800 20165 -2795 20195
rect -2765 20165 -2760 20195
rect -2800 20160 -2760 20165
rect -2720 20195 -2680 20200
rect -2720 20165 -2715 20195
rect -2685 20165 -2680 20195
rect -2720 20160 -2680 20165
rect -2640 20195 -2600 20200
rect -2640 20165 -2635 20195
rect -2605 20165 -2600 20195
rect -2640 20160 -2600 20165
rect -2560 20195 -2520 20200
rect -2560 20165 -2555 20195
rect -2525 20165 -2520 20195
rect -2560 20160 -2520 20165
rect -2480 20195 -2440 20200
rect -2480 20165 -2475 20195
rect -2445 20165 -2440 20195
rect -2480 20160 -2440 20165
rect -2400 20195 -2360 20200
rect -2400 20165 -2395 20195
rect -2365 20165 -2360 20195
rect -2400 20160 -2360 20165
rect -2320 20195 -2280 20200
rect -2320 20165 -2315 20195
rect -2285 20165 -2280 20195
rect -2320 20160 -2280 20165
rect -2240 20195 -2200 20200
rect -2240 20165 -2235 20195
rect -2205 20165 -2200 20195
rect -2240 20160 -2200 20165
rect -2160 20195 -2120 20200
rect -2160 20165 -2155 20195
rect -2125 20165 -2120 20195
rect -2160 20160 -2120 20165
rect -2080 20195 -2040 20200
rect -2080 20165 -2075 20195
rect -2045 20165 -2040 20195
rect -2080 20160 -2040 20165
rect -2000 20195 -1960 20200
rect -2000 20165 -1995 20195
rect -1965 20165 -1960 20195
rect -2000 20160 -1960 20165
rect -1840 20195 -1800 20200
rect -1840 20165 -1835 20195
rect -1805 20165 -1800 20195
rect -1840 20160 -1800 20165
rect -1760 20195 -1720 20200
rect -1760 20165 -1755 20195
rect -1725 20165 -1720 20195
rect -1760 20160 -1720 20165
rect 20520 20035 20560 20040
rect 20520 20005 20525 20035
rect 20555 20005 20560 20035
rect 20520 20000 20560 20005
rect 20600 20035 20640 20040
rect 20600 20005 20605 20035
rect 20635 20005 20640 20035
rect 20600 20000 20640 20005
rect 20680 20035 20720 20040
rect 20680 20005 20685 20035
rect 20715 20005 20720 20035
rect 20680 20000 20720 20005
rect 20760 20035 20800 20040
rect 20760 20005 20765 20035
rect 20795 20005 20800 20035
rect 20760 20000 20800 20005
rect 20840 20035 20880 20040
rect 20840 20005 20845 20035
rect 20875 20005 20880 20035
rect 20840 20000 20880 20005
rect 20920 20035 20960 20040
rect 20920 20005 20925 20035
rect 20955 20005 20960 20035
rect 20920 20000 20960 20005
rect 21000 20035 21040 20040
rect 21000 20005 21005 20035
rect 21035 20005 21040 20035
rect 21000 20000 21040 20005
rect 21080 20035 21120 20040
rect 21080 20005 21085 20035
rect 21115 20005 21120 20035
rect 21080 20000 21120 20005
rect 21160 20035 21200 20040
rect 21160 20005 21165 20035
rect 21195 20005 21200 20035
rect 21160 20000 21200 20005
rect 21240 20035 21280 20040
rect 21240 20005 21245 20035
rect 21275 20005 21280 20035
rect 21240 20000 21280 20005
rect 21320 20035 21360 20040
rect 21320 20005 21325 20035
rect 21355 20005 21360 20035
rect 21320 20000 21360 20005
rect 21400 20035 21440 20040
rect 21400 20005 21405 20035
rect 21435 20005 21440 20035
rect 21400 20000 21440 20005
rect 21480 20035 21520 20040
rect 21480 20005 21485 20035
rect 21515 20005 21520 20035
rect 21480 20000 21520 20005
rect 21560 20035 21600 20040
rect 21560 20005 21565 20035
rect 21595 20005 21600 20035
rect 21560 20000 21600 20005
rect 20520 19875 20560 19880
rect 20520 19845 20525 19875
rect 20555 19845 20560 19875
rect 20520 19840 20560 19845
rect 20600 19875 20640 19880
rect 20600 19845 20605 19875
rect 20635 19845 20640 19875
rect 20600 19840 20640 19845
rect 20680 19875 20720 19880
rect 20680 19845 20685 19875
rect 20715 19845 20720 19875
rect 20680 19840 20720 19845
rect 20760 19875 20800 19880
rect 20760 19845 20765 19875
rect 20795 19845 20800 19875
rect 20760 19840 20800 19845
rect 20840 19875 20880 19880
rect 20840 19845 20845 19875
rect 20875 19845 20880 19875
rect 20840 19840 20880 19845
rect 20920 19875 20960 19880
rect 20920 19845 20925 19875
rect 20955 19845 20960 19875
rect 20920 19840 20960 19845
rect 21000 19875 21040 19880
rect 21000 19845 21005 19875
rect 21035 19845 21040 19875
rect 21000 19840 21040 19845
rect 21080 19875 21120 19880
rect 21080 19845 21085 19875
rect 21115 19845 21120 19875
rect 21080 19840 21120 19845
rect 21160 19875 21200 19880
rect 21160 19845 21165 19875
rect 21195 19845 21200 19875
rect 21160 19840 21200 19845
rect 21240 19875 21280 19880
rect 21240 19845 21245 19875
rect 21275 19845 21280 19875
rect 21240 19840 21280 19845
rect 21320 19875 21360 19880
rect 21320 19845 21325 19875
rect 21355 19845 21360 19875
rect 21320 19840 21360 19845
rect 21400 19875 21440 19880
rect 21400 19845 21405 19875
rect 21435 19845 21440 19875
rect 21400 19840 21440 19845
rect 21480 19875 21520 19880
rect 21480 19845 21485 19875
rect 21515 19845 21520 19875
rect 21480 19840 21520 19845
rect 21560 19875 21600 19880
rect 21560 19845 21565 19875
rect 21595 19845 21600 19875
rect 21560 19840 21600 19845
rect -16560 18875 -16520 18880
rect -16560 18845 -16555 18875
rect -16525 18845 -16520 18875
rect -16560 18840 -16520 18845
rect -16480 18875 -16440 18880
rect -16480 18845 -16475 18875
rect -16445 18845 -16440 18875
rect -16480 18840 -16440 18845
rect -16400 18875 -16360 18880
rect -16400 18845 -16395 18875
rect -16365 18845 -16360 18875
rect -16400 18840 -16360 18845
rect -16320 18875 -16280 18880
rect -16320 18845 -16315 18875
rect -16285 18845 -16280 18875
rect -16320 18840 -16280 18845
rect -16240 18875 -16200 18880
rect -16240 18845 -16235 18875
rect -16205 18845 -16200 18875
rect -16240 18840 -16200 18845
rect -16160 18875 -16120 18880
rect -16160 18845 -16155 18875
rect -16125 18845 -16120 18875
rect -16160 18840 -16120 18845
rect -16080 18875 -16040 18880
rect -16080 18845 -16075 18875
rect -16045 18845 -16040 18875
rect -16080 18840 -16040 18845
rect -16000 18875 -15960 18880
rect -16000 18845 -15995 18875
rect -15965 18845 -15960 18875
rect -16000 18840 -15960 18845
rect -15920 18875 -15880 18880
rect -15920 18845 -15915 18875
rect -15885 18845 -15880 18875
rect -15920 18840 -15880 18845
rect -15840 18875 -15800 18880
rect -15840 18845 -15835 18875
rect -15805 18845 -15800 18875
rect -15840 18840 -15800 18845
rect -15760 18875 -15720 18880
rect -15760 18845 -15755 18875
rect -15725 18845 -15720 18875
rect -15760 18840 -15720 18845
rect -15680 18875 -15640 18880
rect -15680 18845 -15675 18875
rect -15645 18845 -15640 18875
rect -15680 18840 -15640 18845
rect -15600 18875 -15560 18880
rect -15600 18845 -15595 18875
rect -15565 18845 -15560 18875
rect -15600 18840 -15560 18845
rect -16560 18715 -16520 18720
rect -16560 18685 -16555 18715
rect -16525 18685 -16520 18715
rect -16560 18680 -16520 18685
rect -16480 18715 -16440 18720
rect -16480 18685 -16475 18715
rect -16445 18685 -16440 18715
rect -16480 18680 -16440 18685
rect -16400 18715 -16360 18720
rect -16400 18685 -16395 18715
rect -16365 18685 -16360 18715
rect -16400 18680 -16360 18685
rect -16320 18715 -16280 18720
rect -16320 18685 -16315 18715
rect -16285 18685 -16280 18715
rect -16320 18680 -16280 18685
rect -16240 18715 -16200 18720
rect -16240 18685 -16235 18715
rect -16205 18685 -16200 18715
rect -16240 18680 -16200 18685
rect -16160 18715 -16120 18720
rect -16160 18685 -16155 18715
rect -16125 18685 -16120 18715
rect -16160 18680 -16120 18685
rect -16080 18715 -16040 18720
rect -16080 18685 -16075 18715
rect -16045 18685 -16040 18715
rect -16080 18680 -16040 18685
rect -16000 18715 -15960 18720
rect -16000 18685 -15995 18715
rect -15965 18685 -15960 18715
rect -16000 18680 -15960 18685
rect -15920 18715 -15880 18720
rect -15920 18685 -15915 18715
rect -15885 18685 -15880 18715
rect -15920 18680 -15880 18685
rect -15840 18715 -15800 18720
rect -15840 18685 -15835 18715
rect -15805 18685 -15800 18715
rect -15840 18680 -15800 18685
rect -15760 18715 -15720 18720
rect -15760 18685 -15755 18715
rect -15725 18685 -15720 18715
rect -15760 18680 -15720 18685
rect -15680 18715 -15640 18720
rect -15680 18685 -15675 18715
rect -15645 18685 -15640 18715
rect -15680 18680 -15640 18685
rect -15600 18715 -15560 18720
rect -15600 18685 -15595 18715
rect -15565 18685 -15560 18715
rect -15600 18680 -15560 18685
rect -16560 18555 -16520 18560
rect -16560 18525 -16555 18555
rect -16525 18525 -16520 18555
rect -16560 18520 -16520 18525
rect -16480 18555 -16440 18560
rect -16480 18525 -16475 18555
rect -16445 18525 -16440 18555
rect -16480 18520 -16440 18525
rect -16400 18555 -16360 18560
rect -16400 18525 -16395 18555
rect -16365 18525 -16360 18555
rect -16400 18520 -16360 18525
rect -16320 18555 -16280 18560
rect -16320 18525 -16315 18555
rect -16285 18525 -16280 18555
rect -16320 18520 -16280 18525
rect -16240 18555 -16200 18560
rect -16240 18525 -16235 18555
rect -16205 18525 -16200 18555
rect -16240 18520 -16200 18525
rect -16160 18555 -16120 18560
rect -16160 18525 -16155 18555
rect -16125 18525 -16120 18555
rect -16160 18520 -16120 18525
rect -16080 18555 -16040 18560
rect -16080 18525 -16075 18555
rect -16045 18525 -16040 18555
rect -16080 18520 -16040 18525
rect -16000 18555 -15960 18560
rect -16000 18525 -15995 18555
rect -15965 18525 -15960 18555
rect -16000 18520 -15960 18525
rect -15920 18555 -15880 18560
rect -15920 18525 -15915 18555
rect -15885 18525 -15880 18555
rect -15920 18520 -15880 18525
rect -15840 18555 -15800 18560
rect -15840 18525 -15835 18555
rect -15805 18525 -15800 18555
rect -15840 18520 -15800 18525
rect -15760 18555 -15720 18560
rect -15760 18525 -15755 18555
rect -15725 18525 -15720 18555
rect -15760 18520 -15720 18525
rect -15680 18555 -15640 18560
rect -15680 18525 -15675 18555
rect -15645 18525 -15640 18555
rect -15680 18520 -15640 18525
rect -15600 18555 -15560 18560
rect -15600 18525 -15595 18555
rect -15565 18525 -15560 18555
rect -15600 18520 -15560 18525
rect 20520 18035 20560 18040
rect 20520 18005 20525 18035
rect 20555 18005 20560 18035
rect 20520 18000 20560 18005
rect 20600 18035 20640 18040
rect 20600 18005 20605 18035
rect 20635 18005 20640 18035
rect 20600 18000 20640 18005
rect 20680 18035 20720 18040
rect 20680 18005 20685 18035
rect 20715 18005 20720 18035
rect 20680 18000 20720 18005
rect 20760 18035 20800 18040
rect 20760 18005 20765 18035
rect 20795 18005 20800 18035
rect 20760 18000 20800 18005
rect 20840 18035 20880 18040
rect 20840 18005 20845 18035
rect 20875 18005 20880 18035
rect 20840 18000 20880 18005
rect 20920 18035 20960 18040
rect 20920 18005 20925 18035
rect 20955 18005 20960 18035
rect 20920 18000 20960 18005
rect 21000 18035 21040 18040
rect 21000 18005 21005 18035
rect 21035 18005 21040 18035
rect 21000 18000 21040 18005
rect 21080 18035 21120 18040
rect 21080 18005 21085 18035
rect 21115 18005 21120 18035
rect 21080 18000 21120 18005
rect 21160 18035 21200 18040
rect 21160 18005 21165 18035
rect 21195 18005 21200 18035
rect 21160 18000 21200 18005
rect 21240 18035 21280 18040
rect 21240 18005 21245 18035
rect 21275 18005 21280 18035
rect 21240 18000 21280 18005
rect 21320 18035 21360 18040
rect 21320 18005 21325 18035
rect 21355 18005 21360 18035
rect 21320 18000 21360 18005
rect 21400 18035 21440 18040
rect 21400 18005 21405 18035
rect 21435 18005 21440 18035
rect 21400 18000 21440 18005
rect 21480 18035 21520 18040
rect 21480 18005 21485 18035
rect 21515 18005 21520 18035
rect 21480 18000 21520 18005
rect 21560 18035 21600 18040
rect 21560 18005 21565 18035
rect 21595 18005 21600 18035
rect 21560 18000 21600 18005
rect 20520 17875 20560 17880
rect 20520 17845 20525 17875
rect 20555 17845 20560 17875
rect 20520 17840 20560 17845
rect 20600 17875 20640 17880
rect 20600 17845 20605 17875
rect 20635 17845 20640 17875
rect 20600 17840 20640 17845
rect 20680 17875 20720 17880
rect 20680 17845 20685 17875
rect 20715 17845 20720 17875
rect 20680 17840 20720 17845
rect 20760 17875 20800 17880
rect 20760 17845 20765 17875
rect 20795 17845 20800 17875
rect 20760 17840 20800 17845
rect 20840 17875 20880 17880
rect 20840 17845 20845 17875
rect 20875 17845 20880 17875
rect 20840 17840 20880 17845
rect 20920 17875 20960 17880
rect 20920 17845 20925 17875
rect 20955 17845 20960 17875
rect 20920 17840 20960 17845
rect 21000 17875 21040 17880
rect 21000 17845 21005 17875
rect 21035 17845 21040 17875
rect 21000 17840 21040 17845
rect 21080 17875 21120 17880
rect 21080 17845 21085 17875
rect 21115 17845 21120 17875
rect 21080 17840 21120 17845
rect 21160 17875 21200 17880
rect 21160 17845 21165 17875
rect 21195 17845 21200 17875
rect 21160 17840 21200 17845
rect 21240 17875 21280 17880
rect 21240 17845 21245 17875
rect 21275 17845 21280 17875
rect 21240 17840 21280 17845
rect 21320 17875 21360 17880
rect 21320 17845 21325 17875
rect 21355 17845 21360 17875
rect 21320 17840 21360 17845
rect 21400 17875 21440 17880
rect 21400 17845 21405 17875
rect 21435 17845 21440 17875
rect 21400 17840 21440 17845
rect 21480 17875 21520 17880
rect 21480 17845 21485 17875
rect 21515 17845 21520 17875
rect 21480 17840 21520 17845
rect 21560 17875 21600 17880
rect 21560 17845 21565 17875
rect 21595 17845 21600 17875
rect 21560 17840 21600 17845
rect -16560 17355 -16520 17360
rect -16560 17325 -16555 17355
rect -16525 17325 -16520 17355
rect -16560 17320 -16520 17325
rect -16480 17355 -16440 17360
rect -16480 17325 -16475 17355
rect -16445 17325 -16440 17355
rect -16480 17320 -16440 17325
rect -16400 17355 -16360 17360
rect -16400 17325 -16395 17355
rect -16365 17325 -16360 17355
rect -16400 17320 -16360 17325
rect -16320 17355 -16280 17360
rect -16320 17325 -16315 17355
rect -16285 17325 -16280 17355
rect -16320 17320 -16280 17325
rect -16240 17355 -16200 17360
rect -16240 17325 -16235 17355
rect -16205 17325 -16200 17355
rect -16240 17320 -16200 17325
rect -16160 17355 -16120 17360
rect -16160 17325 -16155 17355
rect -16125 17325 -16120 17355
rect -16160 17320 -16120 17325
rect -16080 17355 -16040 17360
rect -16080 17325 -16075 17355
rect -16045 17325 -16040 17355
rect -16080 17320 -16040 17325
rect -16000 17355 -15960 17360
rect -16000 17325 -15995 17355
rect -15965 17325 -15960 17355
rect -16000 17320 -15960 17325
rect -15920 17355 -15880 17360
rect -15920 17325 -15915 17355
rect -15885 17325 -15880 17355
rect -15920 17320 -15880 17325
rect -15840 17355 -15800 17360
rect -15840 17325 -15835 17355
rect -15805 17325 -15800 17355
rect -15840 17320 -15800 17325
rect -15760 17355 -15720 17360
rect -15760 17325 -15755 17355
rect -15725 17325 -15720 17355
rect -15760 17320 -15720 17325
rect -15680 17355 -15640 17360
rect -15680 17325 -15675 17355
rect -15645 17325 -15640 17355
rect -15680 17320 -15640 17325
rect -15600 17355 -15560 17360
rect -15600 17325 -15595 17355
rect -15565 17325 -15560 17355
rect -15600 17320 -15560 17325
rect -14960 17355 -14920 17360
rect -14960 17325 -14955 17355
rect -14925 17325 -14920 17355
rect -14960 17320 -14920 17325
rect -14880 17355 -14840 17360
rect -14880 17325 -14875 17355
rect -14845 17325 -14840 17355
rect -14880 17320 -14840 17325
rect -14800 17355 -14760 17360
rect -14800 17325 -14795 17355
rect -14765 17325 -14760 17355
rect -14800 17320 -14760 17325
rect -14720 17355 -14680 17360
rect -14720 17325 -14715 17355
rect -14685 17325 -14680 17355
rect -14720 17320 -14680 17325
rect -14640 17355 -14600 17360
rect -14640 17325 -14635 17355
rect -14605 17325 -14600 17355
rect -14640 17320 -14600 17325
rect -14560 17355 -14520 17360
rect -14560 17325 -14555 17355
rect -14525 17325 -14520 17355
rect -14560 17320 -14520 17325
rect -14480 17355 -14440 17360
rect -14480 17325 -14475 17355
rect -14445 17325 -14440 17355
rect -14480 17320 -14440 17325
rect -14400 17355 -14360 17360
rect -14400 17325 -14395 17355
rect -14365 17325 -14360 17355
rect -14400 17320 -14360 17325
rect -14320 17355 -14280 17360
rect -14320 17325 -14315 17355
rect -14285 17325 -14280 17355
rect -14320 17320 -14280 17325
rect -14240 17355 -14200 17360
rect -14240 17325 -14235 17355
rect -14205 17325 -14200 17355
rect -14240 17320 -14200 17325
rect -14160 17355 -14120 17360
rect -14160 17325 -14155 17355
rect -14125 17325 -14120 17355
rect -14160 17320 -14120 17325
rect -14080 17355 -14040 17360
rect -14080 17325 -14075 17355
rect -14045 17325 -14040 17355
rect -14080 17320 -14040 17325
rect -14000 17355 -13960 17360
rect -14000 17325 -13995 17355
rect -13965 17325 -13960 17355
rect -14000 17320 -13960 17325
rect -13920 17355 -13880 17360
rect -13920 17325 -13915 17355
rect -13885 17325 -13880 17355
rect -13920 17320 -13880 17325
rect -13840 17355 -13800 17360
rect -13840 17325 -13835 17355
rect -13805 17325 -13800 17355
rect -13840 17320 -13800 17325
rect -13760 17355 -13720 17360
rect -13760 17325 -13755 17355
rect -13725 17325 -13720 17355
rect -13760 17320 -13720 17325
rect -13680 17355 -13640 17360
rect -13680 17325 -13675 17355
rect -13645 17325 -13640 17355
rect -13680 17320 -13640 17325
rect -13600 17355 -13560 17360
rect -13600 17325 -13595 17355
rect -13565 17325 -13560 17355
rect -13600 17320 -13560 17325
rect -13520 17355 -13480 17360
rect -13520 17325 -13515 17355
rect -13485 17325 -13480 17355
rect -13520 17320 -13480 17325
rect -13440 17355 -13400 17360
rect -13440 17325 -13435 17355
rect -13405 17325 -13400 17355
rect -13440 17320 -13400 17325
rect -13360 17355 -13320 17360
rect -13360 17325 -13355 17355
rect -13325 17325 -13320 17355
rect -13360 17320 -13320 17325
rect -13280 17355 -13240 17360
rect -13280 17325 -13275 17355
rect -13245 17325 -13240 17355
rect -13280 17320 -13240 17325
rect -13200 17355 -13160 17360
rect -13200 17325 -13195 17355
rect -13165 17325 -13160 17355
rect -13200 17320 -13160 17325
rect -13120 17355 -13080 17360
rect -13120 17325 -13115 17355
rect -13085 17325 -13080 17355
rect -13120 17320 -13080 17325
rect -13040 17355 -13000 17360
rect -13040 17325 -13035 17355
rect -13005 17325 -13000 17355
rect -13040 17320 -13000 17325
rect -12960 17355 -12920 17360
rect -12960 17325 -12955 17355
rect -12925 17325 -12920 17355
rect -12960 17320 -12920 17325
rect -12880 17355 -12840 17360
rect -12880 17325 -12875 17355
rect -12845 17325 -12840 17355
rect -12880 17320 -12840 17325
rect -12800 17355 -12760 17360
rect -12800 17325 -12795 17355
rect -12765 17325 -12760 17355
rect -12800 17320 -12760 17325
rect -12720 17355 -12680 17360
rect -12720 17325 -12715 17355
rect -12685 17325 -12680 17355
rect -12720 17320 -12680 17325
rect -12640 17355 -12600 17360
rect -12640 17325 -12635 17355
rect -12605 17325 -12600 17355
rect -12640 17320 -12600 17325
rect -12560 17355 -12520 17360
rect -12560 17325 -12555 17355
rect -12525 17325 -12520 17355
rect -12560 17320 -12520 17325
rect -12480 17355 -12440 17360
rect -12480 17325 -12475 17355
rect -12445 17325 -12440 17355
rect -12480 17320 -12440 17325
rect -12400 17355 -12360 17360
rect -12400 17325 -12395 17355
rect -12365 17325 -12360 17355
rect -12400 17320 -12360 17325
rect -12320 17355 -12280 17360
rect -12320 17325 -12315 17355
rect -12285 17325 -12280 17355
rect -12320 17320 -12280 17325
rect -12240 17355 -12200 17360
rect -12240 17325 -12235 17355
rect -12205 17325 -12200 17355
rect -12240 17320 -12200 17325
rect -12160 17355 -12120 17360
rect -12160 17325 -12155 17355
rect -12125 17325 -12120 17355
rect -12160 17320 -12120 17325
rect -12080 17355 -12040 17360
rect -12080 17325 -12075 17355
rect -12045 17325 -12040 17355
rect -12080 17320 -12040 17325
rect -12000 17355 -11960 17360
rect -12000 17325 -11995 17355
rect -11965 17325 -11960 17355
rect -12000 17320 -11960 17325
rect -11920 17355 -11880 17360
rect -11920 17325 -11915 17355
rect -11885 17325 -11880 17355
rect -11920 17320 -11880 17325
rect -11840 17355 -11800 17360
rect -11840 17325 -11835 17355
rect -11805 17325 -11800 17355
rect -11840 17320 -11800 17325
rect -11760 17355 -11720 17360
rect -11760 17325 -11755 17355
rect -11725 17325 -11720 17355
rect -11760 17320 -11720 17325
rect -11680 17355 -11640 17360
rect -11680 17325 -11675 17355
rect -11645 17325 -11640 17355
rect -11680 17320 -11640 17325
rect -11600 17355 -11560 17360
rect -11600 17325 -11595 17355
rect -11565 17325 -11560 17355
rect -11600 17320 -11560 17325
rect -11520 17355 -11480 17360
rect -11520 17325 -11515 17355
rect -11485 17325 -11480 17355
rect -11520 17320 -11480 17325
rect -11440 17355 -11400 17360
rect -11440 17325 -11435 17355
rect -11405 17325 -11400 17355
rect -11440 17320 -11400 17325
rect -11360 17355 -11320 17360
rect -11360 17325 -11355 17355
rect -11325 17325 -11320 17355
rect -11360 17320 -11320 17325
rect -11280 17355 -11240 17360
rect -11280 17325 -11275 17355
rect -11245 17325 -11240 17355
rect -11280 17320 -11240 17325
rect -11200 17355 -11160 17360
rect -11200 17325 -11195 17355
rect -11165 17325 -11160 17355
rect -11200 17320 -11160 17325
rect -11120 17355 -11080 17360
rect -11120 17325 -11115 17355
rect -11085 17325 -11080 17355
rect -11120 17320 -11080 17325
rect -11040 17355 -11000 17360
rect -11040 17325 -11035 17355
rect -11005 17325 -11000 17355
rect -11040 17320 -11000 17325
rect -10960 17355 -10920 17360
rect -10960 17325 -10955 17355
rect -10925 17325 -10920 17355
rect -10960 17320 -10920 17325
rect -10880 17355 -10840 17360
rect -10880 17325 -10875 17355
rect -10845 17325 -10840 17355
rect -10880 17320 -10840 17325
rect -10800 17355 -10760 17360
rect -10800 17325 -10795 17355
rect -10765 17325 -10760 17355
rect -10800 17320 -10760 17325
rect -10720 17355 -10680 17360
rect -10720 17325 -10715 17355
rect -10685 17325 -10680 17355
rect -10720 17320 -10680 17325
rect -10640 17355 -10600 17360
rect -10640 17325 -10635 17355
rect -10605 17325 -10600 17355
rect -10640 17320 -10600 17325
rect -10560 17355 -10520 17360
rect -10560 17325 -10555 17355
rect -10525 17325 -10520 17355
rect -10560 17320 -10520 17325
rect -10480 17355 -10440 17360
rect -10480 17325 -10475 17355
rect -10445 17325 -10440 17355
rect -10480 17320 -10440 17325
rect -10400 17355 -10360 17360
rect -10400 17325 -10395 17355
rect -10365 17325 -10360 17355
rect -10400 17320 -10360 17325
rect -10320 17355 -10280 17360
rect -10320 17325 -10315 17355
rect -10285 17325 -10280 17355
rect -10320 17320 -10280 17325
rect -10240 17355 -10200 17360
rect -10240 17325 -10235 17355
rect -10205 17325 -10200 17355
rect -10240 17320 -10200 17325
rect -10160 17355 -10120 17360
rect -10160 17325 -10155 17355
rect -10125 17325 -10120 17355
rect -10160 17320 -10120 17325
rect -10080 17355 -10040 17360
rect -10080 17325 -10075 17355
rect -10045 17325 -10040 17355
rect -10080 17320 -10040 17325
rect -10000 17355 -9960 17360
rect -10000 17325 -9995 17355
rect -9965 17325 -9960 17355
rect -10000 17320 -9960 17325
rect -9920 17355 -9880 17360
rect -9920 17325 -9915 17355
rect -9885 17325 -9880 17355
rect -9920 17320 -9880 17325
rect -9840 17355 -9800 17360
rect -9840 17325 -9835 17355
rect -9805 17325 -9800 17355
rect -9840 17320 -9800 17325
rect -9760 17355 -9720 17360
rect -9760 17325 -9755 17355
rect -9725 17325 -9720 17355
rect -9760 17320 -9720 17325
rect -9680 17355 -9640 17360
rect -9680 17325 -9675 17355
rect -9645 17325 -9640 17355
rect -9680 17320 -9640 17325
rect -9600 17355 -9560 17360
rect -9600 17325 -9595 17355
rect -9565 17325 -9560 17355
rect -9600 17320 -9560 17325
rect -9520 17355 -9480 17360
rect -9520 17325 -9515 17355
rect -9485 17325 -9480 17355
rect -9520 17320 -9480 17325
rect -9440 17355 -9400 17360
rect -9440 17325 -9435 17355
rect -9405 17325 -9400 17355
rect -9440 17320 -9400 17325
rect -9360 17355 -9320 17360
rect -9360 17325 -9355 17355
rect -9325 17325 -9320 17355
rect -9360 17320 -9320 17325
rect -9280 17355 -9240 17360
rect -9280 17325 -9275 17355
rect -9245 17325 -9240 17355
rect -9280 17320 -9240 17325
rect -9200 17355 -9160 17360
rect -9200 17325 -9195 17355
rect -9165 17325 -9160 17355
rect -9200 17320 -9160 17325
rect -9120 17355 -9080 17360
rect -9120 17325 -9115 17355
rect -9085 17325 -9080 17355
rect -9120 17320 -9080 17325
rect -9040 17355 -9000 17360
rect -9040 17325 -9035 17355
rect -9005 17325 -9000 17355
rect -9040 17320 -9000 17325
rect -8960 17355 -8920 17360
rect -8960 17325 -8955 17355
rect -8925 17325 -8920 17355
rect -8960 17320 -8920 17325
rect -8880 17355 -8840 17360
rect -8880 17325 -8875 17355
rect -8845 17325 -8840 17355
rect -8880 17320 -8840 17325
rect -8800 17355 -8760 17360
rect -8800 17325 -8795 17355
rect -8765 17325 -8760 17355
rect -8800 17320 -8760 17325
rect -8720 17355 -8680 17360
rect -8720 17325 -8715 17355
rect -8685 17325 -8680 17355
rect -8720 17320 -8680 17325
rect -8640 17355 -8600 17360
rect -8640 17325 -8635 17355
rect -8605 17325 -8600 17355
rect -8640 17320 -8600 17325
rect -8560 17355 -8520 17360
rect -8560 17325 -8555 17355
rect -8525 17325 -8520 17355
rect -8560 17320 -8520 17325
rect -8480 17355 -8440 17360
rect -8480 17325 -8475 17355
rect -8445 17325 -8440 17355
rect -8480 17320 -8440 17325
rect -8400 17355 -8360 17360
rect -8400 17325 -8395 17355
rect -8365 17325 -8360 17355
rect -8400 17320 -8360 17325
rect -8320 17355 -8280 17360
rect -8320 17325 -8315 17355
rect -8285 17325 -8280 17355
rect -8320 17320 -8280 17325
rect -8240 17355 -8200 17360
rect -8240 17325 -8235 17355
rect -8205 17325 -8200 17355
rect -8240 17320 -8200 17325
rect -8160 17355 -8120 17360
rect -8160 17325 -8155 17355
rect -8125 17325 -8120 17355
rect -8160 17320 -8120 17325
rect -8080 17355 -8040 17360
rect -8080 17325 -8075 17355
rect -8045 17325 -8040 17355
rect -8080 17320 -8040 17325
rect -8000 17355 -7960 17360
rect -8000 17325 -7995 17355
rect -7965 17325 -7960 17355
rect -8000 17320 -7960 17325
rect -7920 17355 -7880 17360
rect -7920 17325 -7915 17355
rect -7885 17325 -7880 17355
rect -7920 17320 -7880 17325
rect -7840 17355 -7800 17360
rect -7840 17325 -7835 17355
rect -7805 17325 -7800 17355
rect -7840 17320 -7800 17325
rect -7760 17355 -7720 17360
rect -7760 17325 -7755 17355
rect -7725 17325 -7720 17355
rect -7760 17320 -7720 17325
rect -7680 17355 -7640 17360
rect -7680 17325 -7675 17355
rect -7645 17325 -7640 17355
rect -7680 17320 -7640 17325
rect -7600 17355 -7560 17360
rect -7600 17325 -7595 17355
rect -7565 17325 -7560 17355
rect -7600 17320 -7560 17325
rect -7520 17355 -7480 17360
rect -7520 17325 -7515 17355
rect -7485 17325 -7480 17355
rect -7520 17320 -7480 17325
rect -7440 17355 -7400 17360
rect -7440 17325 -7435 17355
rect -7405 17325 -7400 17355
rect -7440 17320 -7400 17325
rect -7360 17355 -7320 17360
rect -7360 17325 -7355 17355
rect -7325 17325 -7320 17355
rect -7360 17320 -7320 17325
rect -7280 17355 -7240 17360
rect -7280 17325 -7275 17355
rect -7245 17325 -7240 17355
rect -7280 17320 -7240 17325
rect -7200 17355 -7160 17360
rect -7200 17325 -7195 17355
rect -7165 17325 -7160 17355
rect -7200 17320 -7160 17325
rect -7120 17355 -7080 17360
rect -7120 17325 -7115 17355
rect -7085 17325 -7080 17355
rect -7120 17320 -7080 17325
rect -7040 17355 -7000 17360
rect -7040 17325 -7035 17355
rect -7005 17325 -7000 17355
rect -7040 17320 -7000 17325
rect -6960 17355 -6920 17360
rect -6960 17325 -6955 17355
rect -6925 17325 -6920 17355
rect -6960 17320 -6920 17325
rect -6880 17355 -6840 17360
rect -6880 17325 -6875 17355
rect -6845 17325 -6840 17355
rect -6880 17320 -6840 17325
rect -6800 17355 -6760 17360
rect -6800 17325 -6795 17355
rect -6765 17325 -6760 17355
rect -6800 17320 -6760 17325
rect -6720 17355 -6680 17360
rect -6720 17325 -6715 17355
rect -6685 17325 -6680 17355
rect -6720 17320 -6680 17325
rect -6640 17355 -6600 17360
rect -6640 17325 -6635 17355
rect -6605 17325 -6600 17355
rect -6640 17320 -6600 17325
rect -6560 17355 -6520 17360
rect -6560 17325 -6555 17355
rect -6525 17325 -6520 17355
rect -6560 17320 -6520 17325
rect -6480 17355 -6440 17360
rect -6480 17325 -6475 17355
rect -6445 17325 -6440 17355
rect -6480 17320 -6440 17325
rect -6400 17355 -6360 17360
rect -6400 17325 -6395 17355
rect -6365 17325 -6360 17355
rect -6400 17320 -6360 17325
rect -6320 17355 -6280 17360
rect -6320 17325 -6315 17355
rect -6285 17325 -6280 17355
rect -6320 17320 -6280 17325
rect -6240 17355 -6200 17360
rect -6240 17325 -6235 17355
rect -6205 17325 -6200 17355
rect -6240 17320 -6200 17325
rect -6160 17355 -6120 17360
rect -6160 17325 -6155 17355
rect -6125 17325 -6120 17355
rect -6160 17320 -6120 17325
rect -6080 17355 -6040 17360
rect -6080 17325 -6075 17355
rect -6045 17325 -6040 17355
rect -6080 17320 -6040 17325
rect -6000 17355 -5960 17360
rect -6000 17325 -5995 17355
rect -5965 17325 -5960 17355
rect -6000 17320 -5960 17325
rect -5920 17355 -5880 17360
rect -5920 17325 -5915 17355
rect -5885 17325 -5880 17355
rect -5920 17320 -5880 17325
rect -5840 17355 -5800 17360
rect -5840 17325 -5835 17355
rect -5805 17325 -5800 17355
rect -5840 17320 -5800 17325
rect -5760 17355 -5720 17360
rect -5760 17325 -5755 17355
rect -5725 17325 -5720 17355
rect -5760 17320 -5720 17325
rect -5440 17355 -5400 17360
rect -5440 17325 -5435 17355
rect -5405 17325 -5400 17355
rect -5440 17320 -5400 17325
rect -5280 17355 -5240 17360
rect -5280 17325 -5275 17355
rect -5245 17325 -5240 17355
rect -5280 17320 -5240 17325
rect -16560 17195 -16520 17200
rect -16560 17165 -16555 17195
rect -16525 17165 -16520 17195
rect -16560 17160 -16520 17165
rect -16480 17195 -16440 17200
rect -16480 17165 -16475 17195
rect -16445 17165 -16440 17195
rect -16480 17160 -16440 17165
rect -16400 17195 -16360 17200
rect -16400 17165 -16395 17195
rect -16365 17165 -16360 17195
rect -16400 17160 -16360 17165
rect -16320 17195 -16280 17200
rect -16320 17165 -16315 17195
rect -16285 17165 -16280 17195
rect -16320 17160 -16280 17165
rect -16240 17195 -16200 17200
rect -16240 17165 -16235 17195
rect -16205 17165 -16200 17195
rect -16240 17160 -16200 17165
rect -16160 17195 -16120 17200
rect -16160 17165 -16155 17195
rect -16125 17165 -16120 17195
rect -16160 17160 -16120 17165
rect -16080 17195 -16040 17200
rect -16080 17165 -16075 17195
rect -16045 17165 -16040 17195
rect -16080 17160 -16040 17165
rect -16000 17195 -15960 17200
rect -16000 17165 -15995 17195
rect -15965 17165 -15960 17195
rect -16000 17160 -15960 17165
rect -15920 17195 -15880 17200
rect -15920 17165 -15915 17195
rect -15885 17165 -15880 17195
rect -15920 17160 -15880 17165
rect -15840 17195 -15800 17200
rect -15840 17165 -15835 17195
rect -15805 17165 -15800 17195
rect -15840 17160 -15800 17165
rect -15760 17195 -15720 17200
rect -15760 17165 -15755 17195
rect -15725 17165 -15720 17195
rect -15760 17160 -15720 17165
rect -15680 17195 -15640 17200
rect -15680 17165 -15675 17195
rect -15645 17165 -15640 17195
rect -15680 17160 -15640 17165
rect -15600 17195 -15560 17200
rect -15600 17165 -15595 17195
rect -15565 17165 -15560 17195
rect -15600 17160 -15560 17165
rect -14960 17195 -14920 17200
rect -14960 17165 -14955 17195
rect -14925 17165 -14920 17195
rect -14960 17160 -14920 17165
rect -14880 17195 -14840 17200
rect -14880 17165 -14875 17195
rect -14845 17165 -14840 17195
rect -14880 17160 -14840 17165
rect -14800 17195 -14760 17200
rect -14800 17165 -14795 17195
rect -14765 17165 -14760 17195
rect -14800 17160 -14760 17165
rect -14720 17195 -14680 17200
rect -14720 17165 -14715 17195
rect -14685 17165 -14680 17195
rect -14720 17160 -14680 17165
rect -14640 17195 -14600 17200
rect -14640 17165 -14635 17195
rect -14605 17165 -14600 17195
rect -14640 17160 -14600 17165
rect -14560 17195 -14520 17200
rect -14560 17165 -14555 17195
rect -14525 17165 -14520 17195
rect -14560 17160 -14520 17165
rect -14480 17195 -14440 17200
rect -14480 17165 -14475 17195
rect -14445 17165 -14440 17195
rect -14480 17160 -14440 17165
rect -14400 17195 -14360 17200
rect -14400 17165 -14395 17195
rect -14365 17165 -14360 17195
rect -14400 17160 -14360 17165
rect -14320 17195 -14280 17200
rect -14320 17165 -14315 17195
rect -14285 17165 -14280 17195
rect -14320 17160 -14280 17165
rect -14240 17195 -14200 17200
rect -14240 17165 -14235 17195
rect -14205 17165 -14200 17195
rect -14240 17160 -14200 17165
rect -14160 17195 -14120 17200
rect -14160 17165 -14155 17195
rect -14125 17165 -14120 17195
rect -14160 17160 -14120 17165
rect -14080 17195 -14040 17200
rect -14080 17165 -14075 17195
rect -14045 17165 -14040 17195
rect -14080 17160 -14040 17165
rect -14000 17195 -13960 17200
rect -14000 17165 -13995 17195
rect -13965 17165 -13960 17195
rect -14000 17160 -13960 17165
rect -13920 17195 -13880 17200
rect -13920 17165 -13915 17195
rect -13885 17165 -13880 17195
rect -13920 17160 -13880 17165
rect -13840 17195 -13800 17200
rect -13840 17165 -13835 17195
rect -13805 17165 -13800 17195
rect -13840 17160 -13800 17165
rect -13760 17195 -13720 17200
rect -13760 17165 -13755 17195
rect -13725 17165 -13720 17195
rect -13760 17160 -13720 17165
rect -13680 17195 -13640 17200
rect -13680 17165 -13675 17195
rect -13645 17165 -13640 17195
rect -13680 17160 -13640 17165
rect -13600 17195 -13560 17200
rect -13600 17165 -13595 17195
rect -13565 17165 -13560 17195
rect -13600 17160 -13560 17165
rect -13520 17195 -13480 17200
rect -13520 17165 -13515 17195
rect -13485 17165 -13480 17195
rect -13520 17160 -13480 17165
rect -13440 17195 -13400 17200
rect -13440 17165 -13435 17195
rect -13405 17165 -13400 17195
rect -13440 17160 -13400 17165
rect -13360 17195 -13320 17200
rect -13360 17165 -13355 17195
rect -13325 17165 -13320 17195
rect -13360 17160 -13320 17165
rect -13280 17195 -13240 17200
rect -13280 17165 -13275 17195
rect -13245 17165 -13240 17195
rect -13280 17160 -13240 17165
rect -13200 17195 -13160 17200
rect -13200 17165 -13195 17195
rect -13165 17165 -13160 17195
rect -13200 17160 -13160 17165
rect -13120 17195 -13080 17200
rect -13120 17165 -13115 17195
rect -13085 17165 -13080 17195
rect -13120 17160 -13080 17165
rect -13040 17195 -13000 17200
rect -13040 17165 -13035 17195
rect -13005 17165 -13000 17195
rect -13040 17160 -13000 17165
rect -12960 17195 -12920 17200
rect -12960 17165 -12955 17195
rect -12925 17165 -12920 17195
rect -12960 17160 -12920 17165
rect -12880 17195 -12840 17200
rect -12880 17165 -12875 17195
rect -12845 17165 -12840 17195
rect -12880 17160 -12840 17165
rect -12800 17195 -12760 17200
rect -12800 17165 -12795 17195
rect -12765 17165 -12760 17195
rect -12800 17160 -12760 17165
rect -12720 17195 -12680 17200
rect -12720 17165 -12715 17195
rect -12685 17165 -12680 17195
rect -12720 17160 -12680 17165
rect -12640 17195 -12600 17200
rect -12640 17165 -12635 17195
rect -12605 17165 -12600 17195
rect -12640 17160 -12600 17165
rect -12560 17195 -12520 17200
rect -12560 17165 -12555 17195
rect -12525 17165 -12520 17195
rect -12560 17160 -12520 17165
rect -12480 17195 -12440 17200
rect -12480 17165 -12475 17195
rect -12445 17165 -12440 17195
rect -12480 17160 -12440 17165
rect -12400 17195 -12360 17200
rect -12400 17165 -12395 17195
rect -12365 17165 -12360 17195
rect -12400 17160 -12360 17165
rect -12320 17195 -12280 17200
rect -12320 17165 -12315 17195
rect -12285 17165 -12280 17195
rect -12320 17160 -12280 17165
rect -12240 17195 -12200 17200
rect -12240 17165 -12235 17195
rect -12205 17165 -12200 17195
rect -12240 17160 -12200 17165
rect -12160 17195 -12120 17200
rect -12160 17165 -12155 17195
rect -12125 17165 -12120 17195
rect -12160 17160 -12120 17165
rect -12080 17195 -12040 17200
rect -12080 17165 -12075 17195
rect -12045 17165 -12040 17195
rect -12080 17160 -12040 17165
rect -12000 17195 -11960 17200
rect -12000 17165 -11995 17195
rect -11965 17165 -11960 17195
rect -12000 17160 -11960 17165
rect -11920 17195 -11880 17200
rect -11920 17165 -11915 17195
rect -11885 17165 -11880 17195
rect -11920 17160 -11880 17165
rect -11840 17195 -11800 17200
rect -11840 17165 -11835 17195
rect -11805 17165 -11800 17195
rect -11840 17160 -11800 17165
rect -11760 17195 -11720 17200
rect -11760 17165 -11755 17195
rect -11725 17165 -11720 17195
rect -11760 17160 -11720 17165
rect -11680 17195 -11640 17200
rect -11680 17165 -11675 17195
rect -11645 17165 -11640 17195
rect -11680 17160 -11640 17165
rect -11600 17195 -11560 17200
rect -11600 17165 -11595 17195
rect -11565 17165 -11560 17195
rect -11600 17160 -11560 17165
rect -11520 17195 -11480 17200
rect -11520 17165 -11515 17195
rect -11485 17165 -11480 17195
rect -11520 17160 -11480 17165
rect -11440 17195 -11400 17200
rect -11440 17165 -11435 17195
rect -11405 17165 -11400 17195
rect -11440 17160 -11400 17165
rect -11360 17195 -11320 17200
rect -11360 17165 -11355 17195
rect -11325 17165 -11320 17195
rect -11360 17160 -11320 17165
rect -11280 17195 -11240 17200
rect -11280 17165 -11275 17195
rect -11245 17165 -11240 17195
rect -11280 17160 -11240 17165
rect -11200 17195 -11160 17200
rect -11200 17165 -11195 17195
rect -11165 17165 -11160 17195
rect -11200 17160 -11160 17165
rect -11120 17195 -11080 17200
rect -11120 17165 -11115 17195
rect -11085 17165 -11080 17195
rect -11120 17160 -11080 17165
rect -11040 17195 -11000 17200
rect -11040 17165 -11035 17195
rect -11005 17165 -11000 17195
rect -11040 17160 -11000 17165
rect -10960 17195 -10920 17200
rect -10960 17165 -10955 17195
rect -10925 17165 -10920 17195
rect -10960 17160 -10920 17165
rect -10880 17195 -10840 17200
rect -10880 17165 -10875 17195
rect -10845 17165 -10840 17195
rect -10880 17160 -10840 17165
rect -10800 17195 -10760 17200
rect -10800 17165 -10795 17195
rect -10765 17165 -10760 17195
rect -10800 17160 -10760 17165
rect -10720 17195 -10680 17200
rect -10720 17165 -10715 17195
rect -10685 17165 -10680 17195
rect -10720 17160 -10680 17165
rect -10640 17195 -10600 17200
rect -10640 17165 -10635 17195
rect -10605 17165 -10600 17195
rect -10640 17160 -10600 17165
rect -10560 17195 -10520 17200
rect -10560 17165 -10555 17195
rect -10525 17165 -10520 17195
rect -10560 17160 -10520 17165
rect -10480 17195 -10440 17200
rect -10480 17165 -10475 17195
rect -10445 17165 -10440 17195
rect -10480 17160 -10440 17165
rect -10400 17195 -10360 17200
rect -10400 17165 -10395 17195
rect -10365 17165 -10360 17195
rect -10400 17160 -10360 17165
rect -10320 17195 -10280 17200
rect -10320 17165 -10315 17195
rect -10285 17165 -10280 17195
rect -10320 17160 -10280 17165
rect -10240 17195 -10200 17200
rect -10240 17165 -10235 17195
rect -10205 17165 -10200 17195
rect -10240 17160 -10200 17165
rect -10160 17195 -10120 17200
rect -10160 17165 -10155 17195
rect -10125 17165 -10120 17195
rect -10160 17160 -10120 17165
rect -10080 17195 -10040 17200
rect -10080 17165 -10075 17195
rect -10045 17165 -10040 17195
rect -10080 17160 -10040 17165
rect -10000 17195 -9960 17200
rect -10000 17165 -9995 17195
rect -9965 17165 -9960 17195
rect -10000 17160 -9960 17165
rect -9920 17195 -9880 17200
rect -9920 17165 -9915 17195
rect -9885 17165 -9880 17195
rect -9920 17160 -9880 17165
rect -9840 17195 -9800 17200
rect -9840 17165 -9835 17195
rect -9805 17165 -9800 17195
rect -9840 17160 -9800 17165
rect -9760 17195 -9720 17200
rect -9760 17165 -9755 17195
rect -9725 17165 -9720 17195
rect -9760 17160 -9720 17165
rect -9680 17195 -9640 17200
rect -9680 17165 -9675 17195
rect -9645 17165 -9640 17195
rect -9680 17160 -9640 17165
rect -9600 17195 -9560 17200
rect -9600 17165 -9595 17195
rect -9565 17165 -9560 17195
rect -9600 17160 -9560 17165
rect -9520 17195 -9480 17200
rect -9520 17165 -9515 17195
rect -9485 17165 -9480 17195
rect -9520 17160 -9480 17165
rect -9440 17195 -9400 17200
rect -9440 17165 -9435 17195
rect -9405 17165 -9400 17195
rect -9440 17160 -9400 17165
rect -9360 17195 -9320 17200
rect -9360 17165 -9355 17195
rect -9325 17165 -9320 17195
rect -9360 17160 -9320 17165
rect -9280 17195 -9240 17200
rect -9280 17165 -9275 17195
rect -9245 17165 -9240 17195
rect -9280 17160 -9240 17165
rect -9200 17195 -9160 17200
rect -9200 17165 -9195 17195
rect -9165 17165 -9160 17195
rect -9200 17160 -9160 17165
rect -9120 17195 -9080 17200
rect -9120 17165 -9115 17195
rect -9085 17165 -9080 17195
rect -9120 17160 -9080 17165
rect -9040 17195 -9000 17200
rect -9040 17165 -9035 17195
rect -9005 17165 -9000 17195
rect -9040 17160 -9000 17165
rect -8960 17195 -8920 17200
rect -8960 17165 -8955 17195
rect -8925 17165 -8920 17195
rect -8960 17160 -8920 17165
rect -8880 17195 -8840 17200
rect -8880 17165 -8875 17195
rect -8845 17165 -8840 17195
rect -8880 17160 -8840 17165
rect -8800 17195 -8760 17200
rect -8800 17165 -8795 17195
rect -8765 17165 -8760 17195
rect -8800 17160 -8760 17165
rect -8720 17195 -8680 17200
rect -8720 17165 -8715 17195
rect -8685 17165 -8680 17195
rect -8720 17160 -8680 17165
rect -8640 17195 -8600 17200
rect -8640 17165 -8635 17195
rect -8605 17165 -8600 17195
rect -8640 17160 -8600 17165
rect -8560 17195 -8520 17200
rect -8560 17165 -8555 17195
rect -8525 17165 -8520 17195
rect -8560 17160 -8520 17165
rect -8480 17195 -8440 17200
rect -8480 17165 -8475 17195
rect -8445 17165 -8440 17195
rect -8480 17160 -8440 17165
rect -8400 17195 -8360 17200
rect -8400 17165 -8395 17195
rect -8365 17165 -8360 17195
rect -8400 17160 -8360 17165
rect -8320 17195 -8280 17200
rect -8320 17165 -8315 17195
rect -8285 17165 -8280 17195
rect -8320 17160 -8280 17165
rect -8240 17195 -8200 17200
rect -8240 17165 -8235 17195
rect -8205 17165 -8200 17195
rect -8240 17160 -8200 17165
rect -8160 17195 -8120 17200
rect -8160 17165 -8155 17195
rect -8125 17165 -8120 17195
rect -8160 17160 -8120 17165
rect -8080 17195 -8040 17200
rect -8080 17165 -8075 17195
rect -8045 17165 -8040 17195
rect -8080 17160 -8040 17165
rect -8000 17195 -7960 17200
rect -8000 17165 -7995 17195
rect -7965 17165 -7960 17195
rect -8000 17160 -7960 17165
rect -7920 17195 -7880 17200
rect -7920 17165 -7915 17195
rect -7885 17165 -7880 17195
rect -7920 17160 -7880 17165
rect -7840 17195 -7800 17200
rect -7840 17165 -7835 17195
rect -7805 17165 -7800 17195
rect -7840 17160 -7800 17165
rect -7760 17195 -7720 17200
rect -7760 17165 -7755 17195
rect -7725 17165 -7720 17195
rect -7760 17160 -7720 17165
rect -7680 17195 -7640 17200
rect -7680 17165 -7675 17195
rect -7645 17165 -7640 17195
rect -7680 17160 -7640 17165
rect -7600 17195 -7560 17200
rect -7600 17165 -7595 17195
rect -7565 17165 -7560 17195
rect -7600 17160 -7560 17165
rect -7520 17195 -7480 17200
rect -7520 17165 -7515 17195
rect -7485 17165 -7480 17195
rect -7520 17160 -7480 17165
rect -7440 17195 -7400 17200
rect -7440 17165 -7435 17195
rect -7405 17165 -7400 17195
rect -7440 17160 -7400 17165
rect -7360 17195 -7320 17200
rect -7360 17165 -7355 17195
rect -7325 17165 -7320 17195
rect -7360 17160 -7320 17165
rect -7280 17195 -7240 17200
rect -7280 17165 -7275 17195
rect -7245 17165 -7240 17195
rect -7280 17160 -7240 17165
rect -7200 17195 -7160 17200
rect -7200 17165 -7195 17195
rect -7165 17165 -7160 17195
rect -7200 17160 -7160 17165
rect -7120 17195 -7080 17200
rect -7120 17165 -7115 17195
rect -7085 17165 -7080 17195
rect -7120 17160 -7080 17165
rect -7040 17195 -7000 17200
rect -7040 17165 -7035 17195
rect -7005 17165 -7000 17195
rect -7040 17160 -7000 17165
rect -6960 17195 -6920 17200
rect -6960 17165 -6955 17195
rect -6925 17165 -6920 17195
rect -6960 17160 -6920 17165
rect -6880 17195 -6840 17200
rect -6880 17165 -6875 17195
rect -6845 17165 -6840 17195
rect -6880 17160 -6840 17165
rect -6800 17195 -6760 17200
rect -6800 17165 -6795 17195
rect -6765 17165 -6760 17195
rect -6800 17160 -6760 17165
rect -6720 17195 -6680 17200
rect -6720 17165 -6715 17195
rect -6685 17165 -6680 17195
rect -6720 17160 -6680 17165
rect -6640 17195 -6600 17200
rect -6640 17165 -6635 17195
rect -6605 17165 -6600 17195
rect -6640 17160 -6600 17165
rect -6560 17195 -6520 17200
rect -6560 17165 -6555 17195
rect -6525 17165 -6520 17195
rect -6560 17160 -6520 17165
rect -6480 17195 -6440 17200
rect -6480 17165 -6475 17195
rect -6445 17165 -6440 17195
rect -6480 17160 -6440 17165
rect -6400 17195 -6360 17200
rect -6400 17165 -6395 17195
rect -6365 17165 -6360 17195
rect -6400 17160 -6360 17165
rect -6320 17195 -6280 17200
rect -6320 17165 -6315 17195
rect -6285 17165 -6280 17195
rect -6320 17160 -6280 17165
rect -6240 17195 -6200 17200
rect -6240 17165 -6235 17195
rect -6205 17165 -6200 17195
rect -6240 17160 -6200 17165
rect -6160 17195 -6120 17200
rect -6160 17165 -6155 17195
rect -6125 17165 -6120 17195
rect -6160 17160 -6120 17165
rect -6080 17195 -6040 17200
rect -6080 17165 -6075 17195
rect -6045 17165 -6040 17195
rect -6080 17160 -6040 17165
rect -6000 17195 -5960 17200
rect -6000 17165 -5995 17195
rect -5965 17165 -5960 17195
rect -6000 17160 -5960 17165
rect -5920 17195 -5880 17200
rect -5920 17165 -5915 17195
rect -5885 17165 -5880 17195
rect -5920 17160 -5880 17165
rect -5840 17195 -5800 17200
rect -5840 17165 -5835 17195
rect -5805 17165 -5800 17195
rect -5840 17160 -5800 17165
rect -5760 17195 -5720 17200
rect -5760 17165 -5755 17195
rect -5725 17165 -5720 17195
rect -5760 17160 -5720 17165
rect -5440 17195 -5400 17200
rect -5440 17165 -5435 17195
rect -5405 17165 -5400 17195
rect -5440 17160 -5400 17165
rect -5280 17195 -5240 17200
rect -5280 17165 -5275 17195
rect -5245 17165 -5240 17195
rect -5280 17160 -5240 17165
rect -14960 16475 -14920 16480
rect -14960 16445 -14955 16475
rect -14925 16445 -14920 16475
rect -14960 16440 -14920 16445
rect -14880 16475 -14840 16480
rect -14880 16445 -14875 16475
rect -14845 16445 -14840 16475
rect -14880 16440 -14840 16445
rect -14800 16475 -14760 16480
rect -14800 16445 -14795 16475
rect -14765 16445 -14760 16475
rect -14800 16440 -14760 16445
rect -14720 16475 -14680 16480
rect -14720 16445 -14715 16475
rect -14685 16445 -14680 16475
rect -14720 16440 -14680 16445
rect -14640 16475 -14600 16480
rect -14640 16445 -14635 16475
rect -14605 16445 -14600 16475
rect -14640 16440 -14600 16445
rect -14560 16475 -14520 16480
rect -14560 16445 -14555 16475
rect -14525 16445 -14520 16475
rect -14560 16440 -14520 16445
rect -14480 16475 -14440 16480
rect -14480 16445 -14475 16475
rect -14445 16445 -14440 16475
rect -14480 16440 -14440 16445
rect -14400 16475 -14360 16480
rect -14400 16445 -14395 16475
rect -14365 16445 -14360 16475
rect -14400 16440 -14360 16445
rect -14320 16475 -14280 16480
rect -14320 16445 -14315 16475
rect -14285 16445 -14280 16475
rect -14320 16440 -14280 16445
rect -14240 16475 -14200 16480
rect -14240 16445 -14235 16475
rect -14205 16445 -14200 16475
rect -14240 16440 -14200 16445
rect -14160 16475 -14120 16480
rect -14160 16445 -14155 16475
rect -14125 16445 -14120 16475
rect -14160 16440 -14120 16445
rect -14080 16475 -14040 16480
rect -14080 16445 -14075 16475
rect -14045 16445 -14040 16475
rect -14080 16440 -14040 16445
rect -14000 16475 -13960 16480
rect -14000 16445 -13995 16475
rect -13965 16445 -13960 16475
rect -14000 16440 -13960 16445
rect -13920 16475 -13880 16480
rect -13920 16445 -13915 16475
rect -13885 16445 -13880 16475
rect -13920 16440 -13880 16445
rect -13840 16475 -13800 16480
rect -13840 16445 -13835 16475
rect -13805 16445 -13800 16475
rect -13840 16440 -13800 16445
rect -13760 16475 -13720 16480
rect -13760 16445 -13755 16475
rect -13725 16445 -13720 16475
rect -13760 16440 -13720 16445
rect -13680 16475 -13640 16480
rect -13680 16445 -13675 16475
rect -13645 16445 -13640 16475
rect -13680 16440 -13640 16445
rect -13600 16475 -13560 16480
rect -13600 16445 -13595 16475
rect -13565 16445 -13560 16475
rect -13600 16440 -13560 16445
rect -13520 16475 -13480 16480
rect -13520 16445 -13515 16475
rect -13485 16445 -13480 16475
rect -13520 16440 -13480 16445
rect -13440 16475 -13400 16480
rect -13440 16445 -13435 16475
rect -13405 16445 -13400 16475
rect -13440 16440 -13400 16445
rect -13360 16475 -13320 16480
rect -13360 16445 -13355 16475
rect -13325 16445 -13320 16475
rect -13360 16440 -13320 16445
rect -13280 16475 -13240 16480
rect -13280 16445 -13275 16475
rect -13245 16445 -13240 16475
rect -13280 16440 -13240 16445
rect -13200 16475 -13160 16480
rect -13200 16445 -13195 16475
rect -13165 16445 -13160 16475
rect -13200 16440 -13160 16445
rect -13120 16475 -13080 16480
rect -13120 16445 -13115 16475
rect -13085 16445 -13080 16475
rect -13120 16440 -13080 16445
rect -13040 16475 -13000 16480
rect -13040 16445 -13035 16475
rect -13005 16445 -13000 16475
rect -13040 16440 -13000 16445
rect -12960 16475 -12920 16480
rect -12960 16445 -12955 16475
rect -12925 16445 -12920 16475
rect -12960 16440 -12920 16445
rect -12880 16475 -12840 16480
rect -12880 16445 -12875 16475
rect -12845 16445 -12840 16475
rect -12880 16440 -12840 16445
rect -12800 16475 -12760 16480
rect -12800 16445 -12795 16475
rect -12765 16445 -12760 16475
rect -12800 16440 -12760 16445
rect -12720 16475 -12680 16480
rect -12720 16445 -12715 16475
rect -12685 16445 -12680 16475
rect -12720 16440 -12680 16445
rect -12640 16475 -12600 16480
rect -12640 16445 -12635 16475
rect -12605 16445 -12600 16475
rect -12640 16440 -12600 16445
rect -12560 16475 -12520 16480
rect -12560 16445 -12555 16475
rect -12525 16445 -12520 16475
rect -12560 16440 -12520 16445
rect -12480 16475 -12440 16480
rect -12480 16445 -12475 16475
rect -12445 16445 -12440 16475
rect -12480 16440 -12440 16445
rect -12400 16475 -12360 16480
rect -12400 16445 -12395 16475
rect -12365 16445 -12360 16475
rect -12400 16440 -12360 16445
rect -12320 16475 -12280 16480
rect -12320 16445 -12315 16475
rect -12285 16445 -12280 16475
rect -12320 16440 -12280 16445
rect -12240 16475 -12200 16480
rect -12240 16445 -12235 16475
rect -12205 16445 -12200 16475
rect -12240 16440 -12200 16445
rect -12160 16475 -12120 16480
rect -12160 16445 -12155 16475
rect -12125 16445 -12120 16475
rect -12160 16440 -12120 16445
rect -12080 16475 -12040 16480
rect -12080 16445 -12075 16475
rect -12045 16445 -12040 16475
rect -12080 16440 -12040 16445
rect -12000 16475 -11960 16480
rect -12000 16445 -11995 16475
rect -11965 16445 -11960 16475
rect -12000 16440 -11960 16445
rect -11920 16475 -11880 16480
rect -11920 16445 -11915 16475
rect -11885 16445 -11880 16475
rect -11920 16440 -11880 16445
rect -11840 16475 -11800 16480
rect -11840 16445 -11835 16475
rect -11805 16445 -11800 16475
rect -11840 16440 -11800 16445
rect -11760 16475 -11720 16480
rect -11760 16445 -11755 16475
rect -11725 16445 -11720 16475
rect -11760 16440 -11720 16445
rect -11680 16475 -11640 16480
rect -11680 16445 -11675 16475
rect -11645 16445 -11640 16475
rect -11680 16440 -11640 16445
rect -11600 16475 -11560 16480
rect -11600 16445 -11595 16475
rect -11565 16445 -11560 16475
rect -11600 16440 -11560 16445
rect -11520 16475 -11480 16480
rect -11520 16445 -11515 16475
rect -11485 16445 -11480 16475
rect -11520 16440 -11480 16445
rect -11440 16475 -11400 16480
rect -11440 16445 -11435 16475
rect -11405 16445 -11400 16475
rect -11440 16440 -11400 16445
rect -11360 16475 -11320 16480
rect -11360 16445 -11355 16475
rect -11325 16445 -11320 16475
rect -11360 16440 -11320 16445
rect -11280 16475 -11240 16480
rect -11280 16445 -11275 16475
rect -11245 16445 -11240 16475
rect -11280 16440 -11240 16445
rect -11200 16475 -11160 16480
rect -11200 16445 -11195 16475
rect -11165 16445 -11160 16475
rect -11200 16440 -11160 16445
rect -11120 16475 -11080 16480
rect -11120 16445 -11115 16475
rect -11085 16445 -11080 16475
rect -11120 16440 -11080 16445
rect -11040 16475 -11000 16480
rect -11040 16445 -11035 16475
rect -11005 16445 -11000 16475
rect -11040 16440 -11000 16445
rect -10960 16475 -10920 16480
rect -10960 16445 -10955 16475
rect -10925 16445 -10920 16475
rect -10960 16440 -10920 16445
rect -10880 16475 -10840 16480
rect -10880 16445 -10875 16475
rect -10845 16445 -10840 16475
rect -10880 16440 -10840 16445
rect -10800 16475 -10760 16480
rect -10800 16445 -10795 16475
rect -10765 16445 -10760 16475
rect -10800 16440 -10760 16445
rect -10720 16475 -10680 16480
rect -10720 16445 -10715 16475
rect -10685 16445 -10680 16475
rect -10720 16440 -10680 16445
rect -10640 16475 -10600 16480
rect -10640 16445 -10635 16475
rect -10605 16445 -10600 16475
rect -10640 16440 -10600 16445
rect -10560 16475 -10520 16480
rect -10560 16445 -10555 16475
rect -10525 16445 -10520 16475
rect -10560 16440 -10520 16445
rect -10480 16475 -10440 16480
rect -10480 16445 -10475 16475
rect -10445 16445 -10440 16475
rect -10480 16440 -10440 16445
rect -10400 16475 -10360 16480
rect -10400 16445 -10395 16475
rect -10365 16445 -10360 16475
rect -10400 16440 -10360 16445
rect -10320 16475 -10280 16480
rect -10320 16445 -10315 16475
rect -10285 16445 -10280 16475
rect -10320 16440 -10280 16445
rect -10240 16475 -10200 16480
rect -10240 16445 -10235 16475
rect -10205 16445 -10200 16475
rect -10240 16440 -10200 16445
rect -10160 16475 -10120 16480
rect -10160 16445 -10155 16475
rect -10125 16445 -10120 16475
rect -10160 16440 -10120 16445
rect -10080 16475 -10040 16480
rect -10080 16445 -10075 16475
rect -10045 16445 -10040 16475
rect -10080 16440 -10040 16445
rect -10000 16475 -9960 16480
rect -10000 16445 -9995 16475
rect -9965 16445 -9960 16475
rect -10000 16440 -9960 16445
rect -9920 16475 -9880 16480
rect -9920 16445 -9915 16475
rect -9885 16445 -9880 16475
rect -9920 16440 -9880 16445
rect -9840 16475 -9800 16480
rect -9840 16445 -9835 16475
rect -9805 16445 -9800 16475
rect -9840 16440 -9800 16445
rect -9760 16475 -9720 16480
rect -9760 16445 -9755 16475
rect -9725 16445 -9720 16475
rect -9760 16440 -9720 16445
rect -9680 16475 -9640 16480
rect -9680 16445 -9675 16475
rect -9645 16445 -9640 16475
rect -9680 16440 -9640 16445
rect -9600 16475 -9560 16480
rect -9600 16445 -9595 16475
rect -9565 16445 -9560 16475
rect -9600 16440 -9560 16445
rect -9520 16475 -9480 16480
rect -9520 16445 -9515 16475
rect -9485 16445 -9480 16475
rect -9520 16440 -9480 16445
rect -9440 16475 -9400 16480
rect -9440 16445 -9435 16475
rect -9405 16445 -9400 16475
rect -9440 16440 -9400 16445
rect -9360 16475 -9320 16480
rect -9360 16445 -9355 16475
rect -9325 16445 -9320 16475
rect -9360 16440 -9320 16445
rect -9280 16475 -9240 16480
rect -9280 16445 -9275 16475
rect -9245 16445 -9240 16475
rect -9280 16440 -9240 16445
rect -9200 16475 -9160 16480
rect -9200 16445 -9195 16475
rect -9165 16445 -9160 16475
rect -9200 16440 -9160 16445
rect -9120 16475 -9080 16480
rect -9120 16445 -9115 16475
rect -9085 16445 -9080 16475
rect -9120 16440 -9080 16445
rect -9040 16475 -9000 16480
rect -9040 16445 -9035 16475
rect -9005 16445 -9000 16475
rect -9040 16440 -9000 16445
rect -8960 16475 -8920 16480
rect -8960 16445 -8955 16475
rect -8925 16445 -8920 16475
rect -8960 16440 -8920 16445
rect -8880 16475 -8840 16480
rect -8880 16445 -8875 16475
rect -8845 16445 -8840 16475
rect -8880 16440 -8840 16445
rect -8800 16475 -8760 16480
rect -8800 16445 -8795 16475
rect -8765 16445 -8760 16475
rect -8800 16440 -8760 16445
rect -8720 16475 -8680 16480
rect -8720 16445 -8715 16475
rect -8685 16445 -8680 16475
rect -8720 16440 -8680 16445
rect -8640 16475 -8600 16480
rect -8640 16445 -8635 16475
rect -8605 16445 -8600 16475
rect -8640 16440 -8600 16445
rect -8560 16475 -8520 16480
rect -8560 16445 -8555 16475
rect -8525 16445 -8520 16475
rect -8560 16440 -8520 16445
rect -8480 16475 -8440 16480
rect -8480 16445 -8475 16475
rect -8445 16445 -8440 16475
rect -8480 16440 -8440 16445
rect -8400 16475 -8360 16480
rect -8400 16445 -8395 16475
rect -8365 16445 -8360 16475
rect -8400 16440 -8360 16445
rect -8320 16475 -8280 16480
rect -8320 16445 -8315 16475
rect -8285 16445 -8280 16475
rect -8320 16440 -8280 16445
rect -8240 16475 -8200 16480
rect -8240 16445 -8235 16475
rect -8205 16445 -8200 16475
rect -8240 16440 -8200 16445
rect -8160 16475 -8120 16480
rect -8160 16445 -8155 16475
rect -8125 16445 -8120 16475
rect -8160 16440 -8120 16445
rect -8080 16475 -8040 16480
rect -8080 16445 -8075 16475
rect -8045 16445 -8040 16475
rect -8080 16440 -8040 16445
rect -8000 16475 -7960 16480
rect -8000 16445 -7995 16475
rect -7965 16445 -7960 16475
rect -8000 16440 -7960 16445
rect -7920 16475 -7880 16480
rect -7920 16445 -7915 16475
rect -7885 16445 -7880 16475
rect -7920 16440 -7880 16445
rect -7840 16475 -7800 16480
rect -7840 16445 -7835 16475
rect -7805 16445 -7800 16475
rect -7840 16440 -7800 16445
rect -7760 16475 -7720 16480
rect -7760 16445 -7755 16475
rect -7725 16445 -7720 16475
rect -7760 16440 -7720 16445
rect -7680 16475 -7640 16480
rect -7680 16445 -7675 16475
rect -7645 16445 -7640 16475
rect -7680 16440 -7640 16445
rect -7600 16475 -7560 16480
rect -7600 16445 -7595 16475
rect -7565 16445 -7560 16475
rect -7600 16440 -7560 16445
rect -7520 16475 -7480 16480
rect -7520 16445 -7515 16475
rect -7485 16445 -7480 16475
rect -7520 16440 -7480 16445
rect -7440 16475 -7400 16480
rect -7440 16445 -7435 16475
rect -7405 16445 -7400 16475
rect -7440 16440 -7400 16445
rect -7360 16475 -7320 16480
rect -7360 16445 -7355 16475
rect -7325 16445 -7320 16475
rect -7360 16440 -7320 16445
rect -7280 16475 -7240 16480
rect -7280 16445 -7275 16475
rect -7245 16445 -7240 16475
rect -7280 16440 -7240 16445
rect -7200 16475 -7160 16480
rect -7200 16445 -7195 16475
rect -7165 16445 -7160 16475
rect -7200 16440 -7160 16445
rect -7120 16475 -7080 16480
rect -7120 16445 -7115 16475
rect -7085 16445 -7080 16475
rect -7120 16440 -7080 16445
rect -7040 16475 -7000 16480
rect -7040 16445 -7035 16475
rect -7005 16445 -7000 16475
rect -7040 16440 -7000 16445
rect -6960 16475 -6920 16480
rect -6960 16445 -6955 16475
rect -6925 16445 -6920 16475
rect -6960 16440 -6920 16445
rect -6880 16475 -6840 16480
rect -6880 16445 -6875 16475
rect -6845 16445 -6840 16475
rect -6880 16440 -6840 16445
rect -6800 16475 -6760 16480
rect -6800 16445 -6795 16475
rect -6765 16445 -6760 16475
rect -6800 16440 -6760 16445
rect -6720 16475 -6680 16480
rect -6720 16445 -6715 16475
rect -6685 16445 -6680 16475
rect -6720 16440 -6680 16445
rect -6640 16475 -6600 16480
rect -6640 16445 -6635 16475
rect -6605 16445 -6600 16475
rect -6640 16440 -6600 16445
rect -6560 16475 -6520 16480
rect -6560 16445 -6555 16475
rect -6525 16445 -6520 16475
rect -6560 16440 -6520 16445
rect -6480 16475 -6440 16480
rect -6480 16445 -6475 16475
rect -6445 16445 -6440 16475
rect -6480 16440 -6440 16445
rect -6400 16475 -6360 16480
rect -6400 16445 -6395 16475
rect -6365 16445 -6360 16475
rect -6400 16440 -6360 16445
rect -6320 16475 -6280 16480
rect -6320 16445 -6315 16475
rect -6285 16445 -6280 16475
rect -6320 16440 -6280 16445
rect -6240 16475 -6200 16480
rect -6240 16445 -6235 16475
rect -6205 16445 -6200 16475
rect -6240 16440 -6200 16445
rect -6160 16475 -6120 16480
rect -6160 16445 -6155 16475
rect -6125 16445 -6120 16475
rect -6160 16440 -6120 16445
rect -6080 16475 -6040 16480
rect -6080 16445 -6075 16475
rect -6045 16445 -6040 16475
rect -6080 16440 -6040 16445
rect -6000 16475 -5960 16480
rect -6000 16445 -5995 16475
rect -5965 16445 -5960 16475
rect -6000 16440 -5960 16445
rect -5920 16475 -5880 16480
rect -5920 16445 -5915 16475
rect -5885 16445 -5880 16475
rect -5920 16440 -5880 16445
rect -5840 16475 -5800 16480
rect -5840 16445 -5835 16475
rect -5805 16445 -5800 16475
rect -5840 16440 -5800 16445
rect -5760 16475 -5720 16480
rect -5760 16445 -5755 16475
rect -5725 16445 -5720 16475
rect -5760 16440 -5720 16445
rect -5600 16475 -5560 16480
rect -5600 16445 -5595 16475
rect -5565 16445 -5560 16475
rect -5600 16440 -5560 16445
rect -5440 16475 -5400 16480
rect -5440 16445 -5435 16475
rect -5405 16445 -5400 16475
rect -5440 16440 -5400 16445
rect -5360 16475 -5320 16480
rect -5360 16445 -5355 16475
rect -5325 16445 -5320 16475
rect -5360 16440 -5320 16445
rect -5280 16475 -5240 16480
rect -5280 16445 -5275 16475
rect -5245 16445 -5240 16475
rect -5280 16440 -5240 16445
rect -5200 16475 -5160 16480
rect -5200 16445 -5195 16475
rect -5165 16445 -5160 16475
rect -5200 16440 -5160 16445
rect -5120 16475 -5080 16480
rect -5120 16445 -5115 16475
rect -5085 16445 -5080 16475
rect -5120 16440 -5080 16445
rect -5040 16475 -5000 16480
rect -5040 16445 -5035 16475
rect -5005 16445 -5000 16475
rect -5040 16440 -5000 16445
rect -4960 16475 -4920 16480
rect -4960 16445 -4955 16475
rect -4925 16445 -4920 16475
rect -4960 16440 -4920 16445
rect -4880 16475 -4840 16480
rect -4880 16445 -4875 16475
rect -4845 16445 -4840 16475
rect -4880 16440 -4840 16445
rect -4800 16475 -4760 16480
rect -4800 16445 -4795 16475
rect -4765 16445 -4760 16475
rect -4800 16440 -4760 16445
rect -4720 16475 -4680 16480
rect -4720 16445 -4715 16475
rect -4685 16445 -4680 16475
rect -4720 16440 -4680 16445
rect -4640 16475 -4600 16480
rect -4640 16445 -4635 16475
rect -4605 16445 -4600 16475
rect -4640 16440 -4600 16445
rect -4560 16475 -4520 16480
rect -4560 16445 -4555 16475
rect -4525 16445 -4520 16475
rect -4560 16440 -4520 16445
rect -4480 16475 -4440 16480
rect -4480 16445 -4475 16475
rect -4445 16445 -4440 16475
rect -4480 16440 -4440 16445
rect -4400 16475 -4360 16480
rect -4400 16445 -4395 16475
rect -4365 16445 -4360 16475
rect -4400 16440 -4360 16445
rect -4320 16475 -4280 16480
rect -4320 16445 -4315 16475
rect -4285 16445 -4280 16475
rect -4320 16440 -4280 16445
rect -4240 16475 -4200 16480
rect -4240 16445 -4235 16475
rect -4205 16445 -4200 16475
rect -4240 16440 -4200 16445
rect -4160 16475 -4120 16480
rect -4160 16445 -4155 16475
rect -4125 16445 -4120 16475
rect -4160 16440 -4120 16445
rect -4080 16475 -4040 16480
rect -4080 16445 -4075 16475
rect -4045 16445 -4040 16475
rect -4080 16440 -4040 16445
rect -4000 16475 -3960 16480
rect -4000 16445 -3995 16475
rect -3965 16445 -3960 16475
rect -4000 16440 -3960 16445
rect -3920 16475 -3880 16480
rect -3920 16445 -3915 16475
rect -3885 16445 -3880 16475
rect -3920 16440 -3880 16445
rect -3840 16475 -3800 16480
rect -3840 16445 -3835 16475
rect -3805 16445 -3800 16475
rect -3840 16440 -3800 16445
rect -3760 16475 -3720 16480
rect -3760 16445 -3755 16475
rect -3725 16445 -3720 16475
rect -3760 16440 -3720 16445
rect -3680 16475 -3640 16480
rect -3680 16445 -3675 16475
rect -3645 16445 -3640 16475
rect -3680 16440 -3640 16445
rect -3600 16475 -3560 16480
rect -3600 16445 -3595 16475
rect -3565 16445 -3560 16475
rect -3600 16440 -3560 16445
rect -3520 16475 -3480 16480
rect -3520 16445 -3515 16475
rect -3485 16445 -3480 16475
rect -3520 16440 -3480 16445
rect -3440 16475 -3400 16480
rect -3440 16445 -3435 16475
rect -3405 16445 -3400 16475
rect -3440 16440 -3400 16445
rect -3360 16475 -3320 16480
rect -3360 16445 -3355 16475
rect -3325 16445 -3320 16475
rect -3360 16440 -3320 16445
rect -3280 16475 -3240 16480
rect -3280 16445 -3275 16475
rect -3245 16445 -3240 16475
rect -3280 16440 -3240 16445
rect -3200 16475 -3160 16480
rect -3200 16445 -3195 16475
rect -3165 16445 -3160 16475
rect -3200 16440 -3160 16445
rect -3120 16475 -3080 16480
rect -3120 16445 -3115 16475
rect -3085 16445 -3080 16475
rect -3120 16440 -3080 16445
rect -3040 16475 -3000 16480
rect -3040 16445 -3035 16475
rect -3005 16445 -3000 16475
rect -3040 16440 -3000 16445
rect -2960 16475 -2920 16480
rect -2960 16445 -2955 16475
rect -2925 16445 -2920 16475
rect -2960 16440 -2920 16445
rect -2880 16475 -2840 16480
rect -2880 16445 -2875 16475
rect -2845 16445 -2840 16475
rect -2880 16440 -2840 16445
rect -2800 16475 -2760 16480
rect -2800 16445 -2795 16475
rect -2765 16445 -2760 16475
rect -2800 16440 -2760 16445
rect -2720 16475 -2680 16480
rect -2720 16445 -2715 16475
rect -2685 16445 -2680 16475
rect -2720 16440 -2680 16445
rect -2640 16475 -2600 16480
rect -2640 16445 -2635 16475
rect -2605 16445 -2600 16475
rect -2640 16440 -2600 16445
rect -2560 16475 -2520 16480
rect -2560 16445 -2555 16475
rect -2525 16445 -2520 16475
rect -2560 16440 -2520 16445
rect -2480 16475 -2440 16480
rect -2480 16445 -2475 16475
rect -2445 16445 -2440 16475
rect -2480 16440 -2440 16445
rect -2400 16475 -2360 16480
rect -2400 16445 -2395 16475
rect -2365 16445 -2360 16475
rect -2400 16440 -2360 16445
rect -2320 16475 -2280 16480
rect -2320 16445 -2315 16475
rect -2285 16445 -2280 16475
rect -2320 16440 -2280 16445
rect -2240 16475 -2200 16480
rect -2240 16445 -2235 16475
rect -2205 16445 -2200 16475
rect -2240 16440 -2200 16445
rect -2160 16475 -2120 16480
rect -2160 16445 -2155 16475
rect -2125 16445 -2120 16475
rect -2160 16440 -2120 16445
rect -2080 16475 -2040 16480
rect -2080 16445 -2075 16475
rect -2045 16445 -2040 16475
rect -2080 16440 -2040 16445
rect -2000 16475 -1960 16480
rect -2000 16445 -1995 16475
rect -1965 16445 -1960 16475
rect -2000 16440 -1960 16445
rect -1840 16475 -1800 16480
rect -1840 16445 -1835 16475
rect -1805 16445 -1800 16475
rect -1840 16440 -1800 16445
rect -1760 16475 -1720 16480
rect -1760 16445 -1755 16475
rect -1725 16445 -1720 16475
rect -1760 16440 -1720 16445
rect -1680 16475 -1640 16480
rect -1680 16445 -1675 16475
rect -1645 16445 -1640 16475
rect -1680 16440 -1640 16445
rect -1600 16475 -1560 16480
rect -1600 16445 -1595 16475
rect -1565 16445 -1560 16475
rect -1600 16440 -1560 16445
rect -1520 16475 -1480 16480
rect -1520 16445 -1515 16475
rect -1485 16445 -1480 16475
rect -1520 16440 -1480 16445
rect -1440 16475 -1400 16480
rect -1440 16445 -1435 16475
rect -1405 16445 -1400 16475
rect -1440 16440 -1400 16445
rect -1360 16475 -1320 16480
rect -1360 16445 -1355 16475
rect -1325 16445 -1320 16475
rect -1360 16440 -1320 16445
rect -1200 16475 -1160 16480
rect -1200 16445 -1195 16475
rect -1165 16445 -1160 16475
rect -1200 16440 -1160 16445
rect -1040 16475 -1000 16480
rect -1040 16445 -1035 16475
rect -1005 16445 -1000 16475
rect -1040 16440 -1000 16445
rect -880 16475 -840 16480
rect -880 16445 -875 16475
rect -845 16445 -840 16475
rect -880 16440 -840 16445
rect -720 16475 -680 16480
rect -720 16445 -715 16475
rect -685 16445 -680 16475
rect -720 16440 -680 16445
rect -560 16475 -520 16480
rect -560 16445 -555 16475
rect -525 16445 -520 16475
rect -560 16440 -520 16445
rect -14960 16315 -14920 16320
rect -14960 16285 -14955 16315
rect -14925 16285 -14920 16315
rect -14960 16280 -14920 16285
rect -14880 16315 -14840 16320
rect -14880 16285 -14875 16315
rect -14845 16285 -14840 16315
rect -14880 16280 -14840 16285
rect -14800 16315 -14760 16320
rect -14800 16285 -14795 16315
rect -14765 16285 -14760 16315
rect -14800 16280 -14760 16285
rect -14720 16315 -14680 16320
rect -14720 16285 -14715 16315
rect -14685 16285 -14680 16315
rect -14720 16280 -14680 16285
rect -14640 16315 -14600 16320
rect -14640 16285 -14635 16315
rect -14605 16285 -14600 16315
rect -14640 16280 -14600 16285
rect -14560 16315 -14520 16320
rect -14560 16285 -14555 16315
rect -14525 16285 -14520 16315
rect -14560 16280 -14520 16285
rect -14480 16315 -14440 16320
rect -14480 16285 -14475 16315
rect -14445 16285 -14440 16315
rect -14480 16280 -14440 16285
rect -14400 16315 -14360 16320
rect -14400 16285 -14395 16315
rect -14365 16285 -14360 16315
rect -14400 16280 -14360 16285
rect -14320 16315 -14280 16320
rect -14320 16285 -14315 16315
rect -14285 16285 -14280 16315
rect -14320 16280 -14280 16285
rect -14240 16315 -14200 16320
rect -14240 16285 -14235 16315
rect -14205 16285 -14200 16315
rect -14240 16280 -14200 16285
rect -14160 16315 -14120 16320
rect -14160 16285 -14155 16315
rect -14125 16285 -14120 16315
rect -14160 16280 -14120 16285
rect -14080 16315 -14040 16320
rect -14080 16285 -14075 16315
rect -14045 16285 -14040 16315
rect -14080 16280 -14040 16285
rect -14000 16315 -13960 16320
rect -14000 16285 -13995 16315
rect -13965 16285 -13960 16315
rect -14000 16280 -13960 16285
rect -13920 16315 -13880 16320
rect -13920 16285 -13915 16315
rect -13885 16285 -13880 16315
rect -13920 16280 -13880 16285
rect -13840 16315 -13800 16320
rect -13840 16285 -13835 16315
rect -13805 16285 -13800 16315
rect -13840 16280 -13800 16285
rect -13760 16315 -13720 16320
rect -13760 16285 -13755 16315
rect -13725 16285 -13720 16315
rect -13760 16280 -13720 16285
rect -13680 16315 -13640 16320
rect -13680 16285 -13675 16315
rect -13645 16285 -13640 16315
rect -13680 16280 -13640 16285
rect -13600 16315 -13560 16320
rect -13600 16285 -13595 16315
rect -13565 16285 -13560 16315
rect -13600 16280 -13560 16285
rect -13520 16315 -13480 16320
rect -13520 16285 -13515 16315
rect -13485 16285 -13480 16315
rect -13520 16280 -13480 16285
rect -13440 16315 -13400 16320
rect -13440 16285 -13435 16315
rect -13405 16285 -13400 16315
rect -13440 16280 -13400 16285
rect -13360 16315 -13320 16320
rect -13360 16285 -13355 16315
rect -13325 16285 -13320 16315
rect -13360 16280 -13320 16285
rect -13280 16315 -13240 16320
rect -13280 16285 -13275 16315
rect -13245 16285 -13240 16315
rect -13280 16280 -13240 16285
rect -13200 16315 -13160 16320
rect -13200 16285 -13195 16315
rect -13165 16285 -13160 16315
rect -13200 16280 -13160 16285
rect -13120 16315 -13080 16320
rect -13120 16285 -13115 16315
rect -13085 16285 -13080 16315
rect -13120 16280 -13080 16285
rect -13040 16315 -13000 16320
rect -13040 16285 -13035 16315
rect -13005 16285 -13000 16315
rect -13040 16280 -13000 16285
rect -12960 16315 -12920 16320
rect -12960 16285 -12955 16315
rect -12925 16285 -12920 16315
rect -12960 16280 -12920 16285
rect -12880 16315 -12840 16320
rect -12880 16285 -12875 16315
rect -12845 16285 -12840 16315
rect -12880 16280 -12840 16285
rect -12800 16315 -12760 16320
rect -12800 16285 -12795 16315
rect -12765 16285 -12760 16315
rect -12800 16280 -12760 16285
rect -12720 16315 -12680 16320
rect -12720 16285 -12715 16315
rect -12685 16285 -12680 16315
rect -12720 16280 -12680 16285
rect -12640 16315 -12600 16320
rect -12640 16285 -12635 16315
rect -12605 16285 -12600 16315
rect -12640 16280 -12600 16285
rect -12560 16315 -12520 16320
rect -12560 16285 -12555 16315
rect -12525 16285 -12520 16315
rect -12560 16280 -12520 16285
rect -12480 16315 -12440 16320
rect -12480 16285 -12475 16315
rect -12445 16285 -12440 16315
rect -12480 16280 -12440 16285
rect -12400 16315 -12360 16320
rect -12400 16285 -12395 16315
rect -12365 16285 -12360 16315
rect -12400 16280 -12360 16285
rect -12320 16315 -12280 16320
rect -12320 16285 -12315 16315
rect -12285 16285 -12280 16315
rect -12320 16280 -12280 16285
rect -12240 16315 -12200 16320
rect -12240 16285 -12235 16315
rect -12205 16285 -12200 16315
rect -12240 16280 -12200 16285
rect -12160 16315 -12120 16320
rect -12160 16285 -12155 16315
rect -12125 16285 -12120 16315
rect -12160 16280 -12120 16285
rect -12080 16315 -12040 16320
rect -12080 16285 -12075 16315
rect -12045 16285 -12040 16315
rect -12080 16280 -12040 16285
rect -12000 16315 -11960 16320
rect -12000 16285 -11995 16315
rect -11965 16285 -11960 16315
rect -12000 16280 -11960 16285
rect -11920 16315 -11880 16320
rect -11920 16285 -11915 16315
rect -11885 16285 -11880 16315
rect -11920 16280 -11880 16285
rect -11840 16315 -11800 16320
rect -11840 16285 -11835 16315
rect -11805 16285 -11800 16315
rect -11840 16280 -11800 16285
rect -11760 16315 -11720 16320
rect -11760 16285 -11755 16315
rect -11725 16285 -11720 16315
rect -11760 16280 -11720 16285
rect -11680 16315 -11640 16320
rect -11680 16285 -11675 16315
rect -11645 16285 -11640 16315
rect -11680 16280 -11640 16285
rect -11600 16315 -11560 16320
rect -11600 16285 -11595 16315
rect -11565 16285 -11560 16315
rect -11600 16280 -11560 16285
rect -11520 16315 -11480 16320
rect -11520 16285 -11515 16315
rect -11485 16285 -11480 16315
rect -11520 16280 -11480 16285
rect -11440 16315 -11400 16320
rect -11440 16285 -11435 16315
rect -11405 16285 -11400 16315
rect -11440 16280 -11400 16285
rect -11360 16315 -11320 16320
rect -11360 16285 -11355 16315
rect -11325 16285 -11320 16315
rect -11360 16280 -11320 16285
rect -11280 16315 -11240 16320
rect -11280 16285 -11275 16315
rect -11245 16285 -11240 16315
rect -11280 16280 -11240 16285
rect -11200 16315 -11160 16320
rect -11200 16285 -11195 16315
rect -11165 16285 -11160 16315
rect -11200 16280 -11160 16285
rect -11120 16315 -11080 16320
rect -11120 16285 -11115 16315
rect -11085 16285 -11080 16315
rect -11120 16280 -11080 16285
rect -11040 16315 -11000 16320
rect -11040 16285 -11035 16315
rect -11005 16285 -11000 16315
rect -11040 16280 -11000 16285
rect -10960 16315 -10920 16320
rect -10960 16285 -10955 16315
rect -10925 16285 -10920 16315
rect -10960 16280 -10920 16285
rect -10880 16315 -10840 16320
rect -10880 16285 -10875 16315
rect -10845 16285 -10840 16315
rect -10880 16280 -10840 16285
rect -10800 16315 -10760 16320
rect -10800 16285 -10795 16315
rect -10765 16285 -10760 16315
rect -10800 16280 -10760 16285
rect -10720 16315 -10680 16320
rect -10720 16285 -10715 16315
rect -10685 16285 -10680 16315
rect -10720 16280 -10680 16285
rect -10640 16315 -10600 16320
rect -10640 16285 -10635 16315
rect -10605 16285 -10600 16315
rect -10640 16280 -10600 16285
rect -10560 16315 -10520 16320
rect -10560 16285 -10555 16315
rect -10525 16285 -10520 16315
rect -10560 16280 -10520 16285
rect -10480 16315 -10440 16320
rect -10480 16285 -10475 16315
rect -10445 16285 -10440 16315
rect -10480 16280 -10440 16285
rect -10400 16315 -10360 16320
rect -10400 16285 -10395 16315
rect -10365 16285 -10360 16315
rect -10400 16280 -10360 16285
rect -10320 16315 -10280 16320
rect -10320 16285 -10315 16315
rect -10285 16285 -10280 16315
rect -10320 16280 -10280 16285
rect -10240 16315 -10200 16320
rect -10240 16285 -10235 16315
rect -10205 16285 -10200 16315
rect -10240 16280 -10200 16285
rect -10160 16315 -10120 16320
rect -10160 16285 -10155 16315
rect -10125 16285 -10120 16315
rect -10160 16280 -10120 16285
rect -10080 16315 -10040 16320
rect -10080 16285 -10075 16315
rect -10045 16285 -10040 16315
rect -10080 16280 -10040 16285
rect -10000 16315 -9960 16320
rect -10000 16285 -9995 16315
rect -9965 16285 -9960 16315
rect -10000 16280 -9960 16285
rect -9920 16315 -9880 16320
rect -9920 16285 -9915 16315
rect -9885 16285 -9880 16315
rect -9920 16280 -9880 16285
rect -9840 16315 -9800 16320
rect -9840 16285 -9835 16315
rect -9805 16285 -9800 16315
rect -9840 16280 -9800 16285
rect -9760 16315 -9720 16320
rect -9760 16285 -9755 16315
rect -9725 16285 -9720 16315
rect -9760 16280 -9720 16285
rect -9680 16315 -9640 16320
rect -9680 16285 -9675 16315
rect -9645 16285 -9640 16315
rect -9680 16280 -9640 16285
rect -9600 16315 -9560 16320
rect -9600 16285 -9595 16315
rect -9565 16285 -9560 16315
rect -9600 16280 -9560 16285
rect -9520 16315 -9480 16320
rect -9520 16285 -9515 16315
rect -9485 16285 -9480 16315
rect -9520 16280 -9480 16285
rect -9440 16315 -9400 16320
rect -9440 16285 -9435 16315
rect -9405 16285 -9400 16315
rect -9440 16280 -9400 16285
rect -9360 16315 -9320 16320
rect -9360 16285 -9355 16315
rect -9325 16285 -9320 16315
rect -9360 16280 -9320 16285
rect -9280 16315 -9240 16320
rect -9280 16285 -9275 16315
rect -9245 16285 -9240 16315
rect -9280 16280 -9240 16285
rect -9200 16315 -9160 16320
rect -9200 16285 -9195 16315
rect -9165 16285 -9160 16315
rect -9200 16280 -9160 16285
rect -9120 16315 -9080 16320
rect -9120 16285 -9115 16315
rect -9085 16285 -9080 16315
rect -9120 16280 -9080 16285
rect -9040 16315 -9000 16320
rect -9040 16285 -9035 16315
rect -9005 16285 -9000 16315
rect -9040 16280 -9000 16285
rect -8960 16315 -8920 16320
rect -8960 16285 -8955 16315
rect -8925 16285 -8920 16315
rect -8960 16280 -8920 16285
rect -8880 16315 -8840 16320
rect -8880 16285 -8875 16315
rect -8845 16285 -8840 16315
rect -8880 16280 -8840 16285
rect -8800 16315 -8760 16320
rect -8800 16285 -8795 16315
rect -8765 16285 -8760 16315
rect -8800 16280 -8760 16285
rect -8720 16315 -8680 16320
rect -8720 16285 -8715 16315
rect -8685 16285 -8680 16315
rect -8720 16280 -8680 16285
rect -8640 16315 -8600 16320
rect -8640 16285 -8635 16315
rect -8605 16285 -8600 16315
rect -8640 16280 -8600 16285
rect -8560 16315 -8520 16320
rect -8560 16285 -8555 16315
rect -8525 16285 -8520 16315
rect -8560 16280 -8520 16285
rect -8480 16315 -8440 16320
rect -8480 16285 -8475 16315
rect -8445 16285 -8440 16315
rect -8480 16280 -8440 16285
rect -8400 16315 -8360 16320
rect -8400 16285 -8395 16315
rect -8365 16285 -8360 16315
rect -8400 16280 -8360 16285
rect -8320 16315 -8280 16320
rect -8320 16285 -8315 16315
rect -8285 16285 -8280 16315
rect -8320 16280 -8280 16285
rect -8240 16315 -8200 16320
rect -8240 16285 -8235 16315
rect -8205 16285 -8200 16315
rect -8240 16280 -8200 16285
rect -8160 16315 -8120 16320
rect -8160 16285 -8155 16315
rect -8125 16285 -8120 16315
rect -8160 16280 -8120 16285
rect -8080 16315 -8040 16320
rect -8080 16285 -8075 16315
rect -8045 16285 -8040 16315
rect -8080 16280 -8040 16285
rect -8000 16315 -7960 16320
rect -8000 16285 -7995 16315
rect -7965 16285 -7960 16315
rect -8000 16280 -7960 16285
rect -7920 16315 -7880 16320
rect -7920 16285 -7915 16315
rect -7885 16285 -7880 16315
rect -7920 16280 -7880 16285
rect -7840 16315 -7800 16320
rect -7840 16285 -7835 16315
rect -7805 16285 -7800 16315
rect -7840 16280 -7800 16285
rect -7760 16315 -7720 16320
rect -7760 16285 -7755 16315
rect -7725 16285 -7720 16315
rect -7760 16280 -7720 16285
rect -7680 16315 -7640 16320
rect -7680 16285 -7675 16315
rect -7645 16285 -7640 16315
rect -7680 16280 -7640 16285
rect -7600 16315 -7560 16320
rect -7600 16285 -7595 16315
rect -7565 16285 -7560 16315
rect -7600 16280 -7560 16285
rect -7520 16315 -7480 16320
rect -7520 16285 -7515 16315
rect -7485 16285 -7480 16315
rect -7520 16280 -7480 16285
rect -7440 16315 -7400 16320
rect -7440 16285 -7435 16315
rect -7405 16285 -7400 16315
rect -7440 16280 -7400 16285
rect -7360 16315 -7320 16320
rect -7360 16285 -7355 16315
rect -7325 16285 -7320 16315
rect -7360 16280 -7320 16285
rect -7280 16315 -7240 16320
rect -7280 16285 -7275 16315
rect -7245 16285 -7240 16315
rect -7280 16280 -7240 16285
rect -7200 16315 -7160 16320
rect -7200 16285 -7195 16315
rect -7165 16285 -7160 16315
rect -7200 16280 -7160 16285
rect -7120 16315 -7080 16320
rect -7120 16285 -7115 16315
rect -7085 16285 -7080 16315
rect -7120 16280 -7080 16285
rect -7040 16315 -7000 16320
rect -7040 16285 -7035 16315
rect -7005 16285 -7000 16315
rect -7040 16280 -7000 16285
rect -6960 16315 -6920 16320
rect -6960 16285 -6955 16315
rect -6925 16285 -6920 16315
rect -6960 16280 -6920 16285
rect -6880 16315 -6840 16320
rect -6880 16285 -6875 16315
rect -6845 16285 -6840 16315
rect -6880 16280 -6840 16285
rect -6800 16315 -6760 16320
rect -6800 16285 -6795 16315
rect -6765 16285 -6760 16315
rect -6800 16280 -6760 16285
rect -6720 16315 -6680 16320
rect -6720 16285 -6715 16315
rect -6685 16285 -6680 16315
rect -6720 16280 -6680 16285
rect -6640 16315 -6600 16320
rect -6640 16285 -6635 16315
rect -6605 16285 -6600 16315
rect -6640 16280 -6600 16285
rect -6560 16315 -6520 16320
rect -6560 16285 -6555 16315
rect -6525 16285 -6520 16315
rect -6560 16280 -6520 16285
rect -6480 16315 -6440 16320
rect -6480 16285 -6475 16315
rect -6445 16285 -6440 16315
rect -6480 16280 -6440 16285
rect -6400 16315 -6360 16320
rect -6400 16285 -6395 16315
rect -6365 16285 -6360 16315
rect -6400 16280 -6360 16285
rect -6320 16315 -6280 16320
rect -6320 16285 -6315 16315
rect -6285 16285 -6280 16315
rect -6320 16280 -6280 16285
rect -6240 16315 -6200 16320
rect -6240 16285 -6235 16315
rect -6205 16285 -6200 16315
rect -6240 16280 -6200 16285
rect -6160 16315 -6120 16320
rect -6160 16285 -6155 16315
rect -6125 16285 -6120 16315
rect -6160 16280 -6120 16285
rect -6080 16315 -6040 16320
rect -6080 16285 -6075 16315
rect -6045 16285 -6040 16315
rect -6080 16280 -6040 16285
rect -6000 16315 -5960 16320
rect -6000 16285 -5995 16315
rect -5965 16285 -5960 16315
rect -6000 16280 -5960 16285
rect -5920 16315 -5880 16320
rect -5920 16285 -5915 16315
rect -5885 16285 -5880 16315
rect -5920 16280 -5880 16285
rect -5840 16315 -5800 16320
rect -5840 16285 -5835 16315
rect -5805 16285 -5800 16315
rect -5840 16280 -5800 16285
rect -5760 16315 -5720 16320
rect -5760 16285 -5755 16315
rect -5725 16285 -5720 16315
rect -5760 16280 -5720 16285
rect -5600 16315 -5560 16320
rect -5600 16285 -5595 16315
rect -5565 16285 -5560 16315
rect -5600 16280 -5560 16285
rect -5440 16315 -5400 16320
rect -5440 16285 -5435 16315
rect -5405 16285 -5400 16315
rect -5440 16280 -5400 16285
rect -5360 16315 -5320 16320
rect -5360 16285 -5355 16315
rect -5325 16285 -5320 16315
rect -5360 16280 -5320 16285
rect -5280 16315 -5240 16320
rect -5280 16285 -5275 16315
rect -5245 16285 -5240 16315
rect -5280 16280 -5240 16285
rect -5200 16315 -5160 16320
rect -5200 16285 -5195 16315
rect -5165 16285 -5160 16315
rect -5200 16280 -5160 16285
rect -5120 16315 -5080 16320
rect -5120 16285 -5115 16315
rect -5085 16285 -5080 16315
rect -5120 16280 -5080 16285
rect -5040 16315 -5000 16320
rect -5040 16285 -5035 16315
rect -5005 16285 -5000 16315
rect -5040 16280 -5000 16285
rect -4960 16315 -4920 16320
rect -4960 16285 -4955 16315
rect -4925 16285 -4920 16315
rect -4960 16280 -4920 16285
rect -4880 16315 -4840 16320
rect -4880 16285 -4875 16315
rect -4845 16285 -4840 16315
rect -4880 16280 -4840 16285
rect -4800 16315 -4760 16320
rect -4800 16285 -4795 16315
rect -4765 16285 -4760 16315
rect -4800 16280 -4760 16285
rect -4720 16315 -4680 16320
rect -4720 16285 -4715 16315
rect -4685 16285 -4680 16315
rect -4720 16280 -4680 16285
rect -4640 16315 -4600 16320
rect -4640 16285 -4635 16315
rect -4605 16285 -4600 16315
rect -4640 16280 -4600 16285
rect -4560 16315 -4520 16320
rect -4560 16285 -4555 16315
rect -4525 16285 -4520 16315
rect -4560 16280 -4520 16285
rect -4480 16315 -4440 16320
rect -4480 16285 -4475 16315
rect -4445 16285 -4440 16315
rect -4480 16280 -4440 16285
rect -4400 16315 -4360 16320
rect -4400 16285 -4395 16315
rect -4365 16285 -4360 16315
rect -4400 16280 -4360 16285
rect -4320 16315 -4280 16320
rect -4320 16285 -4315 16315
rect -4285 16285 -4280 16315
rect -4320 16280 -4280 16285
rect -4240 16315 -4200 16320
rect -4240 16285 -4235 16315
rect -4205 16285 -4200 16315
rect -4240 16280 -4200 16285
rect -4160 16315 -4120 16320
rect -4160 16285 -4155 16315
rect -4125 16285 -4120 16315
rect -4160 16280 -4120 16285
rect -4080 16315 -4040 16320
rect -4080 16285 -4075 16315
rect -4045 16285 -4040 16315
rect -4080 16280 -4040 16285
rect -4000 16315 -3960 16320
rect -4000 16285 -3995 16315
rect -3965 16285 -3960 16315
rect -4000 16280 -3960 16285
rect -3920 16315 -3880 16320
rect -3920 16285 -3915 16315
rect -3885 16285 -3880 16315
rect -3920 16280 -3880 16285
rect -3840 16315 -3800 16320
rect -3840 16285 -3835 16315
rect -3805 16285 -3800 16315
rect -3840 16280 -3800 16285
rect -3760 16315 -3720 16320
rect -3760 16285 -3755 16315
rect -3725 16285 -3720 16315
rect -3760 16280 -3720 16285
rect -3680 16315 -3640 16320
rect -3680 16285 -3675 16315
rect -3645 16285 -3640 16315
rect -3680 16280 -3640 16285
rect -3600 16315 -3560 16320
rect -3600 16285 -3595 16315
rect -3565 16285 -3560 16315
rect -3600 16280 -3560 16285
rect -3520 16315 -3480 16320
rect -3520 16285 -3515 16315
rect -3485 16285 -3480 16315
rect -3520 16280 -3480 16285
rect -3440 16315 -3400 16320
rect -3440 16285 -3435 16315
rect -3405 16285 -3400 16315
rect -3440 16280 -3400 16285
rect -3360 16315 -3320 16320
rect -3360 16285 -3355 16315
rect -3325 16285 -3320 16315
rect -3360 16280 -3320 16285
rect -3280 16315 -3240 16320
rect -3280 16285 -3275 16315
rect -3245 16285 -3240 16315
rect -3280 16280 -3240 16285
rect -3200 16315 -3160 16320
rect -3200 16285 -3195 16315
rect -3165 16285 -3160 16315
rect -3200 16280 -3160 16285
rect -3120 16315 -3080 16320
rect -3120 16285 -3115 16315
rect -3085 16285 -3080 16315
rect -3120 16280 -3080 16285
rect -3040 16315 -3000 16320
rect -3040 16285 -3035 16315
rect -3005 16285 -3000 16315
rect -3040 16280 -3000 16285
rect -2960 16315 -2920 16320
rect -2960 16285 -2955 16315
rect -2925 16285 -2920 16315
rect -2960 16280 -2920 16285
rect -2880 16315 -2840 16320
rect -2880 16285 -2875 16315
rect -2845 16285 -2840 16315
rect -2880 16280 -2840 16285
rect -2800 16315 -2760 16320
rect -2800 16285 -2795 16315
rect -2765 16285 -2760 16315
rect -2800 16280 -2760 16285
rect -2720 16315 -2680 16320
rect -2720 16285 -2715 16315
rect -2685 16285 -2680 16315
rect -2720 16280 -2680 16285
rect -2640 16315 -2600 16320
rect -2640 16285 -2635 16315
rect -2605 16285 -2600 16315
rect -2640 16280 -2600 16285
rect -2560 16315 -2520 16320
rect -2560 16285 -2555 16315
rect -2525 16285 -2520 16315
rect -2560 16280 -2520 16285
rect -2480 16315 -2440 16320
rect -2480 16285 -2475 16315
rect -2445 16285 -2440 16315
rect -2480 16280 -2440 16285
rect -2400 16315 -2360 16320
rect -2400 16285 -2395 16315
rect -2365 16285 -2360 16315
rect -2400 16280 -2360 16285
rect -2320 16315 -2280 16320
rect -2320 16285 -2315 16315
rect -2285 16285 -2280 16315
rect -2320 16280 -2280 16285
rect -2240 16315 -2200 16320
rect -2240 16285 -2235 16315
rect -2205 16285 -2200 16315
rect -2240 16280 -2200 16285
rect -2160 16315 -2120 16320
rect -2160 16285 -2155 16315
rect -2125 16285 -2120 16315
rect -2160 16280 -2120 16285
rect -2080 16315 -2040 16320
rect -2080 16285 -2075 16315
rect -2045 16285 -2040 16315
rect -2080 16280 -2040 16285
rect -2000 16315 -1960 16320
rect -2000 16285 -1995 16315
rect -1965 16285 -1960 16315
rect -2000 16280 -1960 16285
rect -1840 16315 -1800 16320
rect -1840 16285 -1835 16315
rect -1805 16285 -1800 16315
rect -1840 16280 -1800 16285
rect -1760 16315 -1720 16320
rect -1760 16285 -1755 16315
rect -1725 16285 -1720 16315
rect -1760 16280 -1720 16285
rect -1680 16315 -1640 16320
rect -1680 16285 -1675 16315
rect -1645 16285 -1640 16315
rect -1680 16280 -1640 16285
rect -1600 16315 -1560 16320
rect -1600 16285 -1595 16315
rect -1565 16285 -1560 16315
rect -1600 16280 -1560 16285
rect -1520 16315 -1480 16320
rect -1520 16285 -1515 16315
rect -1485 16285 -1480 16315
rect -1520 16280 -1480 16285
rect -1440 16315 -1400 16320
rect -1440 16285 -1435 16315
rect -1405 16285 -1400 16315
rect -1440 16280 -1400 16285
rect -1360 16315 -1320 16320
rect -1360 16285 -1355 16315
rect -1325 16285 -1320 16315
rect -1360 16280 -1320 16285
rect -1200 16315 -1160 16320
rect -1200 16285 -1195 16315
rect -1165 16285 -1160 16315
rect -1200 16280 -1160 16285
rect -1040 16315 -1000 16320
rect -1040 16285 -1035 16315
rect -1005 16285 -1000 16315
rect -1040 16280 -1000 16285
rect -880 16315 -840 16320
rect -880 16285 -875 16315
rect -845 16285 -840 16315
rect -880 16280 -840 16285
rect -720 16315 -680 16320
rect -720 16285 -715 16315
rect -685 16285 -680 16315
rect -720 16280 -680 16285
rect -560 16315 -520 16320
rect -560 16285 -555 16315
rect -525 16285 -520 16315
rect -560 16280 -520 16285
rect -14960 16155 -14920 16160
rect -14960 16125 -14955 16155
rect -14925 16125 -14920 16155
rect -14960 16120 -14920 16125
rect -14880 16155 -14840 16160
rect -14880 16125 -14875 16155
rect -14845 16125 -14840 16155
rect -14880 16120 -14840 16125
rect -14800 16155 -14760 16160
rect -14800 16125 -14795 16155
rect -14765 16125 -14760 16155
rect -14800 16120 -14760 16125
rect -14720 16155 -14680 16160
rect -14720 16125 -14715 16155
rect -14685 16125 -14680 16155
rect -14720 16120 -14680 16125
rect -14640 16155 -14600 16160
rect -14640 16125 -14635 16155
rect -14605 16125 -14600 16155
rect -14640 16120 -14600 16125
rect -14560 16155 -14520 16160
rect -14560 16125 -14555 16155
rect -14525 16125 -14520 16155
rect -14560 16120 -14520 16125
rect -14480 16155 -14440 16160
rect -14480 16125 -14475 16155
rect -14445 16125 -14440 16155
rect -14480 16120 -14440 16125
rect -14400 16155 -14360 16160
rect -14400 16125 -14395 16155
rect -14365 16125 -14360 16155
rect -14400 16120 -14360 16125
rect -14320 16155 -14280 16160
rect -14320 16125 -14315 16155
rect -14285 16125 -14280 16155
rect -14320 16120 -14280 16125
rect -14240 16155 -14200 16160
rect -14240 16125 -14235 16155
rect -14205 16125 -14200 16155
rect -14240 16120 -14200 16125
rect -14160 16155 -14120 16160
rect -14160 16125 -14155 16155
rect -14125 16125 -14120 16155
rect -14160 16120 -14120 16125
rect -14080 16155 -14040 16160
rect -14080 16125 -14075 16155
rect -14045 16125 -14040 16155
rect -14080 16120 -14040 16125
rect -14000 16155 -13960 16160
rect -14000 16125 -13995 16155
rect -13965 16125 -13960 16155
rect -14000 16120 -13960 16125
rect -13920 16155 -13880 16160
rect -13920 16125 -13915 16155
rect -13885 16125 -13880 16155
rect -13920 16120 -13880 16125
rect -13840 16155 -13800 16160
rect -13840 16125 -13835 16155
rect -13805 16125 -13800 16155
rect -13840 16120 -13800 16125
rect -13760 16155 -13720 16160
rect -13760 16125 -13755 16155
rect -13725 16125 -13720 16155
rect -13760 16120 -13720 16125
rect -13680 16155 -13640 16160
rect -13680 16125 -13675 16155
rect -13645 16125 -13640 16155
rect -13680 16120 -13640 16125
rect -13600 16155 -13560 16160
rect -13600 16125 -13595 16155
rect -13565 16125 -13560 16155
rect -13600 16120 -13560 16125
rect -13520 16155 -13480 16160
rect -13520 16125 -13515 16155
rect -13485 16125 -13480 16155
rect -13520 16120 -13480 16125
rect -13440 16155 -13400 16160
rect -13440 16125 -13435 16155
rect -13405 16125 -13400 16155
rect -13440 16120 -13400 16125
rect -13360 16155 -13320 16160
rect -13360 16125 -13355 16155
rect -13325 16125 -13320 16155
rect -13360 16120 -13320 16125
rect -13280 16155 -13240 16160
rect -13280 16125 -13275 16155
rect -13245 16125 -13240 16155
rect -13280 16120 -13240 16125
rect -13200 16155 -13160 16160
rect -13200 16125 -13195 16155
rect -13165 16125 -13160 16155
rect -13200 16120 -13160 16125
rect -13120 16155 -13080 16160
rect -13120 16125 -13115 16155
rect -13085 16125 -13080 16155
rect -13120 16120 -13080 16125
rect -13040 16155 -13000 16160
rect -13040 16125 -13035 16155
rect -13005 16125 -13000 16155
rect -13040 16120 -13000 16125
rect -12960 16155 -12920 16160
rect -12960 16125 -12955 16155
rect -12925 16125 -12920 16155
rect -12960 16120 -12920 16125
rect -12880 16155 -12840 16160
rect -12880 16125 -12875 16155
rect -12845 16125 -12840 16155
rect -12880 16120 -12840 16125
rect -12800 16155 -12760 16160
rect -12800 16125 -12795 16155
rect -12765 16125 -12760 16155
rect -12800 16120 -12760 16125
rect -12720 16155 -12680 16160
rect -12720 16125 -12715 16155
rect -12685 16125 -12680 16155
rect -12720 16120 -12680 16125
rect -12640 16155 -12600 16160
rect -12640 16125 -12635 16155
rect -12605 16125 -12600 16155
rect -12640 16120 -12600 16125
rect -12560 16155 -12520 16160
rect -12560 16125 -12555 16155
rect -12525 16125 -12520 16155
rect -12560 16120 -12520 16125
rect -12480 16155 -12440 16160
rect -12480 16125 -12475 16155
rect -12445 16125 -12440 16155
rect -12480 16120 -12440 16125
rect -12400 16155 -12360 16160
rect -12400 16125 -12395 16155
rect -12365 16125 -12360 16155
rect -12400 16120 -12360 16125
rect -12320 16155 -12280 16160
rect -12320 16125 -12315 16155
rect -12285 16125 -12280 16155
rect -12320 16120 -12280 16125
rect -12240 16155 -12200 16160
rect -12240 16125 -12235 16155
rect -12205 16125 -12200 16155
rect -12240 16120 -12200 16125
rect -12160 16155 -12120 16160
rect -12160 16125 -12155 16155
rect -12125 16125 -12120 16155
rect -12160 16120 -12120 16125
rect -12080 16155 -12040 16160
rect -12080 16125 -12075 16155
rect -12045 16125 -12040 16155
rect -12080 16120 -12040 16125
rect -12000 16155 -11960 16160
rect -12000 16125 -11995 16155
rect -11965 16125 -11960 16155
rect -12000 16120 -11960 16125
rect -11920 16155 -11880 16160
rect -11920 16125 -11915 16155
rect -11885 16125 -11880 16155
rect -11920 16120 -11880 16125
rect -11840 16155 -11800 16160
rect -11840 16125 -11835 16155
rect -11805 16125 -11800 16155
rect -11840 16120 -11800 16125
rect -11760 16155 -11720 16160
rect -11760 16125 -11755 16155
rect -11725 16125 -11720 16155
rect -11760 16120 -11720 16125
rect -11680 16155 -11640 16160
rect -11680 16125 -11675 16155
rect -11645 16125 -11640 16155
rect -11680 16120 -11640 16125
rect -11600 16155 -11560 16160
rect -11600 16125 -11595 16155
rect -11565 16125 -11560 16155
rect -11600 16120 -11560 16125
rect -11520 16155 -11480 16160
rect -11520 16125 -11515 16155
rect -11485 16125 -11480 16155
rect -11520 16120 -11480 16125
rect -11440 16155 -11400 16160
rect -11440 16125 -11435 16155
rect -11405 16125 -11400 16155
rect -11440 16120 -11400 16125
rect -11360 16155 -11320 16160
rect -11360 16125 -11355 16155
rect -11325 16125 -11320 16155
rect -11360 16120 -11320 16125
rect -11280 16155 -11240 16160
rect -11280 16125 -11275 16155
rect -11245 16125 -11240 16155
rect -11280 16120 -11240 16125
rect -11200 16155 -11160 16160
rect -11200 16125 -11195 16155
rect -11165 16125 -11160 16155
rect -11200 16120 -11160 16125
rect -11120 16155 -11080 16160
rect -11120 16125 -11115 16155
rect -11085 16125 -11080 16155
rect -11120 16120 -11080 16125
rect -11040 16155 -11000 16160
rect -11040 16125 -11035 16155
rect -11005 16125 -11000 16155
rect -11040 16120 -11000 16125
rect -10960 16155 -10920 16160
rect -10960 16125 -10955 16155
rect -10925 16125 -10920 16155
rect -10960 16120 -10920 16125
rect -10880 16155 -10840 16160
rect -10880 16125 -10875 16155
rect -10845 16125 -10840 16155
rect -10880 16120 -10840 16125
rect -10800 16155 -10760 16160
rect -10800 16125 -10795 16155
rect -10765 16125 -10760 16155
rect -10800 16120 -10760 16125
rect -10720 16155 -10680 16160
rect -10720 16125 -10715 16155
rect -10685 16125 -10680 16155
rect -10720 16120 -10680 16125
rect -10640 16155 -10600 16160
rect -10640 16125 -10635 16155
rect -10605 16125 -10600 16155
rect -10640 16120 -10600 16125
rect -10560 16155 -10520 16160
rect -10560 16125 -10555 16155
rect -10525 16125 -10520 16155
rect -10560 16120 -10520 16125
rect -10480 16155 -10440 16160
rect -10480 16125 -10475 16155
rect -10445 16125 -10440 16155
rect -10480 16120 -10440 16125
rect -10400 16155 -10360 16160
rect -10400 16125 -10395 16155
rect -10365 16125 -10360 16155
rect -10400 16120 -10360 16125
rect -10320 16155 -10280 16160
rect -10320 16125 -10315 16155
rect -10285 16125 -10280 16155
rect -10320 16120 -10280 16125
rect -10240 16155 -10200 16160
rect -10240 16125 -10235 16155
rect -10205 16125 -10200 16155
rect -10240 16120 -10200 16125
rect -10160 16155 -10120 16160
rect -10160 16125 -10155 16155
rect -10125 16125 -10120 16155
rect -10160 16120 -10120 16125
rect -10080 16155 -10040 16160
rect -10080 16125 -10075 16155
rect -10045 16125 -10040 16155
rect -10080 16120 -10040 16125
rect -10000 16155 -9960 16160
rect -10000 16125 -9995 16155
rect -9965 16125 -9960 16155
rect -10000 16120 -9960 16125
rect -9920 16155 -9880 16160
rect -9920 16125 -9915 16155
rect -9885 16125 -9880 16155
rect -9920 16120 -9880 16125
rect -9840 16155 -9800 16160
rect -9840 16125 -9835 16155
rect -9805 16125 -9800 16155
rect -9840 16120 -9800 16125
rect -9760 16155 -9720 16160
rect -9760 16125 -9755 16155
rect -9725 16125 -9720 16155
rect -9760 16120 -9720 16125
rect -9680 16155 -9640 16160
rect -9680 16125 -9675 16155
rect -9645 16125 -9640 16155
rect -9680 16120 -9640 16125
rect -9600 16155 -9560 16160
rect -9600 16125 -9595 16155
rect -9565 16125 -9560 16155
rect -9600 16120 -9560 16125
rect -9520 16155 -9480 16160
rect -9520 16125 -9515 16155
rect -9485 16125 -9480 16155
rect -9520 16120 -9480 16125
rect -9440 16155 -9400 16160
rect -9440 16125 -9435 16155
rect -9405 16125 -9400 16155
rect -9440 16120 -9400 16125
rect -9360 16155 -9320 16160
rect -9360 16125 -9355 16155
rect -9325 16125 -9320 16155
rect -9360 16120 -9320 16125
rect -9280 16155 -9240 16160
rect -9280 16125 -9275 16155
rect -9245 16125 -9240 16155
rect -9280 16120 -9240 16125
rect -9200 16155 -9160 16160
rect -9200 16125 -9195 16155
rect -9165 16125 -9160 16155
rect -9200 16120 -9160 16125
rect -9120 16155 -9080 16160
rect -9120 16125 -9115 16155
rect -9085 16125 -9080 16155
rect -9120 16120 -9080 16125
rect -9040 16155 -9000 16160
rect -9040 16125 -9035 16155
rect -9005 16125 -9000 16155
rect -9040 16120 -9000 16125
rect -8960 16155 -8920 16160
rect -8960 16125 -8955 16155
rect -8925 16125 -8920 16155
rect -8960 16120 -8920 16125
rect -8880 16155 -8840 16160
rect -8880 16125 -8875 16155
rect -8845 16125 -8840 16155
rect -8880 16120 -8840 16125
rect -8800 16155 -8760 16160
rect -8800 16125 -8795 16155
rect -8765 16125 -8760 16155
rect -8800 16120 -8760 16125
rect -8720 16155 -8680 16160
rect -8720 16125 -8715 16155
rect -8685 16125 -8680 16155
rect -8720 16120 -8680 16125
rect -8640 16155 -8600 16160
rect -8640 16125 -8635 16155
rect -8605 16125 -8600 16155
rect -8640 16120 -8600 16125
rect -8560 16155 -8520 16160
rect -8560 16125 -8555 16155
rect -8525 16125 -8520 16155
rect -8560 16120 -8520 16125
rect -8480 16155 -8440 16160
rect -8480 16125 -8475 16155
rect -8445 16125 -8440 16155
rect -8480 16120 -8440 16125
rect -8400 16155 -8360 16160
rect -8400 16125 -8395 16155
rect -8365 16125 -8360 16155
rect -8400 16120 -8360 16125
rect -8320 16155 -8280 16160
rect -8320 16125 -8315 16155
rect -8285 16125 -8280 16155
rect -8320 16120 -8280 16125
rect -8240 16155 -8200 16160
rect -8240 16125 -8235 16155
rect -8205 16125 -8200 16155
rect -8240 16120 -8200 16125
rect -8160 16155 -8120 16160
rect -8160 16125 -8155 16155
rect -8125 16125 -8120 16155
rect -8160 16120 -8120 16125
rect -8080 16155 -8040 16160
rect -8080 16125 -8075 16155
rect -8045 16125 -8040 16155
rect -8080 16120 -8040 16125
rect -8000 16155 -7960 16160
rect -8000 16125 -7995 16155
rect -7965 16125 -7960 16155
rect -8000 16120 -7960 16125
rect -7920 16155 -7880 16160
rect -7920 16125 -7915 16155
rect -7885 16125 -7880 16155
rect -7920 16120 -7880 16125
rect -7840 16155 -7800 16160
rect -7840 16125 -7835 16155
rect -7805 16125 -7800 16155
rect -7840 16120 -7800 16125
rect -7760 16155 -7720 16160
rect -7760 16125 -7755 16155
rect -7725 16125 -7720 16155
rect -7760 16120 -7720 16125
rect -7680 16155 -7640 16160
rect -7680 16125 -7675 16155
rect -7645 16125 -7640 16155
rect -7680 16120 -7640 16125
rect -7600 16155 -7560 16160
rect -7600 16125 -7595 16155
rect -7565 16125 -7560 16155
rect -7600 16120 -7560 16125
rect -7520 16155 -7480 16160
rect -7520 16125 -7515 16155
rect -7485 16125 -7480 16155
rect -7520 16120 -7480 16125
rect -7440 16155 -7400 16160
rect -7440 16125 -7435 16155
rect -7405 16125 -7400 16155
rect -7440 16120 -7400 16125
rect -7360 16155 -7320 16160
rect -7360 16125 -7355 16155
rect -7325 16125 -7320 16155
rect -7360 16120 -7320 16125
rect -7280 16155 -7240 16160
rect -7280 16125 -7275 16155
rect -7245 16125 -7240 16155
rect -7280 16120 -7240 16125
rect -7200 16155 -7160 16160
rect -7200 16125 -7195 16155
rect -7165 16125 -7160 16155
rect -7200 16120 -7160 16125
rect -7120 16155 -7080 16160
rect -7120 16125 -7115 16155
rect -7085 16125 -7080 16155
rect -7120 16120 -7080 16125
rect -7040 16155 -7000 16160
rect -7040 16125 -7035 16155
rect -7005 16125 -7000 16155
rect -7040 16120 -7000 16125
rect -6960 16155 -6920 16160
rect -6960 16125 -6955 16155
rect -6925 16125 -6920 16155
rect -6960 16120 -6920 16125
rect -6880 16155 -6840 16160
rect -6880 16125 -6875 16155
rect -6845 16125 -6840 16155
rect -6880 16120 -6840 16125
rect -6800 16155 -6760 16160
rect -6800 16125 -6795 16155
rect -6765 16125 -6760 16155
rect -6800 16120 -6760 16125
rect -6720 16155 -6680 16160
rect -6720 16125 -6715 16155
rect -6685 16125 -6680 16155
rect -6720 16120 -6680 16125
rect -6640 16155 -6600 16160
rect -6640 16125 -6635 16155
rect -6605 16125 -6600 16155
rect -6640 16120 -6600 16125
rect -6560 16155 -6520 16160
rect -6560 16125 -6555 16155
rect -6525 16125 -6520 16155
rect -6560 16120 -6520 16125
rect -6480 16155 -6440 16160
rect -6480 16125 -6475 16155
rect -6445 16125 -6440 16155
rect -6480 16120 -6440 16125
rect -6400 16155 -6360 16160
rect -6400 16125 -6395 16155
rect -6365 16125 -6360 16155
rect -6400 16120 -6360 16125
rect -6320 16155 -6280 16160
rect -6320 16125 -6315 16155
rect -6285 16125 -6280 16155
rect -6320 16120 -6280 16125
rect -6240 16155 -6200 16160
rect -6240 16125 -6235 16155
rect -6205 16125 -6200 16155
rect -6240 16120 -6200 16125
rect -6160 16155 -6120 16160
rect -6160 16125 -6155 16155
rect -6125 16125 -6120 16155
rect -6160 16120 -6120 16125
rect -6080 16155 -6040 16160
rect -6080 16125 -6075 16155
rect -6045 16125 -6040 16155
rect -6080 16120 -6040 16125
rect -6000 16155 -5960 16160
rect -6000 16125 -5995 16155
rect -5965 16125 -5960 16155
rect -6000 16120 -5960 16125
rect -5920 16155 -5880 16160
rect -5920 16125 -5915 16155
rect -5885 16125 -5880 16155
rect -5920 16120 -5880 16125
rect -5840 16155 -5800 16160
rect -5840 16125 -5835 16155
rect -5805 16125 -5800 16155
rect -5840 16120 -5800 16125
rect -5760 16155 -5720 16160
rect -5760 16125 -5755 16155
rect -5725 16125 -5720 16155
rect -5760 16120 -5720 16125
rect -5680 16155 -5640 16160
rect -5680 16125 -5675 16155
rect -5645 16125 -5640 16155
rect -5680 16120 -5640 16125
rect -5600 16155 -5560 16160
rect -5600 16125 -5595 16155
rect -5565 16125 -5560 16155
rect -5600 16120 -5560 16125
rect -5440 16155 -5400 16160
rect -5440 16125 -5435 16155
rect -5405 16125 -5400 16155
rect -5440 16120 -5400 16125
rect -5360 16155 -5320 16160
rect -5360 16125 -5355 16155
rect -5325 16125 -5320 16155
rect -5360 16120 -5320 16125
rect -5280 16155 -5240 16160
rect -5280 16125 -5275 16155
rect -5245 16125 -5240 16155
rect -5280 16120 -5240 16125
rect -5200 16155 -5160 16160
rect -5200 16125 -5195 16155
rect -5165 16125 -5160 16155
rect -5200 16120 -5160 16125
rect -5120 16155 -5080 16160
rect -5120 16125 -5115 16155
rect -5085 16125 -5080 16155
rect -5120 16120 -5080 16125
rect -5040 16155 -5000 16160
rect -5040 16125 -5035 16155
rect -5005 16125 -5000 16155
rect -5040 16120 -5000 16125
rect -4960 16155 -4920 16160
rect -4960 16125 -4955 16155
rect -4925 16125 -4920 16155
rect -4960 16120 -4920 16125
rect -4880 16155 -4840 16160
rect -4880 16125 -4875 16155
rect -4845 16125 -4840 16155
rect -4880 16120 -4840 16125
rect -4800 16155 -4760 16160
rect -4800 16125 -4795 16155
rect -4765 16125 -4760 16155
rect -4800 16120 -4760 16125
rect -4720 16155 -4680 16160
rect -4720 16125 -4715 16155
rect -4685 16125 -4680 16155
rect -4720 16120 -4680 16125
rect -4640 16155 -4600 16160
rect -4640 16125 -4635 16155
rect -4605 16125 -4600 16155
rect -4640 16120 -4600 16125
rect -4560 16155 -4520 16160
rect -4560 16125 -4555 16155
rect -4525 16125 -4520 16155
rect -4560 16120 -4520 16125
rect -4480 16155 -4440 16160
rect -4480 16125 -4475 16155
rect -4445 16125 -4440 16155
rect -4480 16120 -4440 16125
rect -4400 16155 -4360 16160
rect -4400 16125 -4395 16155
rect -4365 16125 -4360 16155
rect -4400 16120 -4360 16125
rect -4320 16155 -4280 16160
rect -4320 16125 -4315 16155
rect -4285 16125 -4280 16155
rect -4320 16120 -4280 16125
rect -4240 16155 -4200 16160
rect -4240 16125 -4235 16155
rect -4205 16125 -4200 16155
rect -4240 16120 -4200 16125
rect -4160 16155 -4120 16160
rect -4160 16125 -4155 16155
rect -4125 16125 -4120 16155
rect -4160 16120 -4120 16125
rect -4080 16155 -4040 16160
rect -4080 16125 -4075 16155
rect -4045 16125 -4040 16155
rect -4080 16120 -4040 16125
rect -4000 16155 -3960 16160
rect -4000 16125 -3995 16155
rect -3965 16125 -3960 16155
rect -4000 16120 -3960 16125
rect -3920 16155 -3880 16160
rect -3920 16125 -3915 16155
rect -3885 16125 -3880 16155
rect -3920 16120 -3880 16125
rect -3840 16155 -3800 16160
rect -3840 16125 -3835 16155
rect -3805 16125 -3800 16155
rect -3840 16120 -3800 16125
rect -3760 16155 -3720 16160
rect -3760 16125 -3755 16155
rect -3725 16125 -3720 16155
rect -3760 16120 -3720 16125
rect -3680 16155 -3640 16160
rect -3680 16125 -3675 16155
rect -3645 16125 -3640 16155
rect -3680 16120 -3640 16125
rect -3600 16155 -3560 16160
rect -3600 16125 -3595 16155
rect -3565 16125 -3560 16155
rect -3600 16120 -3560 16125
rect -3520 16155 -3480 16160
rect -3520 16125 -3515 16155
rect -3485 16125 -3480 16155
rect -3520 16120 -3480 16125
rect -3440 16155 -3400 16160
rect -3440 16125 -3435 16155
rect -3405 16125 -3400 16155
rect -3440 16120 -3400 16125
rect -3360 16155 -3320 16160
rect -3360 16125 -3355 16155
rect -3325 16125 -3320 16155
rect -3360 16120 -3320 16125
rect -3280 16155 -3240 16160
rect -3280 16125 -3275 16155
rect -3245 16125 -3240 16155
rect -3280 16120 -3240 16125
rect -3200 16155 -3160 16160
rect -3200 16125 -3195 16155
rect -3165 16125 -3160 16155
rect -3200 16120 -3160 16125
rect -3120 16155 -3080 16160
rect -3120 16125 -3115 16155
rect -3085 16125 -3080 16155
rect -3120 16120 -3080 16125
rect -3040 16155 -3000 16160
rect -3040 16125 -3035 16155
rect -3005 16125 -3000 16155
rect -3040 16120 -3000 16125
rect -2960 16155 -2920 16160
rect -2960 16125 -2955 16155
rect -2925 16125 -2920 16155
rect -2960 16120 -2920 16125
rect -2880 16155 -2840 16160
rect -2880 16125 -2875 16155
rect -2845 16125 -2840 16155
rect -2880 16120 -2840 16125
rect -2800 16155 -2760 16160
rect -2800 16125 -2795 16155
rect -2765 16125 -2760 16155
rect -2800 16120 -2760 16125
rect -2720 16155 -2680 16160
rect -2720 16125 -2715 16155
rect -2685 16125 -2680 16155
rect -2720 16120 -2680 16125
rect -2640 16155 -2600 16160
rect -2640 16125 -2635 16155
rect -2605 16125 -2600 16155
rect -2640 16120 -2600 16125
rect -2560 16155 -2520 16160
rect -2560 16125 -2555 16155
rect -2525 16125 -2520 16155
rect -2560 16120 -2520 16125
rect -2480 16155 -2440 16160
rect -2480 16125 -2475 16155
rect -2445 16125 -2440 16155
rect -2480 16120 -2440 16125
rect -2400 16155 -2360 16160
rect -2400 16125 -2395 16155
rect -2365 16125 -2360 16155
rect -2400 16120 -2360 16125
rect -2320 16155 -2280 16160
rect -2320 16125 -2315 16155
rect -2285 16125 -2280 16155
rect -2320 16120 -2280 16125
rect -2240 16155 -2200 16160
rect -2240 16125 -2235 16155
rect -2205 16125 -2200 16155
rect -2240 16120 -2200 16125
rect -2160 16155 -2120 16160
rect -2160 16125 -2155 16155
rect -2125 16125 -2120 16155
rect -2160 16120 -2120 16125
rect -2080 16155 -2040 16160
rect -2080 16125 -2075 16155
rect -2045 16125 -2040 16155
rect -2080 16120 -2040 16125
rect -2000 16155 -1960 16160
rect -2000 16125 -1995 16155
rect -1965 16125 -1960 16155
rect -2000 16120 -1960 16125
rect -1840 16155 -1800 16160
rect -1840 16125 -1835 16155
rect -1805 16125 -1800 16155
rect -1840 16120 -1800 16125
rect -1760 16155 -1720 16160
rect -1760 16125 -1755 16155
rect -1725 16125 -1720 16155
rect -1760 16120 -1720 16125
rect -1680 16155 -1640 16160
rect -1680 16125 -1675 16155
rect -1645 16125 -1640 16155
rect -1680 16120 -1640 16125
rect -1600 16155 -1560 16160
rect -1600 16125 -1595 16155
rect -1565 16125 -1560 16155
rect -1600 16120 -1560 16125
rect -1520 16155 -1480 16160
rect -1520 16125 -1515 16155
rect -1485 16125 -1480 16155
rect -1520 16120 -1480 16125
rect -1440 16155 -1400 16160
rect -1440 16125 -1435 16155
rect -1405 16125 -1400 16155
rect -1440 16120 -1400 16125
rect -1360 16155 -1320 16160
rect -1360 16125 -1355 16155
rect -1325 16125 -1320 16155
rect -1360 16120 -1320 16125
rect -1200 16155 -1160 16160
rect -1200 16125 -1195 16155
rect -1165 16125 -1160 16155
rect -1200 16120 -1160 16125
rect -1040 16155 -1000 16160
rect -1040 16125 -1035 16155
rect -1005 16125 -1000 16155
rect -1040 16120 -1000 16125
rect -880 16155 -840 16160
rect -880 16125 -875 16155
rect -845 16125 -840 16155
rect -880 16120 -840 16125
rect -720 16155 -680 16160
rect -720 16125 -715 16155
rect -685 16125 -680 16155
rect -720 16120 -680 16125
rect -560 16155 -520 16160
rect -560 16125 -555 16155
rect -525 16125 -520 16155
rect -560 16120 -520 16125
rect -5520 16040 -5480 16080
rect -14960 15995 -14920 16000
rect -14960 15965 -14955 15995
rect -14925 15965 -14920 15995
rect -14960 15960 -14920 15965
rect -14880 15995 -14840 16000
rect -14880 15965 -14875 15995
rect -14845 15965 -14840 15995
rect -14880 15960 -14840 15965
rect -14800 15995 -14760 16000
rect -14800 15965 -14795 15995
rect -14765 15965 -14760 15995
rect -14800 15960 -14760 15965
rect -14720 15995 -14680 16000
rect -14720 15965 -14715 15995
rect -14685 15965 -14680 15995
rect -14720 15960 -14680 15965
rect -14640 15995 -14600 16000
rect -14640 15965 -14635 15995
rect -14605 15965 -14600 15995
rect -14640 15960 -14600 15965
rect -14560 15995 -14520 16000
rect -14560 15965 -14555 15995
rect -14525 15965 -14520 15995
rect -14560 15960 -14520 15965
rect -14480 15995 -14440 16000
rect -14480 15965 -14475 15995
rect -14445 15965 -14440 15995
rect -14480 15960 -14440 15965
rect -14400 15995 -14360 16000
rect -14400 15965 -14395 15995
rect -14365 15965 -14360 15995
rect -14400 15960 -14360 15965
rect -14320 15995 -14280 16000
rect -14320 15965 -14315 15995
rect -14285 15965 -14280 15995
rect -14320 15960 -14280 15965
rect -14240 15995 -14200 16000
rect -14240 15965 -14235 15995
rect -14205 15965 -14200 15995
rect -14240 15960 -14200 15965
rect -14160 15995 -14120 16000
rect -14160 15965 -14155 15995
rect -14125 15965 -14120 15995
rect -14160 15960 -14120 15965
rect -14080 15995 -14040 16000
rect -14080 15965 -14075 15995
rect -14045 15965 -14040 15995
rect -14080 15960 -14040 15965
rect -14000 15995 -13960 16000
rect -14000 15965 -13995 15995
rect -13965 15965 -13960 15995
rect -14000 15960 -13960 15965
rect -13920 15995 -13880 16000
rect -13920 15965 -13915 15995
rect -13885 15965 -13880 15995
rect -13920 15960 -13880 15965
rect -13840 15995 -13800 16000
rect -13840 15965 -13835 15995
rect -13805 15965 -13800 15995
rect -13840 15960 -13800 15965
rect -13760 15995 -13720 16000
rect -13760 15965 -13755 15995
rect -13725 15965 -13720 15995
rect -13760 15960 -13720 15965
rect -13680 15995 -13640 16000
rect -13680 15965 -13675 15995
rect -13645 15965 -13640 15995
rect -13680 15960 -13640 15965
rect -13600 15995 -13560 16000
rect -13600 15965 -13595 15995
rect -13565 15965 -13560 15995
rect -13600 15960 -13560 15965
rect -13520 15995 -13480 16000
rect -13520 15965 -13515 15995
rect -13485 15965 -13480 15995
rect -13520 15960 -13480 15965
rect -13440 15995 -13400 16000
rect -13440 15965 -13435 15995
rect -13405 15965 -13400 15995
rect -13440 15960 -13400 15965
rect -13360 15995 -13320 16000
rect -13360 15965 -13355 15995
rect -13325 15965 -13320 15995
rect -13360 15960 -13320 15965
rect -13280 15995 -13240 16000
rect -13280 15965 -13275 15995
rect -13245 15965 -13240 15995
rect -13280 15960 -13240 15965
rect -13200 15995 -13160 16000
rect -13200 15965 -13195 15995
rect -13165 15965 -13160 15995
rect -13200 15960 -13160 15965
rect -13120 15995 -13080 16000
rect -13120 15965 -13115 15995
rect -13085 15965 -13080 15995
rect -13120 15960 -13080 15965
rect -13040 15995 -13000 16000
rect -13040 15965 -13035 15995
rect -13005 15965 -13000 15995
rect -13040 15960 -13000 15965
rect -12960 15995 -12920 16000
rect -12960 15965 -12955 15995
rect -12925 15965 -12920 15995
rect -12960 15960 -12920 15965
rect -12880 15995 -12840 16000
rect -12880 15965 -12875 15995
rect -12845 15965 -12840 15995
rect -12880 15960 -12840 15965
rect -12800 15995 -12760 16000
rect -12800 15965 -12795 15995
rect -12765 15965 -12760 15995
rect -12800 15960 -12760 15965
rect -12720 15995 -12680 16000
rect -12720 15965 -12715 15995
rect -12685 15965 -12680 15995
rect -12720 15960 -12680 15965
rect -12640 15995 -12600 16000
rect -12640 15965 -12635 15995
rect -12605 15965 -12600 15995
rect -12640 15960 -12600 15965
rect -12560 15995 -12520 16000
rect -12560 15965 -12555 15995
rect -12525 15965 -12520 15995
rect -12560 15960 -12520 15965
rect -12480 15995 -12440 16000
rect -12480 15965 -12475 15995
rect -12445 15965 -12440 15995
rect -12480 15960 -12440 15965
rect -12400 15995 -12360 16000
rect -12400 15965 -12395 15995
rect -12365 15965 -12360 15995
rect -12400 15960 -12360 15965
rect -12320 15995 -12280 16000
rect -12320 15965 -12315 15995
rect -12285 15965 -12280 15995
rect -12320 15960 -12280 15965
rect -12240 15995 -12200 16000
rect -12240 15965 -12235 15995
rect -12205 15965 -12200 15995
rect -12240 15960 -12200 15965
rect -12160 15995 -12120 16000
rect -12160 15965 -12155 15995
rect -12125 15965 -12120 15995
rect -12160 15960 -12120 15965
rect -12080 15995 -12040 16000
rect -12080 15965 -12075 15995
rect -12045 15965 -12040 15995
rect -12080 15960 -12040 15965
rect -12000 15995 -11960 16000
rect -12000 15965 -11995 15995
rect -11965 15965 -11960 15995
rect -12000 15960 -11960 15965
rect -11920 15995 -11880 16000
rect -11920 15965 -11915 15995
rect -11885 15965 -11880 15995
rect -11920 15960 -11880 15965
rect -11840 15995 -11800 16000
rect -11840 15965 -11835 15995
rect -11805 15965 -11800 15995
rect -11840 15960 -11800 15965
rect -11760 15995 -11720 16000
rect -11760 15965 -11755 15995
rect -11725 15965 -11720 15995
rect -11760 15960 -11720 15965
rect -11680 15995 -11640 16000
rect -11680 15965 -11675 15995
rect -11645 15965 -11640 15995
rect -11680 15960 -11640 15965
rect -11600 15995 -11560 16000
rect -11600 15965 -11595 15995
rect -11565 15965 -11560 15995
rect -11600 15960 -11560 15965
rect -11520 15995 -11480 16000
rect -11520 15965 -11515 15995
rect -11485 15965 -11480 15995
rect -11520 15960 -11480 15965
rect -11440 15995 -11400 16000
rect -11440 15965 -11435 15995
rect -11405 15965 -11400 15995
rect -11440 15960 -11400 15965
rect -11360 15995 -11320 16000
rect -11360 15965 -11355 15995
rect -11325 15965 -11320 15995
rect -11360 15960 -11320 15965
rect -11280 15995 -11240 16000
rect -11280 15965 -11275 15995
rect -11245 15965 -11240 15995
rect -11280 15960 -11240 15965
rect -11200 15995 -11160 16000
rect -11200 15965 -11195 15995
rect -11165 15965 -11160 15995
rect -11200 15960 -11160 15965
rect -11120 15995 -11080 16000
rect -11120 15965 -11115 15995
rect -11085 15965 -11080 15995
rect -11120 15960 -11080 15965
rect -11040 15995 -11000 16000
rect -11040 15965 -11035 15995
rect -11005 15965 -11000 15995
rect -11040 15960 -11000 15965
rect -10960 15995 -10920 16000
rect -10960 15965 -10955 15995
rect -10925 15965 -10920 15995
rect -10960 15960 -10920 15965
rect -10880 15995 -10840 16000
rect -10880 15965 -10875 15995
rect -10845 15965 -10840 15995
rect -10880 15960 -10840 15965
rect -10800 15995 -10760 16000
rect -10800 15965 -10795 15995
rect -10765 15965 -10760 15995
rect -10800 15960 -10760 15965
rect -10720 15995 -10680 16000
rect -10720 15965 -10715 15995
rect -10685 15965 -10680 15995
rect -10720 15960 -10680 15965
rect -10640 15995 -10600 16000
rect -10640 15965 -10635 15995
rect -10605 15965 -10600 15995
rect -10640 15960 -10600 15965
rect -10560 15995 -10520 16000
rect -10560 15965 -10555 15995
rect -10525 15965 -10520 15995
rect -10560 15960 -10520 15965
rect -10480 15995 -10440 16000
rect -10480 15965 -10475 15995
rect -10445 15965 -10440 15995
rect -10480 15960 -10440 15965
rect -10400 15995 -10360 16000
rect -10400 15965 -10395 15995
rect -10365 15965 -10360 15995
rect -10400 15960 -10360 15965
rect -10320 15995 -10280 16000
rect -10320 15965 -10315 15995
rect -10285 15965 -10280 15995
rect -10320 15960 -10280 15965
rect -10240 15995 -10200 16000
rect -10240 15965 -10235 15995
rect -10205 15965 -10200 15995
rect -10240 15960 -10200 15965
rect -10160 15995 -10120 16000
rect -10160 15965 -10155 15995
rect -10125 15965 -10120 15995
rect -10160 15960 -10120 15965
rect -10080 15995 -10040 16000
rect -10080 15965 -10075 15995
rect -10045 15965 -10040 15995
rect -10080 15960 -10040 15965
rect -10000 15995 -9960 16000
rect -10000 15965 -9995 15995
rect -9965 15965 -9960 15995
rect -10000 15960 -9960 15965
rect -9920 15995 -9880 16000
rect -9920 15965 -9915 15995
rect -9885 15965 -9880 15995
rect -9920 15960 -9880 15965
rect -9840 15995 -9800 16000
rect -9840 15965 -9835 15995
rect -9805 15965 -9800 15995
rect -9840 15960 -9800 15965
rect -9760 15995 -9720 16000
rect -9760 15965 -9755 15995
rect -9725 15965 -9720 15995
rect -9760 15960 -9720 15965
rect -9680 15995 -9640 16000
rect -9680 15965 -9675 15995
rect -9645 15965 -9640 15995
rect -9680 15960 -9640 15965
rect -9600 15995 -9560 16000
rect -9600 15965 -9595 15995
rect -9565 15965 -9560 15995
rect -9600 15960 -9560 15965
rect -9520 15995 -9480 16000
rect -9520 15965 -9515 15995
rect -9485 15965 -9480 15995
rect -9520 15960 -9480 15965
rect -9440 15995 -9400 16000
rect -9440 15965 -9435 15995
rect -9405 15965 -9400 15995
rect -9440 15960 -9400 15965
rect -9360 15995 -9320 16000
rect -9360 15965 -9355 15995
rect -9325 15965 -9320 15995
rect -9360 15960 -9320 15965
rect -9280 15995 -9240 16000
rect -9280 15965 -9275 15995
rect -9245 15965 -9240 15995
rect -9280 15960 -9240 15965
rect -9200 15995 -9160 16000
rect -9200 15965 -9195 15995
rect -9165 15965 -9160 15995
rect -9200 15960 -9160 15965
rect -9120 15995 -9080 16000
rect -9120 15965 -9115 15995
rect -9085 15965 -9080 15995
rect -9120 15960 -9080 15965
rect -9040 15995 -9000 16000
rect -9040 15965 -9035 15995
rect -9005 15965 -9000 15995
rect -9040 15960 -9000 15965
rect -8960 15995 -8920 16000
rect -8960 15965 -8955 15995
rect -8925 15965 -8920 15995
rect -8960 15960 -8920 15965
rect -8880 15995 -8840 16000
rect -8880 15965 -8875 15995
rect -8845 15965 -8840 15995
rect -8880 15960 -8840 15965
rect -8800 15995 -8760 16000
rect -8800 15965 -8795 15995
rect -8765 15965 -8760 15995
rect -8800 15960 -8760 15965
rect -8720 15995 -8680 16000
rect -8720 15965 -8715 15995
rect -8685 15965 -8680 15995
rect -8720 15960 -8680 15965
rect -8640 15995 -8600 16000
rect -8640 15965 -8635 15995
rect -8605 15965 -8600 15995
rect -8640 15960 -8600 15965
rect -8560 15995 -8520 16000
rect -8560 15965 -8555 15995
rect -8525 15965 -8520 15995
rect -8560 15960 -8520 15965
rect -8480 15995 -8440 16000
rect -8480 15965 -8475 15995
rect -8445 15965 -8440 15995
rect -8480 15960 -8440 15965
rect -8400 15995 -8360 16000
rect -8400 15965 -8395 15995
rect -8365 15965 -8360 15995
rect -8400 15960 -8360 15965
rect -8320 15995 -8280 16000
rect -8320 15965 -8315 15995
rect -8285 15965 -8280 15995
rect -8320 15960 -8280 15965
rect -8240 15995 -8200 16000
rect -8240 15965 -8235 15995
rect -8205 15965 -8200 15995
rect -8240 15960 -8200 15965
rect -8160 15995 -8120 16000
rect -8160 15965 -8155 15995
rect -8125 15965 -8120 15995
rect -8160 15960 -8120 15965
rect -8080 15995 -8040 16000
rect -8080 15965 -8075 15995
rect -8045 15965 -8040 15995
rect -8080 15960 -8040 15965
rect -8000 15995 -7960 16000
rect -8000 15965 -7995 15995
rect -7965 15965 -7960 15995
rect -8000 15960 -7960 15965
rect -7920 15995 -7880 16000
rect -7920 15965 -7915 15995
rect -7885 15965 -7880 15995
rect -7920 15960 -7880 15965
rect -7840 15995 -7800 16000
rect -7840 15965 -7835 15995
rect -7805 15965 -7800 15995
rect -7840 15960 -7800 15965
rect -7760 15995 -7720 16000
rect -7760 15965 -7755 15995
rect -7725 15965 -7720 15995
rect -7760 15960 -7720 15965
rect -7680 15995 -7640 16000
rect -7680 15965 -7675 15995
rect -7645 15965 -7640 15995
rect -7680 15960 -7640 15965
rect -7600 15995 -7560 16000
rect -7600 15965 -7595 15995
rect -7565 15965 -7560 15995
rect -7600 15960 -7560 15965
rect -7520 15995 -7480 16000
rect -7520 15965 -7515 15995
rect -7485 15965 -7480 15995
rect -7520 15960 -7480 15965
rect -7440 15995 -7400 16000
rect -7440 15965 -7435 15995
rect -7405 15965 -7400 15995
rect -7440 15960 -7400 15965
rect -7360 15995 -7320 16000
rect -7360 15965 -7355 15995
rect -7325 15965 -7320 15995
rect -7360 15960 -7320 15965
rect -7280 15995 -7240 16000
rect -7280 15965 -7275 15995
rect -7245 15965 -7240 15995
rect -7280 15960 -7240 15965
rect -7200 15995 -7160 16000
rect -7200 15965 -7195 15995
rect -7165 15965 -7160 15995
rect -7200 15960 -7160 15965
rect -7120 15995 -7080 16000
rect -7120 15965 -7115 15995
rect -7085 15965 -7080 15995
rect -7120 15960 -7080 15965
rect -7040 15995 -7000 16000
rect -7040 15965 -7035 15995
rect -7005 15965 -7000 15995
rect -7040 15960 -7000 15965
rect -6960 15995 -6920 16000
rect -6960 15965 -6955 15995
rect -6925 15965 -6920 15995
rect -6960 15960 -6920 15965
rect -6880 15995 -6840 16000
rect -6880 15965 -6875 15995
rect -6845 15965 -6840 15995
rect -6880 15960 -6840 15965
rect -6800 15995 -6760 16000
rect -6800 15965 -6795 15995
rect -6765 15965 -6760 15995
rect -6800 15960 -6760 15965
rect -6720 15995 -6680 16000
rect -6720 15965 -6715 15995
rect -6685 15965 -6680 15995
rect -6720 15960 -6680 15965
rect -6640 15995 -6600 16000
rect -6640 15965 -6635 15995
rect -6605 15965 -6600 15995
rect -6640 15960 -6600 15965
rect -6560 15995 -6520 16000
rect -6560 15965 -6555 15995
rect -6525 15965 -6520 15995
rect -6560 15960 -6520 15965
rect -6480 15995 -6440 16000
rect -6480 15965 -6475 15995
rect -6445 15965 -6440 15995
rect -6480 15960 -6440 15965
rect -6400 15995 -6360 16000
rect -6400 15965 -6395 15995
rect -6365 15965 -6360 15995
rect -6400 15960 -6360 15965
rect -6320 15995 -6280 16000
rect -6320 15965 -6315 15995
rect -6285 15965 -6280 15995
rect -6320 15960 -6280 15965
rect -6240 15995 -6200 16000
rect -6240 15965 -6235 15995
rect -6205 15965 -6200 15995
rect -6240 15960 -6200 15965
rect -6160 15995 -6120 16000
rect -6160 15965 -6155 15995
rect -6125 15965 -6120 15995
rect -6160 15960 -6120 15965
rect -6080 15995 -6040 16000
rect -6080 15965 -6075 15995
rect -6045 15965 -6040 15995
rect -6080 15960 -6040 15965
rect -6000 15995 -5960 16000
rect -6000 15965 -5995 15995
rect -5965 15965 -5960 15995
rect -6000 15960 -5960 15965
rect -5920 15995 -5880 16000
rect -5920 15965 -5915 15995
rect -5885 15965 -5880 15995
rect -5920 15960 -5880 15965
rect -5840 15995 -5800 16000
rect -5840 15965 -5835 15995
rect -5805 15965 -5800 15995
rect -5840 15960 -5800 15965
rect -5760 15995 -5720 16000
rect -5760 15965 -5755 15995
rect -5725 15965 -5720 15995
rect -5760 15960 -5720 15965
rect -5680 15995 -5640 16000
rect -5680 15965 -5675 15995
rect -5645 15965 -5640 15995
rect -5680 15960 -5640 15965
rect -5600 15995 -5560 16000
rect -5600 15965 -5595 15995
rect -5565 15965 -5560 15995
rect -5600 15960 -5560 15965
rect -5440 15995 -5400 16000
rect -5440 15965 -5435 15995
rect -5405 15965 -5400 15995
rect -5440 15960 -5400 15965
rect -5360 15995 -5320 16000
rect -5360 15965 -5355 15995
rect -5325 15965 -5320 15995
rect -5360 15960 -5320 15965
rect -5280 15995 -5240 16000
rect -5280 15965 -5275 15995
rect -5245 15965 -5240 15995
rect -5280 15960 -5240 15965
rect -5200 15995 -5160 16000
rect -5200 15965 -5195 15995
rect -5165 15965 -5160 15995
rect -5200 15960 -5160 15965
rect -5120 15995 -5080 16000
rect -5120 15965 -5115 15995
rect -5085 15965 -5080 15995
rect -5120 15960 -5080 15965
rect -5040 15995 -5000 16000
rect -5040 15965 -5035 15995
rect -5005 15965 -5000 15995
rect -5040 15960 -5000 15965
rect -4960 15995 -4920 16000
rect -4960 15965 -4955 15995
rect -4925 15965 -4920 15995
rect -4960 15960 -4920 15965
rect -4880 15995 -4840 16000
rect -4880 15965 -4875 15995
rect -4845 15965 -4840 15995
rect -4880 15960 -4840 15965
rect -4800 15995 -4760 16000
rect -4800 15965 -4795 15995
rect -4765 15965 -4760 15995
rect -4800 15960 -4760 15965
rect -4720 15995 -4680 16000
rect -4720 15965 -4715 15995
rect -4685 15965 -4680 15995
rect -4720 15960 -4680 15965
rect -4640 15995 -4600 16000
rect -4640 15965 -4635 15995
rect -4605 15965 -4600 15995
rect -4640 15960 -4600 15965
rect -4560 15995 -4520 16000
rect -4560 15965 -4555 15995
rect -4525 15965 -4520 15995
rect -4560 15960 -4520 15965
rect -4480 15995 -4440 16000
rect -4480 15965 -4475 15995
rect -4445 15965 -4440 15995
rect -4480 15960 -4440 15965
rect -4400 15995 -4360 16000
rect -4400 15965 -4395 15995
rect -4365 15965 -4360 15995
rect -4400 15960 -4360 15965
rect -4320 15995 -4280 16000
rect -4320 15965 -4315 15995
rect -4285 15965 -4280 15995
rect -4320 15960 -4280 15965
rect -4240 15995 -4200 16000
rect -4240 15965 -4235 15995
rect -4205 15965 -4200 15995
rect -4240 15960 -4200 15965
rect -4160 15995 -4120 16000
rect -4160 15965 -4155 15995
rect -4125 15965 -4120 15995
rect -4160 15960 -4120 15965
rect -4080 15995 -4040 16000
rect -4080 15965 -4075 15995
rect -4045 15965 -4040 15995
rect -4080 15960 -4040 15965
rect -4000 15995 -3960 16000
rect -4000 15965 -3995 15995
rect -3965 15965 -3960 15995
rect -4000 15960 -3960 15965
rect -3920 15995 -3880 16000
rect -3920 15965 -3915 15995
rect -3885 15965 -3880 15995
rect -3920 15960 -3880 15965
rect -3840 15995 -3800 16000
rect -3840 15965 -3835 15995
rect -3805 15965 -3800 15995
rect -3840 15960 -3800 15965
rect -3760 15995 -3720 16000
rect -3760 15965 -3755 15995
rect -3725 15965 -3720 15995
rect -3760 15960 -3720 15965
rect -3680 15995 -3640 16000
rect -3680 15965 -3675 15995
rect -3645 15965 -3640 15995
rect -3680 15960 -3640 15965
rect -3600 15995 -3560 16000
rect -3600 15965 -3595 15995
rect -3565 15965 -3560 15995
rect -3600 15960 -3560 15965
rect -3520 15995 -3480 16000
rect -3520 15965 -3515 15995
rect -3485 15965 -3480 15995
rect -3520 15960 -3480 15965
rect -3440 15995 -3400 16000
rect -3440 15965 -3435 15995
rect -3405 15965 -3400 15995
rect -3440 15960 -3400 15965
rect -3360 15995 -3320 16000
rect -3360 15965 -3355 15995
rect -3325 15965 -3320 15995
rect -3360 15960 -3320 15965
rect -3280 15995 -3240 16000
rect -3280 15965 -3275 15995
rect -3245 15965 -3240 15995
rect -3280 15960 -3240 15965
rect -3200 15995 -3160 16000
rect -3200 15965 -3195 15995
rect -3165 15965 -3160 15995
rect -3200 15960 -3160 15965
rect -3120 15995 -3080 16000
rect -3120 15965 -3115 15995
rect -3085 15965 -3080 15995
rect -3120 15960 -3080 15965
rect -3040 15995 -3000 16000
rect -3040 15965 -3035 15995
rect -3005 15965 -3000 15995
rect -3040 15960 -3000 15965
rect -2960 15995 -2920 16000
rect -2960 15965 -2955 15995
rect -2925 15965 -2920 15995
rect -2960 15960 -2920 15965
rect -2880 15995 -2840 16000
rect -2880 15965 -2875 15995
rect -2845 15965 -2840 15995
rect -2880 15960 -2840 15965
rect -2800 15995 -2760 16000
rect -2800 15965 -2795 15995
rect -2765 15965 -2760 15995
rect -2800 15960 -2760 15965
rect -2720 15995 -2680 16000
rect -2720 15965 -2715 15995
rect -2685 15965 -2680 15995
rect -2720 15960 -2680 15965
rect -2640 15995 -2600 16000
rect -2640 15965 -2635 15995
rect -2605 15965 -2600 15995
rect -2640 15960 -2600 15965
rect -2560 15995 -2520 16000
rect -2560 15965 -2555 15995
rect -2525 15965 -2520 15995
rect -2560 15960 -2520 15965
rect -2480 15995 -2440 16000
rect -2480 15965 -2475 15995
rect -2445 15965 -2440 15995
rect -2480 15960 -2440 15965
rect -2400 15995 -2360 16000
rect -2400 15965 -2395 15995
rect -2365 15965 -2360 15995
rect -2400 15960 -2360 15965
rect -2320 15995 -2280 16000
rect -2320 15965 -2315 15995
rect -2285 15965 -2280 15995
rect -2320 15960 -2280 15965
rect -2240 15995 -2200 16000
rect -2240 15965 -2235 15995
rect -2205 15965 -2200 15995
rect -2240 15960 -2200 15965
rect -2160 15995 -2120 16000
rect -2160 15965 -2155 15995
rect -2125 15965 -2120 15995
rect -2160 15960 -2120 15965
rect -2080 15995 -2040 16000
rect -2080 15965 -2075 15995
rect -2045 15965 -2040 15995
rect -2080 15960 -2040 15965
rect -2000 15995 -1960 16000
rect -2000 15965 -1995 15995
rect -1965 15965 -1960 15995
rect -2000 15960 -1960 15965
rect -1840 15995 -1800 16000
rect -1840 15965 -1835 15995
rect -1805 15965 -1800 15995
rect -1840 15960 -1800 15965
rect -1760 15995 -1720 16000
rect -1760 15965 -1755 15995
rect -1725 15965 -1720 15995
rect -1760 15960 -1720 15965
rect -1680 15995 -1640 16000
rect -1680 15965 -1675 15995
rect -1645 15965 -1640 15995
rect -1680 15960 -1640 15965
rect -1600 15995 -1560 16000
rect -1600 15965 -1595 15995
rect -1565 15965 -1560 15995
rect -1600 15960 -1560 15965
rect -1520 15995 -1480 16000
rect -1520 15965 -1515 15995
rect -1485 15965 -1480 15995
rect -1520 15960 -1480 15965
rect -1440 15995 -1400 16000
rect -1440 15965 -1435 15995
rect -1405 15965 -1400 15995
rect -1440 15960 -1400 15965
rect -1360 15995 -1320 16000
rect -1360 15965 -1355 15995
rect -1325 15965 -1320 15995
rect -1360 15960 -1320 15965
rect -1200 15995 -1160 16000
rect -1200 15965 -1195 15995
rect -1165 15965 -1160 15995
rect -1200 15960 -1160 15965
rect -1040 15995 -1000 16000
rect -1040 15965 -1035 15995
rect -1005 15965 -1000 15995
rect -1040 15960 -1000 15965
rect -880 15995 -840 16000
rect -880 15965 -875 15995
rect -845 15965 -840 15995
rect -880 15960 -840 15965
rect -720 15995 -680 16000
rect -720 15965 -715 15995
rect -685 15965 -680 15995
rect -720 15960 -680 15965
rect -560 15995 -520 16000
rect -560 15965 -555 15995
rect -525 15965 -520 15995
rect -560 15960 -520 15965
<< via1 >>
rect -14955 21430 -14925 21435
rect -14955 21410 -14950 21430
rect -14950 21410 -14930 21430
rect -14930 21410 -14925 21430
rect -14955 21405 -14925 21410
rect -14875 21430 -14845 21435
rect -14875 21410 -14870 21430
rect -14870 21410 -14850 21430
rect -14850 21410 -14845 21430
rect -14875 21405 -14845 21410
rect -14795 21430 -14765 21435
rect -14795 21410 -14790 21430
rect -14790 21410 -14770 21430
rect -14770 21410 -14765 21430
rect -14795 21405 -14765 21410
rect -14715 21430 -14685 21435
rect -14715 21410 -14710 21430
rect -14710 21410 -14690 21430
rect -14690 21410 -14685 21430
rect -14715 21405 -14685 21410
rect -14635 21430 -14605 21435
rect -14635 21410 -14630 21430
rect -14630 21410 -14610 21430
rect -14610 21410 -14605 21430
rect -14635 21405 -14605 21410
rect -14555 21430 -14525 21435
rect -14555 21410 -14550 21430
rect -14550 21410 -14530 21430
rect -14530 21410 -14525 21430
rect -14555 21405 -14525 21410
rect -14475 21430 -14445 21435
rect -14475 21410 -14470 21430
rect -14470 21410 -14450 21430
rect -14450 21410 -14445 21430
rect -14475 21405 -14445 21410
rect -14395 21430 -14365 21435
rect -14395 21410 -14390 21430
rect -14390 21410 -14370 21430
rect -14370 21410 -14365 21430
rect -14395 21405 -14365 21410
rect -14315 21430 -14285 21435
rect -14315 21410 -14310 21430
rect -14310 21410 -14290 21430
rect -14290 21410 -14285 21430
rect -14315 21405 -14285 21410
rect -14235 21430 -14205 21435
rect -14235 21410 -14230 21430
rect -14230 21410 -14210 21430
rect -14210 21410 -14205 21430
rect -14235 21405 -14205 21410
rect -14155 21430 -14125 21435
rect -14155 21410 -14150 21430
rect -14150 21410 -14130 21430
rect -14130 21410 -14125 21430
rect -14155 21405 -14125 21410
rect -14075 21430 -14045 21435
rect -14075 21410 -14070 21430
rect -14070 21410 -14050 21430
rect -14050 21410 -14045 21430
rect -14075 21405 -14045 21410
rect -13995 21430 -13965 21435
rect -13995 21410 -13990 21430
rect -13990 21410 -13970 21430
rect -13970 21410 -13965 21430
rect -13995 21405 -13965 21410
rect -13915 21430 -13885 21435
rect -13915 21410 -13910 21430
rect -13910 21410 -13890 21430
rect -13890 21410 -13885 21430
rect -13915 21405 -13885 21410
rect -13835 21430 -13805 21435
rect -13835 21410 -13830 21430
rect -13830 21410 -13810 21430
rect -13810 21410 -13805 21430
rect -13835 21405 -13805 21410
rect -13755 21430 -13725 21435
rect -13755 21410 -13750 21430
rect -13750 21410 -13730 21430
rect -13730 21410 -13725 21430
rect -13755 21405 -13725 21410
rect -13675 21430 -13645 21435
rect -13675 21410 -13670 21430
rect -13670 21410 -13650 21430
rect -13650 21410 -13645 21430
rect -13675 21405 -13645 21410
rect -13595 21430 -13565 21435
rect -13595 21410 -13590 21430
rect -13590 21410 -13570 21430
rect -13570 21410 -13565 21430
rect -13595 21405 -13565 21410
rect -13515 21430 -13485 21435
rect -13515 21410 -13510 21430
rect -13510 21410 -13490 21430
rect -13490 21410 -13485 21430
rect -13515 21405 -13485 21410
rect -13435 21430 -13405 21435
rect -13435 21410 -13430 21430
rect -13430 21410 -13410 21430
rect -13410 21410 -13405 21430
rect -13435 21405 -13405 21410
rect -13355 21430 -13325 21435
rect -13355 21410 -13350 21430
rect -13350 21410 -13330 21430
rect -13330 21410 -13325 21430
rect -13355 21405 -13325 21410
rect -13275 21430 -13245 21435
rect -13275 21410 -13270 21430
rect -13270 21410 -13250 21430
rect -13250 21410 -13245 21430
rect -13275 21405 -13245 21410
rect -13195 21430 -13165 21435
rect -13195 21410 -13190 21430
rect -13190 21410 -13170 21430
rect -13170 21410 -13165 21430
rect -13195 21405 -13165 21410
rect -13115 21430 -13085 21435
rect -13115 21410 -13110 21430
rect -13110 21410 -13090 21430
rect -13090 21410 -13085 21430
rect -13115 21405 -13085 21410
rect -13035 21430 -13005 21435
rect -13035 21410 -13030 21430
rect -13030 21410 -13010 21430
rect -13010 21410 -13005 21430
rect -13035 21405 -13005 21410
rect -12955 21430 -12925 21435
rect -12955 21410 -12950 21430
rect -12950 21410 -12930 21430
rect -12930 21410 -12925 21430
rect -12955 21405 -12925 21410
rect -12875 21430 -12845 21435
rect -12875 21410 -12870 21430
rect -12870 21410 -12850 21430
rect -12850 21410 -12845 21430
rect -12875 21405 -12845 21410
rect -12795 21430 -12765 21435
rect -12795 21410 -12790 21430
rect -12790 21410 -12770 21430
rect -12770 21410 -12765 21430
rect -12795 21405 -12765 21410
rect -12715 21430 -12685 21435
rect -12715 21410 -12710 21430
rect -12710 21410 -12690 21430
rect -12690 21410 -12685 21430
rect -12715 21405 -12685 21410
rect -12635 21430 -12605 21435
rect -12635 21410 -12630 21430
rect -12630 21410 -12610 21430
rect -12610 21410 -12605 21430
rect -12635 21405 -12605 21410
rect -12555 21430 -12525 21435
rect -12555 21410 -12550 21430
rect -12550 21410 -12530 21430
rect -12530 21410 -12525 21430
rect -12555 21405 -12525 21410
rect -12475 21430 -12445 21435
rect -12475 21410 -12470 21430
rect -12470 21410 -12450 21430
rect -12450 21410 -12445 21430
rect -12475 21405 -12445 21410
rect -12395 21430 -12365 21435
rect -12395 21410 -12390 21430
rect -12390 21410 -12370 21430
rect -12370 21410 -12365 21430
rect -12395 21405 -12365 21410
rect -12315 21430 -12285 21435
rect -12315 21410 -12310 21430
rect -12310 21410 -12290 21430
rect -12290 21410 -12285 21430
rect -12315 21405 -12285 21410
rect -12235 21430 -12205 21435
rect -12235 21410 -12230 21430
rect -12230 21410 -12210 21430
rect -12210 21410 -12205 21430
rect -12235 21405 -12205 21410
rect -12155 21430 -12125 21435
rect -12155 21410 -12150 21430
rect -12150 21410 -12130 21430
rect -12130 21410 -12125 21430
rect -12155 21405 -12125 21410
rect -12075 21430 -12045 21435
rect -12075 21410 -12070 21430
rect -12070 21410 -12050 21430
rect -12050 21410 -12045 21430
rect -12075 21405 -12045 21410
rect -11995 21430 -11965 21435
rect -11995 21410 -11990 21430
rect -11990 21410 -11970 21430
rect -11970 21410 -11965 21430
rect -11995 21405 -11965 21410
rect -11915 21430 -11885 21435
rect -11915 21410 -11910 21430
rect -11910 21410 -11890 21430
rect -11890 21410 -11885 21430
rect -11915 21405 -11885 21410
rect -11835 21430 -11805 21435
rect -11835 21410 -11830 21430
rect -11830 21410 -11810 21430
rect -11810 21410 -11805 21430
rect -11835 21405 -11805 21410
rect -11755 21430 -11725 21435
rect -11755 21410 -11750 21430
rect -11750 21410 -11730 21430
rect -11730 21410 -11725 21430
rect -11755 21405 -11725 21410
rect -11675 21430 -11645 21435
rect -11675 21410 -11670 21430
rect -11670 21410 -11650 21430
rect -11650 21410 -11645 21430
rect -11675 21405 -11645 21410
rect -11595 21430 -11565 21435
rect -11595 21410 -11590 21430
rect -11590 21410 -11570 21430
rect -11570 21410 -11565 21430
rect -11595 21405 -11565 21410
rect -11515 21430 -11485 21435
rect -11515 21410 -11510 21430
rect -11510 21410 -11490 21430
rect -11490 21410 -11485 21430
rect -11515 21405 -11485 21410
rect -11435 21430 -11405 21435
rect -11435 21410 -11430 21430
rect -11430 21410 -11410 21430
rect -11410 21410 -11405 21430
rect -11435 21405 -11405 21410
rect -11355 21430 -11325 21435
rect -11355 21410 -11350 21430
rect -11350 21410 -11330 21430
rect -11330 21410 -11325 21430
rect -11355 21405 -11325 21410
rect -11275 21430 -11245 21435
rect -11275 21410 -11270 21430
rect -11270 21410 -11250 21430
rect -11250 21410 -11245 21430
rect -11275 21405 -11245 21410
rect -11195 21430 -11165 21435
rect -11195 21410 -11190 21430
rect -11190 21410 -11170 21430
rect -11170 21410 -11165 21430
rect -11195 21405 -11165 21410
rect -11115 21430 -11085 21435
rect -11115 21410 -11110 21430
rect -11110 21410 -11090 21430
rect -11090 21410 -11085 21430
rect -11115 21405 -11085 21410
rect -11035 21430 -11005 21435
rect -11035 21410 -11030 21430
rect -11030 21410 -11010 21430
rect -11010 21410 -11005 21430
rect -11035 21405 -11005 21410
rect -10955 21430 -10925 21435
rect -10955 21410 -10950 21430
rect -10950 21410 -10930 21430
rect -10930 21410 -10925 21430
rect -10955 21405 -10925 21410
rect -10875 21430 -10845 21435
rect -10875 21410 -10870 21430
rect -10870 21410 -10850 21430
rect -10850 21410 -10845 21430
rect -10875 21405 -10845 21410
rect -10795 21430 -10765 21435
rect -10795 21410 -10790 21430
rect -10790 21410 -10770 21430
rect -10770 21410 -10765 21430
rect -10795 21405 -10765 21410
rect -10715 21430 -10685 21435
rect -10715 21410 -10710 21430
rect -10710 21410 -10690 21430
rect -10690 21410 -10685 21430
rect -10715 21405 -10685 21410
rect -10635 21430 -10605 21435
rect -10635 21410 -10630 21430
rect -10630 21410 -10610 21430
rect -10610 21410 -10605 21430
rect -10635 21405 -10605 21410
rect -10555 21430 -10525 21435
rect -10555 21410 -10550 21430
rect -10550 21410 -10530 21430
rect -10530 21410 -10525 21430
rect -10555 21405 -10525 21410
rect -10475 21430 -10445 21435
rect -10475 21410 -10470 21430
rect -10470 21410 -10450 21430
rect -10450 21410 -10445 21430
rect -10475 21405 -10445 21410
rect -10395 21430 -10365 21435
rect -10395 21410 -10390 21430
rect -10390 21410 -10370 21430
rect -10370 21410 -10365 21430
rect -10395 21405 -10365 21410
rect -10315 21430 -10285 21435
rect -10315 21410 -10310 21430
rect -10310 21410 -10290 21430
rect -10290 21410 -10285 21430
rect -10315 21405 -10285 21410
rect -10235 21430 -10205 21435
rect -10235 21410 -10230 21430
rect -10230 21410 -10210 21430
rect -10210 21410 -10205 21430
rect -10235 21405 -10205 21410
rect -10155 21430 -10125 21435
rect -10155 21410 -10150 21430
rect -10150 21410 -10130 21430
rect -10130 21410 -10125 21430
rect -10155 21405 -10125 21410
rect -10075 21430 -10045 21435
rect -10075 21410 -10070 21430
rect -10070 21410 -10050 21430
rect -10050 21410 -10045 21430
rect -10075 21405 -10045 21410
rect -9995 21430 -9965 21435
rect -9995 21410 -9990 21430
rect -9990 21410 -9970 21430
rect -9970 21410 -9965 21430
rect -9995 21405 -9965 21410
rect -9915 21430 -9885 21435
rect -9915 21410 -9910 21430
rect -9910 21410 -9890 21430
rect -9890 21410 -9885 21430
rect -9915 21405 -9885 21410
rect -9835 21430 -9805 21435
rect -9835 21410 -9830 21430
rect -9830 21410 -9810 21430
rect -9810 21410 -9805 21430
rect -9835 21405 -9805 21410
rect -9755 21430 -9725 21435
rect -9755 21410 -9750 21430
rect -9750 21410 -9730 21430
rect -9730 21410 -9725 21430
rect -9755 21405 -9725 21410
rect -9675 21430 -9645 21435
rect -9675 21410 -9670 21430
rect -9670 21410 -9650 21430
rect -9650 21410 -9645 21430
rect -9675 21405 -9645 21410
rect -9595 21430 -9565 21435
rect -9595 21410 -9590 21430
rect -9590 21410 -9570 21430
rect -9570 21410 -9565 21430
rect -9595 21405 -9565 21410
rect -9515 21430 -9485 21435
rect -9515 21410 -9510 21430
rect -9510 21410 -9490 21430
rect -9490 21410 -9485 21430
rect -9515 21405 -9485 21410
rect -9435 21430 -9405 21435
rect -9435 21410 -9430 21430
rect -9430 21410 -9410 21430
rect -9410 21410 -9405 21430
rect -9435 21405 -9405 21410
rect -9355 21430 -9325 21435
rect -9355 21410 -9350 21430
rect -9350 21410 -9330 21430
rect -9330 21410 -9325 21430
rect -9355 21405 -9325 21410
rect -9275 21430 -9245 21435
rect -9275 21410 -9270 21430
rect -9270 21410 -9250 21430
rect -9250 21410 -9245 21430
rect -9275 21405 -9245 21410
rect -9195 21430 -9165 21435
rect -9195 21410 -9190 21430
rect -9190 21410 -9170 21430
rect -9170 21410 -9165 21430
rect -9195 21405 -9165 21410
rect -9115 21430 -9085 21435
rect -9115 21410 -9110 21430
rect -9110 21410 -9090 21430
rect -9090 21410 -9085 21430
rect -9115 21405 -9085 21410
rect -9035 21430 -9005 21435
rect -9035 21410 -9030 21430
rect -9030 21410 -9010 21430
rect -9010 21410 -9005 21430
rect -9035 21405 -9005 21410
rect -8955 21430 -8925 21435
rect -8955 21410 -8950 21430
rect -8950 21410 -8930 21430
rect -8930 21410 -8925 21430
rect -8955 21405 -8925 21410
rect -8875 21430 -8845 21435
rect -8875 21410 -8870 21430
rect -8870 21410 -8850 21430
rect -8850 21410 -8845 21430
rect -8875 21405 -8845 21410
rect -8795 21430 -8765 21435
rect -8795 21410 -8790 21430
rect -8790 21410 -8770 21430
rect -8770 21410 -8765 21430
rect -8795 21405 -8765 21410
rect -8715 21430 -8685 21435
rect -8715 21410 -8710 21430
rect -8710 21410 -8690 21430
rect -8690 21410 -8685 21430
rect -8715 21405 -8685 21410
rect -8635 21430 -8605 21435
rect -8635 21410 -8630 21430
rect -8630 21410 -8610 21430
rect -8610 21410 -8605 21430
rect -8635 21405 -8605 21410
rect -8555 21430 -8525 21435
rect -8555 21410 -8550 21430
rect -8550 21410 -8530 21430
rect -8530 21410 -8525 21430
rect -8555 21405 -8525 21410
rect -8475 21430 -8445 21435
rect -8475 21410 -8470 21430
rect -8470 21410 -8450 21430
rect -8450 21410 -8445 21430
rect -8475 21405 -8445 21410
rect -8395 21430 -8365 21435
rect -8395 21410 -8390 21430
rect -8390 21410 -8370 21430
rect -8370 21410 -8365 21430
rect -8395 21405 -8365 21410
rect -8315 21430 -8285 21435
rect -8315 21410 -8310 21430
rect -8310 21410 -8290 21430
rect -8290 21410 -8285 21430
rect -8315 21405 -8285 21410
rect -8235 21430 -8205 21435
rect -8235 21410 -8230 21430
rect -8230 21410 -8210 21430
rect -8210 21410 -8205 21430
rect -8235 21405 -8205 21410
rect -8155 21430 -8125 21435
rect -8155 21410 -8150 21430
rect -8150 21410 -8130 21430
rect -8130 21410 -8125 21430
rect -8155 21405 -8125 21410
rect -8075 21430 -8045 21435
rect -8075 21410 -8070 21430
rect -8070 21410 -8050 21430
rect -8050 21410 -8045 21430
rect -8075 21405 -8045 21410
rect -7995 21430 -7965 21435
rect -7995 21410 -7990 21430
rect -7990 21410 -7970 21430
rect -7970 21410 -7965 21430
rect -7995 21405 -7965 21410
rect -7915 21430 -7885 21435
rect -7915 21410 -7910 21430
rect -7910 21410 -7890 21430
rect -7890 21410 -7885 21430
rect -7915 21405 -7885 21410
rect -7835 21430 -7805 21435
rect -7835 21410 -7830 21430
rect -7830 21410 -7810 21430
rect -7810 21410 -7805 21430
rect -7835 21405 -7805 21410
rect -7755 21430 -7725 21435
rect -7755 21410 -7750 21430
rect -7750 21410 -7730 21430
rect -7730 21410 -7725 21430
rect -7755 21405 -7725 21410
rect -7675 21430 -7645 21435
rect -7675 21410 -7670 21430
rect -7670 21410 -7650 21430
rect -7650 21410 -7645 21430
rect -7675 21405 -7645 21410
rect -7595 21430 -7565 21435
rect -7595 21410 -7590 21430
rect -7590 21410 -7570 21430
rect -7570 21410 -7565 21430
rect -7595 21405 -7565 21410
rect -7515 21430 -7485 21435
rect -7515 21410 -7510 21430
rect -7510 21410 -7490 21430
rect -7490 21410 -7485 21430
rect -7515 21405 -7485 21410
rect -7435 21430 -7405 21435
rect -7435 21410 -7430 21430
rect -7430 21410 -7410 21430
rect -7410 21410 -7405 21430
rect -7435 21405 -7405 21410
rect -7355 21430 -7325 21435
rect -7355 21410 -7350 21430
rect -7350 21410 -7330 21430
rect -7330 21410 -7325 21430
rect -7355 21405 -7325 21410
rect -7275 21430 -7245 21435
rect -7275 21410 -7270 21430
rect -7270 21410 -7250 21430
rect -7250 21410 -7245 21430
rect -7275 21405 -7245 21410
rect -7195 21430 -7165 21435
rect -7195 21410 -7190 21430
rect -7190 21410 -7170 21430
rect -7170 21410 -7165 21430
rect -7195 21405 -7165 21410
rect -7115 21430 -7085 21435
rect -7115 21410 -7110 21430
rect -7110 21410 -7090 21430
rect -7090 21410 -7085 21430
rect -7115 21405 -7085 21410
rect -7035 21430 -7005 21435
rect -7035 21410 -7030 21430
rect -7030 21410 -7010 21430
rect -7010 21410 -7005 21430
rect -7035 21405 -7005 21410
rect -6955 21430 -6925 21435
rect -6955 21410 -6950 21430
rect -6950 21410 -6930 21430
rect -6930 21410 -6925 21430
rect -6955 21405 -6925 21410
rect -6875 21430 -6845 21435
rect -6875 21410 -6870 21430
rect -6870 21410 -6850 21430
rect -6850 21410 -6845 21430
rect -6875 21405 -6845 21410
rect -6795 21430 -6765 21435
rect -6795 21410 -6790 21430
rect -6790 21410 -6770 21430
rect -6770 21410 -6765 21430
rect -6795 21405 -6765 21410
rect -6715 21430 -6685 21435
rect -6715 21410 -6710 21430
rect -6710 21410 -6690 21430
rect -6690 21410 -6685 21430
rect -6715 21405 -6685 21410
rect -6635 21430 -6605 21435
rect -6635 21410 -6630 21430
rect -6630 21410 -6610 21430
rect -6610 21410 -6605 21430
rect -6635 21405 -6605 21410
rect -6555 21430 -6525 21435
rect -6555 21410 -6550 21430
rect -6550 21410 -6530 21430
rect -6530 21410 -6525 21430
rect -6555 21405 -6525 21410
rect -6475 21430 -6445 21435
rect -6475 21410 -6470 21430
rect -6470 21410 -6450 21430
rect -6450 21410 -6445 21430
rect -6475 21405 -6445 21410
rect -6395 21430 -6365 21435
rect -6395 21410 -6390 21430
rect -6390 21410 -6370 21430
rect -6370 21410 -6365 21430
rect -6395 21405 -6365 21410
rect -6315 21430 -6285 21435
rect -6315 21410 -6310 21430
rect -6310 21410 -6290 21430
rect -6290 21410 -6285 21430
rect -6315 21405 -6285 21410
rect -6235 21430 -6205 21435
rect -6235 21410 -6230 21430
rect -6230 21410 -6210 21430
rect -6210 21410 -6205 21430
rect -6235 21405 -6205 21410
rect -6155 21430 -6125 21435
rect -6155 21410 -6150 21430
rect -6150 21410 -6130 21430
rect -6130 21410 -6125 21430
rect -6155 21405 -6125 21410
rect -5675 21430 -5645 21435
rect -5675 21410 -5670 21430
rect -5670 21410 -5650 21430
rect -5650 21410 -5645 21430
rect -5675 21405 -5645 21410
rect -5595 21430 -5565 21435
rect -5595 21410 -5590 21430
rect -5590 21410 -5570 21430
rect -5570 21410 -5565 21430
rect -5595 21405 -5565 21410
rect -5515 21430 -5485 21435
rect -5515 21410 -5510 21430
rect -5510 21410 -5490 21430
rect -5490 21410 -5485 21430
rect -5515 21405 -5485 21410
rect -5435 21430 -5405 21435
rect -5435 21410 -5430 21430
rect -5430 21410 -5410 21430
rect -5410 21410 -5405 21430
rect -5435 21405 -5405 21410
rect -5355 21430 -5325 21435
rect -5355 21410 -5350 21430
rect -5350 21410 -5330 21430
rect -5330 21410 -5325 21430
rect -5355 21405 -5325 21410
rect -5275 21430 -5245 21435
rect -5275 21410 -5270 21430
rect -5270 21410 -5250 21430
rect -5250 21410 -5245 21430
rect -5275 21405 -5245 21410
rect -5195 21430 -5165 21435
rect -5195 21410 -5190 21430
rect -5190 21410 -5170 21430
rect -5170 21410 -5165 21430
rect -5195 21405 -5165 21410
rect -5115 21430 -5085 21435
rect -5115 21410 -5110 21430
rect -5110 21410 -5090 21430
rect -5090 21410 -5085 21430
rect -5115 21405 -5085 21410
rect -5035 21430 -5005 21435
rect -5035 21410 -5030 21430
rect -5030 21410 -5010 21430
rect -5010 21410 -5005 21430
rect -5035 21405 -5005 21410
rect -4955 21430 -4925 21435
rect -4955 21410 -4950 21430
rect -4950 21410 -4930 21430
rect -4930 21410 -4925 21430
rect -4955 21405 -4925 21410
rect -4875 21430 -4845 21435
rect -4875 21410 -4870 21430
rect -4870 21410 -4850 21430
rect -4850 21410 -4845 21430
rect -4875 21405 -4845 21410
rect -4795 21430 -4765 21435
rect -4795 21410 -4790 21430
rect -4790 21410 -4770 21430
rect -4770 21410 -4765 21430
rect -4795 21405 -4765 21410
rect -4715 21430 -4685 21435
rect -4715 21410 -4710 21430
rect -4710 21410 -4690 21430
rect -4690 21410 -4685 21430
rect -4715 21405 -4685 21410
rect -4635 21430 -4605 21435
rect -4635 21410 -4630 21430
rect -4630 21410 -4610 21430
rect -4610 21410 -4605 21430
rect -4635 21405 -4605 21410
rect -4555 21430 -4525 21435
rect -4555 21410 -4550 21430
rect -4550 21410 -4530 21430
rect -4530 21410 -4525 21430
rect -4555 21405 -4525 21410
rect -4475 21430 -4445 21435
rect -4475 21410 -4470 21430
rect -4470 21410 -4450 21430
rect -4450 21410 -4445 21430
rect -4475 21405 -4445 21410
rect -4395 21430 -4365 21435
rect -4395 21410 -4390 21430
rect -4390 21410 -4370 21430
rect -4370 21410 -4365 21430
rect -4395 21405 -4365 21410
rect -4315 21430 -4285 21435
rect -4315 21410 -4310 21430
rect -4310 21410 -4290 21430
rect -4290 21410 -4285 21430
rect -4315 21405 -4285 21410
rect -4235 21430 -4205 21435
rect -4235 21410 -4230 21430
rect -4230 21410 -4210 21430
rect -4210 21410 -4205 21430
rect -4235 21405 -4205 21410
rect -4155 21430 -4125 21435
rect -4155 21410 -4150 21430
rect -4150 21410 -4130 21430
rect -4130 21410 -4125 21430
rect -4155 21405 -4125 21410
rect -4075 21430 -4045 21435
rect -4075 21410 -4070 21430
rect -4070 21410 -4050 21430
rect -4050 21410 -4045 21430
rect -4075 21405 -4045 21410
rect -3995 21430 -3965 21435
rect -3995 21410 -3990 21430
rect -3990 21410 -3970 21430
rect -3970 21410 -3965 21430
rect -3995 21405 -3965 21410
rect -3915 21430 -3885 21435
rect -3915 21410 -3910 21430
rect -3910 21410 -3890 21430
rect -3890 21410 -3885 21430
rect -3915 21405 -3885 21410
rect -3835 21430 -3805 21435
rect -3835 21410 -3830 21430
rect -3830 21410 -3810 21430
rect -3810 21410 -3805 21430
rect -3835 21405 -3805 21410
rect -3755 21430 -3725 21435
rect -3755 21410 -3750 21430
rect -3750 21410 -3730 21430
rect -3730 21410 -3725 21430
rect -3755 21405 -3725 21410
rect -3675 21430 -3645 21435
rect -3675 21410 -3670 21430
rect -3670 21410 -3650 21430
rect -3650 21410 -3645 21430
rect -3675 21405 -3645 21410
rect -3595 21430 -3565 21435
rect -3595 21410 -3590 21430
rect -3590 21410 -3570 21430
rect -3570 21410 -3565 21430
rect -3595 21405 -3565 21410
rect -3515 21430 -3485 21435
rect -3515 21410 -3510 21430
rect -3510 21410 -3490 21430
rect -3490 21410 -3485 21430
rect -3515 21405 -3485 21410
rect -3435 21430 -3405 21435
rect -3435 21410 -3430 21430
rect -3430 21410 -3410 21430
rect -3410 21410 -3405 21430
rect -3435 21405 -3405 21410
rect -3355 21430 -3325 21435
rect -3355 21410 -3350 21430
rect -3350 21410 -3330 21430
rect -3330 21410 -3325 21430
rect -3355 21405 -3325 21410
rect -3275 21430 -3245 21435
rect -3275 21410 -3270 21430
rect -3270 21410 -3250 21430
rect -3250 21410 -3245 21430
rect -3275 21405 -3245 21410
rect -3195 21430 -3165 21435
rect -3195 21410 -3190 21430
rect -3190 21410 -3170 21430
rect -3170 21410 -3165 21430
rect -3195 21405 -3165 21410
rect -3115 21430 -3085 21435
rect -3115 21410 -3110 21430
rect -3110 21410 -3090 21430
rect -3090 21410 -3085 21430
rect -3115 21405 -3085 21410
rect -3035 21430 -3005 21435
rect -3035 21410 -3030 21430
rect -3030 21410 -3010 21430
rect -3010 21410 -3005 21430
rect -3035 21405 -3005 21410
rect -2955 21430 -2925 21435
rect -2955 21410 -2950 21430
rect -2950 21410 -2930 21430
rect -2930 21410 -2925 21430
rect -2955 21405 -2925 21410
rect -2875 21430 -2845 21435
rect -2875 21410 -2870 21430
rect -2870 21410 -2850 21430
rect -2850 21410 -2845 21430
rect -2875 21405 -2845 21410
rect -2795 21430 -2765 21435
rect -2795 21410 -2790 21430
rect -2790 21410 -2770 21430
rect -2770 21410 -2765 21430
rect -2795 21405 -2765 21410
rect -2715 21430 -2685 21435
rect -2715 21410 -2710 21430
rect -2710 21410 -2690 21430
rect -2690 21410 -2685 21430
rect -2715 21405 -2685 21410
rect -2635 21430 -2605 21435
rect -2635 21410 -2630 21430
rect -2630 21410 -2610 21430
rect -2610 21410 -2605 21430
rect -2635 21405 -2605 21410
rect -2555 21430 -2525 21435
rect -2555 21410 -2550 21430
rect -2550 21410 -2530 21430
rect -2530 21410 -2525 21430
rect -2555 21405 -2525 21410
rect -2475 21430 -2445 21435
rect -2475 21410 -2470 21430
rect -2470 21410 -2450 21430
rect -2450 21410 -2445 21430
rect -2475 21405 -2445 21410
rect -2395 21430 -2365 21435
rect -2395 21410 -2390 21430
rect -2390 21410 -2370 21430
rect -2370 21410 -2365 21430
rect -2395 21405 -2365 21410
rect -2315 21430 -2285 21435
rect -2315 21410 -2310 21430
rect -2310 21410 -2290 21430
rect -2290 21410 -2285 21430
rect -2315 21405 -2285 21410
rect -2235 21430 -2205 21435
rect -2235 21410 -2230 21430
rect -2230 21410 -2210 21430
rect -2210 21410 -2205 21430
rect -2235 21405 -2205 21410
rect -2155 21430 -2125 21435
rect -2155 21410 -2150 21430
rect -2150 21410 -2130 21430
rect -2130 21410 -2125 21430
rect -2155 21405 -2125 21410
rect -2075 21430 -2045 21435
rect -2075 21410 -2070 21430
rect -2070 21410 -2050 21430
rect -2050 21410 -2045 21430
rect -2075 21405 -2045 21410
rect -1995 21430 -1965 21435
rect -1995 21410 -1990 21430
rect -1990 21410 -1970 21430
rect -1970 21410 -1965 21430
rect -1995 21405 -1965 21410
rect -1835 21430 -1805 21435
rect -1835 21410 -1830 21430
rect -1830 21410 -1810 21430
rect -1810 21410 -1805 21430
rect -1835 21405 -1805 21410
rect -1755 21430 -1725 21435
rect -1755 21410 -1750 21430
rect -1750 21410 -1730 21430
rect -1730 21410 -1725 21430
rect -1755 21405 -1725 21410
rect -1675 21430 -1645 21435
rect -1675 21410 -1670 21430
rect -1670 21410 -1650 21430
rect -1650 21410 -1645 21430
rect -1675 21405 -1645 21410
rect -1515 21430 -1485 21435
rect -1515 21410 -1510 21430
rect -1510 21410 -1490 21430
rect -1490 21410 -1485 21430
rect -1515 21405 -1485 21410
rect -1355 21430 -1325 21435
rect -1355 21410 -1350 21430
rect -1350 21410 -1330 21430
rect -1330 21410 -1325 21430
rect -1355 21405 -1325 21410
rect -1275 21430 -1245 21435
rect -1275 21410 -1270 21430
rect -1270 21410 -1250 21430
rect -1250 21410 -1245 21430
rect -1275 21405 -1245 21410
rect -1195 21430 -1165 21435
rect -1195 21410 -1190 21430
rect -1190 21410 -1170 21430
rect -1170 21410 -1165 21430
rect -1195 21405 -1165 21410
rect -1115 21430 -1085 21435
rect -1115 21410 -1110 21430
rect -1110 21410 -1090 21430
rect -1090 21410 -1085 21430
rect -1115 21405 -1085 21410
rect -1035 21430 -1005 21435
rect -1035 21410 -1030 21430
rect -1030 21410 -1010 21430
rect -1010 21410 -1005 21430
rect -1035 21405 -1005 21410
rect -875 21430 -845 21435
rect -875 21410 -870 21430
rect -870 21410 -850 21430
rect -850 21410 -845 21430
rect -875 21405 -845 21410
rect -715 21430 -685 21435
rect -715 21410 -710 21430
rect -710 21410 -690 21430
rect -690 21410 -685 21430
rect -715 21405 -685 21410
rect -555 21430 -525 21435
rect -555 21410 -550 21430
rect -550 21410 -530 21430
rect -530 21410 -525 21430
rect -555 21405 -525 21410
rect -14955 21270 -14925 21275
rect -14955 21250 -14950 21270
rect -14950 21250 -14930 21270
rect -14930 21250 -14925 21270
rect -14955 21245 -14925 21250
rect -14875 21270 -14845 21275
rect -14875 21250 -14870 21270
rect -14870 21250 -14850 21270
rect -14850 21250 -14845 21270
rect -14875 21245 -14845 21250
rect -14795 21270 -14765 21275
rect -14795 21250 -14790 21270
rect -14790 21250 -14770 21270
rect -14770 21250 -14765 21270
rect -14795 21245 -14765 21250
rect -14715 21270 -14685 21275
rect -14715 21250 -14710 21270
rect -14710 21250 -14690 21270
rect -14690 21250 -14685 21270
rect -14715 21245 -14685 21250
rect -14635 21270 -14605 21275
rect -14635 21250 -14630 21270
rect -14630 21250 -14610 21270
rect -14610 21250 -14605 21270
rect -14635 21245 -14605 21250
rect -14555 21270 -14525 21275
rect -14555 21250 -14550 21270
rect -14550 21250 -14530 21270
rect -14530 21250 -14525 21270
rect -14555 21245 -14525 21250
rect -14475 21270 -14445 21275
rect -14475 21250 -14470 21270
rect -14470 21250 -14450 21270
rect -14450 21250 -14445 21270
rect -14475 21245 -14445 21250
rect -14395 21270 -14365 21275
rect -14395 21250 -14390 21270
rect -14390 21250 -14370 21270
rect -14370 21250 -14365 21270
rect -14395 21245 -14365 21250
rect -14315 21270 -14285 21275
rect -14315 21250 -14310 21270
rect -14310 21250 -14290 21270
rect -14290 21250 -14285 21270
rect -14315 21245 -14285 21250
rect -14235 21270 -14205 21275
rect -14235 21250 -14230 21270
rect -14230 21250 -14210 21270
rect -14210 21250 -14205 21270
rect -14235 21245 -14205 21250
rect -14155 21270 -14125 21275
rect -14155 21250 -14150 21270
rect -14150 21250 -14130 21270
rect -14130 21250 -14125 21270
rect -14155 21245 -14125 21250
rect -14075 21270 -14045 21275
rect -14075 21250 -14070 21270
rect -14070 21250 -14050 21270
rect -14050 21250 -14045 21270
rect -14075 21245 -14045 21250
rect -13995 21270 -13965 21275
rect -13995 21250 -13990 21270
rect -13990 21250 -13970 21270
rect -13970 21250 -13965 21270
rect -13995 21245 -13965 21250
rect -13915 21270 -13885 21275
rect -13915 21250 -13910 21270
rect -13910 21250 -13890 21270
rect -13890 21250 -13885 21270
rect -13915 21245 -13885 21250
rect -13835 21270 -13805 21275
rect -13835 21250 -13830 21270
rect -13830 21250 -13810 21270
rect -13810 21250 -13805 21270
rect -13835 21245 -13805 21250
rect -13755 21270 -13725 21275
rect -13755 21250 -13750 21270
rect -13750 21250 -13730 21270
rect -13730 21250 -13725 21270
rect -13755 21245 -13725 21250
rect -13675 21270 -13645 21275
rect -13675 21250 -13670 21270
rect -13670 21250 -13650 21270
rect -13650 21250 -13645 21270
rect -13675 21245 -13645 21250
rect -13595 21270 -13565 21275
rect -13595 21250 -13590 21270
rect -13590 21250 -13570 21270
rect -13570 21250 -13565 21270
rect -13595 21245 -13565 21250
rect -13515 21270 -13485 21275
rect -13515 21250 -13510 21270
rect -13510 21250 -13490 21270
rect -13490 21250 -13485 21270
rect -13515 21245 -13485 21250
rect -13435 21270 -13405 21275
rect -13435 21250 -13430 21270
rect -13430 21250 -13410 21270
rect -13410 21250 -13405 21270
rect -13435 21245 -13405 21250
rect -13355 21270 -13325 21275
rect -13355 21250 -13350 21270
rect -13350 21250 -13330 21270
rect -13330 21250 -13325 21270
rect -13355 21245 -13325 21250
rect -13275 21270 -13245 21275
rect -13275 21250 -13270 21270
rect -13270 21250 -13250 21270
rect -13250 21250 -13245 21270
rect -13275 21245 -13245 21250
rect -13195 21270 -13165 21275
rect -13195 21250 -13190 21270
rect -13190 21250 -13170 21270
rect -13170 21250 -13165 21270
rect -13195 21245 -13165 21250
rect -13115 21270 -13085 21275
rect -13115 21250 -13110 21270
rect -13110 21250 -13090 21270
rect -13090 21250 -13085 21270
rect -13115 21245 -13085 21250
rect -13035 21270 -13005 21275
rect -13035 21250 -13030 21270
rect -13030 21250 -13010 21270
rect -13010 21250 -13005 21270
rect -13035 21245 -13005 21250
rect -12955 21270 -12925 21275
rect -12955 21250 -12950 21270
rect -12950 21250 -12930 21270
rect -12930 21250 -12925 21270
rect -12955 21245 -12925 21250
rect -12875 21270 -12845 21275
rect -12875 21250 -12870 21270
rect -12870 21250 -12850 21270
rect -12850 21250 -12845 21270
rect -12875 21245 -12845 21250
rect -12795 21270 -12765 21275
rect -12795 21250 -12790 21270
rect -12790 21250 -12770 21270
rect -12770 21250 -12765 21270
rect -12795 21245 -12765 21250
rect -12715 21270 -12685 21275
rect -12715 21250 -12710 21270
rect -12710 21250 -12690 21270
rect -12690 21250 -12685 21270
rect -12715 21245 -12685 21250
rect -12635 21270 -12605 21275
rect -12635 21250 -12630 21270
rect -12630 21250 -12610 21270
rect -12610 21250 -12605 21270
rect -12635 21245 -12605 21250
rect -12555 21270 -12525 21275
rect -12555 21250 -12550 21270
rect -12550 21250 -12530 21270
rect -12530 21250 -12525 21270
rect -12555 21245 -12525 21250
rect -12475 21270 -12445 21275
rect -12475 21250 -12470 21270
rect -12470 21250 -12450 21270
rect -12450 21250 -12445 21270
rect -12475 21245 -12445 21250
rect -12395 21270 -12365 21275
rect -12395 21250 -12390 21270
rect -12390 21250 -12370 21270
rect -12370 21250 -12365 21270
rect -12395 21245 -12365 21250
rect -12315 21270 -12285 21275
rect -12315 21250 -12310 21270
rect -12310 21250 -12290 21270
rect -12290 21250 -12285 21270
rect -12315 21245 -12285 21250
rect -12235 21270 -12205 21275
rect -12235 21250 -12230 21270
rect -12230 21250 -12210 21270
rect -12210 21250 -12205 21270
rect -12235 21245 -12205 21250
rect -12155 21270 -12125 21275
rect -12155 21250 -12150 21270
rect -12150 21250 -12130 21270
rect -12130 21250 -12125 21270
rect -12155 21245 -12125 21250
rect -12075 21270 -12045 21275
rect -12075 21250 -12070 21270
rect -12070 21250 -12050 21270
rect -12050 21250 -12045 21270
rect -12075 21245 -12045 21250
rect -11995 21270 -11965 21275
rect -11995 21250 -11990 21270
rect -11990 21250 -11970 21270
rect -11970 21250 -11965 21270
rect -11995 21245 -11965 21250
rect -11915 21270 -11885 21275
rect -11915 21250 -11910 21270
rect -11910 21250 -11890 21270
rect -11890 21250 -11885 21270
rect -11915 21245 -11885 21250
rect -11835 21270 -11805 21275
rect -11835 21250 -11830 21270
rect -11830 21250 -11810 21270
rect -11810 21250 -11805 21270
rect -11835 21245 -11805 21250
rect -11755 21270 -11725 21275
rect -11755 21250 -11750 21270
rect -11750 21250 -11730 21270
rect -11730 21250 -11725 21270
rect -11755 21245 -11725 21250
rect -11675 21270 -11645 21275
rect -11675 21250 -11670 21270
rect -11670 21250 -11650 21270
rect -11650 21250 -11645 21270
rect -11675 21245 -11645 21250
rect -11595 21270 -11565 21275
rect -11595 21250 -11590 21270
rect -11590 21250 -11570 21270
rect -11570 21250 -11565 21270
rect -11595 21245 -11565 21250
rect -11515 21270 -11485 21275
rect -11515 21250 -11510 21270
rect -11510 21250 -11490 21270
rect -11490 21250 -11485 21270
rect -11515 21245 -11485 21250
rect -11435 21270 -11405 21275
rect -11435 21250 -11430 21270
rect -11430 21250 -11410 21270
rect -11410 21250 -11405 21270
rect -11435 21245 -11405 21250
rect -11355 21270 -11325 21275
rect -11355 21250 -11350 21270
rect -11350 21250 -11330 21270
rect -11330 21250 -11325 21270
rect -11355 21245 -11325 21250
rect -11275 21270 -11245 21275
rect -11275 21250 -11270 21270
rect -11270 21250 -11250 21270
rect -11250 21250 -11245 21270
rect -11275 21245 -11245 21250
rect -11195 21270 -11165 21275
rect -11195 21250 -11190 21270
rect -11190 21250 -11170 21270
rect -11170 21250 -11165 21270
rect -11195 21245 -11165 21250
rect -11115 21270 -11085 21275
rect -11115 21250 -11110 21270
rect -11110 21250 -11090 21270
rect -11090 21250 -11085 21270
rect -11115 21245 -11085 21250
rect -11035 21270 -11005 21275
rect -11035 21250 -11030 21270
rect -11030 21250 -11010 21270
rect -11010 21250 -11005 21270
rect -11035 21245 -11005 21250
rect -10955 21270 -10925 21275
rect -10955 21250 -10950 21270
rect -10950 21250 -10930 21270
rect -10930 21250 -10925 21270
rect -10955 21245 -10925 21250
rect -10875 21270 -10845 21275
rect -10875 21250 -10870 21270
rect -10870 21250 -10850 21270
rect -10850 21250 -10845 21270
rect -10875 21245 -10845 21250
rect -10795 21270 -10765 21275
rect -10795 21250 -10790 21270
rect -10790 21250 -10770 21270
rect -10770 21250 -10765 21270
rect -10795 21245 -10765 21250
rect -10715 21270 -10685 21275
rect -10715 21250 -10710 21270
rect -10710 21250 -10690 21270
rect -10690 21250 -10685 21270
rect -10715 21245 -10685 21250
rect -10635 21270 -10605 21275
rect -10635 21250 -10630 21270
rect -10630 21250 -10610 21270
rect -10610 21250 -10605 21270
rect -10635 21245 -10605 21250
rect -10555 21270 -10525 21275
rect -10555 21250 -10550 21270
rect -10550 21250 -10530 21270
rect -10530 21250 -10525 21270
rect -10555 21245 -10525 21250
rect -10475 21270 -10445 21275
rect -10475 21250 -10470 21270
rect -10470 21250 -10450 21270
rect -10450 21250 -10445 21270
rect -10475 21245 -10445 21250
rect -10395 21270 -10365 21275
rect -10395 21250 -10390 21270
rect -10390 21250 -10370 21270
rect -10370 21250 -10365 21270
rect -10395 21245 -10365 21250
rect -10315 21270 -10285 21275
rect -10315 21250 -10310 21270
rect -10310 21250 -10290 21270
rect -10290 21250 -10285 21270
rect -10315 21245 -10285 21250
rect -10235 21270 -10205 21275
rect -10235 21250 -10230 21270
rect -10230 21250 -10210 21270
rect -10210 21250 -10205 21270
rect -10235 21245 -10205 21250
rect -10155 21270 -10125 21275
rect -10155 21250 -10150 21270
rect -10150 21250 -10130 21270
rect -10130 21250 -10125 21270
rect -10155 21245 -10125 21250
rect -10075 21270 -10045 21275
rect -10075 21250 -10070 21270
rect -10070 21250 -10050 21270
rect -10050 21250 -10045 21270
rect -10075 21245 -10045 21250
rect -9995 21270 -9965 21275
rect -9995 21250 -9990 21270
rect -9990 21250 -9970 21270
rect -9970 21250 -9965 21270
rect -9995 21245 -9965 21250
rect -9915 21270 -9885 21275
rect -9915 21250 -9910 21270
rect -9910 21250 -9890 21270
rect -9890 21250 -9885 21270
rect -9915 21245 -9885 21250
rect -9835 21270 -9805 21275
rect -9835 21250 -9830 21270
rect -9830 21250 -9810 21270
rect -9810 21250 -9805 21270
rect -9835 21245 -9805 21250
rect -9755 21270 -9725 21275
rect -9755 21250 -9750 21270
rect -9750 21250 -9730 21270
rect -9730 21250 -9725 21270
rect -9755 21245 -9725 21250
rect -9675 21270 -9645 21275
rect -9675 21250 -9670 21270
rect -9670 21250 -9650 21270
rect -9650 21250 -9645 21270
rect -9675 21245 -9645 21250
rect -9595 21270 -9565 21275
rect -9595 21250 -9590 21270
rect -9590 21250 -9570 21270
rect -9570 21250 -9565 21270
rect -9595 21245 -9565 21250
rect -9515 21270 -9485 21275
rect -9515 21250 -9510 21270
rect -9510 21250 -9490 21270
rect -9490 21250 -9485 21270
rect -9515 21245 -9485 21250
rect -9435 21270 -9405 21275
rect -9435 21250 -9430 21270
rect -9430 21250 -9410 21270
rect -9410 21250 -9405 21270
rect -9435 21245 -9405 21250
rect -9355 21270 -9325 21275
rect -9355 21250 -9350 21270
rect -9350 21250 -9330 21270
rect -9330 21250 -9325 21270
rect -9355 21245 -9325 21250
rect -9275 21270 -9245 21275
rect -9275 21250 -9270 21270
rect -9270 21250 -9250 21270
rect -9250 21250 -9245 21270
rect -9275 21245 -9245 21250
rect -9195 21270 -9165 21275
rect -9195 21250 -9190 21270
rect -9190 21250 -9170 21270
rect -9170 21250 -9165 21270
rect -9195 21245 -9165 21250
rect -9115 21270 -9085 21275
rect -9115 21250 -9110 21270
rect -9110 21250 -9090 21270
rect -9090 21250 -9085 21270
rect -9115 21245 -9085 21250
rect -9035 21270 -9005 21275
rect -9035 21250 -9030 21270
rect -9030 21250 -9010 21270
rect -9010 21250 -9005 21270
rect -9035 21245 -9005 21250
rect -8955 21270 -8925 21275
rect -8955 21250 -8950 21270
rect -8950 21250 -8930 21270
rect -8930 21250 -8925 21270
rect -8955 21245 -8925 21250
rect -8875 21270 -8845 21275
rect -8875 21250 -8870 21270
rect -8870 21250 -8850 21270
rect -8850 21250 -8845 21270
rect -8875 21245 -8845 21250
rect -8795 21270 -8765 21275
rect -8795 21250 -8790 21270
rect -8790 21250 -8770 21270
rect -8770 21250 -8765 21270
rect -8795 21245 -8765 21250
rect -8715 21270 -8685 21275
rect -8715 21250 -8710 21270
rect -8710 21250 -8690 21270
rect -8690 21250 -8685 21270
rect -8715 21245 -8685 21250
rect -8635 21270 -8605 21275
rect -8635 21250 -8630 21270
rect -8630 21250 -8610 21270
rect -8610 21250 -8605 21270
rect -8635 21245 -8605 21250
rect -8555 21270 -8525 21275
rect -8555 21250 -8550 21270
rect -8550 21250 -8530 21270
rect -8530 21250 -8525 21270
rect -8555 21245 -8525 21250
rect -8475 21270 -8445 21275
rect -8475 21250 -8470 21270
rect -8470 21250 -8450 21270
rect -8450 21250 -8445 21270
rect -8475 21245 -8445 21250
rect -8395 21270 -8365 21275
rect -8395 21250 -8390 21270
rect -8390 21250 -8370 21270
rect -8370 21250 -8365 21270
rect -8395 21245 -8365 21250
rect -8315 21270 -8285 21275
rect -8315 21250 -8310 21270
rect -8310 21250 -8290 21270
rect -8290 21250 -8285 21270
rect -8315 21245 -8285 21250
rect -8235 21270 -8205 21275
rect -8235 21250 -8230 21270
rect -8230 21250 -8210 21270
rect -8210 21250 -8205 21270
rect -8235 21245 -8205 21250
rect -8155 21270 -8125 21275
rect -8155 21250 -8150 21270
rect -8150 21250 -8130 21270
rect -8130 21250 -8125 21270
rect -8155 21245 -8125 21250
rect -8075 21270 -8045 21275
rect -8075 21250 -8070 21270
rect -8070 21250 -8050 21270
rect -8050 21250 -8045 21270
rect -8075 21245 -8045 21250
rect -7995 21270 -7965 21275
rect -7995 21250 -7990 21270
rect -7990 21250 -7970 21270
rect -7970 21250 -7965 21270
rect -7995 21245 -7965 21250
rect -7915 21270 -7885 21275
rect -7915 21250 -7910 21270
rect -7910 21250 -7890 21270
rect -7890 21250 -7885 21270
rect -7915 21245 -7885 21250
rect -7835 21270 -7805 21275
rect -7835 21250 -7830 21270
rect -7830 21250 -7810 21270
rect -7810 21250 -7805 21270
rect -7835 21245 -7805 21250
rect -7755 21270 -7725 21275
rect -7755 21250 -7750 21270
rect -7750 21250 -7730 21270
rect -7730 21250 -7725 21270
rect -7755 21245 -7725 21250
rect -7675 21270 -7645 21275
rect -7675 21250 -7670 21270
rect -7670 21250 -7650 21270
rect -7650 21250 -7645 21270
rect -7675 21245 -7645 21250
rect -7595 21270 -7565 21275
rect -7595 21250 -7590 21270
rect -7590 21250 -7570 21270
rect -7570 21250 -7565 21270
rect -7595 21245 -7565 21250
rect -7515 21270 -7485 21275
rect -7515 21250 -7510 21270
rect -7510 21250 -7490 21270
rect -7490 21250 -7485 21270
rect -7515 21245 -7485 21250
rect -7435 21270 -7405 21275
rect -7435 21250 -7430 21270
rect -7430 21250 -7410 21270
rect -7410 21250 -7405 21270
rect -7435 21245 -7405 21250
rect -7355 21270 -7325 21275
rect -7355 21250 -7350 21270
rect -7350 21250 -7330 21270
rect -7330 21250 -7325 21270
rect -7355 21245 -7325 21250
rect -7275 21270 -7245 21275
rect -7275 21250 -7270 21270
rect -7270 21250 -7250 21270
rect -7250 21250 -7245 21270
rect -7275 21245 -7245 21250
rect -7195 21270 -7165 21275
rect -7195 21250 -7190 21270
rect -7190 21250 -7170 21270
rect -7170 21250 -7165 21270
rect -7195 21245 -7165 21250
rect -7115 21270 -7085 21275
rect -7115 21250 -7110 21270
rect -7110 21250 -7090 21270
rect -7090 21250 -7085 21270
rect -7115 21245 -7085 21250
rect -7035 21270 -7005 21275
rect -7035 21250 -7030 21270
rect -7030 21250 -7010 21270
rect -7010 21250 -7005 21270
rect -7035 21245 -7005 21250
rect -6955 21270 -6925 21275
rect -6955 21250 -6950 21270
rect -6950 21250 -6930 21270
rect -6930 21250 -6925 21270
rect -6955 21245 -6925 21250
rect -6875 21270 -6845 21275
rect -6875 21250 -6870 21270
rect -6870 21250 -6850 21270
rect -6850 21250 -6845 21270
rect -6875 21245 -6845 21250
rect -6795 21270 -6765 21275
rect -6795 21250 -6790 21270
rect -6790 21250 -6770 21270
rect -6770 21250 -6765 21270
rect -6795 21245 -6765 21250
rect -6715 21270 -6685 21275
rect -6715 21250 -6710 21270
rect -6710 21250 -6690 21270
rect -6690 21250 -6685 21270
rect -6715 21245 -6685 21250
rect -6635 21270 -6605 21275
rect -6635 21250 -6630 21270
rect -6630 21250 -6610 21270
rect -6610 21250 -6605 21270
rect -6635 21245 -6605 21250
rect -6555 21270 -6525 21275
rect -6555 21250 -6550 21270
rect -6550 21250 -6530 21270
rect -6530 21250 -6525 21270
rect -6555 21245 -6525 21250
rect -6475 21270 -6445 21275
rect -6475 21250 -6470 21270
rect -6470 21250 -6450 21270
rect -6450 21250 -6445 21270
rect -6475 21245 -6445 21250
rect -6395 21270 -6365 21275
rect -6395 21250 -6390 21270
rect -6390 21250 -6370 21270
rect -6370 21250 -6365 21270
rect -6395 21245 -6365 21250
rect -6315 21270 -6285 21275
rect -6315 21250 -6310 21270
rect -6310 21250 -6290 21270
rect -6290 21250 -6285 21270
rect -6315 21245 -6285 21250
rect -6235 21270 -6205 21275
rect -6235 21250 -6230 21270
rect -6230 21250 -6210 21270
rect -6210 21250 -6205 21270
rect -6235 21245 -6205 21250
rect -6155 21270 -6125 21275
rect -6155 21250 -6150 21270
rect -6150 21250 -6130 21270
rect -6130 21250 -6125 21270
rect -6155 21245 -6125 21250
rect -5675 21270 -5645 21275
rect -5675 21250 -5670 21270
rect -5670 21250 -5650 21270
rect -5650 21250 -5645 21270
rect -5675 21245 -5645 21250
rect -5595 21270 -5565 21275
rect -5595 21250 -5590 21270
rect -5590 21250 -5570 21270
rect -5570 21250 -5565 21270
rect -5595 21245 -5565 21250
rect -5515 21270 -5485 21275
rect -5515 21250 -5510 21270
rect -5510 21250 -5490 21270
rect -5490 21250 -5485 21270
rect -5515 21245 -5485 21250
rect -5435 21270 -5405 21275
rect -5435 21250 -5430 21270
rect -5430 21250 -5410 21270
rect -5410 21250 -5405 21270
rect -5435 21245 -5405 21250
rect -5355 21270 -5325 21275
rect -5355 21250 -5350 21270
rect -5350 21250 -5330 21270
rect -5330 21250 -5325 21270
rect -5355 21245 -5325 21250
rect -5275 21270 -5245 21275
rect -5275 21250 -5270 21270
rect -5270 21250 -5250 21270
rect -5250 21250 -5245 21270
rect -5275 21245 -5245 21250
rect -5195 21270 -5165 21275
rect -5195 21250 -5190 21270
rect -5190 21250 -5170 21270
rect -5170 21250 -5165 21270
rect -5195 21245 -5165 21250
rect -5115 21270 -5085 21275
rect -5115 21250 -5110 21270
rect -5110 21250 -5090 21270
rect -5090 21250 -5085 21270
rect -5115 21245 -5085 21250
rect -5035 21270 -5005 21275
rect -5035 21250 -5030 21270
rect -5030 21250 -5010 21270
rect -5010 21250 -5005 21270
rect -5035 21245 -5005 21250
rect -4955 21270 -4925 21275
rect -4955 21250 -4950 21270
rect -4950 21250 -4930 21270
rect -4930 21250 -4925 21270
rect -4955 21245 -4925 21250
rect -4875 21270 -4845 21275
rect -4875 21250 -4870 21270
rect -4870 21250 -4850 21270
rect -4850 21250 -4845 21270
rect -4875 21245 -4845 21250
rect -4795 21270 -4765 21275
rect -4795 21250 -4790 21270
rect -4790 21250 -4770 21270
rect -4770 21250 -4765 21270
rect -4795 21245 -4765 21250
rect -4715 21270 -4685 21275
rect -4715 21250 -4710 21270
rect -4710 21250 -4690 21270
rect -4690 21250 -4685 21270
rect -4715 21245 -4685 21250
rect -4635 21270 -4605 21275
rect -4635 21250 -4630 21270
rect -4630 21250 -4610 21270
rect -4610 21250 -4605 21270
rect -4635 21245 -4605 21250
rect -4555 21270 -4525 21275
rect -4555 21250 -4550 21270
rect -4550 21250 -4530 21270
rect -4530 21250 -4525 21270
rect -4555 21245 -4525 21250
rect -4475 21270 -4445 21275
rect -4475 21250 -4470 21270
rect -4470 21250 -4450 21270
rect -4450 21250 -4445 21270
rect -4475 21245 -4445 21250
rect -4395 21270 -4365 21275
rect -4395 21250 -4390 21270
rect -4390 21250 -4370 21270
rect -4370 21250 -4365 21270
rect -4395 21245 -4365 21250
rect -4315 21270 -4285 21275
rect -4315 21250 -4310 21270
rect -4310 21250 -4290 21270
rect -4290 21250 -4285 21270
rect -4315 21245 -4285 21250
rect -4235 21270 -4205 21275
rect -4235 21250 -4230 21270
rect -4230 21250 -4210 21270
rect -4210 21250 -4205 21270
rect -4235 21245 -4205 21250
rect -4155 21270 -4125 21275
rect -4155 21250 -4150 21270
rect -4150 21250 -4130 21270
rect -4130 21250 -4125 21270
rect -4155 21245 -4125 21250
rect -4075 21270 -4045 21275
rect -4075 21250 -4070 21270
rect -4070 21250 -4050 21270
rect -4050 21250 -4045 21270
rect -4075 21245 -4045 21250
rect -3995 21270 -3965 21275
rect -3995 21250 -3990 21270
rect -3990 21250 -3970 21270
rect -3970 21250 -3965 21270
rect -3995 21245 -3965 21250
rect -3915 21270 -3885 21275
rect -3915 21250 -3910 21270
rect -3910 21250 -3890 21270
rect -3890 21250 -3885 21270
rect -3915 21245 -3885 21250
rect -3835 21270 -3805 21275
rect -3835 21250 -3830 21270
rect -3830 21250 -3810 21270
rect -3810 21250 -3805 21270
rect -3835 21245 -3805 21250
rect -3755 21270 -3725 21275
rect -3755 21250 -3750 21270
rect -3750 21250 -3730 21270
rect -3730 21250 -3725 21270
rect -3755 21245 -3725 21250
rect -3675 21270 -3645 21275
rect -3675 21250 -3670 21270
rect -3670 21250 -3650 21270
rect -3650 21250 -3645 21270
rect -3675 21245 -3645 21250
rect -3595 21270 -3565 21275
rect -3595 21250 -3590 21270
rect -3590 21250 -3570 21270
rect -3570 21250 -3565 21270
rect -3595 21245 -3565 21250
rect -3515 21270 -3485 21275
rect -3515 21250 -3510 21270
rect -3510 21250 -3490 21270
rect -3490 21250 -3485 21270
rect -3515 21245 -3485 21250
rect -3435 21270 -3405 21275
rect -3435 21250 -3430 21270
rect -3430 21250 -3410 21270
rect -3410 21250 -3405 21270
rect -3435 21245 -3405 21250
rect -3355 21270 -3325 21275
rect -3355 21250 -3350 21270
rect -3350 21250 -3330 21270
rect -3330 21250 -3325 21270
rect -3355 21245 -3325 21250
rect -3275 21270 -3245 21275
rect -3275 21250 -3270 21270
rect -3270 21250 -3250 21270
rect -3250 21250 -3245 21270
rect -3275 21245 -3245 21250
rect -3195 21270 -3165 21275
rect -3195 21250 -3190 21270
rect -3190 21250 -3170 21270
rect -3170 21250 -3165 21270
rect -3195 21245 -3165 21250
rect -3115 21270 -3085 21275
rect -3115 21250 -3110 21270
rect -3110 21250 -3090 21270
rect -3090 21250 -3085 21270
rect -3115 21245 -3085 21250
rect -3035 21270 -3005 21275
rect -3035 21250 -3030 21270
rect -3030 21250 -3010 21270
rect -3010 21250 -3005 21270
rect -3035 21245 -3005 21250
rect -2955 21270 -2925 21275
rect -2955 21250 -2950 21270
rect -2950 21250 -2930 21270
rect -2930 21250 -2925 21270
rect -2955 21245 -2925 21250
rect -2875 21270 -2845 21275
rect -2875 21250 -2870 21270
rect -2870 21250 -2850 21270
rect -2850 21250 -2845 21270
rect -2875 21245 -2845 21250
rect -2795 21270 -2765 21275
rect -2795 21250 -2790 21270
rect -2790 21250 -2770 21270
rect -2770 21250 -2765 21270
rect -2795 21245 -2765 21250
rect -2715 21270 -2685 21275
rect -2715 21250 -2710 21270
rect -2710 21250 -2690 21270
rect -2690 21250 -2685 21270
rect -2715 21245 -2685 21250
rect -2635 21270 -2605 21275
rect -2635 21250 -2630 21270
rect -2630 21250 -2610 21270
rect -2610 21250 -2605 21270
rect -2635 21245 -2605 21250
rect -2555 21270 -2525 21275
rect -2555 21250 -2550 21270
rect -2550 21250 -2530 21270
rect -2530 21250 -2525 21270
rect -2555 21245 -2525 21250
rect -2475 21270 -2445 21275
rect -2475 21250 -2470 21270
rect -2470 21250 -2450 21270
rect -2450 21250 -2445 21270
rect -2475 21245 -2445 21250
rect -2395 21270 -2365 21275
rect -2395 21250 -2390 21270
rect -2390 21250 -2370 21270
rect -2370 21250 -2365 21270
rect -2395 21245 -2365 21250
rect -2315 21270 -2285 21275
rect -2315 21250 -2310 21270
rect -2310 21250 -2290 21270
rect -2290 21250 -2285 21270
rect -2315 21245 -2285 21250
rect -2235 21270 -2205 21275
rect -2235 21250 -2230 21270
rect -2230 21250 -2210 21270
rect -2210 21250 -2205 21270
rect -2235 21245 -2205 21250
rect -2155 21270 -2125 21275
rect -2155 21250 -2150 21270
rect -2150 21250 -2130 21270
rect -2130 21250 -2125 21270
rect -2155 21245 -2125 21250
rect -2075 21270 -2045 21275
rect -2075 21250 -2070 21270
rect -2070 21250 -2050 21270
rect -2050 21250 -2045 21270
rect -2075 21245 -2045 21250
rect -1995 21270 -1965 21275
rect -1995 21250 -1990 21270
rect -1990 21250 -1970 21270
rect -1970 21250 -1965 21270
rect -1995 21245 -1965 21250
rect -1835 21270 -1805 21275
rect -1835 21250 -1830 21270
rect -1830 21250 -1810 21270
rect -1810 21250 -1805 21270
rect -1835 21245 -1805 21250
rect -1755 21270 -1725 21275
rect -1755 21250 -1750 21270
rect -1750 21250 -1730 21270
rect -1730 21250 -1725 21270
rect -1755 21245 -1725 21250
rect -1675 21270 -1645 21275
rect -1675 21250 -1670 21270
rect -1670 21250 -1650 21270
rect -1650 21250 -1645 21270
rect -1675 21245 -1645 21250
rect -1515 21270 -1485 21275
rect -1515 21250 -1510 21270
rect -1510 21250 -1490 21270
rect -1490 21250 -1485 21270
rect -1515 21245 -1485 21250
rect -1355 21270 -1325 21275
rect -1355 21250 -1350 21270
rect -1350 21250 -1330 21270
rect -1330 21250 -1325 21270
rect -1355 21245 -1325 21250
rect -1275 21270 -1245 21275
rect -1275 21250 -1270 21270
rect -1270 21250 -1250 21270
rect -1250 21250 -1245 21270
rect -1275 21245 -1245 21250
rect -1195 21270 -1165 21275
rect -1195 21250 -1190 21270
rect -1190 21250 -1170 21270
rect -1170 21250 -1165 21270
rect -1195 21245 -1165 21250
rect -1115 21270 -1085 21275
rect -1115 21250 -1110 21270
rect -1110 21250 -1090 21270
rect -1090 21250 -1085 21270
rect -1115 21245 -1085 21250
rect -1035 21270 -1005 21275
rect -1035 21250 -1030 21270
rect -1030 21250 -1010 21270
rect -1010 21250 -1005 21270
rect -1035 21245 -1005 21250
rect -875 21270 -845 21275
rect -875 21250 -870 21270
rect -870 21250 -850 21270
rect -850 21250 -845 21270
rect -875 21245 -845 21250
rect -715 21270 -685 21275
rect -715 21250 -710 21270
rect -710 21250 -690 21270
rect -690 21250 -685 21270
rect -715 21245 -685 21250
rect -555 21270 -525 21275
rect -555 21250 -550 21270
rect -550 21250 -530 21270
rect -530 21250 -525 21270
rect -555 21245 -525 21250
rect -14955 21110 -14925 21115
rect -14955 21090 -14950 21110
rect -14950 21090 -14930 21110
rect -14930 21090 -14925 21110
rect -14955 21085 -14925 21090
rect -14875 21110 -14845 21115
rect -14875 21090 -14870 21110
rect -14870 21090 -14850 21110
rect -14850 21090 -14845 21110
rect -14875 21085 -14845 21090
rect -14795 21110 -14765 21115
rect -14795 21090 -14790 21110
rect -14790 21090 -14770 21110
rect -14770 21090 -14765 21110
rect -14795 21085 -14765 21090
rect -14715 21110 -14685 21115
rect -14715 21090 -14710 21110
rect -14710 21090 -14690 21110
rect -14690 21090 -14685 21110
rect -14715 21085 -14685 21090
rect -14635 21110 -14605 21115
rect -14635 21090 -14630 21110
rect -14630 21090 -14610 21110
rect -14610 21090 -14605 21110
rect -14635 21085 -14605 21090
rect -14555 21110 -14525 21115
rect -14555 21090 -14550 21110
rect -14550 21090 -14530 21110
rect -14530 21090 -14525 21110
rect -14555 21085 -14525 21090
rect -14475 21110 -14445 21115
rect -14475 21090 -14470 21110
rect -14470 21090 -14450 21110
rect -14450 21090 -14445 21110
rect -14475 21085 -14445 21090
rect -14395 21110 -14365 21115
rect -14395 21090 -14390 21110
rect -14390 21090 -14370 21110
rect -14370 21090 -14365 21110
rect -14395 21085 -14365 21090
rect -14315 21110 -14285 21115
rect -14315 21090 -14310 21110
rect -14310 21090 -14290 21110
rect -14290 21090 -14285 21110
rect -14315 21085 -14285 21090
rect -14235 21110 -14205 21115
rect -14235 21090 -14230 21110
rect -14230 21090 -14210 21110
rect -14210 21090 -14205 21110
rect -14235 21085 -14205 21090
rect -14155 21110 -14125 21115
rect -14155 21090 -14150 21110
rect -14150 21090 -14130 21110
rect -14130 21090 -14125 21110
rect -14155 21085 -14125 21090
rect -14075 21110 -14045 21115
rect -14075 21090 -14070 21110
rect -14070 21090 -14050 21110
rect -14050 21090 -14045 21110
rect -14075 21085 -14045 21090
rect -13995 21110 -13965 21115
rect -13995 21090 -13990 21110
rect -13990 21090 -13970 21110
rect -13970 21090 -13965 21110
rect -13995 21085 -13965 21090
rect -13915 21110 -13885 21115
rect -13915 21090 -13910 21110
rect -13910 21090 -13890 21110
rect -13890 21090 -13885 21110
rect -13915 21085 -13885 21090
rect -13835 21110 -13805 21115
rect -13835 21090 -13830 21110
rect -13830 21090 -13810 21110
rect -13810 21090 -13805 21110
rect -13835 21085 -13805 21090
rect -13755 21110 -13725 21115
rect -13755 21090 -13750 21110
rect -13750 21090 -13730 21110
rect -13730 21090 -13725 21110
rect -13755 21085 -13725 21090
rect -13675 21110 -13645 21115
rect -13675 21090 -13670 21110
rect -13670 21090 -13650 21110
rect -13650 21090 -13645 21110
rect -13675 21085 -13645 21090
rect -13595 21110 -13565 21115
rect -13595 21090 -13590 21110
rect -13590 21090 -13570 21110
rect -13570 21090 -13565 21110
rect -13595 21085 -13565 21090
rect -13515 21110 -13485 21115
rect -13515 21090 -13510 21110
rect -13510 21090 -13490 21110
rect -13490 21090 -13485 21110
rect -13515 21085 -13485 21090
rect -13435 21110 -13405 21115
rect -13435 21090 -13430 21110
rect -13430 21090 -13410 21110
rect -13410 21090 -13405 21110
rect -13435 21085 -13405 21090
rect -13355 21110 -13325 21115
rect -13355 21090 -13350 21110
rect -13350 21090 -13330 21110
rect -13330 21090 -13325 21110
rect -13355 21085 -13325 21090
rect -13275 21110 -13245 21115
rect -13275 21090 -13270 21110
rect -13270 21090 -13250 21110
rect -13250 21090 -13245 21110
rect -13275 21085 -13245 21090
rect -13195 21110 -13165 21115
rect -13195 21090 -13190 21110
rect -13190 21090 -13170 21110
rect -13170 21090 -13165 21110
rect -13195 21085 -13165 21090
rect -13115 21110 -13085 21115
rect -13115 21090 -13110 21110
rect -13110 21090 -13090 21110
rect -13090 21090 -13085 21110
rect -13115 21085 -13085 21090
rect -13035 21110 -13005 21115
rect -13035 21090 -13030 21110
rect -13030 21090 -13010 21110
rect -13010 21090 -13005 21110
rect -13035 21085 -13005 21090
rect -12955 21110 -12925 21115
rect -12955 21090 -12950 21110
rect -12950 21090 -12930 21110
rect -12930 21090 -12925 21110
rect -12955 21085 -12925 21090
rect -12875 21110 -12845 21115
rect -12875 21090 -12870 21110
rect -12870 21090 -12850 21110
rect -12850 21090 -12845 21110
rect -12875 21085 -12845 21090
rect -12795 21110 -12765 21115
rect -12795 21090 -12790 21110
rect -12790 21090 -12770 21110
rect -12770 21090 -12765 21110
rect -12795 21085 -12765 21090
rect -12715 21110 -12685 21115
rect -12715 21090 -12710 21110
rect -12710 21090 -12690 21110
rect -12690 21090 -12685 21110
rect -12715 21085 -12685 21090
rect -12635 21110 -12605 21115
rect -12635 21090 -12630 21110
rect -12630 21090 -12610 21110
rect -12610 21090 -12605 21110
rect -12635 21085 -12605 21090
rect -12555 21110 -12525 21115
rect -12555 21090 -12550 21110
rect -12550 21090 -12530 21110
rect -12530 21090 -12525 21110
rect -12555 21085 -12525 21090
rect -12475 21110 -12445 21115
rect -12475 21090 -12470 21110
rect -12470 21090 -12450 21110
rect -12450 21090 -12445 21110
rect -12475 21085 -12445 21090
rect -12395 21110 -12365 21115
rect -12395 21090 -12390 21110
rect -12390 21090 -12370 21110
rect -12370 21090 -12365 21110
rect -12395 21085 -12365 21090
rect -12315 21110 -12285 21115
rect -12315 21090 -12310 21110
rect -12310 21090 -12290 21110
rect -12290 21090 -12285 21110
rect -12315 21085 -12285 21090
rect -12235 21110 -12205 21115
rect -12235 21090 -12230 21110
rect -12230 21090 -12210 21110
rect -12210 21090 -12205 21110
rect -12235 21085 -12205 21090
rect -12155 21110 -12125 21115
rect -12155 21090 -12150 21110
rect -12150 21090 -12130 21110
rect -12130 21090 -12125 21110
rect -12155 21085 -12125 21090
rect -12075 21110 -12045 21115
rect -12075 21090 -12070 21110
rect -12070 21090 -12050 21110
rect -12050 21090 -12045 21110
rect -12075 21085 -12045 21090
rect -11995 21110 -11965 21115
rect -11995 21090 -11990 21110
rect -11990 21090 -11970 21110
rect -11970 21090 -11965 21110
rect -11995 21085 -11965 21090
rect -11915 21110 -11885 21115
rect -11915 21090 -11910 21110
rect -11910 21090 -11890 21110
rect -11890 21090 -11885 21110
rect -11915 21085 -11885 21090
rect -11835 21110 -11805 21115
rect -11835 21090 -11830 21110
rect -11830 21090 -11810 21110
rect -11810 21090 -11805 21110
rect -11835 21085 -11805 21090
rect -11755 21110 -11725 21115
rect -11755 21090 -11750 21110
rect -11750 21090 -11730 21110
rect -11730 21090 -11725 21110
rect -11755 21085 -11725 21090
rect -11675 21110 -11645 21115
rect -11675 21090 -11670 21110
rect -11670 21090 -11650 21110
rect -11650 21090 -11645 21110
rect -11675 21085 -11645 21090
rect -11595 21110 -11565 21115
rect -11595 21090 -11590 21110
rect -11590 21090 -11570 21110
rect -11570 21090 -11565 21110
rect -11595 21085 -11565 21090
rect -11515 21110 -11485 21115
rect -11515 21090 -11510 21110
rect -11510 21090 -11490 21110
rect -11490 21090 -11485 21110
rect -11515 21085 -11485 21090
rect -11435 21110 -11405 21115
rect -11435 21090 -11430 21110
rect -11430 21090 -11410 21110
rect -11410 21090 -11405 21110
rect -11435 21085 -11405 21090
rect -11355 21110 -11325 21115
rect -11355 21090 -11350 21110
rect -11350 21090 -11330 21110
rect -11330 21090 -11325 21110
rect -11355 21085 -11325 21090
rect -11275 21110 -11245 21115
rect -11275 21090 -11270 21110
rect -11270 21090 -11250 21110
rect -11250 21090 -11245 21110
rect -11275 21085 -11245 21090
rect -11195 21110 -11165 21115
rect -11195 21090 -11190 21110
rect -11190 21090 -11170 21110
rect -11170 21090 -11165 21110
rect -11195 21085 -11165 21090
rect -11115 21110 -11085 21115
rect -11115 21090 -11110 21110
rect -11110 21090 -11090 21110
rect -11090 21090 -11085 21110
rect -11115 21085 -11085 21090
rect -11035 21110 -11005 21115
rect -11035 21090 -11030 21110
rect -11030 21090 -11010 21110
rect -11010 21090 -11005 21110
rect -11035 21085 -11005 21090
rect -10955 21110 -10925 21115
rect -10955 21090 -10950 21110
rect -10950 21090 -10930 21110
rect -10930 21090 -10925 21110
rect -10955 21085 -10925 21090
rect -10875 21110 -10845 21115
rect -10875 21090 -10870 21110
rect -10870 21090 -10850 21110
rect -10850 21090 -10845 21110
rect -10875 21085 -10845 21090
rect -10795 21110 -10765 21115
rect -10795 21090 -10790 21110
rect -10790 21090 -10770 21110
rect -10770 21090 -10765 21110
rect -10795 21085 -10765 21090
rect -10715 21110 -10685 21115
rect -10715 21090 -10710 21110
rect -10710 21090 -10690 21110
rect -10690 21090 -10685 21110
rect -10715 21085 -10685 21090
rect -10635 21110 -10605 21115
rect -10635 21090 -10630 21110
rect -10630 21090 -10610 21110
rect -10610 21090 -10605 21110
rect -10635 21085 -10605 21090
rect -10555 21110 -10525 21115
rect -10555 21090 -10550 21110
rect -10550 21090 -10530 21110
rect -10530 21090 -10525 21110
rect -10555 21085 -10525 21090
rect -10475 21110 -10445 21115
rect -10475 21090 -10470 21110
rect -10470 21090 -10450 21110
rect -10450 21090 -10445 21110
rect -10475 21085 -10445 21090
rect -10395 21110 -10365 21115
rect -10395 21090 -10390 21110
rect -10390 21090 -10370 21110
rect -10370 21090 -10365 21110
rect -10395 21085 -10365 21090
rect -10315 21110 -10285 21115
rect -10315 21090 -10310 21110
rect -10310 21090 -10290 21110
rect -10290 21090 -10285 21110
rect -10315 21085 -10285 21090
rect -10235 21110 -10205 21115
rect -10235 21090 -10230 21110
rect -10230 21090 -10210 21110
rect -10210 21090 -10205 21110
rect -10235 21085 -10205 21090
rect -10155 21110 -10125 21115
rect -10155 21090 -10150 21110
rect -10150 21090 -10130 21110
rect -10130 21090 -10125 21110
rect -10155 21085 -10125 21090
rect -10075 21110 -10045 21115
rect -10075 21090 -10070 21110
rect -10070 21090 -10050 21110
rect -10050 21090 -10045 21110
rect -10075 21085 -10045 21090
rect -9995 21110 -9965 21115
rect -9995 21090 -9990 21110
rect -9990 21090 -9970 21110
rect -9970 21090 -9965 21110
rect -9995 21085 -9965 21090
rect -9915 21110 -9885 21115
rect -9915 21090 -9910 21110
rect -9910 21090 -9890 21110
rect -9890 21090 -9885 21110
rect -9915 21085 -9885 21090
rect -9835 21110 -9805 21115
rect -9835 21090 -9830 21110
rect -9830 21090 -9810 21110
rect -9810 21090 -9805 21110
rect -9835 21085 -9805 21090
rect -9755 21110 -9725 21115
rect -9755 21090 -9750 21110
rect -9750 21090 -9730 21110
rect -9730 21090 -9725 21110
rect -9755 21085 -9725 21090
rect -9675 21110 -9645 21115
rect -9675 21090 -9670 21110
rect -9670 21090 -9650 21110
rect -9650 21090 -9645 21110
rect -9675 21085 -9645 21090
rect -9595 21110 -9565 21115
rect -9595 21090 -9590 21110
rect -9590 21090 -9570 21110
rect -9570 21090 -9565 21110
rect -9595 21085 -9565 21090
rect -9515 21110 -9485 21115
rect -9515 21090 -9510 21110
rect -9510 21090 -9490 21110
rect -9490 21090 -9485 21110
rect -9515 21085 -9485 21090
rect -9435 21110 -9405 21115
rect -9435 21090 -9430 21110
rect -9430 21090 -9410 21110
rect -9410 21090 -9405 21110
rect -9435 21085 -9405 21090
rect -9355 21110 -9325 21115
rect -9355 21090 -9350 21110
rect -9350 21090 -9330 21110
rect -9330 21090 -9325 21110
rect -9355 21085 -9325 21090
rect -9275 21110 -9245 21115
rect -9275 21090 -9270 21110
rect -9270 21090 -9250 21110
rect -9250 21090 -9245 21110
rect -9275 21085 -9245 21090
rect -9195 21110 -9165 21115
rect -9195 21090 -9190 21110
rect -9190 21090 -9170 21110
rect -9170 21090 -9165 21110
rect -9195 21085 -9165 21090
rect -9115 21110 -9085 21115
rect -9115 21090 -9110 21110
rect -9110 21090 -9090 21110
rect -9090 21090 -9085 21110
rect -9115 21085 -9085 21090
rect -9035 21110 -9005 21115
rect -9035 21090 -9030 21110
rect -9030 21090 -9010 21110
rect -9010 21090 -9005 21110
rect -9035 21085 -9005 21090
rect -8955 21110 -8925 21115
rect -8955 21090 -8950 21110
rect -8950 21090 -8930 21110
rect -8930 21090 -8925 21110
rect -8955 21085 -8925 21090
rect -8875 21110 -8845 21115
rect -8875 21090 -8870 21110
rect -8870 21090 -8850 21110
rect -8850 21090 -8845 21110
rect -8875 21085 -8845 21090
rect -8795 21110 -8765 21115
rect -8795 21090 -8790 21110
rect -8790 21090 -8770 21110
rect -8770 21090 -8765 21110
rect -8795 21085 -8765 21090
rect -8715 21110 -8685 21115
rect -8715 21090 -8710 21110
rect -8710 21090 -8690 21110
rect -8690 21090 -8685 21110
rect -8715 21085 -8685 21090
rect -8635 21110 -8605 21115
rect -8635 21090 -8630 21110
rect -8630 21090 -8610 21110
rect -8610 21090 -8605 21110
rect -8635 21085 -8605 21090
rect -8555 21110 -8525 21115
rect -8555 21090 -8550 21110
rect -8550 21090 -8530 21110
rect -8530 21090 -8525 21110
rect -8555 21085 -8525 21090
rect -8475 21110 -8445 21115
rect -8475 21090 -8470 21110
rect -8470 21090 -8450 21110
rect -8450 21090 -8445 21110
rect -8475 21085 -8445 21090
rect -8395 21110 -8365 21115
rect -8395 21090 -8390 21110
rect -8390 21090 -8370 21110
rect -8370 21090 -8365 21110
rect -8395 21085 -8365 21090
rect -8315 21110 -8285 21115
rect -8315 21090 -8310 21110
rect -8310 21090 -8290 21110
rect -8290 21090 -8285 21110
rect -8315 21085 -8285 21090
rect -8235 21110 -8205 21115
rect -8235 21090 -8230 21110
rect -8230 21090 -8210 21110
rect -8210 21090 -8205 21110
rect -8235 21085 -8205 21090
rect -8155 21110 -8125 21115
rect -8155 21090 -8150 21110
rect -8150 21090 -8130 21110
rect -8130 21090 -8125 21110
rect -8155 21085 -8125 21090
rect -8075 21110 -8045 21115
rect -8075 21090 -8070 21110
rect -8070 21090 -8050 21110
rect -8050 21090 -8045 21110
rect -8075 21085 -8045 21090
rect -7995 21110 -7965 21115
rect -7995 21090 -7990 21110
rect -7990 21090 -7970 21110
rect -7970 21090 -7965 21110
rect -7995 21085 -7965 21090
rect -7915 21110 -7885 21115
rect -7915 21090 -7910 21110
rect -7910 21090 -7890 21110
rect -7890 21090 -7885 21110
rect -7915 21085 -7885 21090
rect -7835 21110 -7805 21115
rect -7835 21090 -7830 21110
rect -7830 21090 -7810 21110
rect -7810 21090 -7805 21110
rect -7835 21085 -7805 21090
rect -7755 21110 -7725 21115
rect -7755 21090 -7750 21110
rect -7750 21090 -7730 21110
rect -7730 21090 -7725 21110
rect -7755 21085 -7725 21090
rect -7675 21110 -7645 21115
rect -7675 21090 -7670 21110
rect -7670 21090 -7650 21110
rect -7650 21090 -7645 21110
rect -7675 21085 -7645 21090
rect -7595 21110 -7565 21115
rect -7595 21090 -7590 21110
rect -7590 21090 -7570 21110
rect -7570 21090 -7565 21110
rect -7595 21085 -7565 21090
rect -7515 21110 -7485 21115
rect -7515 21090 -7510 21110
rect -7510 21090 -7490 21110
rect -7490 21090 -7485 21110
rect -7515 21085 -7485 21090
rect -7435 21110 -7405 21115
rect -7435 21090 -7430 21110
rect -7430 21090 -7410 21110
rect -7410 21090 -7405 21110
rect -7435 21085 -7405 21090
rect -7355 21110 -7325 21115
rect -7355 21090 -7350 21110
rect -7350 21090 -7330 21110
rect -7330 21090 -7325 21110
rect -7355 21085 -7325 21090
rect -7275 21110 -7245 21115
rect -7275 21090 -7270 21110
rect -7270 21090 -7250 21110
rect -7250 21090 -7245 21110
rect -7275 21085 -7245 21090
rect -7195 21110 -7165 21115
rect -7195 21090 -7190 21110
rect -7190 21090 -7170 21110
rect -7170 21090 -7165 21110
rect -7195 21085 -7165 21090
rect -7115 21110 -7085 21115
rect -7115 21090 -7110 21110
rect -7110 21090 -7090 21110
rect -7090 21090 -7085 21110
rect -7115 21085 -7085 21090
rect -7035 21110 -7005 21115
rect -7035 21090 -7030 21110
rect -7030 21090 -7010 21110
rect -7010 21090 -7005 21110
rect -7035 21085 -7005 21090
rect -6955 21110 -6925 21115
rect -6955 21090 -6950 21110
rect -6950 21090 -6930 21110
rect -6930 21090 -6925 21110
rect -6955 21085 -6925 21090
rect -6875 21110 -6845 21115
rect -6875 21090 -6870 21110
rect -6870 21090 -6850 21110
rect -6850 21090 -6845 21110
rect -6875 21085 -6845 21090
rect -6795 21110 -6765 21115
rect -6795 21090 -6790 21110
rect -6790 21090 -6770 21110
rect -6770 21090 -6765 21110
rect -6795 21085 -6765 21090
rect -6715 21110 -6685 21115
rect -6715 21090 -6710 21110
rect -6710 21090 -6690 21110
rect -6690 21090 -6685 21110
rect -6715 21085 -6685 21090
rect -6635 21110 -6605 21115
rect -6635 21090 -6630 21110
rect -6630 21090 -6610 21110
rect -6610 21090 -6605 21110
rect -6635 21085 -6605 21090
rect -6555 21110 -6525 21115
rect -6555 21090 -6550 21110
rect -6550 21090 -6530 21110
rect -6530 21090 -6525 21110
rect -6555 21085 -6525 21090
rect -6475 21110 -6445 21115
rect -6475 21090 -6470 21110
rect -6470 21090 -6450 21110
rect -6450 21090 -6445 21110
rect -6475 21085 -6445 21090
rect -6395 21110 -6365 21115
rect -6395 21090 -6390 21110
rect -6390 21090 -6370 21110
rect -6370 21090 -6365 21110
rect -6395 21085 -6365 21090
rect -6315 21110 -6285 21115
rect -6315 21090 -6310 21110
rect -6310 21090 -6290 21110
rect -6290 21090 -6285 21110
rect -6315 21085 -6285 21090
rect -6235 21110 -6205 21115
rect -6235 21090 -6230 21110
rect -6230 21090 -6210 21110
rect -6210 21090 -6205 21110
rect -6235 21085 -6205 21090
rect -6155 21110 -6125 21115
rect -6155 21090 -6150 21110
rect -6150 21090 -6130 21110
rect -6130 21090 -6125 21110
rect -6155 21085 -6125 21090
rect -5675 21110 -5645 21115
rect -5675 21090 -5670 21110
rect -5670 21090 -5650 21110
rect -5650 21090 -5645 21110
rect -5675 21085 -5645 21090
rect -5595 21110 -5565 21115
rect -5595 21090 -5590 21110
rect -5590 21090 -5570 21110
rect -5570 21090 -5565 21110
rect -5595 21085 -5565 21090
rect -5515 21110 -5485 21115
rect -5515 21090 -5510 21110
rect -5510 21090 -5490 21110
rect -5490 21090 -5485 21110
rect -5515 21085 -5485 21090
rect -5435 21110 -5405 21115
rect -5435 21090 -5430 21110
rect -5430 21090 -5410 21110
rect -5410 21090 -5405 21110
rect -5435 21085 -5405 21090
rect -5355 21110 -5325 21115
rect -5355 21090 -5350 21110
rect -5350 21090 -5330 21110
rect -5330 21090 -5325 21110
rect -5355 21085 -5325 21090
rect -5275 21110 -5245 21115
rect -5275 21090 -5270 21110
rect -5270 21090 -5250 21110
rect -5250 21090 -5245 21110
rect -5275 21085 -5245 21090
rect -5195 21110 -5165 21115
rect -5195 21090 -5190 21110
rect -5190 21090 -5170 21110
rect -5170 21090 -5165 21110
rect -5195 21085 -5165 21090
rect -5115 21110 -5085 21115
rect -5115 21090 -5110 21110
rect -5110 21090 -5090 21110
rect -5090 21090 -5085 21110
rect -5115 21085 -5085 21090
rect -5035 21110 -5005 21115
rect -5035 21090 -5030 21110
rect -5030 21090 -5010 21110
rect -5010 21090 -5005 21110
rect -5035 21085 -5005 21090
rect -4955 21110 -4925 21115
rect -4955 21090 -4950 21110
rect -4950 21090 -4930 21110
rect -4930 21090 -4925 21110
rect -4955 21085 -4925 21090
rect -4875 21110 -4845 21115
rect -4875 21090 -4870 21110
rect -4870 21090 -4850 21110
rect -4850 21090 -4845 21110
rect -4875 21085 -4845 21090
rect -4795 21110 -4765 21115
rect -4795 21090 -4790 21110
rect -4790 21090 -4770 21110
rect -4770 21090 -4765 21110
rect -4795 21085 -4765 21090
rect -4715 21110 -4685 21115
rect -4715 21090 -4710 21110
rect -4710 21090 -4690 21110
rect -4690 21090 -4685 21110
rect -4715 21085 -4685 21090
rect -4635 21110 -4605 21115
rect -4635 21090 -4630 21110
rect -4630 21090 -4610 21110
rect -4610 21090 -4605 21110
rect -4635 21085 -4605 21090
rect -4555 21110 -4525 21115
rect -4555 21090 -4550 21110
rect -4550 21090 -4530 21110
rect -4530 21090 -4525 21110
rect -4555 21085 -4525 21090
rect -4475 21110 -4445 21115
rect -4475 21090 -4470 21110
rect -4470 21090 -4450 21110
rect -4450 21090 -4445 21110
rect -4475 21085 -4445 21090
rect -4395 21110 -4365 21115
rect -4395 21090 -4390 21110
rect -4390 21090 -4370 21110
rect -4370 21090 -4365 21110
rect -4395 21085 -4365 21090
rect -4315 21110 -4285 21115
rect -4315 21090 -4310 21110
rect -4310 21090 -4290 21110
rect -4290 21090 -4285 21110
rect -4315 21085 -4285 21090
rect -4235 21110 -4205 21115
rect -4235 21090 -4230 21110
rect -4230 21090 -4210 21110
rect -4210 21090 -4205 21110
rect -4235 21085 -4205 21090
rect -4155 21110 -4125 21115
rect -4155 21090 -4150 21110
rect -4150 21090 -4130 21110
rect -4130 21090 -4125 21110
rect -4155 21085 -4125 21090
rect -4075 21110 -4045 21115
rect -4075 21090 -4070 21110
rect -4070 21090 -4050 21110
rect -4050 21090 -4045 21110
rect -4075 21085 -4045 21090
rect -3995 21110 -3965 21115
rect -3995 21090 -3990 21110
rect -3990 21090 -3970 21110
rect -3970 21090 -3965 21110
rect -3995 21085 -3965 21090
rect -3915 21110 -3885 21115
rect -3915 21090 -3910 21110
rect -3910 21090 -3890 21110
rect -3890 21090 -3885 21110
rect -3915 21085 -3885 21090
rect -3835 21110 -3805 21115
rect -3835 21090 -3830 21110
rect -3830 21090 -3810 21110
rect -3810 21090 -3805 21110
rect -3835 21085 -3805 21090
rect -3755 21110 -3725 21115
rect -3755 21090 -3750 21110
rect -3750 21090 -3730 21110
rect -3730 21090 -3725 21110
rect -3755 21085 -3725 21090
rect -3675 21110 -3645 21115
rect -3675 21090 -3670 21110
rect -3670 21090 -3650 21110
rect -3650 21090 -3645 21110
rect -3675 21085 -3645 21090
rect -3595 21110 -3565 21115
rect -3595 21090 -3590 21110
rect -3590 21090 -3570 21110
rect -3570 21090 -3565 21110
rect -3595 21085 -3565 21090
rect -3515 21110 -3485 21115
rect -3515 21090 -3510 21110
rect -3510 21090 -3490 21110
rect -3490 21090 -3485 21110
rect -3515 21085 -3485 21090
rect -3435 21110 -3405 21115
rect -3435 21090 -3430 21110
rect -3430 21090 -3410 21110
rect -3410 21090 -3405 21110
rect -3435 21085 -3405 21090
rect -3355 21110 -3325 21115
rect -3355 21090 -3350 21110
rect -3350 21090 -3330 21110
rect -3330 21090 -3325 21110
rect -3355 21085 -3325 21090
rect -3275 21110 -3245 21115
rect -3275 21090 -3270 21110
rect -3270 21090 -3250 21110
rect -3250 21090 -3245 21110
rect -3275 21085 -3245 21090
rect -3195 21110 -3165 21115
rect -3195 21090 -3190 21110
rect -3190 21090 -3170 21110
rect -3170 21090 -3165 21110
rect -3195 21085 -3165 21090
rect -3115 21110 -3085 21115
rect -3115 21090 -3110 21110
rect -3110 21090 -3090 21110
rect -3090 21090 -3085 21110
rect -3115 21085 -3085 21090
rect -3035 21110 -3005 21115
rect -3035 21090 -3030 21110
rect -3030 21090 -3010 21110
rect -3010 21090 -3005 21110
rect -3035 21085 -3005 21090
rect -2955 21110 -2925 21115
rect -2955 21090 -2950 21110
rect -2950 21090 -2930 21110
rect -2930 21090 -2925 21110
rect -2955 21085 -2925 21090
rect -2875 21110 -2845 21115
rect -2875 21090 -2870 21110
rect -2870 21090 -2850 21110
rect -2850 21090 -2845 21110
rect -2875 21085 -2845 21090
rect -2795 21110 -2765 21115
rect -2795 21090 -2790 21110
rect -2790 21090 -2770 21110
rect -2770 21090 -2765 21110
rect -2795 21085 -2765 21090
rect -2715 21110 -2685 21115
rect -2715 21090 -2710 21110
rect -2710 21090 -2690 21110
rect -2690 21090 -2685 21110
rect -2715 21085 -2685 21090
rect -2635 21110 -2605 21115
rect -2635 21090 -2630 21110
rect -2630 21090 -2610 21110
rect -2610 21090 -2605 21110
rect -2635 21085 -2605 21090
rect -2555 21110 -2525 21115
rect -2555 21090 -2550 21110
rect -2550 21090 -2530 21110
rect -2530 21090 -2525 21110
rect -2555 21085 -2525 21090
rect -2475 21110 -2445 21115
rect -2475 21090 -2470 21110
rect -2470 21090 -2450 21110
rect -2450 21090 -2445 21110
rect -2475 21085 -2445 21090
rect -2395 21110 -2365 21115
rect -2395 21090 -2390 21110
rect -2390 21090 -2370 21110
rect -2370 21090 -2365 21110
rect -2395 21085 -2365 21090
rect -2315 21110 -2285 21115
rect -2315 21090 -2310 21110
rect -2310 21090 -2290 21110
rect -2290 21090 -2285 21110
rect -2315 21085 -2285 21090
rect -2235 21110 -2205 21115
rect -2235 21090 -2230 21110
rect -2230 21090 -2210 21110
rect -2210 21090 -2205 21110
rect -2235 21085 -2205 21090
rect -2155 21110 -2125 21115
rect -2155 21090 -2150 21110
rect -2150 21090 -2130 21110
rect -2130 21090 -2125 21110
rect -2155 21085 -2125 21090
rect -2075 21110 -2045 21115
rect -2075 21090 -2070 21110
rect -2070 21090 -2050 21110
rect -2050 21090 -2045 21110
rect -2075 21085 -2045 21090
rect -1995 21110 -1965 21115
rect -1995 21090 -1990 21110
rect -1990 21090 -1970 21110
rect -1970 21090 -1965 21110
rect -1995 21085 -1965 21090
rect -1835 21110 -1805 21115
rect -1835 21090 -1830 21110
rect -1830 21090 -1810 21110
rect -1810 21090 -1805 21110
rect -1835 21085 -1805 21090
rect -1755 21110 -1725 21115
rect -1755 21090 -1750 21110
rect -1750 21090 -1730 21110
rect -1730 21090 -1725 21110
rect -1755 21085 -1725 21090
rect -1675 21110 -1645 21115
rect -1675 21090 -1670 21110
rect -1670 21090 -1650 21110
rect -1650 21090 -1645 21110
rect -1675 21085 -1645 21090
rect -1515 21110 -1485 21115
rect -1515 21090 -1510 21110
rect -1510 21090 -1490 21110
rect -1490 21090 -1485 21110
rect -1515 21085 -1485 21090
rect -1355 21110 -1325 21115
rect -1355 21090 -1350 21110
rect -1350 21090 -1330 21110
rect -1330 21090 -1325 21110
rect -1355 21085 -1325 21090
rect -1275 21110 -1245 21115
rect -1275 21090 -1270 21110
rect -1270 21090 -1250 21110
rect -1250 21090 -1245 21110
rect -1275 21085 -1245 21090
rect -1195 21110 -1165 21115
rect -1195 21090 -1190 21110
rect -1190 21090 -1170 21110
rect -1170 21090 -1165 21110
rect -1195 21085 -1165 21090
rect -1115 21110 -1085 21115
rect -1115 21090 -1110 21110
rect -1110 21090 -1090 21110
rect -1090 21090 -1085 21110
rect -1115 21085 -1085 21090
rect -1035 21110 -1005 21115
rect -1035 21090 -1030 21110
rect -1030 21090 -1010 21110
rect -1010 21090 -1005 21110
rect -1035 21085 -1005 21090
rect -875 21110 -845 21115
rect -875 21090 -870 21110
rect -870 21090 -850 21110
rect -850 21090 -845 21110
rect -875 21085 -845 21090
rect -715 21110 -685 21115
rect -715 21090 -710 21110
rect -710 21090 -690 21110
rect -690 21090 -685 21110
rect -715 21085 -685 21090
rect -555 21110 -525 21115
rect -555 21090 -550 21110
rect -550 21090 -530 21110
rect -530 21090 -525 21110
rect -555 21085 -525 21090
rect -14955 20950 -14925 20955
rect -14955 20930 -14950 20950
rect -14950 20930 -14930 20950
rect -14930 20930 -14925 20950
rect -14955 20925 -14925 20930
rect -14875 20950 -14845 20955
rect -14875 20930 -14870 20950
rect -14870 20930 -14850 20950
rect -14850 20930 -14845 20950
rect -14875 20925 -14845 20930
rect -14795 20950 -14765 20955
rect -14795 20930 -14790 20950
rect -14790 20930 -14770 20950
rect -14770 20930 -14765 20950
rect -14795 20925 -14765 20930
rect -14715 20950 -14685 20955
rect -14715 20930 -14710 20950
rect -14710 20930 -14690 20950
rect -14690 20930 -14685 20950
rect -14715 20925 -14685 20930
rect -14635 20950 -14605 20955
rect -14635 20930 -14630 20950
rect -14630 20930 -14610 20950
rect -14610 20930 -14605 20950
rect -14635 20925 -14605 20930
rect -14555 20950 -14525 20955
rect -14555 20930 -14550 20950
rect -14550 20930 -14530 20950
rect -14530 20930 -14525 20950
rect -14555 20925 -14525 20930
rect -14475 20950 -14445 20955
rect -14475 20930 -14470 20950
rect -14470 20930 -14450 20950
rect -14450 20930 -14445 20950
rect -14475 20925 -14445 20930
rect -14395 20950 -14365 20955
rect -14395 20930 -14390 20950
rect -14390 20930 -14370 20950
rect -14370 20930 -14365 20950
rect -14395 20925 -14365 20930
rect -14315 20950 -14285 20955
rect -14315 20930 -14310 20950
rect -14310 20930 -14290 20950
rect -14290 20930 -14285 20950
rect -14315 20925 -14285 20930
rect -14235 20950 -14205 20955
rect -14235 20930 -14230 20950
rect -14230 20930 -14210 20950
rect -14210 20930 -14205 20950
rect -14235 20925 -14205 20930
rect -14155 20950 -14125 20955
rect -14155 20930 -14150 20950
rect -14150 20930 -14130 20950
rect -14130 20930 -14125 20950
rect -14155 20925 -14125 20930
rect -14075 20950 -14045 20955
rect -14075 20930 -14070 20950
rect -14070 20930 -14050 20950
rect -14050 20930 -14045 20950
rect -14075 20925 -14045 20930
rect -13995 20950 -13965 20955
rect -13995 20930 -13990 20950
rect -13990 20930 -13970 20950
rect -13970 20930 -13965 20950
rect -13995 20925 -13965 20930
rect -13915 20950 -13885 20955
rect -13915 20930 -13910 20950
rect -13910 20930 -13890 20950
rect -13890 20930 -13885 20950
rect -13915 20925 -13885 20930
rect -13835 20950 -13805 20955
rect -13835 20930 -13830 20950
rect -13830 20930 -13810 20950
rect -13810 20930 -13805 20950
rect -13835 20925 -13805 20930
rect -13755 20950 -13725 20955
rect -13755 20930 -13750 20950
rect -13750 20930 -13730 20950
rect -13730 20930 -13725 20950
rect -13755 20925 -13725 20930
rect -13675 20950 -13645 20955
rect -13675 20930 -13670 20950
rect -13670 20930 -13650 20950
rect -13650 20930 -13645 20950
rect -13675 20925 -13645 20930
rect -13595 20950 -13565 20955
rect -13595 20930 -13590 20950
rect -13590 20930 -13570 20950
rect -13570 20930 -13565 20950
rect -13595 20925 -13565 20930
rect -13515 20950 -13485 20955
rect -13515 20930 -13510 20950
rect -13510 20930 -13490 20950
rect -13490 20930 -13485 20950
rect -13515 20925 -13485 20930
rect -13435 20950 -13405 20955
rect -13435 20930 -13430 20950
rect -13430 20930 -13410 20950
rect -13410 20930 -13405 20950
rect -13435 20925 -13405 20930
rect -13355 20950 -13325 20955
rect -13355 20930 -13350 20950
rect -13350 20930 -13330 20950
rect -13330 20930 -13325 20950
rect -13355 20925 -13325 20930
rect -13275 20950 -13245 20955
rect -13275 20930 -13270 20950
rect -13270 20930 -13250 20950
rect -13250 20930 -13245 20950
rect -13275 20925 -13245 20930
rect -13195 20950 -13165 20955
rect -13195 20930 -13190 20950
rect -13190 20930 -13170 20950
rect -13170 20930 -13165 20950
rect -13195 20925 -13165 20930
rect -13115 20950 -13085 20955
rect -13115 20930 -13110 20950
rect -13110 20930 -13090 20950
rect -13090 20930 -13085 20950
rect -13115 20925 -13085 20930
rect -13035 20950 -13005 20955
rect -13035 20930 -13030 20950
rect -13030 20930 -13010 20950
rect -13010 20930 -13005 20950
rect -13035 20925 -13005 20930
rect -12955 20950 -12925 20955
rect -12955 20930 -12950 20950
rect -12950 20930 -12930 20950
rect -12930 20930 -12925 20950
rect -12955 20925 -12925 20930
rect -12875 20950 -12845 20955
rect -12875 20930 -12870 20950
rect -12870 20930 -12850 20950
rect -12850 20930 -12845 20950
rect -12875 20925 -12845 20930
rect -12795 20950 -12765 20955
rect -12795 20930 -12790 20950
rect -12790 20930 -12770 20950
rect -12770 20930 -12765 20950
rect -12795 20925 -12765 20930
rect -12715 20950 -12685 20955
rect -12715 20930 -12710 20950
rect -12710 20930 -12690 20950
rect -12690 20930 -12685 20950
rect -12715 20925 -12685 20930
rect -12635 20950 -12605 20955
rect -12635 20930 -12630 20950
rect -12630 20930 -12610 20950
rect -12610 20930 -12605 20950
rect -12635 20925 -12605 20930
rect -12555 20950 -12525 20955
rect -12555 20930 -12550 20950
rect -12550 20930 -12530 20950
rect -12530 20930 -12525 20950
rect -12555 20925 -12525 20930
rect -12475 20950 -12445 20955
rect -12475 20930 -12470 20950
rect -12470 20930 -12450 20950
rect -12450 20930 -12445 20950
rect -12475 20925 -12445 20930
rect -12395 20950 -12365 20955
rect -12395 20930 -12390 20950
rect -12390 20930 -12370 20950
rect -12370 20930 -12365 20950
rect -12395 20925 -12365 20930
rect -12315 20950 -12285 20955
rect -12315 20930 -12310 20950
rect -12310 20930 -12290 20950
rect -12290 20930 -12285 20950
rect -12315 20925 -12285 20930
rect -12235 20950 -12205 20955
rect -12235 20930 -12230 20950
rect -12230 20930 -12210 20950
rect -12210 20930 -12205 20950
rect -12235 20925 -12205 20930
rect -12155 20950 -12125 20955
rect -12155 20930 -12150 20950
rect -12150 20930 -12130 20950
rect -12130 20930 -12125 20950
rect -12155 20925 -12125 20930
rect -12075 20950 -12045 20955
rect -12075 20930 -12070 20950
rect -12070 20930 -12050 20950
rect -12050 20930 -12045 20950
rect -12075 20925 -12045 20930
rect -11995 20950 -11965 20955
rect -11995 20930 -11990 20950
rect -11990 20930 -11970 20950
rect -11970 20930 -11965 20950
rect -11995 20925 -11965 20930
rect -11915 20950 -11885 20955
rect -11915 20930 -11910 20950
rect -11910 20930 -11890 20950
rect -11890 20930 -11885 20950
rect -11915 20925 -11885 20930
rect -11835 20950 -11805 20955
rect -11835 20930 -11830 20950
rect -11830 20930 -11810 20950
rect -11810 20930 -11805 20950
rect -11835 20925 -11805 20930
rect -11755 20950 -11725 20955
rect -11755 20930 -11750 20950
rect -11750 20930 -11730 20950
rect -11730 20930 -11725 20950
rect -11755 20925 -11725 20930
rect -11675 20950 -11645 20955
rect -11675 20930 -11670 20950
rect -11670 20930 -11650 20950
rect -11650 20930 -11645 20950
rect -11675 20925 -11645 20930
rect -11595 20950 -11565 20955
rect -11595 20930 -11590 20950
rect -11590 20930 -11570 20950
rect -11570 20930 -11565 20950
rect -11595 20925 -11565 20930
rect -11515 20950 -11485 20955
rect -11515 20930 -11510 20950
rect -11510 20930 -11490 20950
rect -11490 20930 -11485 20950
rect -11515 20925 -11485 20930
rect -11435 20950 -11405 20955
rect -11435 20930 -11430 20950
rect -11430 20930 -11410 20950
rect -11410 20930 -11405 20950
rect -11435 20925 -11405 20930
rect -11355 20950 -11325 20955
rect -11355 20930 -11350 20950
rect -11350 20930 -11330 20950
rect -11330 20930 -11325 20950
rect -11355 20925 -11325 20930
rect -11275 20950 -11245 20955
rect -11275 20930 -11270 20950
rect -11270 20930 -11250 20950
rect -11250 20930 -11245 20950
rect -11275 20925 -11245 20930
rect -11195 20950 -11165 20955
rect -11195 20930 -11190 20950
rect -11190 20930 -11170 20950
rect -11170 20930 -11165 20950
rect -11195 20925 -11165 20930
rect -11115 20950 -11085 20955
rect -11115 20930 -11110 20950
rect -11110 20930 -11090 20950
rect -11090 20930 -11085 20950
rect -11115 20925 -11085 20930
rect -11035 20950 -11005 20955
rect -11035 20930 -11030 20950
rect -11030 20930 -11010 20950
rect -11010 20930 -11005 20950
rect -11035 20925 -11005 20930
rect -10955 20950 -10925 20955
rect -10955 20930 -10950 20950
rect -10950 20930 -10930 20950
rect -10930 20930 -10925 20950
rect -10955 20925 -10925 20930
rect -10875 20950 -10845 20955
rect -10875 20930 -10870 20950
rect -10870 20930 -10850 20950
rect -10850 20930 -10845 20950
rect -10875 20925 -10845 20930
rect -10795 20950 -10765 20955
rect -10795 20930 -10790 20950
rect -10790 20930 -10770 20950
rect -10770 20930 -10765 20950
rect -10795 20925 -10765 20930
rect -10715 20950 -10685 20955
rect -10715 20930 -10710 20950
rect -10710 20930 -10690 20950
rect -10690 20930 -10685 20950
rect -10715 20925 -10685 20930
rect -10635 20950 -10605 20955
rect -10635 20930 -10630 20950
rect -10630 20930 -10610 20950
rect -10610 20930 -10605 20950
rect -10635 20925 -10605 20930
rect -10555 20950 -10525 20955
rect -10555 20930 -10550 20950
rect -10550 20930 -10530 20950
rect -10530 20930 -10525 20950
rect -10555 20925 -10525 20930
rect -10475 20950 -10445 20955
rect -10475 20930 -10470 20950
rect -10470 20930 -10450 20950
rect -10450 20930 -10445 20950
rect -10475 20925 -10445 20930
rect -10395 20950 -10365 20955
rect -10395 20930 -10390 20950
rect -10390 20930 -10370 20950
rect -10370 20930 -10365 20950
rect -10395 20925 -10365 20930
rect -10315 20950 -10285 20955
rect -10315 20930 -10310 20950
rect -10310 20930 -10290 20950
rect -10290 20930 -10285 20950
rect -10315 20925 -10285 20930
rect -10235 20950 -10205 20955
rect -10235 20930 -10230 20950
rect -10230 20930 -10210 20950
rect -10210 20930 -10205 20950
rect -10235 20925 -10205 20930
rect -10155 20950 -10125 20955
rect -10155 20930 -10150 20950
rect -10150 20930 -10130 20950
rect -10130 20930 -10125 20950
rect -10155 20925 -10125 20930
rect -10075 20950 -10045 20955
rect -10075 20930 -10070 20950
rect -10070 20930 -10050 20950
rect -10050 20930 -10045 20950
rect -10075 20925 -10045 20930
rect -9995 20950 -9965 20955
rect -9995 20930 -9990 20950
rect -9990 20930 -9970 20950
rect -9970 20930 -9965 20950
rect -9995 20925 -9965 20930
rect -9915 20950 -9885 20955
rect -9915 20930 -9910 20950
rect -9910 20930 -9890 20950
rect -9890 20930 -9885 20950
rect -9915 20925 -9885 20930
rect -9835 20950 -9805 20955
rect -9835 20930 -9830 20950
rect -9830 20930 -9810 20950
rect -9810 20930 -9805 20950
rect -9835 20925 -9805 20930
rect -9755 20950 -9725 20955
rect -9755 20930 -9750 20950
rect -9750 20930 -9730 20950
rect -9730 20930 -9725 20950
rect -9755 20925 -9725 20930
rect -9675 20950 -9645 20955
rect -9675 20930 -9670 20950
rect -9670 20930 -9650 20950
rect -9650 20930 -9645 20950
rect -9675 20925 -9645 20930
rect -9595 20950 -9565 20955
rect -9595 20930 -9590 20950
rect -9590 20930 -9570 20950
rect -9570 20930 -9565 20950
rect -9595 20925 -9565 20930
rect -9515 20950 -9485 20955
rect -9515 20930 -9510 20950
rect -9510 20930 -9490 20950
rect -9490 20930 -9485 20950
rect -9515 20925 -9485 20930
rect -9435 20950 -9405 20955
rect -9435 20930 -9430 20950
rect -9430 20930 -9410 20950
rect -9410 20930 -9405 20950
rect -9435 20925 -9405 20930
rect -9355 20950 -9325 20955
rect -9355 20930 -9350 20950
rect -9350 20930 -9330 20950
rect -9330 20930 -9325 20950
rect -9355 20925 -9325 20930
rect -9275 20950 -9245 20955
rect -9275 20930 -9270 20950
rect -9270 20930 -9250 20950
rect -9250 20930 -9245 20950
rect -9275 20925 -9245 20930
rect -9195 20950 -9165 20955
rect -9195 20930 -9190 20950
rect -9190 20930 -9170 20950
rect -9170 20930 -9165 20950
rect -9195 20925 -9165 20930
rect -9115 20950 -9085 20955
rect -9115 20930 -9110 20950
rect -9110 20930 -9090 20950
rect -9090 20930 -9085 20950
rect -9115 20925 -9085 20930
rect -9035 20950 -9005 20955
rect -9035 20930 -9030 20950
rect -9030 20930 -9010 20950
rect -9010 20930 -9005 20950
rect -9035 20925 -9005 20930
rect -8955 20950 -8925 20955
rect -8955 20930 -8950 20950
rect -8950 20930 -8930 20950
rect -8930 20930 -8925 20950
rect -8955 20925 -8925 20930
rect -8875 20950 -8845 20955
rect -8875 20930 -8870 20950
rect -8870 20930 -8850 20950
rect -8850 20930 -8845 20950
rect -8875 20925 -8845 20930
rect -8795 20950 -8765 20955
rect -8795 20930 -8790 20950
rect -8790 20930 -8770 20950
rect -8770 20930 -8765 20950
rect -8795 20925 -8765 20930
rect -8715 20950 -8685 20955
rect -8715 20930 -8710 20950
rect -8710 20930 -8690 20950
rect -8690 20930 -8685 20950
rect -8715 20925 -8685 20930
rect -8635 20950 -8605 20955
rect -8635 20930 -8630 20950
rect -8630 20930 -8610 20950
rect -8610 20930 -8605 20950
rect -8635 20925 -8605 20930
rect -8555 20950 -8525 20955
rect -8555 20930 -8550 20950
rect -8550 20930 -8530 20950
rect -8530 20930 -8525 20950
rect -8555 20925 -8525 20930
rect -8475 20950 -8445 20955
rect -8475 20930 -8470 20950
rect -8470 20930 -8450 20950
rect -8450 20930 -8445 20950
rect -8475 20925 -8445 20930
rect -8395 20950 -8365 20955
rect -8395 20930 -8390 20950
rect -8390 20930 -8370 20950
rect -8370 20930 -8365 20950
rect -8395 20925 -8365 20930
rect -8315 20950 -8285 20955
rect -8315 20930 -8310 20950
rect -8310 20930 -8290 20950
rect -8290 20930 -8285 20950
rect -8315 20925 -8285 20930
rect -8235 20950 -8205 20955
rect -8235 20930 -8230 20950
rect -8230 20930 -8210 20950
rect -8210 20930 -8205 20950
rect -8235 20925 -8205 20930
rect -8155 20950 -8125 20955
rect -8155 20930 -8150 20950
rect -8150 20930 -8130 20950
rect -8130 20930 -8125 20950
rect -8155 20925 -8125 20930
rect -8075 20950 -8045 20955
rect -8075 20930 -8070 20950
rect -8070 20930 -8050 20950
rect -8050 20930 -8045 20950
rect -8075 20925 -8045 20930
rect -7995 20950 -7965 20955
rect -7995 20930 -7990 20950
rect -7990 20930 -7970 20950
rect -7970 20930 -7965 20950
rect -7995 20925 -7965 20930
rect -7915 20950 -7885 20955
rect -7915 20930 -7910 20950
rect -7910 20930 -7890 20950
rect -7890 20930 -7885 20950
rect -7915 20925 -7885 20930
rect -7835 20950 -7805 20955
rect -7835 20930 -7830 20950
rect -7830 20930 -7810 20950
rect -7810 20930 -7805 20950
rect -7835 20925 -7805 20930
rect -7755 20950 -7725 20955
rect -7755 20930 -7750 20950
rect -7750 20930 -7730 20950
rect -7730 20930 -7725 20950
rect -7755 20925 -7725 20930
rect -7675 20950 -7645 20955
rect -7675 20930 -7670 20950
rect -7670 20930 -7650 20950
rect -7650 20930 -7645 20950
rect -7675 20925 -7645 20930
rect -7595 20950 -7565 20955
rect -7595 20930 -7590 20950
rect -7590 20930 -7570 20950
rect -7570 20930 -7565 20950
rect -7595 20925 -7565 20930
rect -7515 20950 -7485 20955
rect -7515 20930 -7510 20950
rect -7510 20930 -7490 20950
rect -7490 20930 -7485 20950
rect -7515 20925 -7485 20930
rect -7435 20950 -7405 20955
rect -7435 20930 -7430 20950
rect -7430 20930 -7410 20950
rect -7410 20930 -7405 20950
rect -7435 20925 -7405 20930
rect -7355 20950 -7325 20955
rect -7355 20930 -7350 20950
rect -7350 20930 -7330 20950
rect -7330 20930 -7325 20950
rect -7355 20925 -7325 20930
rect -7275 20950 -7245 20955
rect -7275 20930 -7270 20950
rect -7270 20930 -7250 20950
rect -7250 20930 -7245 20950
rect -7275 20925 -7245 20930
rect -7195 20950 -7165 20955
rect -7195 20930 -7190 20950
rect -7190 20930 -7170 20950
rect -7170 20930 -7165 20950
rect -7195 20925 -7165 20930
rect -7115 20950 -7085 20955
rect -7115 20930 -7110 20950
rect -7110 20930 -7090 20950
rect -7090 20930 -7085 20950
rect -7115 20925 -7085 20930
rect -7035 20950 -7005 20955
rect -7035 20930 -7030 20950
rect -7030 20930 -7010 20950
rect -7010 20930 -7005 20950
rect -7035 20925 -7005 20930
rect -6955 20950 -6925 20955
rect -6955 20930 -6950 20950
rect -6950 20930 -6930 20950
rect -6930 20930 -6925 20950
rect -6955 20925 -6925 20930
rect -6875 20950 -6845 20955
rect -6875 20930 -6870 20950
rect -6870 20930 -6850 20950
rect -6850 20930 -6845 20950
rect -6875 20925 -6845 20930
rect -6795 20950 -6765 20955
rect -6795 20930 -6790 20950
rect -6790 20930 -6770 20950
rect -6770 20930 -6765 20950
rect -6795 20925 -6765 20930
rect -6715 20950 -6685 20955
rect -6715 20930 -6710 20950
rect -6710 20930 -6690 20950
rect -6690 20930 -6685 20950
rect -6715 20925 -6685 20930
rect -6635 20950 -6605 20955
rect -6635 20930 -6630 20950
rect -6630 20930 -6610 20950
rect -6610 20930 -6605 20950
rect -6635 20925 -6605 20930
rect -6555 20950 -6525 20955
rect -6555 20930 -6550 20950
rect -6550 20930 -6530 20950
rect -6530 20930 -6525 20950
rect -6555 20925 -6525 20930
rect -6475 20950 -6445 20955
rect -6475 20930 -6470 20950
rect -6470 20930 -6450 20950
rect -6450 20930 -6445 20950
rect -6475 20925 -6445 20930
rect -6395 20950 -6365 20955
rect -6395 20930 -6390 20950
rect -6390 20930 -6370 20950
rect -6370 20930 -6365 20950
rect -6395 20925 -6365 20930
rect -6315 20950 -6285 20955
rect -6315 20930 -6310 20950
rect -6310 20930 -6290 20950
rect -6290 20930 -6285 20950
rect -6315 20925 -6285 20930
rect -6235 20950 -6205 20955
rect -6235 20930 -6230 20950
rect -6230 20930 -6210 20950
rect -6210 20930 -6205 20950
rect -6235 20925 -6205 20930
rect -6155 20950 -6125 20955
rect -6155 20930 -6150 20950
rect -6150 20930 -6130 20950
rect -6130 20930 -6125 20950
rect -6155 20925 -6125 20930
rect -5675 20950 -5645 20955
rect -5675 20930 -5670 20950
rect -5670 20930 -5650 20950
rect -5650 20930 -5645 20950
rect -5675 20925 -5645 20930
rect -5595 20950 -5565 20955
rect -5595 20930 -5590 20950
rect -5590 20930 -5570 20950
rect -5570 20930 -5565 20950
rect -5595 20925 -5565 20930
rect -5515 20950 -5485 20955
rect -5515 20930 -5510 20950
rect -5510 20930 -5490 20950
rect -5490 20930 -5485 20950
rect -5515 20925 -5485 20930
rect -5435 20950 -5405 20955
rect -5435 20930 -5430 20950
rect -5430 20930 -5410 20950
rect -5410 20930 -5405 20950
rect -5435 20925 -5405 20930
rect -5355 20950 -5325 20955
rect -5355 20930 -5350 20950
rect -5350 20930 -5330 20950
rect -5330 20930 -5325 20950
rect -5355 20925 -5325 20930
rect -5275 20950 -5245 20955
rect -5275 20930 -5270 20950
rect -5270 20930 -5250 20950
rect -5250 20930 -5245 20950
rect -5275 20925 -5245 20930
rect -5195 20950 -5165 20955
rect -5195 20930 -5190 20950
rect -5190 20930 -5170 20950
rect -5170 20930 -5165 20950
rect -5195 20925 -5165 20930
rect -5115 20950 -5085 20955
rect -5115 20930 -5110 20950
rect -5110 20930 -5090 20950
rect -5090 20930 -5085 20950
rect -5115 20925 -5085 20930
rect -5035 20950 -5005 20955
rect -5035 20930 -5030 20950
rect -5030 20930 -5010 20950
rect -5010 20930 -5005 20950
rect -5035 20925 -5005 20930
rect -4955 20950 -4925 20955
rect -4955 20930 -4950 20950
rect -4950 20930 -4930 20950
rect -4930 20930 -4925 20950
rect -4955 20925 -4925 20930
rect -4875 20950 -4845 20955
rect -4875 20930 -4870 20950
rect -4870 20930 -4850 20950
rect -4850 20930 -4845 20950
rect -4875 20925 -4845 20930
rect -4795 20950 -4765 20955
rect -4795 20930 -4790 20950
rect -4790 20930 -4770 20950
rect -4770 20930 -4765 20950
rect -4795 20925 -4765 20930
rect -4715 20950 -4685 20955
rect -4715 20930 -4710 20950
rect -4710 20930 -4690 20950
rect -4690 20930 -4685 20950
rect -4715 20925 -4685 20930
rect -4635 20950 -4605 20955
rect -4635 20930 -4630 20950
rect -4630 20930 -4610 20950
rect -4610 20930 -4605 20950
rect -4635 20925 -4605 20930
rect -4555 20950 -4525 20955
rect -4555 20930 -4550 20950
rect -4550 20930 -4530 20950
rect -4530 20930 -4525 20950
rect -4555 20925 -4525 20930
rect -4475 20950 -4445 20955
rect -4475 20930 -4470 20950
rect -4470 20930 -4450 20950
rect -4450 20930 -4445 20950
rect -4475 20925 -4445 20930
rect -4395 20950 -4365 20955
rect -4395 20930 -4390 20950
rect -4390 20930 -4370 20950
rect -4370 20930 -4365 20950
rect -4395 20925 -4365 20930
rect -4315 20950 -4285 20955
rect -4315 20930 -4310 20950
rect -4310 20930 -4290 20950
rect -4290 20930 -4285 20950
rect -4315 20925 -4285 20930
rect -4235 20950 -4205 20955
rect -4235 20930 -4230 20950
rect -4230 20930 -4210 20950
rect -4210 20930 -4205 20950
rect -4235 20925 -4205 20930
rect -4155 20950 -4125 20955
rect -4155 20930 -4150 20950
rect -4150 20930 -4130 20950
rect -4130 20930 -4125 20950
rect -4155 20925 -4125 20930
rect -4075 20950 -4045 20955
rect -4075 20930 -4070 20950
rect -4070 20930 -4050 20950
rect -4050 20930 -4045 20950
rect -4075 20925 -4045 20930
rect -3995 20950 -3965 20955
rect -3995 20930 -3990 20950
rect -3990 20930 -3970 20950
rect -3970 20930 -3965 20950
rect -3995 20925 -3965 20930
rect -3915 20950 -3885 20955
rect -3915 20930 -3910 20950
rect -3910 20930 -3890 20950
rect -3890 20930 -3885 20950
rect -3915 20925 -3885 20930
rect -3835 20950 -3805 20955
rect -3835 20930 -3830 20950
rect -3830 20930 -3810 20950
rect -3810 20930 -3805 20950
rect -3835 20925 -3805 20930
rect -3755 20950 -3725 20955
rect -3755 20930 -3750 20950
rect -3750 20930 -3730 20950
rect -3730 20930 -3725 20950
rect -3755 20925 -3725 20930
rect -3675 20950 -3645 20955
rect -3675 20930 -3670 20950
rect -3670 20930 -3650 20950
rect -3650 20930 -3645 20950
rect -3675 20925 -3645 20930
rect -3595 20950 -3565 20955
rect -3595 20930 -3590 20950
rect -3590 20930 -3570 20950
rect -3570 20930 -3565 20950
rect -3595 20925 -3565 20930
rect -3515 20950 -3485 20955
rect -3515 20930 -3510 20950
rect -3510 20930 -3490 20950
rect -3490 20930 -3485 20950
rect -3515 20925 -3485 20930
rect -3435 20950 -3405 20955
rect -3435 20930 -3430 20950
rect -3430 20930 -3410 20950
rect -3410 20930 -3405 20950
rect -3435 20925 -3405 20930
rect -3355 20950 -3325 20955
rect -3355 20930 -3350 20950
rect -3350 20930 -3330 20950
rect -3330 20930 -3325 20950
rect -3355 20925 -3325 20930
rect -3275 20950 -3245 20955
rect -3275 20930 -3270 20950
rect -3270 20930 -3250 20950
rect -3250 20930 -3245 20950
rect -3275 20925 -3245 20930
rect -3195 20950 -3165 20955
rect -3195 20930 -3190 20950
rect -3190 20930 -3170 20950
rect -3170 20930 -3165 20950
rect -3195 20925 -3165 20930
rect -3115 20950 -3085 20955
rect -3115 20930 -3110 20950
rect -3110 20930 -3090 20950
rect -3090 20930 -3085 20950
rect -3115 20925 -3085 20930
rect -3035 20950 -3005 20955
rect -3035 20930 -3030 20950
rect -3030 20930 -3010 20950
rect -3010 20930 -3005 20950
rect -3035 20925 -3005 20930
rect -2955 20950 -2925 20955
rect -2955 20930 -2950 20950
rect -2950 20930 -2930 20950
rect -2930 20930 -2925 20950
rect -2955 20925 -2925 20930
rect -2875 20950 -2845 20955
rect -2875 20930 -2870 20950
rect -2870 20930 -2850 20950
rect -2850 20930 -2845 20950
rect -2875 20925 -2845 20930
rect -2795 20950 -2765 20955
rect -2795 20930 -2790 20950
rect -2790 20930 -2770 20950
rect -2770 20930 -2765 20950
rect -2795 20925 -2765 20930
rect -2715 20950 -2685 20955
rect -2715 20930 -2710 20950
rect -2710 20930 -2690 20950
rect -2690 20930 -2685 20950
rect -2715 20925 -2685 20930
rect -2635 20950 -2605 20955
rect -2635 20930 -2630 20950
rect -2630 20930 -2610 20950
rect -2610 20930 -2605 20950
rect -2635 20925 -2605 20930
rect -2555 20950 -2525 20955
rect -2555 20930 -2550 20950
rect -2550 20930 -2530 20950
rect -2530 20930 -2525 20950
rect -2555 20925 -2525 20930
rect -2475 20950 -2445 20955
rect -2475 20930 -2470 20950
rect -2470 20930 -2450 20950
rect -2450 20930 -2445 20950
rect -2475 20925 -2445 20930
rect -2395 20950 -2365 20955
rect -2395 20930 -2390 20950
rect -2390 20930 -2370 20950
rect -2370 20930 -2365 20950
rect -2395 20925 -2365 20930
rect -2315 20950 -2285 20955
rect -2315 20930 -2310 20950
rect -2310 20930 -2290 20950
rect -2290 20930 -2285 20950
rect -2315 20925 -2285 20930
rect -2235 20950 -2205 20955
rect -2235 20930 -2230 20950
rect -2230 20930 -2210 20950
rect -2210 20930 -2205 20950
rect -2235 20925 -2205 20930
rect -2155 20950 -2125 20955
rect -2155 20930 -2150 20950
rect -2150 20930 -2130 20950
rect -2130 20930 -2125 20950
rect -2155 20925 -2125 20930
rect -2075 20950 -2045 20955
rect -2075 20930 -2070 20950
rect -2070 20930 -2050 20950
rect -2050 20930 -2045 20950
rect -2075 20925 -2045 20930
rect -1995 20950 -1965 20955
rect -1995 20930 -1990 20950
rect -1990 20930 -1970 20950
rect -1970 20930 -1965 20950
rect -1995 20925 -1965 20930
rect -1835 20950 -1805 20955
rect -1835 20930 -1830 20950
rect -1830 20930 -1810 20950
rect -1810 20930 -1805 20950
rect -1835 20925 -1805 20930
rect -1755 20950 -1725 20955
rect -1755 20930 -1750 20950
rect -1750 20930 -1730 20950
rect -1730 20930 -1725 20950
rect -1755 20925 -1725 20930
rect -1675 20950 -1645 20955
rect -1675 20930 -1670 20950
rect -1670 20930 -1650 20950
rect -1650 20930 -1645 20950
rect -1675 20925 -1645 20930
rect -1515 20950 -1485 20955
rect -1515 20930 -1510 20950
rect -1510 20930 -1490 20950
rect -1490 20930 -1485 20950
rect -1515 20925 -1485 20930
rect -1355 20950 -1325 20955
rect -1355 20930 -1350 20950
rect -1350 20930 -1330 20950
rect -1330 20930 -1325 20950
rect -1355 20925 -1325 20930
rect -1275 20950 -1245 20955
rect -1275 20930 -1270 20950
rect -1270 20930 -1250 20950
rect -1250 20930 -1245 20950
rect -1275 20925 -1245 20930
rect -1195 20950 -1165 20955
rect -1195 20930 -1190 20950
rect -1190 20930 -1170 20950
rect -1170 20930 -1165 20950
rect -1195 20925 -1165 20930
rect -1115 20950 -1085 20955
rect -1115 20930 -1110 20950
rect -1110 20930 -1090 20950
rect -1090 20930 -1085 20950
rect -1115 20925 -1085 20930
rect -1035 20950 -1005 20955
rect -1035 20930 -1030 20950
rect -1030 20930 -1010 20950
rect -1010 20930 -1005 20950
rect -1035 20925 -1005 20930
rect -875 20950 -845 20955
rect -875 20930 -870 20950
rect -870 20930 -850 20950
rect -850 20930 -845 20950
rect -875 20925 -845 20930
rect -715 20950 -685 20955
rect -715 20930 -710 20950
rect -710 20930 -690 20950
rect -690 20930 -685 20950
rect -715 20925 -685 20930
rect -555 20950 -525 20955
rect -555 20930 -550 20950
rect -550 20930 -530 20950
rect -530 20930 -525 20950
rect -555 20925 -525 20930
rect -16555 20670 -16525 20675
rect -16555 20650 -16550 20670
rect -16550 20650 -16530 20670
rect -16530 20650 -16525 20670
rect -16555 20645 -16525 20650
rect -16475 20670 -16445 20675
rect -16475 20650 -16470 20670
rect -16470 20650 -16450 20670
rect -16450 20650 -16445 20670
rect -16475 20645 -16445 20650
rect -16395 20670 -16365 20675
rect -16395 20650 -16390 20670
rect -16390 20650 -16370 20670
rect -16370 20650 -16365 20670
rect -16395 20645 -16365 20650
rect -16315 20670 -16285 20675
rect -16315 20650 -16310 20670
rect -16310 20650 -16290 20670
rect -16290 20650 -16285 20670
rect -16315 20645 -16285 20650
rect -16235 20670 -16205 20675
rect -16235 20650 -16230 20670
rect -16230 20650 -16210 20670
rect -16210 20650 -16205 20670
rect -16235 20645 -16205 20650
rect -16155 20670 -16125 20675
rect -16155 20650 -16150 20670
rect -16150 20650 -16130 20670
rect -16130 20650 -16125 20670
rect -16155 20645 -16125 20650
rect -16075 20670 -16045 20675
rect -16075 20650 -16070 20670
rect -16070 20650 -16050 20670
rect -16050 20650 -16045 20670
rect -16075 20645 -16045 20650
rect -15995 20670 -15965 20675
rect -15995 20650 -15990 20670
rect -15990 20650 -15970 20670
rect -15970 20650 -15965 20670
rect -15995 20645 -15965 20650
rect -15915 20670 -15885 20675
rect -15915 20650 -15910 20670
rect -15910 20650 -15890 20670
rect -15890 20650 -15885 20670
rect -15915 20645 -15885 20650
rect -15835 20670 -15805 20675
rect -15835 20650 -15830 20670
rect -15830 20650 -15810 20670
rect -15810 20650 -15805 20670
rect -15835 20645 -15805 20650
rect -15755 20670 -15725 20675
rect -15755 20650 -15750 20670
rect -15750 20650 -15730 20670
rect -15730 20650 -15725 20670
rect -15755 20645 -15725 20650
rect -15675 20670 -15645 20675
rect -15675 20650 -15670 20670
rect -15670 20650 -15650 20670
rect -15650 20650 -15645 20670
rect -15675 20645 -15645 20650
rect -15595 20670 -15565 20675
rect -15595 20650 -15590 20670
rect -15590 20650 -15570 20670
rect -15570 20650 -15565 20670
rect -15595 20645 -15565 20650
rect -14955 20670 -14925 20675
rect -14955 20650 -14950 20670
rect -14950 20650 -14930 20670
rect -14930 20650 -14925 20670
rect -14955 20645 -14925 20650
rect -14875 20670 -14845 20675
rect -14875 20650 -14870 20670
rect -14870 20650 -14850 20670
rect -14850 20650 -14845 20670
rect -14875 20645 -14845 20650
rect -14795 20670 -14765 20675
rect -14795 20650 -14790 20670
rect -14790 20650 -14770 20670
rect -14770 20650 -14765 20670
rect -14795 20645 -14765 20650
rect -14715 20670 -14685 20675
rect -14715 20650 -14710 20670
rect -14710 20650 -14690 20670
rect -14690 20650 -14685 20670
rect -14715 20645 -14685 20650
rect -14635 20670 -14605 20675
rect -14635 20650 -14630 20670
rect -14630 20650 -14610 20670
rect -14610 20650 -14605 20670
rect -14635 20645 -14605 20650
rect -14555 20670 -14525 20675
rect -14555 20650 -14550 20670
rect -14550 20650 -14530 20670
rect -14530 20650 -14525 20670
rect -14555 20645 -14525 20650
rect -14475 20670 -14445 20675
rect -14475 20650 -14470 20670
rect -14470 20650 -14450 20670
rect -14450 20650 -14445 20670
rect -14475 20645 -14445 20650
rect -14395 20670 -14365 20675
rect -14395 20650 -14390 20670
rect -14390 20650 -14370 20670
rect -14370 20650 -14365 20670
rect -14395 20645 -14365 20650
rect -14315 20670 -14285 20675
rect -14315 20650 -14310 20670
rect -14310 20650 -14290 20670
rect -14290 20650 -14285 20670
rect -14315 20645 -14285 20650
rect -14235 20670 -14205 20675
rect -14235 20650 -14230 20670
rect -14230 20650 -14210 20670
rect -14210 20650 -14205 20670
rect -14235 20645 -14205 20650
rect -14155 20670 -14125 20675
rect -14155 20650 -14150 20670
rect -14150 20650 -14130 20670
rect -14130 20650 -14125 20670
rect -14155 20645 -14125 20650
rect -14075 20670 -14045 20675
rect -14075 20650 -14070 20670
rect -14070 20650 -14050 20670
rect -14050 20650 -14045 20670
rect -14075 20645 -14045 20650
rect -13995 20670 -13965 20675
rect -13995 20650 -13990 20670
rect -13990 20650 -13970 20670
rect -13970 20650 -13965 20670
rect -13995 20645 -13965 20650
rect -13915 20670 -13885 20675
rect -13915 20650 -13910 20670
rect -13910 20650 -13890 20670
rect -13890 20650 -13885 20670
rect -13915 20645 -13885 20650
rect -13835 20670 -13805 20675
rect -13835 20650 -13830 20670
rect -13830 20650 -13810 20670
rect -13810 20650 -13805 20670
rect -13835 20645 -13805 20650
rect -13755 20670 -13725 20675
rect -13755 20650 -13750 20670
rect -13750 20650 -13730 20670
rect -13730 20650 -13725 20670
rect -13755 20645 -13725 20650
rect -13675 20670 -13645 20675
rect -13675 20650 -13670 20670
rect -13670 20650 -13650 20670
rect -13650 20650 -13645 20670
rect -13675 20645 -13645 20650
rect -13595 20670 -13565 20675
rect -13595 20650 -13590 20670
rect -13590 20650 -13570 20670
rect -13570 20650 -13565 20670
rect -13595 20645 -13565 20650
rect -13515 20670 -13485 20675
rect -13515 20650 -13510 20670
rect -13510 20650 -13490 20670
rect -13490 20650 -13485 20670
rect -13515 20645 -13485 20650
rect -13435 20670 -13405 20675
rect -13435 20650 -13430 20670
rect -13430 20650 -13410 20670
rect -13410 20650 -13405 20670
rect -13435 20645 -13405 20650
rect -13355 20670 -13325 20675
rect -13355 20650 -13350 20670
rect -13350 20650 -13330 20670
rect -13330 20650 -13325 20670
rect -13355 20645 -13325 20650
rect -13275 20670 -13245 20675
rect -13275 20650 -13270 20670
rect -13270 20650 -13250 20670
rect -13250 20650 -13245 20670
rect -13275 20645 -13245 20650
rect -13195 20670 -13165 20675
rect -13195 20650 -13190 20670
rect -13190 20650 -13170 20670
rect -13170 20650 -13165 20670
rect -13195 20645 -13165 20650
rect -13115 20670 -13085 20675
rect -13115 20650 -13110 20670
rect -13110 20650 -13090 20670
rect -13090 20650 -13085 20670
rect -13115 20645 -13085 20650
rect -13035 20670 -13005 20675
rect -13035 20650 -13030 20670
rect -13030 20650 -13010 20670
rect -13010 20650 -13005 20670
rect -13035 20645 -13005 20650
rect -12955 20670 -12925 20675
rect -12955 20650 -12950 20670
rect -12950 20650 -12930 20670
rect -12930 20650 -12925 20670
rect -12955 20645 -12925 20650
rect -12875 20670 -12845 20675
rect -12875 20650 -12870 20670
rect -12870 20650 -12850 20670
rect -12850 20650 -12845 20670
rect -12875 20645 -12845 20650
rect -12795 20670 -12765 20675
rect -12795 20650 -12790 20670
rect -12790 20650 -12770 20670
rect -12770 20650 -12765 20670
rect -12795 20645 -12765 20650
rect -12715 20670 -12685 20675
rect -12715 20650 -12710 20670
rect -12710 20650 -12690 20670
rect -12690 20650 -12685 20670
rect -12715 20645 -12685 20650
rect -12635 20670 -12605 20675
rect -12635 20650 -12630 20670
rect -12630 20650 -12610 20670
rect -12610 20650 -12605 20670
rect -12635 20645 -12605 20650
rect -12555 20670 -12525 20675
rect -12555 20650 -12550 20670
rect -12550 20650 -12530 20670
rect -12530 20650 -12525 20670
rect -12555 20645 -12525 20650
rect -12475 20670 -12445 20675
rect -12475 20650 -12470 20670
rect -12470 20650 -12450 20670
rect -12450 20650 -12445 20670
rect -12475 20645 -12445 20650
rect -12395 20670 -12365 20675
rect -12395 20650 -12390 20670
rect -12390 20650 -12370 20670
rect -12370 20650 -12365 20670
rect -12395 20645 -12365 20650
rect -12315 20670 -12285 20675
rect -12315 20650 -12310 20670
rect -12310 20650 -12290 20670
rect -12290 20650 -12285 20670
rect -12315 20645 -12285 20650
rect -12235 20670 -12205 20675
rect -12235 20650 -12230 20670
rect -12230 20650 -12210 20670
rect -12210 20650 -12205 20670
rect -12235 20645 -12205 20650
rect -12155 20670 -12125 20675
rect -12155 20650 -12150 20670
rect -12150 20650 -12130 20670
rect -12130 20650 -12125 20670
rect -12155 20645 -12125 20650
rect -12075 20670 -12045 20675
rect -12075 20650 -12070 20670
rect -12070 20650 -12050 20670
rect -12050 20650 -12045 20670
rect -12075 20645 -12045 20650
rect -11995 20670 -11965 20675
rect -11995 20650 -11990 20670
rect -11990 20650 -11970 20670
rect -11970 20650 -11965 20670
rect -11995 20645 -11965 20650
rect -11915 20670 -11885 20675
rect -11915 20650 -11910 20670
rect -11910 20650 -11890 20670
rect -11890 20650 -11885 20670
rect -11915 20645 -11885 20650
rect -11835 20670 -11805 20675
rect -11835 20650 -11830 20670
rect -11830 20650 -11810 20670
rect -11810 20650 -11805 20670
rect -11835 20645 -11805 20650
rect -11755 20670 -11725 20675
rect -11755 20650 -11750 20670
rect -11750 20650 -11730 20670
rect -11730 20650 -11725 20670
rect -11755 20645 -11725 20650
rect -11675 20670 -11645 20675
rect -11675 20650 -11670 20670
rect -11670 20650 -11650 20670
rect -11650 20650 -11645 20670
rect -11675 20645 -11645 20650
rect -11595 20670 -11565 20675
rect -11595 20650 -11590 20670
rect -11590 20650 -11570 20670
rect -11570 20650 -11565 20670
rect -11595 20645 -11565 20650
rect -11515 20670 -11485 20675
rect -11515 20650 -11510 20670
rect -11510 20650 -11490 20670
rect -11490 20650 -11485 20670
rect -11515 20645 -11485 20650
rect -11435 20670 -11405 20675
rect -11435 20650 -11430 20670
rect -11430 20650 -11410 20670
rect -11410 20650 -11405 20670
rect -11435 20645 -11405 20650
rect -11355 20670 -11325 20675
rect -11355 20650 -11350 20670
rect -11350 20650 -11330 20670
rect -11330 20650 -11325 20670
rect -11355 20645 -11325 20650
rect -11275 20670 -11245 20675
rect -11275 20650 -11270 20670
rect -11270 20650 -11250 20670
rect -11250 20650 -11245 20670
rect -11275 20645 -11245 20650
rect -11195 20670 -11165 20675
rect -11195 20650 -11190 20670
rect -11190 20650 -11170 20670
rect -11170 20650 -11165 20670
rect -11195 20645 -11165 20650
rect -11115 20670 -11085 20675
rect -11115 20650 -11110 20670
rect -11110 20650 -11090 20670
rect -11090 20650 -11085 20670
rect -11115 20645 -11085 20650
rect -11035 20670 -11005 20675
rect -11035 20650 -11030 20670
rect -11030 20650 -11010 20670
rect -11010 20650 -11005 20670
rect -11035 20645 -11005 20650
rect -10955 20670 -10925 20675
rect -10955 20650 -10950 20670
rect -10950 20650 -10930 20670
rect -10930 20650 -10925 20670
rect -10955 20645 -10925 20650
rect -10875 20670 -10845 20675
rect -10875 20650 -10870 20670
rect -10870 20650 -10850 20670
rect -10850 20650 -10845 20670
rect -10875 20645 -10845 20650
rect -10795 20670 -10765 20675
rect -10795 20650 -10790 20670
rect -10790 20650 -10770 20670
rect -10770 20650 -10765 20670
rect -10795 20645 -10765 20650
rect -10715 20670 -10685 20675
rect -10715 20650 -10710 20670
rect -10710 20650 -10690 20670
rect -10690 20650 -10685 20670
rect -10715 20645 -10685 20650
rect -10635 20670 -10605 20675
rect -10635 20650 -10630 20670
rect -10630 20650 -10610 20670
rect -10610 20650 -10605 20670
rect -10635 20645 -10605 20650
rect -10555 20670 -10525 20675
rect -10555 20650 -10550 20670
rect -10550 20650 -10530 20670
rect -10530 20650 -10525 20670
rect -10555 20645 -10525 20650
rect -10475 20670 -10445 20675
rect -10475 20650 -10470 20670
rect -10470 20650 -10450 20670
rect -10450 20650 -10445 20670
rect -10475 20645 -10445 20650
rect -10395 20670 -10365 20675
rect -10395 20650 -10390 20670
rect -10390 20650 -10370 20670
rect -10370 20650 -10365 20670
rect -10395 20645 -10365 20650
rect -10315 20670 -10285 20675
rect -10315 20650 -10310 20670
rect -10310 20650 -10290 20670
rect -10290 20650 -10285 20670
rect -10315 20645 -10285 20650
rect -10235 20670 -10205 20675
rect -10235 20650 -10230 20670
rect -10230 20650 -10210 20670
rect -10210 20650 -10205 20670
rect -10235 20645 -10205 20650
rect -10155 20670 -10125 20675
rect -10155 20650 -10150 20670
rect -10150 20650 -10130 20670
rect -10130 20650 -10125 20670
rect -10155 20645 -10125 20650
rect -10075 20670 -10045 20675
rect -10075 20650 -10070 20670
rect -10070 20650 -10050 20670
rect -10050 20650 -10045 20670
rect -10075 20645 -10045 20650
rect -9995 20670 -9965 20675
rect -9995 20650 -9990 20670
rect -9990 20650 -9970 20670
rect -9970 20650 -9965 20670
rect -9995 20645 -9965 20650
rect -9915 20670 -9885 20675
rect -9915 20650 -9910 20670
rect -9910 20650 -9890 20670
rect -9890 20650 -9885 20670
rect -9915 20645 -9885 20650
rect -9835 20670 -9805 20675
rect -9835 20650 -9830 20670
rect -9830 20650 -9810 20670
rect -9810 20650 -9805 20670
rect -9835 20645 -9805 20650
rect -9755 20670 -9725 20675
rect -9755 20650 -9750 20670
rect -9750 20650 -9730 20670
rect -9730 20650 -9725 20670
rect -9755 20645 -9725 20650
rect -9675 20670 -9645 20675
rect -9675 20650 -9670 20670
rect -9670 20650 -9650 20670
rect -9650 20650 -9645 20670
rect -9675 20645 -9645 20650
rect -9595 20670 -9565 20675
rect -9595 20650 -9590 20670
rect -9590 20650 -9570 20670
rect -9570 20650 -9565 20670
rect -9595 20645 -9565 20650
rect -9515 20670 -9485 20675
rect -9515 20650 -9510 20670
rect -9510 20650 -9490 20670
rect -9490 20650 -9485 20670
rect -9515 20645 -9485 20650
rect -9435 20670 -9405 20675
rect -9435 20650 -9430 20670
rect -9430 20650 -9410 20670
rect -9410 20650 -9405 20670
rect -9435 20645 -9405 20650
rect -9355 20670 -9325 20675
rect -9355 20650 -9350 20670
rect -9350 20650 -9330 20670
rect -9330 20650 -9325 20670
rect -9355 20645 -9325 20650
rect -9275 20670 -9245 20675
rect -9275 20650 -9270 20670
rect -9270 20650 -9250 20670
rect -9250 20650 -9245 20670
rect -9275 20645 -9245 20650
rect -9195 20670 -9165 20675
rect -9195 20650 -9190 20670
rect -9190 20650 -9170 20670
rect -9170 20650 -9165 20670
rect -9195 20645 -9165 20650
rect -9115 20670 -9085 20675
rect -9115 20650 -9110 20670
rect -9110 20650 -9090 20670
rect -9090 20650 -9085 20670
rect -9115 20645 -9085 20650
rect -9035 20670 -9005 20675
rect -9035 20650 -9030 20670
rect -9030 20650 -9010 20670
rect -9010 20650 -9005 20670
rect -9035 20645 -9005 20650
rect -8955 20670 -8925 20675
rect -8955 20650 -8950 20670
rect -8950 20650 -8930 20670
rect -8930 20650 -8925 20670
rect -8955 20645 -8925 20650
rect -8875 20670 -8845 20675
rect -8875 20650 -8870 20670
rect -8870 20650 -8850 20670
rect -8850 20650 -8845 20670
rect -8875 20645 -8845 20650
rect -8795 20670 -8765 20675
rect -8795 20650 -8790 20670
rect -8790 20650 -8770 20670
rect -8770 20650 -8765 20670
rect -8795 20645 -8765 20650
rect -8715 20670 -8685 20675
rect -8715 20650 -8710 20670
rect -8710 20650 -8690 20670
rect -8690 20650 -8685 20670
rect -8715 20645 -8685 20650
rect -8635 20670 -8605 20675
rect -8635 20650 -8630 20670
rect -8630 20650 -8610 20670
rect -8610 20650 -8605 20670
rect -8635 20645 -8605 20650
rect -8555 20670 -8525 20675
rect -8555 20650 -8550 20670
rect -8550 20650 -8530 20670
rect -8530 20650 -8525 20670
rect -8555 20645 -8525 20650
rect -8475 20670 -8445 20675
rect -8475 20650 -8470 20670
rect -8470 20650 -8450 20670
rect -8450 20650 -8445 20670
rect -8475 20645 -8445 20650
rect -8395 20670 -8365 20675
rect -8395 20650 -8390 20670
rect -8390 20650 -8370 20670
rect -8370 20650 -8365 20670
rect -8395 20645 -8365 20650
rect -8315 20670 -8285 20675
rect -8315 20650 -8310 20670
rect -8310 20650 -8290 20670
rect -8290 20650 -8285 20670
rect -8315 20645 -8285 20650
rect -8235 20670 -8205 20675
rect -8235 20650 -8230 20670
rect -8230 20650 -8210 20670
rect -8210 20650 -8205 20670
rect -8235 20645 -8205 20650
rect -8155 20670 -8125 20675
rect -8155 20650 -8150 20670
rect -8150 20650 -8130 20670
rect -8130 20650 -8125 20670
rect -8155 20645 -8125 20650
rect -8075 20670 -8045 20675
rect -8075 20650 -8070 20670
rect -8070 20650 -8050 20670
rect -8050 20650 -8045 20670
rect -8075 20645 -8045 20650
rect -7995 20670 -7965 20675
rect -7995 20650 -7990 20670
rect -7990 20650 -7970 20670
rect -7970 20650 -7965 20670
rect -7995 20645 -7965 20650
rect -7915 20670 -7885 20675
rect -7915 20650 -7910 20670
rect -7910 20650 -7890 20670
rect -7890 20650 -7885 20670
rect -7915 20645 -7885 20650
rect -7835 20670 -7805 20675
rect -7835 20650 -7830 20670
rect -7830 20650 -7810 20670
rect -7810 20650 -7805 20670
rect -7835 20645 -7805 20650
rect -7755 20670 -7725 20675
rect -7755 20650 -7750 20670
rect -7750 20650 -7730 20670
rect -7730 20650 -7725 20670
rect -7755 20645 -7725 20650
rect -7675 20670 -7645 20675
rect -7675 20650 -7670 20670
rect -7670 20650 -7650 20670
rect -7650 20650 -7645 20670
rect -7675 20645 -7645 20650
rect -7595 20670 -7565 20675
rect -7595 20650 -7590 20670
rect -7590 20650 -7570 20670
rect -7570 20650 -7565 20670
rect -7595 20645 -7565 20650
rect -7515 20670 -7485 20675
rect -7515 20650 -7510 20670
rect -7510 20650 -7490 20670
rect -7490 20650 -7485 20670
rect -7515 20645 -7485 20650
rect -7435 20670 -7405 20675
rect -7435 20650 -7430 20670
rect -7430 20650 -7410 20670
rect -7410 20650 -7405 20670
rect -7435 20645 -7405 20650
rect -7355 20670 -7325 20675
rect -7355 20650 -7350 20670
rect -7350 20650 -7330 20670
rect -7330 20650 -7325 20670
rect -7355 20645 -7325 20650
rect -7275 20670 -7245 20675
rect -7275 20650 -7270 20670
rect -7270 20650 -7250 20670
rect -7250 20650 -7245 20670
rect -7275 20645 -7245 20650
rect -7195 20670 -7165 20675
rect -7195 20650 -7190 20670
rect -7190 20650 -7170 20670
rect -7170 20650 -7165 20670
rect -7195 20645 -7165 20650
rect -7115 20670 -7085 20675
rect -7115 20650 -7110 20670
rect -7110 20650 -7090 20670
rect -7090 20650 -7085 20670
rect -7115 20645 -7085 20650
rect -7035 20670 -7005 20675
rect -7035 20650 -7030 20670
rect -7030 20650 -7010 20670
rect -7010 20650 -7005 20670
rect -7035 20645 -7005 20650
rect -6955 20670 -6925 20675
rect -6955 20650 -6950 20670
rect -6950 20650 -6930 20670
rect -6930 20650 -6925 20670
rect -6955 20645 -6925 20650
rect -6875 20670 -6845 20675
rect -6875 20650 -6870 20670
rect -6870 20650 -6850 20670
rect -6850 20650 -6845 20670
rect -6875 20645 -6845 20650
rect -6795 20670 -6765 20675
rect -6795 20650 -6790 20670
rect -6790 20650 -6770 20670
rect -6770 20650 -6765 20670
rect -6795 20645 -6765 20650
rect -6715 20670 -6685 20675
rect -6715 20650 -6710 20670
rect -6710 20650 -6690 20670
rect -6690 20650 -6685 20670
rect -6715 20645 -6685 20650
rect -6635 20670 -6605 20675
rect -6635 20650 -6630 20670
rect -6630 20650 -6610 20670
rect -6610 20650 -6605 20670
rect -6635 20645 -6605 20650
rect -6555 20670 -6525 20675
rect -6555 20650 -6550 20670
rect -6550 20650 -6530 20670
rect -6530 20650 -6525 20670
rect -6555 20645 -6525 20650
rect -6475 20670 -6445 20675
rect -6475 20650 -6470 20670
rect -6470 20650 -6450 20670
rect -6450 20650 -6445 20670
rect -6475 20645 -6445 20650
rect -6395 20670 -6365 20675
rect -6395 20650 -6390 20670
rect -6390 20650 -6370 20670
rect -6370 20650 -6365 20670
rect -6395 20645 -6365 20650
rect -6315 20670 -6285 20675
rect -6315 20650 -6310 20670
rect -6310 20650 -6290 20670
rect -6290 20650 -6285 20670
rect -6315 20645 -6285 20650
rect -6235 20670 -6205 20675
rect -6235 20650 -6230 20670
rect -6230 20650 -6210 20670
rect -6210 20650 -6205 20670
rect -6235 20645 -6205 20650
rect -6155 20670 -6125 20675
rect -6155 20650 -6150 20670
rect -6150 20650 -6130 20670
rect -6130 20650 -6125 20670
rect -6155 20645 -6125 20650
rect -5675 20670 -5645 20675
rect -5675 20650 -5670 20670
rect -5670 20650 -5650 20670
rect -5650 20650 -5645 20670
rect -5675 20645 -5645 20650
rect -5595 20670 -5565 20675
rect -5595 20650 -5590 20670
rect -5590 20650 -5570 20670
rect -5570 20650 -5565 20670
rect -5595 20645 -5565 20650
rect -5515 20670 -5485 20675
rect -5515 20650 -5510 20670
rect -5510 20650 -5490 20670
rect -5490 20650 -5485 20670
rect -5515 20645 -5485 20650
rect -5435 20670 -5405 20675
rect -5435 20650 -5430 20670
rect -5430 20650 -5410 20670
rect -5410 20650 -5405 20670
rect -5435 20645 -5405 20650
rect -5355 20670 -5325 20675
rect -5355 20650 -5350 20670
rect -5350 20650 -5330 20670
rect -5330 20650 -5325 20670
rect -5355 20645 -5325 20650
rect -5275 20670 -5245 20675
rect -5275 20650 -5270 20670
rect -5270 20650 -5250 20670
rect -5250 20650 -5245 20670
rect -5275 20645 -5245 20650
rect -5195 20670 -5165 20675
rect -5195 20650 -5190 20670
rect -5190 20650 -5170 20670
rect -5170 20650 -5165 20670
rect -5195 20645 -5165 20650
rect -5115 20670 -5085 20675
rect -5115 20650 -5110 20670
rect -5110 20650 -5090 20670
rect -5090 20650 -5085 20670
rect -5115 20645 -5085 20650
rect -5035 20670 -5005 20675
rect -5035 20650 -5030 20670
rect -5030 20650 -5010 20670
rect -5010 20650 -5005 20670
rect -5035 20645 -5005 20650
rect -4955 20670 -4925 20675
rect -4955 20650 -4950 20670
rect -4950 20650 -4930 20670
rect -4930 20650 -4925 20670
rect -4955 20645 -4925 20650
rect -4875 20670 -4845 20675
rect -4875 20650 -4870 20670
rect -4870 20650 -4850 20670
rect -4850 20650 -4845 20670
rect -4875 20645 -4845 20650
rect -4795 20670 -4765 20675
rect -4795 20650 -4790 20670
rect -4790 20650 -4770 20670
rect -4770 20650 -4765 20670
rect -4795 20645 -4765 20650
rect -4715 20670 -4685 20675
rect -4715 20650 -4710 20670
rect -4710 20650 -4690 20670
rect -4690 20650 -4685 20670
rect -4715 20645 -4685 20650
rect -4635 20670 -4605 20675
rect -4635 20650 -4630 20670
rect -4630 20650 -4610 20670
rect -4610 20650 -4605 20670
rect -4635 20645 -4605 20650
rect -4555 20670 -4525 20675
rect -4555 20650 -4550 20670
rect -4550 20650 -4530 20670
rect -4530 20650 -4525 20670
rect -4555 20645 -4525 20650
rect -4475 20670 -4445 20675
rect -4475 20650 -4470 20670
rect -4470 20650 -4450 20670
rect -4450 20650 -4445 20670
rect -4475 20645 -4445 20650
rect -4395 20670 -4365 20675
rect -4395 20650 -4390 20670
rect -4390 20650 -4370 20670
rect -4370 20650 -4365 20670
rect -4395 20645 -4365 20650
rect -4315 20670 -4285 20675
rect -4315 20650 -4310 20670
rect -4310 20650 -4290 20670
rect -4290 20650 -4285 20670
rect -4315 20645 -4285 20650
rect -4235 20670 -4205 20675
rect -4235 20650 -4230 20670
rect -4230 20650 -4210 20670
rect -4210 20650 -4205 20670
rect -4235 20645 -4205 20650
rect -4155 20670 -4125 20675
rect -4155 20650 -4150 20670
rect -4150 20650 -4130 20670
rect -4130 20650 -4125 20670
rect -4155 20645 -4125 20650
rect -4075 20670 -4045 20675
rect -4075 20650 -4070 20670
rect -4070 20650 -4050 20670
rect -4050 20650 -4045 20670
rect -4075 20645 -4045 20650
rect -3995 20670 -3965 20675
rect -3995 20650 -3990 20670
rect -3990 20650 -3970 20670
rect -3970 20650 -3965 20670
rect -3995 20645 -3965 20650
rect -3915 20670 -3885 20675
rect -3915 20650 -3910 20670
rect -3910 20650 -3890 20670
rect -3890 20650 -3885 20670
rect -3915 20645 -3885 20650
rect -3835 20670 -3805 20675
rect -3835 20650 -3830 20670
rect -3830 20650 -3810 20670
rect -3810 20650 -3805 20670
rect -3835 20645 -3805 20650
rect -3755 20670 -3725 20675
rect -3755 20650 -3750 20670
rect -3750 20650 -3730 20670
rect -3730 20650 -3725 20670
rect -3755 20645 -3725 20650
rect -3675 20670 -3645 20675
rect -3675 20650 -3670 20670
rect -3670 20650 -3650 20670
rect -3650 20650 -3645 20670
rect -3675 20645 -3645 20650
rect -3595 20670 -3565 20675
rect -3595 20650 -3590 20670
rect -3590 20650 -3570 20670
rect -3570 20650 -3565 20670
rect -3595 20645 -3565 20650
rect -3515 20670 -3485 20675
rect -3515 20650 -3510 20670
rect -3510 20650 -3490 20670
rect -3490 20650 -3485 20670
rect -3515 20645 -3485 20650
rect -3435 20670 -3405 20675
rect -3435 20650 -3430 20670
rect -3430 20650 -3410 20670
rect -3410 20650 -3405 20670
rect -3435 20645 -3405 20650
rect -3355 20670 -3325 20675
rect -3355 20650 -3350 20670
rect -3350 20650 -3330 20670
rect -3330 20650 -3325 20670
rect -3355 20645 -3325 20650
rect -3275 20670 -3245 20675
rect -3275 20650 -3270 20670
rect -3270 20650 -3250 20670
rect -3250 20650 -3245 20670
rect -3275 20645 -3245 20650
rect -3195 20670 -3165 20675
rect -3195 20650 -3190 20670
rect -3190 20650 -3170 20670
rect -3170 20650 -3165 20670
rect -3195 20645 -3165 20650
rect -3115 20670 -3085 20675
rect -3115 20650 -3110 20670
rect -3110 20650 -3090 20670
rect -3090 20650 -3085 20670
rect -3115 20645 -3085 20650
rect -3035 20670 -3005 20675
rect -3035 20650 -3030 20670
rect -3030 20650 -3010 20670
rect -3010 20650 -3005 20670
rect -3035 20645 -3005 20650
rect -2955 20670 -2925 20675
rect -2955 20650 -2950 20670
rect -2950 20650 -2930 20670
rect -2930 20650 -2925 20670
rect -2955 20645 -2925 20650
rect -2875 20670 -2845 20675
rect -2875 20650 -2870 20670
rect -2870 20650 -2850 20670
rect -2850 20650 -2845 20670
rect -2875 20645 -2845 20650
rect -2795 20670 -2765 20675
rect -2795 20650 -2790 20670
rect -2790 20650 -2770 20670
rect -2770 20650 -2765 20670
rect -2795 20645 -2765 20650
rect -2715 20670 -2685 20675
rect -2715 20650 -2710 20670
rect -2710 20650 -2690 20670
rect -2690 20650 -2685 20670
rect -2715 20645 -2685 20650
rect -2635 20670 -2605 20675
rect -2635 20650 -2630 20670
rect -2630 20650 -2610 20670
rect -2610 20650 -2605 20670
rect -2635 20645 -2605 20650
rect -2555 20670 -2525 20675
rect -2555 20650 -2550 20670
rect -2550 20650 -2530 20670
rect -2530 20650 -2525 20670
rect -2555 20645 -2525 20650
rect -2475 20670 -2445 20675
rect -2475 20650 -2470 20670
rect -2470 20650 -2450 20670
rect -2450 20650 -2445 20670
rect -2475 20645 -2445 20650
rect -2395 20670 -2365 20675
rect -2395 20650 -2390 20670
rect -2390 20650 -2370 20670
rect -2370 20650 -2365 20670
rect -2395 20645 -2365 20650
rect -2315 20670 -2285 20675
rect -2315 20650 -2310 20670
rect -2310 20650 -2290 20670
rect -2290 20650 -2285 20670
rect -2315 20645 -2285 20650
rect -2235 20670 -2205 20675
rect -2235 20650 -2230 20670
rect -2230 20650 -2210 20670
rect -2210 20650 -2205 20670
rect -2235 20645 -2205 20650
rect -2155 20670 -2125 20675
rect -2155 20650 -2150 20670
rect -2150 20650 -2130 20670
rect -2130 20650 -2125 20670
rect -2155 20645 -2125 20650
rect -2075 20670 -2045 20675
rect -2075 20650 -2070 20670
rect -2070 20650 -2050 20670
rect -2050 20650 -2045 20670
rect -2075 20645 -2045 20650
rect -1995 20670 -1965 20675
rect -1995 20650 -1990 20670
rect -1990 20650 -1970 20670
rect -1970 20650 -1965 20670
rect -1995 20645 -1965 20650
rect -1835 20670 -1805 20675
rect -1835 20650 -1830 20670
rect -1830 20650 -1810 20670
rect -1810 20650 -1805 20670
rect -1835 20645 -1805 20650
rect -1755 20670 -1725 20675
rect -1755 20650 -1750 20670
rect -1750 20650 -1730 20670
rect -1730 20650 -1725 20670
rect -1755 20645 -1725 20650
rect 20525 20670 20555 20675
rect 20525 20650 20530 20670
rect 20530 20650 20550 20670
rect 20550 20650 20555 20670
rect 20525 20645 20555 20650
rect 20605 20670 20635 20675
rect 20605 20650 20610 20670
rect 20610 20650 20630 20670
rect 20630 20650 20635 20670
rect 20605 20645 20635 20650
rect 20685 20670 20715 20675
rect 20685 20650 20690 20670
rect 20690 20650 20710 20670
rect 20710 20650 20715 20670
rect 20685 20645 20715 20650
rect 20765 20670 20795 20675
rect 20765 20650 20770 20670
rect 20770 20650 20790 20670
rect 20790 20650 20795 20670
rect 20765 20645 20795 20650
rect 20845 20670 20875 20675
rect 20845 20650 20850 20670
rect 20850 20650 20870 20670
rect 20870 20650 20875 20670
rect 20845 20645 20875 20650
rect 20925 20670 20955 20675
rect 20925 20650 20930 20670
rect 20930 20650 20950 20670
rect 20950 20650 20955 20670
rect 20925 20645 20955 20650
rect 21005 20670 21035 20675
rect 21005 20650 21010 20670
rect 21010 20650 21030 20670
rect 21030 20650 21035 20670
rect 21005 20645 21035 20650
rect 21085 20670 21115 20675
rect 21085 20650 21090 20670
rect 21090 20650 21110 20670
rect 21110 20650 21115 20670
rect 21085 20645 21115 20650
rect 21165 20670 21195 20675
rect 21165 20650 21170 20670
rect 21170 20650 21190 20670
rect 21190 20650 21195 20670
rect 21165 20645 21195 20650
rect 21245 20670 21275 20675
rect 21245 20650 21250 20670
rect 21250 20650 21270 20670
rect 21270 20650 21275 20670
rect 21245 20645 21275 20650
rect 21325 20670 21355 20675
rect 21325 20650 21330 20670
rect 21330 20650 21350 20670
rect 21350 20650 21355 20670
rect 21325 20645 21355 20650
rect 21405 20670 21435 20675
rect 21405 20650 21410 20670
rect 21410 20650 21430 20670
rect 21430 20650 21435 20670
rect 21405 20645 21435 20650
rect 21485 20670 21515 20675
rect 21485 20650 21490 20670
rect 21490 20650 21510 20670
rect 21510 20650 21515 20670
rect 21485 20645 21515 20650
rect 21565 20670 21595 20675
rect 21565 20650 21570 20670
rect 21570 20650 21590 20670
rect 21590 20650 21595 20670
rect 21565 20645 21595 20650
rect -16555 20510 -16525 20515
rect -16555 20490 -16550 20510
rect -16550 20490 -16530 20510
rect -16530 20490 -16525 20510
rect -16555 20485 -16525 20490
rect -16475 20510 -16445 20515
rect -16475 20490 -16470 20510
rect -16470 20490 -16450 20510
rect -16450 20490 -16445 20510
rect -16475 20485 -16445 20490
rect -16395 20510 -16365 20515
rect -16395 20490 -16390 20510
rect -16390 20490 -16370 20510
rect -16370 20490 -16365 20510
rect -16395 20485 -16365 20490
rect -16315 20510 -16285 20515
rect -16315 20490 -16310 20510
rect -16310 20490 -16290 20510
rect -16290 20490 -16285 20510
rect -16315 20485 -16285 20490
rect -16235 20510 -16205 20515
rect -16235 20490 -16230 20510
rect -16230 20490 -16210 20510
rect -16210 20490 -16205 20510
rect -16235 20485 -16205 20490
rect -16155 20510 -16125 20515
rect -16155 20490 -16150 20510
rect -16150 20490 -16130 20510
rect -16130 20490 -16125 20510
rect -16155 20485 -16125 20490
rect -16075 20510 -16045 20515
rect -16075 20490 -16070 20510
rect -16070 20490 -16050 20510
rect -16050 20490 -16045 20510
rect -16075 20485 -16045 20490
rect -15995 20510 -15965 20515
rect -15995 20490 -15990 20510
rect -15990 20490 -15970 20510
rect -15970 20490 -15965 20510
rect -15995 20485 -15965 20490
rect -15915 20510 -15885 20515
rect -15915 20490 -15910 20510
rect -15910 20490 -15890 20510
rect -15890 20490 -15885 20510
rect -15915 20485 -15885 20490
rect -15835 20510 -15805 20515
rect -15835 20490 -15830 20510
rect -15830 20490 -15810 20510
rect -15810 20490 -15805 20510
rect -15835 20485 -15805 20490
rect -15755 20510 -15725 20515
rect -15755 20490 -15750 20510
rect -15750 20490 -15730 20510
rect -15730 20490 -15725 20510
rect -15755 20485 -15725 20490
rect -15675 20510 -15645 20515
rect -15675 20490 -15670 20510
rect -15670 20490 -15650 20510
rect -15650 20490 -15645 20510
rect -15675 20485 -15645 20490
rect -15595 20510 -15565 20515
rect -15595 20490 -15590 20510
rect -15590 20490 -15570 20510
rect -15570 20490 -15565 20510
rect -15595 20485 -15565 20490
rect -14955 20510 -14925 20515
rect -14955 20490 -14950 20510
rect -14950 20490 -14930 20510
rect -14930 20490 -14925 20510
rect -14955 20485 -14925 20490
rect -14875 20510 -14845 20515
rect -14875 20490 -14870 20510
rect -14870 20490 -14850 20510
rect -14850 20490 -14845 20510
rect -14875 20485 -14845 20490
rect -14795 20510 -14765 20515
rect -14795 20490 -14790 20510
rect -14790 20490 -14770 20510
rect -14770 20490 -14765 20510
rect -14795 20485 -14765 20490
rect -14715 20510 -14685 20515
rect -14715 20490 -14710 20510
rect -14710 20490 -14690 20510
rect -14690 20490 -14685 20510
rect -14715 20485 -14685 20490
rect -14635 20510 -14605 20515
rect -14635 20490 -14630 20510
rect -14630 20490 -14610 20510
rect -14610 20490 -14605 20510
rect -14635 20485 -14605 20490
rect -14555 20510 -14525 20515
rect -14555 20490 -14550 20510
rect -14550 20490 -14530 20510
rect -14530 20490 -14525 20510
rect -14555 20485 -14525 20490
rect -14475 20510 -14445 20515
rect -14475 20490 -14470 20510
rect -14470 20490 -14450 20510
rect -14450 20490 -14445 20510
rect -14475 20485 -14445 20490
rect -14395 20510 -14365 20515
rect -14395 20490 -14390 20510
rect -14390 20490 -14370 20510
rect -14370 20490 -14365 20510
rect -14395 20485 -14365 20490
rect -14315 20510 -14285 20515
rect -14315 20490 -14310 20510
rect -14310 20490 -14290 20510
rect -14290 20490 -14285 20510
rect -14315 20485 -14285 20490
rect -14235 20510 -14205 20515
rect -14235 20490 -14230 20510
rect -14230 20490 -14210 20510
rect -14210 20490 -14205 20510
rect -14235 20485 -14205 20490
rect -14155 20510 -14125 20515
rect -14155 20490 -14150 20510
rect -14150 20490 -14130 20510
rect -14130 20490 -14125 20510
rect -14155 20485 -14125 20490
rect -14075 20510 -14045 20515
rect -14075 20490 -14070 20510
rect -14070 20490 -14050 20510
rect -14050 20490 -14045 20510
rect -14075 20485 -14045 20490
rect -13995 20510 -13965 20515
rect -13995 20490 -13990 20510
rect -13990 20490 -13970 20510
rect -13970 20490 -13965 20510
rect -13995 20485 -13965 20490
rect -13915 20510 -13885 20515
rect -13915 20490 -13910 20510
rect -13910 20490 -13890 20510
rect -13890 20490 -13885 20510
rect -13915 20485 -13885 20490
rect -13835 20510 -13805 20515
rect -13835 20490 -13830 20510
rect -13830 20490 -13810 20510
rect -13810 20490 -13805 20510
rect -13835 20485 -13805 20490
rect -13755 20510 -13725 20515
rect -13755 20490 -13750 20510
rect -13750 20490 -13730 20510
rect -13730 20490 -13725 20510
rect -13755 20485 -13725 20490
rect -13675 20510 -13645 20515
rect -13675 20490 -13670 20510
rect -13670 20490 -13650 20510
rect -13650 20490 -13645 20510
rect -13675 20485 -13645 20490
rect -13595 20510 -13565 20515
rect -13595 20490 -13590 20510
rect -13590 20490 -13570 20510
rect -13570 20490 -13565 20510
rect -13595 20485 -13565 20490
rect -13515 20510 -13485 20515
rect -13515 20490 -13510 20510
rect -13510 20490 -13490 20510
rect -13490 20490 -13485 20510
rect -13515 20485 -13485 20490
rect -13435 20510 -13405 20515
rect -13435 20490 -13430 20510
rect -13430 20490 -13410 20510
rect -13410 20490 -13405 20510
rect -13435 20485 -13405 20490
rect -13355 20510 -13325 20515
rect -13355 20490 -13350 20510
rect -13350 20490 -13330 20510
rect -13330 20490 -13325 20510
rect -13355 20485 -13325 20490
rect -13275 20510 -13245 20515
rect -13275 20490 -13270 20510
rect -13270 20490 -13250 20510
rect -13250 20490 -13245 20510
rect -13275 20485 -13245 20490
rect -13195 20510 -13165 20515
rect -13195 20490 -13190 20510
rect -13190 20490 -13170 20510
rect -13170 20490 -13165 20510
rect -13195 20485 -13165 20490
rect -13115 20510 -13085 20515
rect -13115 20490 -13110 20510
rect -13110 20490 -13090 20510
rect -13090 20490 -13085 20510
rect -13115 20485 -13085 20490
rect -13035 20510 -13005 20515
rect -13035 20490 -13030 20510
rect -13030 20490 -13010 20510
rect -13010 20490 -13005 20510
rect -13035 20485 -13005 20490
rect -12955 20510 -12925 20515
rect -12955 20490 -12950 20510
rect -12950 20490 -12930 20510
rect -12930 20490 -12925 20510
rect -12955 20485 -12925 20490
rect -12875 20510 -12845 20515
rect -12875 20490 -12870 20510
rect -12870 20490 -12850 20510
rect -12850 20490 -12845 20510
rect -12875 20485 -12845 20490
rect -12795 20510 -12765 20515
rect -12795 20490 -12790 20510
rect -12790 20490 -12770 20510
rect -12770 20490 -12765 20510
rect -12795 20485 -12765 20490
rect -12715 20510 -12685 20515
rect -12715 20490 -12710 20510
rect -12710 20490 -12690 20510
rect -12690 20490 -12685 20510
rect -12715 20485 -12685 20490
rect -12635 20510 -12605 20515
rect -12635 20490 -12630 20510
rect -12630 20490 -12610 20510
rect -12610 20490 -12605 20510
rect -12635 20485 -12605 20490
rect -12555 20510 -12525 20515
rect -12555 20490 -12550 20510
rect -12550 20490 -12530 20510
rect -12530 20490 -12525 20510
rect -12555 20485 -12525 20490
rect -12475 20510 -12445 20515
rect -12475 20490 -12470 20510
rect -12470 20490 -12450 20510
rect -12450 20490 -12445 20510
rect -12475 20485 -12445 20490
rect -12395 20510 -12365 20515
rect -12395 20490 -12390 20510
rect -12390 20490 -12370 20510
rect -12370 20490 -12365 20510
rect -12395 20485 -12365 20490
rect -12315 20510 -12285 20515
rect -12315 20490 -12310 20510
rect -12310 20490 -12290 20510
rect -12290 20490 -12285 20510
rect -12315 20485 -12285 20490
rect -12235 20510 -12205 20515
rect -12235 20490 -12230 20510
rect -12230 20490 -12210 20510
rect -12210 20490 -12205 20510
rect -12235 20485 -12205 20490
rect -12155 20510 -12125 20515
rect -12155 20490 -12150 20510
rect -12150 20490 -12130 20510
rect -12130 20490 -12125 20510
rect -12155 20485 -12125 20490
rect -12075 20510 -12045 20515
rect -12075 20490 -12070 20510
rect -12070 20490 -12050 20510
rect -12050 20490 -12045 20510
rect -12075 20485 -12045 20490
rect -11995 20510 -11965 20515
rect -11995 20490 -11990 20510
rect -11990 20490 -11970 20510
rect -11970 20490 -11965 20510
rect -11995 20485 -11965 20490
rect -11915 20510 -11885 20515
rect -11915 20490 -11910 20510
rect -11910 20490 -11890 20510
rect -11890 20490 -11885 20510
rect -11915 20485 -11885 20490
rect -11835 20510 -11805 20515
rect -11835 20490 -11830 20510
rect -11830 20490 -11810 20510
rect -11810 20490 -11805 20510
rect -11835 20485 -11805 20490
rect -11755 20510 -11725 20515
rect -11755 20490 -11750 20510
rect -11750 20490 -11730 20510
rect -11730 20490 -11725 20510
rect -11755 20485 -11725 20490
rect -11675 20510 -11645 20515
rect -11675 20490 -11670 20510
rect -11670 20490 -11650 20510
rect -11650 20490 -11645 20510
rect -11675 20485 -11645 20490
rect -11595 20510 -11565 20515
rect -11595 20490 -11590 20510
rect -11590 20490 -11570 20510
rect -11570 20490 -11565 20510
rect -11595 20485 -11565 20490
rect -11515 20510 -11485 20515
rect -11515 20490 -11510 20510
rect -11510 20490 -11490 20510
rect -11490 20490 -11485 20510
rect -11515 20485 -11485 20490
rect -11435 20510 -11405 20515
rect -11435 20490 -11430 20510
rect -11430 20490 -11410 20510
rect -11410 20490 -11405 20510
rect -11435 20485 -11405 20490
rect -11355 20510 -11325 20515
rect -11355 20490 -11350 20510
rect -11350 20490 -11330 20510
rect -11330 20490 -11325 20510
rect -11355 20485 -11325 20490
rect -11275 20510 -11245 20515
rect -11275 20490 -11270 20510
rect -11270 20490 -11250 20510
rect -11250 20490 -11245 20510
rect -11275 20485 -11245 20490
rect -11195 20510 -11165 20515
rect -11195 20490 -11190 20510
rect -11190 20490 -11170 20510
rect -11170 20490 -11165 20510
rect -11195 20485 -11165 20490
rect -11115 20510 -11085 20515
rect -11115 20490 -11110 20510
rect -11110 20490 -11090 20510
rect -11090 20490 -11085 20510
rect -11115 20485 -11085 20490
rect -11035 20510 -11005 20515
rect -11035 20490 -11030 20510
rect -11030 20490 -11010 20510
rect -11010 20490 -11005 20510
rect -11035 20485 -11005 20490
rect -10955 20510 -10925 20515
rect -10955 20490 -10950 20510
rect -10950 20490 -10930 20510
rect -10930 20490 -10925 20510
rect -10955 20485 -10925 20490
rect -10875 20510 -10845 20515
rect -10875 20490 -10870 20510
rect -10870 20490 -10850 20510
rect -10850 20490 -10845 20510
rect -10875 20485 -10845 20490
rect -10795 20510 -10765 20515
rect -10795 20490 -10790 20510
rect -10790 20490 -10770 20510
rect -10770 20490 -10765 20510
rect -10795 20485 -10765 20490
rect -10715 20510 -10685 20515
rect -10715 20490 -10710 20510
rect -10710 20490 -10690 20510
rect -10690 20490 -10685 20510
rect -10715 20485 -10685 20490
rect -10635 20510 -10605 20515
rect -10635 20490 -10630 20510
rect -10630 20490 -10610 20510
rect -10610 20490 -10605 20510
rect -10635 20485 -10605 20490
rect -10555 20510 -10525 20515
rect -10555 20490 -10550 20510
rect -10550 20490 -10530 20510
rect -10530 20490 -10525 20510
rect -10555 20485 -10525 20490
rect -10475 20510 -10445 20515
rect -10475 20490 -10470 20510
rect -10470 20490 -10450 20510
rect -10450 20490 -10445 20510
rect -10475 20485 -10445 20490
rect -10395 20510 -10365 20515
rect -10395 20490 -10390 20510
rect -10390 20490 -10370 20510
rect -10370 20490 -10365 20510
rect -10395 20485 -10365 20490
rect -10315 20510 -10285 20515
rect -10315 20490 -10310 20510
rect -10310 20490 -10290 20510
rect -10290 20490 -10285 20510
rect -10315 20485 -10285 20490
rect -10235 20510 -10205 20515
rect -10235 20490 -10230 20510
rect -10230 20490 -10210 20510
rect -10210 20490 -10205 20510
rect -10235 20485 -10205 20490
rect -10155 20510 -10125 20515
rect -10155 20490 -10150 20510
rect -10150 20490 -10130 20510
rect -10130 20490 -10125 20510
rect -10155 20485 -10125 20490
rect -10075 20510 -10045 20515
rect -10075 20490 -10070 20510
rect -10070 20490 -10050 20510
rect -10050 20490 -10045 20510
rect -10075 20485 -10045 20490
rect -9995 20510 -9965 20515
rect -9995 20490 -9990 20510
rect -9990 20490 -9970 20510
rect -9970 20490 -9965 20510
rect -9995 20485 -9965 20490
rect -9915 20510 -9885 20515
rect -9915 20490 -9910 20510
rect -9910 20490 -9890 20510
rect -9890 20490 -9885 20510
rect -9915 20485 -9885 20490
rect -9835 20510 -9805 20515
rect -9835 20490 -9830 20510
rect -9830 20490 -9810 20510
rect -9810 20490 -9805 20510
rect -9835 20485 -9805 20490
rect -9755 20510 -9725 20515
rect -9755 20490 -9750 20510
rect -9750 20490 -9730 20510
rect -9730 20490 -9725 20510
rect -9755 20485 -9725 20490
rect -9675 20510 -9645 20515
rect -9675 20490 -9670 20510
rect -9670 20490 -9650 20510
rect -9650 20490 -9645 20510
rect -9675 20485 -9645 20490
rect -9595 20510 -9565 20515
rect -9595 20490 -9590 20510
rect -9590 20490 -9570 20510
rect -9570 20490 -9565 20510
rect -9595 20485 -9565 20490
rect -9515 20510 -9485 20515
rect -9515 20490 -9510 20510
rect -9510 20490 -9490 20510
rect -9490 20490 -9485 20510
rect -9515 20485 -9485 20490
rect -9435 20510 -9405 20515
rect -9435 20490 -9430 20510
rect -9430 20490 -9410 20510
rect -9410 20490 -9405 20510
rect -9435 20485 -9405 20490
rect -9355 20510 -9325 20515
rect -9355 20490 -9350 20510
rect -9350 20490 -9330 20510
rect -9330 20490 -9325 20510
rect -9355 20485 -9325 20490
rect -9275 20510 -9245 20515
rect -9275 20490 -9270 20510
rect -9270 20490 -9250 20510
rect -9250 20490 -9245 20510
rect -9275 20485 -9245 20490
rect -9195 20510 -9165 20515
rect -9195 20490 -9190 20510
rect -9190 20490 -9170 20510
rect -9170 20490 -9165 20510
rect -9195 20485 -9165 20490
rect -9115 20510 -9085 20515
rect -9115 20490 -9110 20510
rect -9110 20490 -9090 20510
rect -9090 20490 -9085 20510
rect -9115 20485 -9085 20490
rect -9035 20510 -9005 20515
rect -9035 20490 -9030 20510
rect -9030 20490 -9010 20510
rect -9010 20490 -9005 20510
rect -9035 20485 -9005 20490
rect -8955 20510 -8925 20515
rect -8955 20490 -8950 20510
rect -8950 20490 -8930 20510
rect -8930 20490 -8925 20510
rect -8955 20485 -8925 20490
rect -8875 20510 -8845 20515
rect -8875 20490 -8870 20510
rect -8870 20490 -8850 20510
rect -8850 20490 -8845 20510
rect -8875 20485 -8845 20490
rect -8795 20510 -8765 20515
rect -8795 20490 -8790 20510
rect -8790 20490 -8770 20510
rect -8770 20490 -8765 20510
rect -8795 20485 -8765 20490
rect -8715 20510 -8685 20515
rect -8715 20490 -8710 20510
rect -8710 20490 -8690 20510
rect -8690 20490 -8685 20510
rect -8715 20485 -8685 20490
rect -8635 20510 -8605 20515
rect -8635 20490 -8630 20510
rect -8630 20490 -8610 20510
rect -8610 20490 -8605 20510
rect -8635 20485 -8605 20490
rect -8555 20510 -8525 20515
rect -8555 20490 -8550 20510
rect -8550 20490 -8530 20510
rect -8530 20490 -8525 20510
rect -8555 20485 -8525 20490
rect -8475 20510 -8445 20515
rect -8475 20490 -8470 20510
rect -8470 20490 -8450 20510
rect -8450 20490 -8445 20510
rect -8475 20485 -8445 20490
rect -8395 20510 -8365 20515
rect -8395 20490 -8390 20510
rect -8390 20490 -8370 20510
rect -8370 20490 -8365 20510
rect -8395 20485 -8365 20490
rect -8315 20510 -8285 20515
rect -8315 20490 -8310 20510
rect -8310 20490 -8290 20510
rect -8290 20490 -8285 20510
rect -8315 20485 -8285 20490
rect -8235 20510 -8205 20515
rect -8235 20490 -8230 20510
rect -8230 20490 -8210 20510
rect -8210 20490 -8205 20510
rect -8235 20485 -8205 20490
rect -8155 20510 -8125 20515
rect -8155 20490 -8150 20510
rect -8150 20490 -8130 20510
rect -8130 20490 -8125 20510
rect -8155 20485 -8125 20490
rect -8075 20510 -8045 20515
rect -8075 20490 -8070 20510
rect -8070 20490 -8050 20510
rect -8050 20490 -8045 20510
rect -8075 20485 -8045 20490
rect -7995 20510 -7965 20515
rect -7995 20490 -7990 20510
rect -7990 20490 -7970 20510
rect -7970 20490 -7965 20510
rect -7995 20485 -7965 20490
rect -7915 20510 -7885 20515
rect -7915 20490 -7910 20510
rect -7910 20490 -7890 20510
rect -7890 20490 -7885 20510
rect -7915 20485 -7885 20490
rect -7835 20510 -7805 20515
rect -7835 20490 -7830 20510
rect -7830 20490 -7810 20510
rect -7810 20490 -7805 20510
rect -7835 20485 -7805 20490
rect -7755 20510 -7725 20515
rect -7755 20490 -7750 20510
rect -7750 20490 -7730 20510
rect -7730 20490 -7725 20510
rect -7755 20485 -7725 20490
rect -7675 20510 -7645 20515
rect -7675 20490 -7670 20510
rect -7670 20490 -7650 20510
rect -7650 20490 -7645 20510
rect -7675 20485 -7645 20490
rect -7595 20510 -7565 20515
rect -7595 20490 -7590 20510
rect -7590 20490 -7570 20510
rect -7570 20490 -7565 20510
rect -7595 20485 -7565 20490
rect -7515 20510 -7485 20515
rect -7515 20490 -7510 20510
rect -7510 20490 -7490 20510
rect -7490 20490 -7485 20510
rect -7515 20485 -7485 20490
rect -7435 20510 -7405 20515
rect -7435 20490 -7430 20510
rect -7430 20490 -7410 20510
rect -7410 20490 -7405 20510
rect -7435 20485 -7405 20490
rect -7355 20510 -7325 20515
rect -7355 20490 -7350 20510
rect -7350 20490 -7330 20510
rect -7330 20490 -7325 20510
rect -7355 20485 -7325 20490
rect -7275 20510 -7245 20515
rect -7275 20490 -7270 20510
rect -7270 20490 -7250 20510
rect -7250 20490 -7245 20510
rect -7275 20485 -7245 20490
rect -7195 20510 -7165 20515
rect -7195 20490 -7190 20510
rect -7190 20490 -7170 20510
rect -7170 20490 -7165 20510
rect -7195 20485 -7165 20490
rect -7115 20510 -7085 20515
rect -7115 20490 -7110 20510
rect -7110 20490 -7090 20510
rect -7090 20490 -7085 20510
rect -7115 20485 -7085 20490
rect -7035 20510 -7005 20515
rect -7035 20490 -7030 20510
rect -7030 20490 -7010 20510
rect -7010 20490 -7005 20510
rect -7035 20485 -7005 20490
rect -6955 20510 -6925 20515
rect -6955 20490 -6950 20510
rect -6950 20490 -6930 20510
rect -6930 20490 -6925 20510
rect -6955 20485 -6925 20490
rect -6875 20510 -6845 20515
rect -6875 20490 -6870 20510
rect -6870 20490 -6850 20510
rect -6850 20490 -6845 20510
rect -6875 20485 -6845 20490
rect -6795 20510 -6765 20515
rect -6795 20490 -6790 20510
rect -6790 20490 -6770 20510
rect -6770 20490 -6765 20510
rect -6795 20485 -6765 20490
rect -6715 20510 -6685 20515
rect -6715 20490 -6710 20510
rect -6710 20490 -6690 20510
rect -6690 20490 -6685 20510
rect -6715 20485 -6685 20490
rect -6635 20510 -6605 20515
rect -6635 20490 -6630 20510
rect -6630 20490 -6610 20510
rect -6610 20490 -6605 20510
rect -6635 20485 -6605 20490
rect -6555 20510 -6525 20515
rect -6555 20490 -6550 20510
rect -6550 20490 -6530 20510
rect -6530 20490 -6525 20510
rect -6555 20485 -6525 20490
rect -6475 20510 -6445 20515
rect -6475 20490 -6470 20510
rect -6470 20490 -6450 20510
rect -6450 20490 -6445 20510
rect -6475 20485 -6445 20490
rect -6395 20510 -6365 20515
rect -6395 20490 -6390 20510
rect -6390 20490 -6370 20510
rect -6370 20490 -6365 20510
rect -6395 20485 -6365 20490
rect -6315 20510 -6285 20515
rect -6315 20490 -6310 20510
rect -6310 20490 -6290 20510
rect -6290 20490 -6285 20510
rect -6315 20485 -6285 20490
rect -6235 20510 -6205 20515
rect -6235 20490 -6230 20510
rect -6230 20490 -6210 20510
rect -6210 20490 -6205 20510
rect -6235 20485 -6205 20490
rect -6155 20510 -6125 20515
rect -6155 20490 -6150 20510
rect -6150 20490 -6130 20510
rect -6130 20490 -6125 20510
rect -6155 20485 -6125 20490
rect -5675 20510 -5645 20515
rect -5675 20490 -5670 20510
rect -5670 20490 -5650 20510
rect -5650 20490 -5645 20510
rect -5675 20485 -5645 20490
rect -5595 20510 -5565 20515
rect -5595 20490 -5590 20510
rect -5590 20490 -5570 20510
rect -5570 20490 -5565 20510
rect -5595 20485 -5565 20490
rect -5515 20510 -5485 20515
rect -5515 20490 -5510 20510
rect -5510 20490 -5490 20510
rect -5490 20490 -5485 20510
rect -5515 20485 -5485 20490
rect -5435 20510 -5405 20515
rect -5435 20490 -5430 20510
rect -5430 20490 -5410 20510
rect -5410 20490 -5405 20510
rect -5435 20485 -5405 20490
rect -5355 20510 -5325 20515
rect -5355 20490 -5350 20510
rect -5350 20490 -5330 20510
rect -5330 20490 -5325 20510
rect -5355 20485 -5325 20490
rect -5275 20510 -5245 20515
rect -5275 20490 -5270 20510
rect -5270 20490 -5250 20510
rect -5250 20490 -5245 20510
rect -5275 20485 -5245 20490
rect -5195 20510 -5165 20515
rect -5195 20490 -5190 20510
rect -5190 20490 -5170 20510
rect -5170 20490 -5165 20510
rect -5195 20485 -5165 20490
rect -5115 20510 -5085 20515
rect -5115 20490 -5110 20510
rect -5110 20490 -5090 20510
rect -5090 20490 -5085 20510
rect -5115 20485 -5085 20490
rect -5035 20510 -5005 20515
rect -5035 20490 -5030 20510
rect -5030 20490 -5010 20510
rect -5010 20490 -5005 20510
rect -5035 20485 -5005 20490
rect -4955 20510 -4925 20515
rect -4955 20490 -4950 20510
rect -4950 20490 -4930 20510
rect -4930 20490 -4925 20510
rect -4955 20485 -4925 20490
rect -4875 20510 -4845 20515
rect -4875 20490 -4870 20510
rect -4870 20490 -4850 20510
rect -4850 20490 -4845 20510
rect -4875 20485 -4845 20490
rect -4795 20510 -4765 20515
rect -4795 20490 -4790 20510
rect -4790 20490 -4770 20510
rect -4770 20490 -4765 20510
rect -4795 20485 -4765 20490
rect -4715 20510 -4685 20515
rect -4715 20490 -4710 20510
rect -4710 20490 -4690 20510
rect -4690 20490 -4685 20510
rect -4715 20485 -4685 20490
rect -4635 20510 -4605 20515
rect -4635 20490 -4630 20510
rect -4630 20490 -4610 20510
rect -4610 20490 -4605 20510
rect -4635 20485 -4605 20490
rect -4555 20510 -4525 20515
rect -4555 20490 -4550 20510
rect -4550 20490 -4530 20510
rect -4530 20490 -4525 20510
rect -4555 20485 -4525 20490
rect -4475 20510 -4445 20515
rect -4475 20490 -4470 20510
rect -4470 20490 -4450 20510
rect -4450 20490 -4445 20510
rect -4475 20485 -4445 20490
rect -4395 20510 -4365 20515
rect -4395 20490 -4390 20510
rect -4390 20490 -4370 20510
rect -4370 20490 -4365 20510
rect -4395 20485 -4365 20490
rect -4315 20510 -4285 20515
rect -4315 20490 -4310 20510
rect -4310 20490 -4290 20510
rect -4290 20490 -4285 20510
rect -4315 20485 -4285 20490
rect -4235 20510 -4205 20515
rect -4235 20490 -4230 20510
rect -4230 20490 -4210 20510
rect -4210 20490 -4205 20510
rect -4235 20485 -4205 20490
rect -4155 20510 -4125 20515
rect -4155 20490 -4150 20510
rect -4150 20490 -4130 20510
rect -4130 20490 -4125 20510
rect -4155 20485 -4125 20490
rect -4075 20510 -4045 20515
rect -4075 20490 -4070 20510
rect -4070 20490 -4050 20510
rect -4050 20490 -4045 20510
rect -4075 20485 -4045 20490
rect -3995 20510 -3965 20515
rect -3995 20490 -3990 20510
rect -3990 20490 -3970 20510
rect -3970 20490 -3965 20510
rect -3995 20485 -3965 20490
rect -3915 20510 -3885 20515
rect -3915 20490 -3910 20510
rect -3910 20490 -3890 20510
rect -3890 20490 -3885 20510
rect -3915 20485 -3885 20490
rect -3835 20510 -3805 20515
rect -3835 20490 -3830 20510
rect -3830 20490 -3810 20510
rect -3810 20490 -3805 20510
rect -3835 20485 -3805 20490
rect -3755 20510 -3725 20515
rect -3755 20490 -3750 20510
rect -3750 20490 -3730 20510
rect -3730 20490 -3725 20510
rect -3755 20485 -3725 20490
rect -3675 20510 -3645 20515
rect -3675 20490 -3670 20510
rect -3670 20490 -3650 20510
rect -3650 20490 -3645 20510
rect -3675 20485 -3645 20490
rect -3595 20510 -3565 20515
rect -3595 20490 -3590 20510
rect -3590 20490 -3570 20510
rect -3570 20490 -3565 20510
rect -3595 20485 -3565 20490
rect -3515 20510 -3485 20515
rect -3515 20490 -3510 20510
rect -3510 20490 -3490 20510
rect -3490 20490 -3485 20510
rect -3515 20485 -3485 20490
rect -3435 20510 -3405 20515
rect -3435 20490 -3430 20510
rect -3430 20490 -3410 20510
rect -3410 20490 -3405 20510
rect -3435 20485 -3405 20490
rect -3355 20510 -3325 20515
rect -3355 20490 -3350 20510
rect -3350 20490 -3330 20510
rect -3330 20490 -3325 20510
rect -3355 20485 -3325 20490
rect -3275 20510 -3245 20515
rect -3275 20490 -3270 20510
rect -3270 20490 -3250 20510
rect -3250 20490 -3245 20510
rect -3275 20485 -3245 20490
rect -3195 20510 -3165 20515
rect -3195 20490 -3190 20510
rect -3190 20490 -3170 20510
rect -3170 20490 -3165 20510
rect -3195 20485 -3165 20490
rect -3115 20510 -3085 20515
rect -3115 20490 -3110 20510
rect -3110 20490 -3090 20510
rect -3090 20490 -3085 20510
rect -3115 20485 -3085 20490
rect -3035 20510 -3005 20515
rect -3035 20490 -3030 20510
rect -3030 20490 -3010 20510
rect -3010 20490 -3005 20510
rect -3035 20485 -3005 20490
rect -2955 20510 -2925 20515
rect -2955 20490 -2950 20510
rect -2950 20490 -2930 20510
rect -2930 20490 -2925 20510
rect -2955 20485 -2925 20490
rect -2875 20510 -2845 20515
rect -2875 20490 -2870 20510
rect -2870 20490 -2850 20510
rect -2850 20490 -2845 20510
rect -2875 20485 -2845 20490
rect -2795 20510 -2765 20515
rect -2795 20490 -2790 20510
rect -2790 20490 -2770 20510
rect -2770 20490 -2765 20510
rect -2795 20485 -2765 20490
rect -2715 20510 -2685 20515
rect -2715 20490 -2710 20510
rect -2710 20490 -2690 20510
rect -2690 20490 -2685 20510
rect -2715 20485 -2685 20490
rect -2635 20510 -2605 20515
rect -2635 20490 -2630 20510
rect -2630 20490 -2610 20510
rect -2610 20490 -2605 20510
rect -2635 20485 -2605 20490
rect -2555 20510 -2525 20515
rect -2555 20490 -2550 20510
rect -2550 20490 -2530 20510
rect -2530 20490 -2525 20510
rect -2555 20485 -2525 20490
rect -2475 20510 -2445 20515
rect -2475 20490 -2470 20510
rect -2470 20490 -2450 20510
rect -2450 20490 -2445 20510
rect -2475 20485 -2445 20490
rect -2395 20510 -2365 20515
rect -2395 20490 -2390 20510
rect -2390 20490 -2370 20510
rect -2370 20490 -2365 20510
rect -2395 20485 -2365 20490
rect -2315 20510 -2285 20515
rect -2315 20490 -2310 20510
rect -2310 20490 -2290 20510
rect -2290 20490 -2285 20510
rect -2315 20485 -2285 20490
rect -2235 20510 -2205 20515
rect -2235 20490 -2230 20510
rect -2230 20490 -2210 20510
rect -2210 20490 -2205 20510
rect -2235 20485 -2205 20490
rect -2155 20510 -2125 20515
rect -2155 20490 -2150 20510
rect -2150 20490 -2130 20510
rect -2130 20490 -2125 20510
rect -2155 20485 -2125 20490
rect -2075 20510 -2045 20515
rect -2075 20490 -2070 20510
rect -2070 20490 -2050 20510
rect -2050 20490 -2045 20510
rect -2075 20485 -2045 20490
rect -1995 20510 -1965 20515
rect -1995 20490 -1990 20510
rect -1990 20490 -1970 20510
rect -1970 20490 -1965 20510
rect -1995 20485 -1965 20490
rect -1835 20510 -1805 20515
rect -1835 20490 -1830 20510
rect -1830 20490 -1810 20510
rect -1810 20490 -1805 20510
rect -1835 20485 -1805 20490
rect -1755 20510 -1725 20515
rect -1755 20490 -1750 20510
rect -1750 20490 -1730 20510
rect -1730 20490 -1725 20510
rect -1755 20485 -1725 20490
rect 20525 20510 20555 20515
rect 20525 20490 20530 20510
rect 20530 20490 20550 20510
rect 20550 20490 20555 20510
rect 20525 20485 20555 20490
rect 20605 20510 20635 20515
rect 20605 20490 20610 20510
rect 20610 20490 20630 20510
rect 20630 20490 20635 20510
rect 20605 20485 20635 20490
rect 20685 20510 20715 20515
rect 20685 20490 20690 20510
rect 20690 20490 20710 20510
rect 20710 20490 20715 20510
rect 20685 20485 20715 20490
rect 20765 20510 20795 20515
rect 20765 20490 20770 20510
rect 20770 20490 20790 20510
rect 20790 20490 20795 20510
rect 20765 20485 20795 20490
rect 20845 20510 20875 20515
rect 20845 20490 20850 20510
rect 20850 20490 20870 20510
rect 20870 20490 20875 20510
rect 20845 20485 20875 20490
rect 20925 20510 20955 20515
rect 20925 20490 20930 20510
rect 20930 20490 20950 20510
rect 20950 20490 20955 20510
rect 20925 20485 20955 20490
rect 21005 20510 21035 20515
rect 21005 20490 21010 20510
rect 21010 20490 21030 20510
rect 21030 20490 21035 20510
rect 21005 20485 21035 20490
rect 21085 20510 21115 20515
rect 21085 20490 21090 20510
rect 21090 20490 21110 20510
rect 21110 20490 21115 20510
rect 21085 20485 21115 20490
rect 21165 20510 21195 20515
rect 21165 20490 21170 20510
rect 21170 20490 21190 20510
rect 21190 20490 21195 20510
rect 21165 20485 21195 20490
rect 21245 20510 21275 20515
rect 21245 20490 21250 20510
rect 21250 20490 21270 20510
rect 21270 20490 21275 20510
rect 21245 20485 21275 20490
rect 21325 20510 21355 20515
rect 21325 20490 21330 20510
rect 21330 20490 21350 20510
rect 21350 20490 21355 20510
rect 21325 20485 21355 20490
rect 21405 20510 21435 20515
rect 21405 20490 21410 20510
rect 21410 20490 21430 20510
rect 21430 20490 21435 20510
rect 21405 20485 21435 20490
rect 21485 20510 21515 20515
rect 21485 20490 21490 20510
rect 21490 20490 21510 20510
rect 21510 20490 21515 20510
rect 21485 20485 21515 20490
rect 21565 20510 21595 20515
rect 21565 20490 21570 20510
rect 21570 20490 21590 20510
rect 21590 20490 21595 20510
rect 21565 20485 21595 20490
rect -5275 20350 -5245 20355
rect -5275 20330 -5270 20350
rect -5270 20330 -5250 20350
rect -5250 20330 -5245 20350
rect -5275 20325 -5245 20330
rect -5115 20350 -5085 20355
rect -5115 20330 -5110 20350
rect -5110 20330 -5090 20350
rect -5090 20330 -5085 20350
rect -5115 20325 -5085 20330
rect -5035 20350 -5005 20355
rect -5035 20330 -5030 20350
rect -5030 20330 -5010 20350
rect -5010 20330 -5005 20350
rect -5035 20325 -5005 20330
rect -4955 20350 -4925 20355
rect -4955 20330 -4950 20350
rect -4950 20330 -4930 20350
rect -4930 20330 -4925 20350
rect -4955 20325 -4925 20330
rect -4875 20350 -4845 20355
rect -4875 20330 -4870 20350
rect -4870 20330 -4850 20350
rect -4850 20330 -4845 20350
rect -4875 20325 -4845 20330
rect -4795 20350 -4765 20355
rect -4795 20330 -4790 20350
rect -4790 20330 -4770 20350
rect -4770 20330 -4765 20350
rect -4795 20325 -4765 20330
rect -4715 20350 -4685 20355
rect -4715 20330 -4710 20350
rect -4710 20330 -4690 20350
rect -4690 20330 -4685 20350
rect -4715 20325 -4685 20330
rect -4635 20350 -4605 20355
rect -4635 20330 -4630 20350
rect -4630 20330 -4610 20350
rect -4610 20330 -4605 20350
rect -4635 20325 -4605 20330
rect -4555 20350 -4525 20355
rect -4555 20330 -4550 20350
rect -4550 20330 -4530 20350
rect -4530 20330 -4525 20350
rect -4555 20325 -4525 20330
rect -4475 20350 -4445 20355
rect -4475 20330 -4470 20350
rect -4470 20330 -4450 20350
rect -4450 20330 -4445 20350
rect -4475 20325 -4445 20330
rect -4395 20350 -4365 20355
rect -4395 20330 -4390 20350
rect -4390 20330 -4370 20350
rect -4370 20330 -4365 20350
rect -4395 20325 -4365 20330
rect -4315 20350 -4285 20355
rect -4315 20330 -4310 20350
rect -4310 20330 -4290 20350
rect -4290 20330 -4285 20350
rect -4315 20325 -4285 20330
rect -4235 20350 -4205 20355
rect -4235 20330 -4230 20350
rect -4230 20330 -4210 20350
rect -4210 20330 -4205 20350
rect -4235 20325 -4205 20330
rect -4155 20350 -4125 20355
rect -4155 20330 -4150 20350
rect -4150 20330 -4130 20350
rect -4130 20330 -4125 20350
rect -4155 20325 -4125 20330
rect -4075 20350 -4045 20355
rect -4075 20330 -4070 20350
rect -4070 20330 -4050 20350
rect -4050 20330 -4045 20350
rect -4075 20325 -4045 20330
rect -3995 20350 -3965 20355
rect -3995 20330 -3990 20350
rect -3990 20330 -3970 20350
rect -3970 20330 -3965 20350
rect -3995 20325 -3965 20330
rect -3915 20350 -3885 20355
rect -3915 20330 -3910 20350
rect -3910 20330 -3890 20350
rect -3890 20330 -3885 20350
rect -3915 20325 -3885 20330
rect -3835 20350 -3805 20355
rect -3835 20330 -3830 20350
rect -3830 20330 -3810 20350
rect -3810 20330 -3805 20350
rect -3835 20325 -3805 20330
rect -3755 20350 -3725 20355
rect -3755 20330 -3750 20350
rect -3750 20330 -3730 20350
rect -3730 20330 -3725 20350
rect -3755 20325 -3725 20330
rect -3675 20350 -3645 20355
rect -3675 20330 -3670 20350
rect -3670 20330 -3650 20350
rect -3650 20330 -3645 20350
rect -3675 20325 -3645 20330
rect -3595 20350 -3565 20355
rect -3595 20330 -3590 20350
rect -3590 20330 -3570 20350
rect -3570 20330 -3565 20350
rect -3595 20325 -3565 20330
rect -3515 20350 -3485 20355
rect -3515 20330 -3510 20350
rect -3510 20330 -3490 20350
rect -3490 20330 -3485 20350
rect -3515 20325 -3485 20330
rect -3435 20350 -3405 20355
rect -3435 20330 -3430 20350
rect -3430 20330 -3410 20350
rect -3410 20330 -3405 20350
rect -3435 20325 -3405 20330
rect -3355 20350 -3325 20355
rect -3355 20330 -3350 20350
rect -3350 20330 -3330 20350
rect -3330 20330 -3325 20350
rect -3355 20325 -3325 20330
rect -3275 20350 -3245 20355
rect -3275 20330 -3270 20350
rect -3270 20330 -3250 20350
rect -3250 20330 -3245 20350
rect -3275 20325 -3245 20330
rect -3195 20350 -3165 20355
rect -3195 20330 -3190 20350
rect -3190 20330 -3170 20350
rect -3170 20330 -3165 20350
rect -3195 20325 -3165 20330
rect -3115 20350 -3085 20355
rect -3115 20330 -3110 20350
rect -3110 20330 -3090 20350
rect -3090 20330 -3085 20350
rect -3115 20325 -3085 20330
rect -3035 20350 -3005 20355
rect -3035 20330 -3030 20350
rect -3030 20330 -3010 20350
rect -3010 20330 -3005 20350
rect -3035 20325 -3005 20330
rect -2955 20350 -2925 20355
rect -2955 20330 -2950 20350
rect -2950 20330 -2930 20350
rect -2930 20330 -2925 20350
rect -2955 20325 -2925 20330
rect -2875 20350 -2845 20355
rect -2875 20330 -2870 20350
rect -2870 20330 -2850 20350
rect -2850 20330 -2845 20350
rect -2875 20325 -2845 20330
rect -2795 20350 -2765 20355
rect -2795 20330 -2790 20350
rect -2790 20330 -2770 20350
rect -2770 20330 -2765 20350
rect -2795 20325 -2765 20330
rect -2715 20350 -2685 20355
rect -2715 20330 -2710 20350
rect -2710 20330 -2690 20350
rect -2690 20330 -2685 20350
rect -2715 20325 -2685 20330
rect -2635 20350 -2605 20355
rect -2635 20330 -2630 20350
rect -2630 20330 -2610 20350
rect -2610 20330 -2605 20350
rect -2635 20325 -2605 20330
rect -2555 20350 -2525 20355
rect -2555 20330 -2550 20350
rect -2550 20330 -2530 20350
rect -2530 20330 -2525 20350
rect -2555 20325 -2525 20330
rect -2475 20350 -2445 20355
rect -2475 20330 -2470 20350
rect -2470 20330 -2450 20350
rect -2450 20330 -2445 20350
rect -2475 20325 -2445 20330
rect -2395 20350 -2365 20355
rect -2395 20330 -2390 20350
rect -2390 20330 -2370 20350
rect -2370 20330 -2365 20350
rect -2395 20325 -2365 20330
rect -2315 20350 -2285 20355
rect -2315 20330 -2310 20350
rect -2310 20330 -2290 20350
rect -2290 20330 -2285 20350
rect -2315 20325 -2285 20330
rect -2235 20350 -2205 20355
rect -2235 20330 -2230 20350
rect -2230 20330 -2210 20350
rect -2210 20330 -2205 20350
rect -2235 20325 -2205 20330
rect -2155 20350 -2125 20355
rect -2155 20330 -2150 20350
rect -2150 20330 -2130 20350
rect -2130 20330 -2125 20350
rect -2155 20325 -2125 20330
rect -2075 20350 -2045 20355
rect -2075 20330 -2070 20350
rect -2070 20330 -2050 20350
rect -2050 20330 -2045 20350
rect -2075 20325 -2045 20330
rect -1995 20350 -1965 20355
rect -1995 20330 -1990 20350
rect -1990 20330 -1970 20350
rect -1970 20330 -1965 20350
rect -1995 20325 -1965 20330
rect -1835 20350 -1805 20355
rect -1835 20330 -1830 20350
rect -1830 20330 -1810 20350
rect -1810 20330 -1805 20350
rect -1835 20325 -1805 20330
rect -1755 20350 -1725 20355
rect -1755 20330 -1750 20350
rect -1750 20330 -1730 20350
rect -1730 20330 -1725 20350
rect -1755 20325 -1725 20330
rect -5275 20190 -5245 20195
rect -5275 20170 -5270 20190
rect -5270 20170 -5250 20190
rect -5250 20170 -5245 20190
rect -5275 20165 -5245 20170
rect -5115 20190 -5085 20195
rect -5115 20170 -5110 20190
rect -5110 20170 -5090 20190
rect -5090 20170 -5085 20190
rect -5115 20165 -5085 20170
rect -5035 20190 -5005 20195
rect -5035 20170 -5030 20190
rect -5030 20170 -5010 20190
rect -5010 20170 -5005 20190
rect -5035 20165 -5005 20170
rect -4955 20190 -4925 20195
rect -4955 20170 -4950 20190
rect -4950 20170 -4930 20190
rect -4930 20170 -4925 20190
rect -4955 20165 -4925 20170
rect -4875 20190 -4845 20195
rect -4875 20170 -4870 20190
rect -4870 20170 -4850 20190
rect -4850 20170 -4845 20190
rect -4875 20165 -4845 20170
rect -4795 20190 -4765 20195
rect -4795 20170 -4790 20190
rect -4790 20170 -4770 20190
rect -4770 20170 -4765 20190
rect -4795 20165 -4765 20170
rect -4715 20190 -4685 20195
rect -4715 20170 -4710 20190
rect -4710 20170 -4690 20190
rect -4690 20170 -4685 20190
rect -4715 20165 -4685 20170
rect -4635 20190 -4605 20195
rect -4635 20170 -4630 20190
rect -4630 20170 -4610 20190
rect -4610 20170 -4605 20190
rect -4635 20165 -4605 20170
rect -4555 20190 -4525 20195
rect -4555 20170 -4550 20190
rect -4550 20170 -4530 20190
rect -4530 20170 -4525 20190
rect -4555 20165 -4525 20170
rect -4475 20190 -4445 20195
rect -4475 20170 -4470 20190
rect -4470 20170 -4450 20190
rect -4450 20170 -4445 20190
rect -4475 20165 -4445 20170
rect -4395 20190 -4365 20195
rect -4395 20170 -4390 20190
rect -4390 20170 -4370 20190
rect -4370 20170 -4365 20190
rect -4395 20165 -4365 20170
rect -4315 20190 -4285 20195
rect -4315 20170 -4310 20190
rect -4310 20170 -4290 20190
rect -4290 20170 -4285 20190
rect -4315 20165 -4285 20170
rect -4235 20190 -4205 20195
rect -4235 20170 -4230 20190
rect -4230 20170 -4210 20190
rect -4210 20170 -4205 20190
rect -4235 20165 -4205 20170
rect -4155 20190 -4125 20195
rect -4155 20170 -4150 20190
rect -4150 20170 -4130 20190
rect -4130 20170 -4125 20190
rect -4155 20165 -4125 20170
rect -4075 20190 -4045 20195
rect -4075 20170 -4070 20190
rect -4070 20170 -4050 20190
rect -4050 20170 -4045 20190
rect -4075 20165 -4045 20170
rect -3995 20190 -3965 20195
rect -3995 20170 -3990 20190
rect -3990 20170 -3970 20190
rect -3970 20170 -3965 20190
rect -3995 20165 -3965 20170
rect -3915 20190 -3885 20195
rect -3915 20170 -3910 20190
rect -3910 20170 -3890 20190
rect -3890 20170 -3885 20190
rect -3915 20165 -3885 20170
rect -3835 20190 -3805 20195
rect -3835 20170 -3830 20190
rect -3830 20170 -3810 20190
rect -3810 20170 -3805 20190
rect -3835 20165 -3805 20170
rect -3755 20190 -3725 20195
rect -3755 20170 -3750 20190
rect -3750 20170 -3730 20190
rect -3730 20170 -3725 20190
rect -3755 20165 -3725 20170
rect -3675 20190 -3645 20195
rect -3675 20170 -3670 20190
rect -3670 20170 -3650 20190
rect -3650 20170 -3645 20190
rect -3675 20165 -3645 20170
rect -3595 20190 -3565 20195
rect -3595 20170 -3590 20190
rect -3590 20170 -3570 20190
rect -3570 20170 -3565 20190
rect -3595 20165 -3565 20170
rect -3515 20190 -3485 20195
rect -3515 20170 -3510 20190
rect -3510 20170 -3490 20190
rect -3490 20170 -3485 20190
rect -3515 20165 -3485 20170
rect -3435 20190 -3405 20195
rect -3435 20170 -3430 20190
rect -3430 20170 -3410 20190
rect -3410 20170 -3405 20190
rect -3435 20165 -3405 20170
rect -3355 20190 -3325 20195
rect -3355 20170 -3350 20190
rect -3350 20170 -3330 20190
rect -3330 20170 -3325 20190
rect -3355 20165 -3325 20170
rect -3275 20190 -3245 20195
rect -3275 20170 -3270 20190
rect -3270 20170 -3250 20190
rect -3250 20170 -3245 20190
rect -3275 20165 -3245 20170
rect -3195 20190 -3165 20195
rect -3195 20170 -3190 20190
rect -3190 20170 -3170 20190
rect -3170 20170 -3165 20190
rect -3195 20165 -3165 20170
rect -3115 20190 -3085 20195
rect -3115 20170 -3110 20190
rect -3110 20170 -3090 20190
rect -3090 20170 -3085 20190
rect -3115 20165 -3085 20170
rect -3035 20190 -3005 20195
rect -3035 20170 -3030 20190
rect -3030 20170 -3010 20190
rect -3010 20170 -3005 20190
rect -3035 20165 -3005 20170
rect -2955 20190 -2925 20195
rect -2955 20170 -2950 20190
rect -2950 20170 -2930 20190
rect -2930 20170 -2925 20190
rect -2955 20165 -2925 20170
rect -2875 20190 -2845 20195
rect -2875 20170 -2870 20190
rect -2870 20170 -2850 20190
rect -2850 20170 -2845 20190
rect -2875 20165 -2845 20170
rect -2795 20190 -2765 20195
rect -2795 20170 -2790 20190
rect -2790 20170 -2770 20190
rect -2770 20170 -2765 20190
rect -2795 20165 -2765 20170
rect -2715 20190 -2685 20195
rect -2715 20170 -2710 20190
rect -2710 20170 -2690 20190
rect -2690 20170 -2685 20190
rect -2715 20165 -2685 20170
rect -2635 20190 -2605 20195
rect -2635 20170 -2630 20190
rect -2630 20170 -2610 20190
rect -2610 20170 -2605 20190
rect -2635 20165 -2605 20170
rect -2555 20190 -2525 20195
rect -2555 20170 -2550 20190
rect -2550 20170 -2530 20190
rect -2530 20170 -2525 20190
rect -2555 20165 -2525 20170
rect -2475 20190 -2445 20195
rect -2475 20170 -2470 20190
rect -2470 20170 -2450 20190
rect -2450 20170 -2445 20190
rect -2475 20165 -2445 20170
rect -2395 20190 -2365 20195
rect -2395 20170 -2390 20190
rect -2390 20170 -2370 20190
rect -2370 20170 -2365 20190
rect -2395 20165 -2365 20170
rect -2315 20190 -2285 20195
rect -2315 20170 -2310 20190
rect -2310 20170 -2290 20190
rect -2290 20170 -2285 20190
rect -2315 20165 -2285 20170
rect -2235 20190 -2205 20195
rect -2235 20170 -2230 20190
rect -2230 20170 -2210 20190
rect -2210 20170 -2205 20190
rect -2235 20165 -2205 20170
rect -2155 20190 -2125 20195
rect -2155 20170 -2150 20190
rect -2150 20170 -2130 20190
rect -2130 20170 -2125 20190
rect -2155 20165 -2125 20170
rect -2075 20190 -2045 20195
rect -2075 20170 -2070 20190
rect -2070 20170 -2050 20190
rect -2050 20170 -2045 20190
rect -2075 20165 -2045 20170
rect -1995 20190 -1965 20195
rect -1995 20170 -1990 20190
rect -1990 20170 -1970 20190
rect -1970 20170 -1965 20190
rect -1995 20165 -1965 20170
rect -1835 20190 -1805 20195
rect -1835 20170 -1830 20190
rect -1830 20170 -1810 20190
rect -1810 20170 -1805 20190
rect -1835 20165 -1805 20170
rect -1755 20190 -1725 20195
rect -1755 20170 -1750 20190
rect -1750 20170 -1730 20190
rect -1730 20170 -1725 20190
rect -1755 20165 -1725 20170
rect 20525 20030 20555 20035
rect 20525 20010 20530 20030
rect 20530 20010 20550 20030
rect 20550 20010 20555 20030
rect 20525 20005 20555 20010
rect 20605 20030 20635 20035
rect 20605 20010 20610 20030
rect 20610 20010 20630 20030
rect 20630 20010 20635 20030
rect 20605 20005 20635 20010
rect 20685 20030 20715 20035
rect 20685 20010 20690 20030
rect 20690 20010 20710 20030
rect 20710 20010 20715 20030
rect 20685 20005 20715 20010
rect 20765 20030 20795 20035
rect 20765 20010 20770 20030
rect 20770 20010 20790 20030
rect 20790 20010 20795 20030
rect 20765 20005 20795 20010
rect 20845 20030 20875 20035
rect 20845 20010 20850 20030
rect 20850 20010 20870 20030
rect 20870 20010 20875 20030
rect 20845 20005 20875 20010
rect 20925 20030 20955 20035
rect 20925 20010 20930 20030
rect 20930 20010 20950 20030
rect 20950 20010 20955 20030
rect 20925 20005 20955 20010
rect 21005 20030 21035 20035
rect 21005 20010 21010 20030
rect 21010 20010 21030 20030
rect 21030 20010 21035 20030
rect 21005 20005 21035 20010
rect 21085 20030 21115 20035
rect 21085 20010 21090 20030
rect 21090 20010 21110 20030
rect 21110 20010 21115 20030
rect 21085 20005 21115 20010
rect 21165 20030 21195 20035
rect 21165 20010 21170 20030
rect 21170 20010 21190 20030
rect 21190 20010 21195 20030
rect 21165 20005 21195 20010
rect 21245 20030 21275 20035
rect 21245 20010 21250 20030
rect 21250 20010 21270 20030
rect 21270 20010 21275 20030
rect 21245 20005 21275 20010
rect 21325 20030 21355 20035
rect 21325 20010 21330 20030
rect 21330 20010 21350 20030
rect 21350 20010 21355 20030
rect 21325 20005 21355 20010
rect 21405 20030 21435 20035
rect 21405 20010 21410 20030
rect 21410 20010 21430 20030
rect 21430 20010 21435 20030
rect 21405 20005 21435 20010
rect 21485 20030 21515 20035
rect 21485 20010 21490 20030
rect 21490 20010 21510 20030
rect 21510 20010 21515 20030
rect 21485 20005 21515 20010
rect 21565 20030 21595 20035
rect 21565 20010 21570 20030
rect 21570 20010 21590 20030
rect 21590 20010 21595 20030
rect 21565 20005 21595 20010
rect 20525 19870 20555 19875
rect 20525 19850 20530 19870
rect 20530 19850 20550 19870
rect 20550 19850 20555 19870
rect 20525 19845 20555 19850
rect 20605 19870 20635 19875
rect 20605 19850 20610 19870
rect 20610 19850 20630 19870
rect 20630 19850 20635 19870
rect 20605 19845 20635 19850
rect 20685 19870 20715 19875
rect 20685 19850 20690 19870
rect 20690 19850 20710 19870
rect 20710 19850 20715 19870
rect 20685 19845 20715 19850
rect 20765 19870 20795 19875
rect 20765 19850 20770 19870
rect 20770 19850 20790 19870
rect 20790 19850 20795 19870
rect 20765 19845 20795 19850
rect 20845 19870 20875 19875
rect 20845 19850 20850 19870
rect 20850 19850 20870 19870
rect 20870 19850 20875 19870
rect 20845 19845 20875 19850
rect 20925 19870 20955 19875
rect 20925 19850 20930 19870
rect 20930 19850 20950 19870
rect 20950 19850 20955 19870
rect 20925 19845 20955 19850
rect 21005 19870 21035 19875
rect 21005 19850 21010 19870
rect 21010 19850 21030 19870
rect 21030 19850 21035 19870
rect 21005 19845 21035 19850
rect 21085 19870 21115 19875
rect 21085 19850 21090 19870
rect 21090 19850 21110 19870
rect 21110 19850 21115 19870
rect 21085 19845 21115 19850
rect 21165 19870 21195 19875
rect 21165 19850 21170 19870
rect 21170 19850 21190 19870
rect 21190 19850 21195 19870
rect 21165 19845 21195 19850
rect 21245 19870 21275 19875
rect 21245 19850 21250 19870
rect 21250 19850 21270 19870
rect 21270 19850 21275 19870
rect 21245 19845 21275 19850
rect 21325 19870 21355 19875
rect 21325 19850 21330 19870
rect 21330 19850 21350 19870
rect 21350 19850 21355 19870
rect 21325 19845 21355 19850
rect 21405 19870 21435 19875
rect 21405 19850 21410 19870
rect 21410 19850 21430 19870
rect 21430 19850 21435 19870
rect 21405 19845 21435 19850
rect 21485 19870 21515 19875
rect 21485 19850 21490 19870
rect 21490 19850 21510 19870
rect 21510 19850 21515 19870
rect 21485 19845 21515 19850
rect 21565 19870 21595 19875
rect 21565 19850 21570 19870
rect 21570 19850 21590 19870
rect 21590 19850 21595 19870
rect 21565 19845 21595 19850
rect -16555 18870 -16525 18875
rect -16555 18850 -16550 18870
rect -16550 18850 -16530 18870
rect -16530 18850 -16525 18870
rect -16555 18845 -16525 18850
rect -16475 18870 -16445 18875
rect -16475 18850 -16470 18870
rect -16470 18850 -16450 18870
rect -16450 18850 -16445 18870
rect -16475 18845 -16445 18850
rect -16395 18870 -16365 18875
rect -16395 18850 -16390 18870
rect -16390 18850 -16370 18870
rect -16370 18850 -16365 18870
rect -16395 18845 -16365 18850
rect -16315 18870 -16285 18875
rect -16315 18850 -16310 18870
rect -16310 18850 -16290 18870
rect -16290 18850 -16285 18870
rect -16315 18845 -16285 18850
rect -16235 18870 -16205 18875
rect -16235 18850 -16230 18870
rect -16230 18850 -16210 18870
rect -16210 18850 -16205 18870
rect -16235 18845 -16205 18850
rect -16155 18870 -16125 18875
rect -16155 18850 -16150 18870
rect -16150 18850 -16130 18870
rect -16130 18850 -16125 18870
rect -16155 18845 -16125 18850
rect -16075 18870 -16045 18875
rect -16075 18850 -16070 18870
rect -16070 18850 -16050 18870
rect -16050 18850 -16045 18870
rect -16075 18845 -16045 18850
rect -15995 18870 -15965 18875
rect -15995 18850 -15990 18870
rect -15990 18850 -15970 18870
rect -15970 18850 -15965 18870
rect -15995 18845 -15965 18850
rect -15915 18870 -15885 18875
rect -15915 18850 -15910 18870
rect -15910 18850 -15890 18870
rect -15890 18850 -15885 18870
rect -15915 18845 -15885 18850
rect -15835 18870 -15805 18875
rect -15835 18850 -15830 18870
rect -15830 18850 -15810 18870
rect -15810 18850 -15805 18870
rect -15835 18845 -15805 18850
rect -15755 18870 -15725 18875
rect -15755 18850 -15750 18870
rect -15750 18850 -15730 18870
rect -15730 18850 -15725 18870
rect -15755 18845 -15725 18850
rect -15675 18870 -15645 18875
rect -15675 18850 -15670 18870
rect -15670 18850 -15650 18870
rect -15650 18850 -15645 18870
rect -15675 18845 -15645 18850
rect -15595 18870 -15565 18875
rect -15595 18850 -15590 18870
rect -15590 18850 -15570 18870
rect -15570 18850 -15565 18870
rect -15595 18845 -15565 18850
rect -16555 18710 -16525 18715
rect -16555 18690 -16550 18710
rect -16550 18690 -16530 18710
rect -16530 18690 -16525 18710
rect -16555 18685 -16525 18690
rect -16475 18710 -16445 18715
rect -16475 18690 -16470 18710
rect -16470 18690 -16450 18710
rect -16450 18690 -16445 18710
rect -16475 18685 -16445 18690
rect -16395 18710 -16365 18715
rect -16395 18690 -16390 18710
rect -16390 18690 -16370 18710
rect -16370 18690 -16365 18710
rect -16395 18685 -16365 18690
rect -16315 18710 -16285 18715
rect -16315 18690 -16310 18710
rect -16310 18690 -16290 18710
rect -16290 18690 -16285 18710
rect -16315 18685 -16285 18690
rect -16235 18710 -16205 18715
rect -16235 18690 -16230 18710
rect -16230 18690 -16210 18710
rect -16210 18690 -16205 18710
rect -16235 18685 -16205 18690
rect -16155 18710 -16125 18715
rect -16155 18690 -16150 18710
rect -16150 18690 -16130 18710
rect -16130 18690 -16125 18710
rect -16155 18685 -16125 18690
rect -16075 18710 -16045 18715
rect -16075 18690 -16070 18710
rect -16070 18690 -16050 18710
rect -16050 18690 -16045 18710
rect -16075 18685 -16045 18690
rect -15995 18710 -15965 18715
rect -15995 18690 -15990 18710
rect -15990 18690 -15970 18710
rect -15970 18690 -15965 18710
rect -15995 18685 -15965 18690
rect -15915 18710 -15885 18715
rect -15915 18690 -15910 18710
rect -15910 18690 -15890 18710
rect -15890 18690 -15885 18710
rect -15915 18685 -15885 18690
rect -15835 18710 -15805 18715
rect -15835 18690 -15830 18710
rect -15830 18690 -15810 18710
rect -15810 18690 -15805 18710
rect -15835 18685 -15805 18690
rect -15755 18710 -15725 18715
rect -15755 18690 -15750 18710
rect -15750 18690 -15730 18710
rect -15730 18690 -15725 18710
rect -15755 18685 -15725 18690
rect -15675 18710 -15645 18715
rect -15675 18690 -15670 18710
rect -15670 18690 -15650 18710
rect -15650 18690 -15645 18710
rect -15675 18685 -15645 18690
rect -15595 18710 -15565 18715
rect -15595 18690 -15590 18710
rect -15590 18690 -15570 18710
rect -15570 18690 -15565 18710
rect -15595 18685 -15565 18690
rect -16555 18550 -16525 18555
rect -16555 18530 -16550 18550
rect -16550 18530 -16530 18550
rect -16530 18530 -16525 18550
rect -16555 18525 -16525 18530
rect -16475 18550 -16445 18555
rect -16475 18530 -16470 18550
rect -16470 18530 -16450 18550
rect -16450 18530 -16445 18550
rect -16475 18525 -16445 18530
rect -16395 18550 -16365 18555
rect -16395 18530 -16390 18550
rect -16390 18530 -16370 18550
rect -16370 18530 -16365 18550
rect -16395 18525 -16365 18530
rect -16315 18550 -16285 18555
rect -16315 18530 -16310 18550
rect -16310 18530 -16290 18550
rect -16290 18530 -16285 18550
rect -16315 18525 -16285 18530
rect -16235 18550 -16205 18555
rect -16235 18530 -16230 18550
rect -16230 18530 -16210 18550
rect -16210 18530 -16205 18550
rect -16235 18525 -16205 18530
rect -16155 18550 -16125 18555
rect -16155 18530 -16150 18550
rect -16150 18530 -16130 18550
rect -16130 18530 -16125 18550
rect -16155 18525 -16125 18530
rect -16075 18550 -16045 18555
rect -16075 18530 -16070 18550
rect -16070 18530 -16050 18550
rect -16050 18530 -16045 18550
rect -16075 18525 -16045 18530
rect -15995 18550 -15965 18555
rect -15995 18530 -15990 18550
rect -15990 18530 -15970 18550
rect -15970 18530 -15965 18550
rect -15995 18525 -15965 18530
rect -15915 18550 -15885 18555
rect -15915 18530 -15910 18550
rect -15910 18530 -15890 18550
rect -15890 18530 -15885 18550
rect -15915 18525 -15885 18530
rect -15835 18550 -15805 18555
rect -15835 18530 -15830 18550
rect -15830 18530 -15810 18550
rect -15810 18530 -15805 18550
rect -15835 18525 -15805 18530
rect -15755 18550 -15725 18555
rect -15755 18530 -15750 18550
rect -15750 18530 -15730 18550
rect -15730 18530 -15725 18550
rect -15755 18525 -15725 18530
rect -15675 18550 -15645 18555
rect -15675 18530 -15670 18550
rect -15670 18530 -15650 18550
rect -15650 18530 -15645 18550
rect -15675 18525 -15645 18530
rect -15595 18550 -15565 18555
rect -15595 18530 -15590 18550
rect -15590 18530 -15570 18550
rect -15570 18530 -15565 18550
rect -15595 18525 -15565 18530
rect 20525 18030 20555 18035
rect 20525 18010 20530 18030
rect 20530 18010 20550 18030
rect 20550 18010 20555 18030
rect 20525 18005 20555 18010
rect 20605 18030 20635 18035
rect 20605 18010 20610 18030
rect 20610 18010 20630 18030
rect 20630 18010 20635 18030
rect 20605 18005 20635 18010
rect 20685 18030 20715 18035
rect 20685 18010 20690 18030
rect 20690 18010 20710 18030
rect 20710 18010 20715 18030
rect 20685 18005 20715 18010
rect 20765 18030 20795 18035
rect 20765 18010 20770 18030
rect 20770 18010 20790 18030
rect 20790 18010 20795 18030
rect 20765 18005 20795 18010
rect 20845 18030 20875 18035
rect 20845 18010 20850 18030
rect 20850 18010 20870 18030
rect 20870 18010 20875 18030
rect 20845 18005 20875 18010
rect 20925 18030 20955 18035
rect 20925 18010 20930 18030
rect 20930 18010 20950 18030
rect 20950 18010 20955 18030
rect 20925 18005 20955 18010
rect 21005 18030 21035 18035
rect 21005 18010 21010 18030
rect 21010 18010 21030 18030
rect 21030 18010 21035 18030
rect 21005 18005 21035 18010
rect 21085 18030 21115 18035
rect 21085 18010 21090 18030
rect 21090 18010 21110 18030
rect 21110 18010 21115 18030
rect 21085 18005 21115 18010
rect 21165 18030 21195 18035
rect 21165 18010 21170 18030
rect 21170 18010 21190 18030
rect 21190 18010 21195 18030
rect 21165 18005 21195 18010
rect 21245 18030 21275 18035
rect 21245 18010 21250 18030
rect 21250 18010 21270 18030
rect 21270 18010 21275 18030
rect 21245 18005 21275 18010
rect 21325 18030 21355 18035
rect 21325 18010 21330 18030
rect 21330 18010 21350 18030
rect 21350 18010 21355 18030
rect 21325 18005 21355 18010
rect 21405 18030 21435 18035
rect 21405 18010 21410 18030
rect 21410 18010 21430 18030
rect 21430 18010 21435 18030
rect 21405 18005 21435 18010
rect 21485 18030 21515 18035
rect 21485 18010 21490 18030
rect 21490 18010 21510 18030
rect 21510 18010 21515 18030
rect 21485 18005 21515 18010
rect 21565 18030 21595 18035
rect 21565 18010 21570 18030
rect 21570 18010 21590 18030
rect 21590 18010 21595 18030
rect 21565 18005 21595 18010
rect 20525 17870 20555 17875
rect 20525 17850 20530 17870
rect 20530 17850 20550 17870
rect 20550 17850 20555 17870
rect 20525 17845 20555 17850
rect 20605 17870 20635 17875
rect 20605 17850 20610 17870
rect 20610 17850 20630 17870
rect 20630 17850 20635 17870
rect 20605 17845 20635 17850
rect 20685 17870 20715 17875
rect 20685 17850 20690 17870
rect 20690 17850 20710 17870
rect 20710 17850 20715 17870
rect 20685 17845 20715 17850
rect 20765 17870 20795 17875
rect 20765 17850 20770 17870
rect 20770 17850 20790 17870
rect 20790 17850 20795 17870
rect 20765 17845 20795 17850
rect 20845 17870 20875 17875
rect 20845 17850 20850 17870
rect 20850 17850 20870 17870
rect 20870 17850 20875 17870
rect 20845 17845 20875 17850
rect 20925 17870 20955 17875
rect 20925 17850 20930 17870
rect 20930 17850 20950 17870
rect 20950 17850 20955 17870
rect 20925 17845 20955 17850
rect 21005 17870 21035 17875
rect 21005 17850 21010 17870
rect 21010 17850 21030 17870
rect 21030 17850 21035 17870
rect 21005 17845 21035 17850
rect 21085 17870 21115 17875
rect 21085 17850 21090 17870
rect 21090 17850 21110 17870
rect 21110 17850 21115 17870
rect 21085 17845 21115 17850
rect 21165 17870 21195 17875
rect 21165 17850 21170 17870
rect 21170 17850 21190 17870
rect 21190 17850 21195 17870
rect 21165 17845 21195 17850
rect 21245 17870 21275 17875
rect 21245 17850 21250 17870
rect 21250 17850 21270 17870
rect 21270 17850 21275 17870
rect 21245 17845 21275 17850
rect 21325 17870 21355 17875
rect 21325 17850 21330 17870
rect 21330 17850 21350 17870
rect 21350 17850 21355 17870
rect 21325 17845 21355 17850
rect 21405 17870 21435 17875
rect 21405 17850 21410 17870
rect 21410 17850 21430 17870
rect 21430 17850 21435 17870
rect 21405 17845 21435 17850
rect 21485 17870 21515 17875
rect 21485 17850 21490 17870
rect 21490 17850 21510 17870
rect 21510 17850 21515 17870
rect 21485 17845 21515 17850
rect 21565 17870 21595 17875
rect 21565 17850 21570 17870
rect 21570 17850 21590 17870
rect 21590 17850 21595 17870
rect 21565 17845 21595 17850
rect -16555 17350 -16525 17355
rect -16555 17330 -16550 17350
rect -16550 17330 -16530 17350
rect -16530 17330 -16525 17350
rect -16555 17325 -16525 17330
rect -16475 17350 -16445 17355
rect -16475 17330 -16470 17350
rect -16470 17330 -16450 17350
rect -16450 17330 -16445 17350
rect -16475 17325 -16445 17330
rect -16395 17350 -16365 17355
rect -16395 17330 -16390 17350
rect -16390 17330 -16370 17350
rect -16370 17330 -16365 17350
rect -16395 17325 -16365 17330
rect -16315 17350 -16285 17355
rect -16315 17330 -16310 17350
rect -16310 17330 -16290 17350
rect -16290 17330 -16285 17350
rect -16315 17325 -16285 17330
rect -16235 17350 -16205 17355
rect -16235 17330 -16230 17350
rect -16230 17330 -16210 17350
rect -16210 17330 -16205 17350
rect -16235 17325 -16205 17330
rect -16155 17350 -16125 17355
rect -16155 17330 -16150 17350
rect -16150 17330 -16130 17350
rect -16130 17330 -16125 17350
rect -16155 17325 -16125 17330
rect -16075 17350 -16045 17355
rect -16075 17330 -16070 17350
rect -16070 17330 -16050 17350
rect -16050 17330 -16045 17350
rect -16075 17325 -16045 17330
rect -15995 17350 -15965 17355
rect -15995 17330 -15990 17350
rect -15990 17330 -15970 17350
rect -15970 17330 -15965 17350
rect -15995 17325 -15965 17330
rect -15915 17350 -15885 17355
rect -15915 17330 -15910 17350
rect -15910 17330 -15890 17350
rect -15890 17330 -15885 17350
rect -15915 17325 -15885 17330
rect -15835 17350 -15805 17355
rect -15835 17330 -15830 17350
rect -15830 17330 -15810 17350
rect -15810 17330 -15805 17350
rect -15835 17325 -15805 17330
rect -15755 17350 -15725 17355
rect -15755 17330 -15750 17350
rect -15750 17330 -15730 17350
rect -15730 17330 -15725 17350
rect -15755 17325 -15725 17330
rect -15675 17350 -15645 17355
rect -15675 17330 -15670 17350
rect -15670 17330 -15650 17350
rect -15650 17330 -15645 17350
rect -15675 17325 -15645 17330
rect -15595 17350 -15565 17355
rect -15595 17330 -15590 17350
rect -15590 17330 -15570 17350
rect -15570 17330 -15565 17350
rect -15595 17325 -15565 17330
rect -14955 17350 -14925 17355
rect -14955 17330 -14950 17350
rect -14950 17330 -14930 17350
rect -14930 17330 -14925 17350
rect -14955 17325 -14925 17330
rect -14875 17350 -14845 17355
rect -14875 17330 -14870 17350
rect -14870 17330 -14850 17350
rect -14850 17330 -14845 17350
rect -14875 17325 -14845 17330
rect -14795 17350 -14765 17355
rect -14795 17330 -14790 17350
rect -14790 17330 -14770 17350
rect -14770 17330 -14765 17350
rect -14795 17325 -14765 17330
rect -14715 17350 -14685 17355
rect -14715 17330 -14710 17350
rect -14710 17330 -14690 17350
rect -14690 17330 -14685 17350
rect -14715 17325 -14685 17330
rect -14635 17350 -14605 17355
rect -14635 17330 -14630 17350
rect -14630 17330 -14610 17350
rect -14610 17330 -14605 17350
rect -14635 17325 -14605 17330
rect -14555 17350 -14525 17355
rect -14555 17330 -14550 17350
rect -14550 17330 -14530 17350
rect -14530 17330 -14525 17350
rect -14555 17325 -14525 17330
rect -14475 17350 -14445 17355
rect -14475 17330 -14470 17350
rect -14470 17330 -14450 17350
rect -14450 17330 -14445 17350
rect -14475 17325 -14445 17330
rect -14395 17350 -14365 17355
rect -14395 17330 -14390 17350
rect -14390 17330 -14370 17350
rect -14370 17330 -14365 17350
rect -14395 17325 -14365 17330
rect -14315 17350 -14285 17355
rect -14315 17330 -14310 17350
rect -14310 17330 -14290 17350
rect -14290 17330 -14285 17350
rect -14315 17325 -14285 17330
rect -14235 17350 -14205 17355
rect -14235 17330 -14230 17350
rect -14230 17330 -14210 17350
rect -14210 17330 -14205 17350
rect -14235 17325 -14205 17330
rect -14155 17350 -14125 17355
rect -14155 17330 -14150 17350
rect -14150 17330 -14130 17350
rect -14130 17330 -14125 17350
rect -14155 17325 -14125 17330
rect -14075 17350 -14045 17355
rect -14075 17330 -14070 17350
rect -14070 17330 -14050 17350
rect -14050 17330 -14045 17350
rect -14075 17325 -14045 17330
rect -13995 17350 -13965 17355
rect -13995 17330 -13990 17350
rect -13990 17330 -13970 17350
rect -13970 17330 -13965 17350
rect -13995 17325 -13965 17330
rect -13915 17350 -13885 17355
rect -13915 17330 -13910 17350
rect -13910 17330 -13890 17350
rect -13890 17330 -13885 17350
rect -13915 17325 -13885 17330
rect -13835 17350 -13805 17355
rect -13835 17330 -13830 17350
rect -13830 17330 -13810 17350
rect -13810 17330 -13805 17350
rect -13835 17325 -13805 17330
rect -13755 17350 -13725 17355
rect -13755 17330 -13750 17350
rect -13750 17330 -13730 17350
rect -13730 17330 -13725 17350
rect -13755 17325 -13725 17330
rect -13675 17350 -13645 17355
rect -13675 17330 -13670 17350
rect -13670 17330 -13650 17350
rect -13650 17330 -13645 17350
rect -13675 17325 -13645 17330
rect -13595 17350 -13565 17355
rect -13595 17330 -13590 17350
rect -13590 17330 -13570 17350
rect -13570 17330 -13565 17350
rect -13595 17325 -13565 17330
rect -13515 17350 -13485 17355
rect -13515 17330 -13510 17350
rect -13510 17330 -13490 17350
rect -13490 17330 -13485 17350
rect -13515 17325 -13485 17330
rect -13435 17350 -13405 17355
rect -13435 17330 -13430 17350
rect -13430 17330 -13410 17350
rect -13410 17330 -13405 17350
rect -13435 17325 -13405 17330
rect -13355 17350 -13325 17355
rect -13355 17330 -13350 17350
rect -13350 17330 -13330 17350
rect -13330 17330 -13325 17350
rect -13355 17325 -13325 17330
rect -13275 17350 -13245 17355
rect -13275 17330 -13270 17350
rect -13270 17330 -13250 17350
rect -13250 17330 -13245 17350
rect -13275 17325 -13245 17330
rect -13195 17350 -13165 17355
rect -13195 17330 -13190 17350
rect -13190 17330 -13170 17350
rect -13170 17330 -13165 17350
rect -13195 17325 -13165 17330
rect -13115 17350 -13085 17355
rect -13115 17330 -13110 17350
rect -13110 17330 -13090 17350
rect -13090 17330 -13085 17350
rect -13115 17325 -13085 17330
rect -13035 17350 -13005 17355
rect -13035 17330 -13030 17350
rect -13030 17330 -13010 17350
rect -13010 17330 -13005 17350
rect -13035 17325 -13005 17330
rect -12955 17350 -12925 17355
rect -12955 17330 -12950 17350
rect -12950 17330 -12930 17350
rect -12930 17330 -12925 17350
rect -12955 17325 -12925 17330
rect -12875 17350 -12845 17355
rect -12875 17330 -12870 17350
rect -12870 17330 -12850 17350
rect -12850 17330 -12845 17350
rect -12875 17325 -12845 17330
rect -12795 17350 -12765 17355
rect -12795 17330 -12790 17350
rect -12790 17330 -12770 17350
rect -12770 17330 -12765 17350
rect -12795 17325 -12765 17330
rect -12715 17350 -12685 17355
rect -12715 17330 -12710 17350
rect -12710 17330 -12690 17350
rect -12690 17330 -12685 17350
rect -12715 17325 -12685 17330
rect -12635 17350 -12605 17355
rect -12635 17330 -12630 17350
rect -12630 17330 -12610 17350
rect -12610 17330 -12605 17350
rect -12635 17325 -12605 17330
rect -12555 17350 -12525 17355
rect -12555 17330 -12550 17350
rect -12550 17330 -12530 17350
rect -12530 17330 -12525 17350
rect -12555 17325 -12525 17330
rect -12475 17350 -12445 17355
rect -12475 17330 -12470 17350
rect -12470 17330 -12450 17350
rect -12450 17330 -12445 17350
rect -12475 17325 -12445 17330
rect -12395 17350 -12365 17355
rect -12395 17330 -12390 17350
rect -12390 17330 -12370 17350
rect -12370 17330 -12365 17350
rect -12395 17325 -12365 17330
rect -12315 17350 -12285 17355
rect -12315 17330 -12310 17350
rect -12310 17330 -12290 17350
rect -12290 17330 -12285 17350
rect -12315 17325 -12285 17330
rect -12235 17350 -12205 17355
rect -12235 17330 -12230 17350
rect -12230 17330 -12210 17350
rect -12210 17330 -12205 17350
rect -12235 17325 -12205 17330
rect -12155 17350 -12125 17355
rect -12155 17330 -12150 17350
rect -12150 17330 -12130 17350
rect -12130 17330 -12125 17350
rect -12155 17325 -12125 17330
rect -12075 17350 -12045 17355
rect -12075 17330 -12070 17350
rect -12070 17330 -12050 17350
rect -12050 17330 -12045 17350
rect -12075 17325 -12045 17330
rect -11995 17350 -11965 17355
rect -11995 17330 -11990 17350
rect -11990 17330 -11970 17350
rect -11970 17330 -11965 17350
rect -11995 17325 -11965 17330
rect -11915 17350 -11885 17355
rect -11915 17330 -11910 17350
rect -11910 17330 -11890 17350
rect -11890 17330 -11885 17350
rect -11915 17325 -11885 17330
rect -11835 17350 -11805 17355
rect -11835 17330 -11830 17350
rect -11830 17330 -11810 17350
rect -11810 17330 -11805 17350
rect -11835 17325 -11805 17330
rect -11755 17350 -11725 17355
rect -11755 17330 -11750 17350
rect -11750 17330 -11730 17350
rect -11730 17330 -11725 17350
rect -11755 17325 -11725 17330
rect -11675 17350 -11645 17355
rect -11675 17330 -11670 17350
rect -11670 17330 -11650 17350
rect -11650 17330 -11645 17350
rect -11675 17325 -11645 17330
rect -11595 17350 -11565 17355
rect -11595 17330 -11590 17350
rect -11590 17330 -11570 17350
rect -11570 17330 -11565 17350
rect -11595 17325 -11565 17330
rect -11515 17350 -11485 17355
rect -11515 17330 -11510 17350
rect -11510 17330 -11490 17350
rect -11490 17330 -11485 17350
rect -11515 17325 -11485 17330
rect -11435 17350 -11405 17355
rect -11435 17330 -11430 17350
rect -11430 17330 -11410 17350
rect -11410 17330 -11405 17350
rect -11435 17325 -11405 17330
rect -11355 17350 -11325 17355
rect -11355 17330 -11350 17350
rect -11350 17330 -11330 17350
rect -11330 17330 -11325 17350
rect -11355 17325 -11325 17330
rect -11275 17350 -11245 17355
rect -11275 17330 -11270 17350
rect -11270 17330 -11250 17350
rect -11250 17330 -11245 17350
rect -11275 17325 -11245 17330
rect -11195 17350 -11165 17355
rect -11195 17330 -11190 17350
rect -11190 17330 -11170 17350
rect -11170 17330 -11165 17350
rect -11195 17325 -11165 17330
rect -11115 17350 -11085 17355
rect -11115 17330 -11110 17350
rect -11110 17330 -11090 17350
rect -11090 17330 -11085 17350
rect -11115 17325 -11085 17330
rect -11035 17350 -11005 17355
rect -11035 17330 -11030 17350
rect -11030 17330 -11010 17350
rect -11010 17330 -11005 17350
rect -11035 17325 -11005 17330
rect -10955 17350 -10925 17355
rect -10955 17330 -10950 17350
rect -10950 17330 -10930 17350
rect -10930 17330 -10925 17350
rect -10955 17325 -10925 17330
rect -10875 17350 -10845 17355
rect -10875 17330 -10870 17350
rect -10870 17330 -10850 17350
rect -10850 17330 -10845 17350
rect -10875 17325 -10845 17330
rect -10795 17350 -10765 17355
rect -10795 17330 -10790 17350
rect -10790 17330 -10770 17350
rect -10770 17330 -10765 17350
rect -10795 17325 -10765 17330
rect -10715 17350 -10685 17355
rect -10715 17330 -10710 17350
rect -10710 17330 -10690 17350
rect -10690 17330 -10685 17350
rect -10715 17325 -10685 17330
rect -10635 17350 -10605 17355
rect -10635 17330 -10630 17350
rect -10630 17330 -10610 17350
rect -10610 17330 -10605 17350
rect -10635 17325 -10605 17330
rect -10555 17350 -10525 17355
rect -10555 17330 -10550 17350
rect -10550 17330 -10530 17350
rect -10530 17330 -10525 17350
rect -10555 17325 -10525 17330
rect -10475 17350 -10445 17355
rect -10475 17330 -10470 17350
rect -10470 17330 -10450 17350
rect -10450 17330 -10445 17350
rect -10475 17325 -10445 17330
rect -10395 17350 -10365 17355
rect -10395 17330 -10390 17350
rect -10390 17330 -10370 17350
rect -10370 17330 -10365 17350
rect -10395 17325 -10365 17330
rect -10315 17350 -10285 17355
rect -10315 17330 -10310 17350
rect -10310 17330 -10290 17350
rect -10290 17330 -10285 17350
rect -10315 17325 -10285 17330
rect -10235 17350 -10205 17355
rect -10235 17330 -10230 17350
rect -10230 17330 -10210 17350
rect -10210 17330 -10205 17350
rect -10235 17325 -10205 17330
rect -10155 17350 -10125 17355
rect -10155 17330 -10150 17350
rect -10150 17330 -10130 17350
rect -10130 17330 -10125 17350
rect -10155 17325 -10125 17330
rect -10075 17350 -10045 17355
rect -10075 17330 -10070 17350
rect -10070 17330 -10050 17350
rect -10050 17330 -10045 17350
rect -10075 17325 -10045 17330
rect -9995 17350 -9965 17355
rect -9995 17330 -9990 17350
rect -9990 17330 -9970 17350
rect -9970 17330 -9965 17350
rect -9995 17325 -9965 17330
rect -9915 17350 -9885 17355
rect -9915 17330 -9910 17350
rect -9910 17330 -9890 17350
rect -9890 17330 -9885 17350
rect -9915 17325 -9885 17330
rect -9835 17350 -9805 17355
rect -9835 17330 -9830 17350
rect -9830 17330 -9810 17350
rect -9810 17330 -9805 17350
rect -9835 17325 -9805 17330
rect -9755 17350 -9725 17355
rect -9755 17330 -9750 17350
rect -9750 17330 -9730 17350
rect -9730 17330 -9725 17350
rect -9755 17325 -9725 17330
rect -9675 17350 -9645 17355
rect -9675 17330 -9670 17350
rect -9670 17330 -9650 17350
rect -9650 17330 -9645 17350
rect -9675 17325 -9645 17330
rect -9595 17350 -9565 17355
rect -9595 17330 -9590 17350
rect -9590 17330 -9570 17350
rect -9570 17330 -9565 17350
rect -9595 17325 -9565 17330
rect -9515 17350 -9485 17355
rect -9515 17330 -9510 17350
rect -9510 17330 -9490 17350
rect -9490 17330 -9485 17350
rect -9515 17325 -9485 17330
rect -9435 17350 -9405 17355
rect -9435 17330 -9430 17350
rect -9430 17330 -9410 17350
rect -9410 17330 -9405 17350
rect -9435 17325 -9405 17330
rect -9355 17350 -9325 17355
rect -9355 17330 -9350 17350
rect -9350 17330 -9330 17350
rect -9330 17330 -9325 17350
rect -9355 17325 -9325 17330
rect -9275 17350 -9245 17355
rect -9275 17330 -9270 17350
rect -9270 17330 -9250 17350
rect -9250 17330 -9245 17350
rect -9275 17325 -9245 17330
rect -9195 17350 -9165 17355
rect -9195 17330 -9190 17350
rect -9190 17330 -9170 17350
rect -9170 17330 -9165 17350
rect -9195 17325 -9165 17330
rect -9115 17350 -9085 17355
rect -9115 17330 -9110 17350
rect -9110 17330 -9090 17350
rect -9090 17330 -9085 17350
rect -9115 17325 -9085 17330
rect -9035 17350 -9005 17355
rect -9035 17330 -9030 17350
rect -9030 17330 -9010 17350
rect -9010 17330 -9005 17350
rect -9035 17325 -9005 17330
rect -8955 17350 -8925 17355
rect -8955 17330 -8950 17350
rect -8950 17330 -8930 17350
rect -8930 17330 -8925 17350
rect -8955 17325 -8925 17330
rect -8875 17350 -8845 17355
rect -8875 17330 -8870 17350
rect -8870 17330 -8850 17350
rect -8850 17330 -8845 17350
rect -8875 17325 -8845 17330
rect -8795 17350 -8765 17355
rect -8795 17330 -8790 17350
rect -8790 17330 -8770 17350
rect -8770 17330 -8765 17350
rect -8795 17325 -8765 17330
rect -8715 17350 -8685 17355
rect -8715 17330 -8710 17350
rect -8710 17330 -8690 17350
rect -8690 17330 -8685 17350
rect -8715 17325 -8685 17330
rect -8635 17350 -8605 17355
rect -8635 17330 -8630 17350
rect -8630 17330 -8610 17350
rect -8610 17330 -8605 17350
rect -8635 17325 -8605 17330
rect -8555 17350 -8525 17355
rect -8555 17330 -8550 17350
rect -8550 17330 -8530 17350
rect -8530 17330 -8525 17350
rect -8555 17325 -8525 17330
rect -8475 17350 -8445 17355
rect -8475 17330 -8470 17350
rect -8470 17330 -8450 17350
rect -8450 17330 -8445 17350
rect -8475 17325 -8445 17330
rect -8395 17350 -8365 17355
rect -8395 17330 -8390 17350
rect -8390 17330 -8370 17350
rect -8370 17330 -8365 17350
rect -8395 17325 -8365 17330
rect -8315 17350 -8285 17355
rect -8315 17330 -8310 17350
rect -8310 17330 -8290 17350
rect -8290 17330 -8285 17350
rect -8315 17325 -8285 17330
rect -8235 17350 -8205 17355
rect -8235 17330 -8230 17350
rect -8230 17330 -8210 17350
rect -8210 17330 -8205 17350
rect -8235 17325 -8205 17330
rect -8155 17350 -8125 17355
rect -8155 17330 -8150 17350
rect -8150 17330 -8130 17350
rect -8130 17330 -8125 17350
rect -8155 17325 -8125 17330
rect -8075 17350 -8045 17355
rect -8075 17330 -8070 17350
rect -8070 17330 -8050 17350
rect -8050 17330 -8045 17350
rect -8075 17325 -8045 17330
rect -7995 17350 -7965 17355
rect -7995 17330 -7990 17350
rect -7990 17330 -7970 17350
rect -7970 17330 -7965 17350
rect -7995 17325 -7965 17330
rect -7915 17350 -7885 17355
rect -7915 17330 -7910 17350
rect -7910 17330 -7890 17350
rect -7890 17330 -7885 17350
rect -7915 17325 -7885 17330
rect -7835 17350 -7805 17355
rect -7835 17330 -7830 17350
rect -7830 17330 -7810 17350
rect -7810 17330 -7805 17350
rect -7835 17325 -7805 17330
rect -7755 17350 -7725 17355
rect -7755 17330 -7750 17350
rect -7750 17330 -7730 17350
rect -7730 17330 -7725 17350
rect -7755 17325 -7725 17330
rect -7675 17350 -7645 17355
rect -7675 17330 -7670 17350
rect -7670 17330 -7650 17350
rect -7650 17330 -7645 17350
rect -7675 17325 -7645 17330
rect -7595 17350 -7565 17355
rect -7595 17330 -7590 17350
rect -7590 17330 -7570 17350
rect -7570 17330 -7565 17350
rect -7595 17325 -7565 17330
rect -7515 17350 -7485 17355
rect -7515 17330 -7510 17350
rect -7510 17330 -7490 17350
rect -7490 17330 -7485 17350
rect -7515 17325 -7485 17330
rect -7435 17350 -7405 17355
rect -7435 17330 -7430 17350
rect -7430 17330 -7410 17350
rect -7410 17330 -7405 17350
rect -7435 17325 -7405 17330
rect -7355 17350 -7325 17355
rect -7355 17330 -7350 17350
rect -7350 17330 -7330 17350
rect -7330 17330 -7325 17350
rect -7355 17325 -7325 17330
rect -7275 17350 -7245 17355
rect -7275 17330 -7270 17350
rect -7270 17330 -7250 17350
rect -7250 17330 -7245 17350
rect -7275 17325 -7245 17330
rect -7195 17350 -7165 17355
rect -7195 17330 -7190 17350
rect -7190 17330 -7170 17350
rect -7170 17330 -7165 17350
rect -7195 17325 -7165 17330
rect -7115 17350 -7085 17355
rect -7115 17330 -7110 17350
rect -7110 17330 -7090 17350
rect -7090 17330 -7085 17350
rect -7115 17325 -7085 17330
rect -7035 17350 -7005 17355
rect -7035 17330 -7030 17350
rect -7030 17330 -7010 17350
rect -7010 17330 -7005 17350
rect -7035 17325 -7005 17330
rect -6955 17350 -6925 17355
rect -6955 17330 -6950 17350
rect -6950 17330 -6930 17350
rect -6930 17330 -6925 17350
rect -6955 17325 -6925 17330
rect -6875 17350 -6845 17355
rect -6875 17330 -6870 17350
rect -6870 17330 -6850 17350
rect -6850 17330 -6845 17350
rect -6875 17325 -6845 17330
rect -6795 17350 -6765 17355
rect -6795 17330 -6790 17350
rect -6790 17330 -6770 17350
rect -6770 17330 -6765 17350
rect -6795 17325 -6765 17330
rect -6715 17350 -6685 17355
rect -6715 17330 -6710 17350
rect -6710 17330 -6690 17350
rect -6690 17330 -6685 17350
rect -6715 17325 -6685 17330
rect -6635 17350 -6605 17355
rect -6635 17330 -6630 17350
rect -6630 17330 -6610 17350
rect -6610 17330 -6605 17350
rect -6635 17325 -6605 17330
rect -6555 17350 -6525 17355
rect -6555 17330 -6550 17350
rect -6550 17330 -6530 17350
rect -6530 17330 -6525 17350
rect -6555 17325 -6525 17330
rect -6475 17350 -6445 17355
rect -6475 17330 -6470 17350
rect -6470 17330 -6450 17350
rect -6450 17330 -6445 17350
rect -6475 17325 -6445 17330
rect -6395 17350 -6365 17355
rect -6395 17330 -6390 17350
rect -6390 17330 -6370 17350
rect -6370 17330 -6365 17350
rect -6395 17325 -6365 17330
rect -6315 17350 -6285 17355
rect -6315 17330 -6310 17350
rect -6310 17330 -6290 17350
rect -6290 17330 -6285 17350
rect -6315 17325 -6285 17330
rect -6235 17350 -6205 17355
rect -6235 17330 -6230 17350
rect -6230 17330 -6210 17350
rect -6210 17330 -6205 17350
rect -6235 17325 -6205 17330
rect -6155 17350 -6125 17355
rect -6155 17330 -6150 17350
rect -6150 17330 -6130 17350
rect -6130 17330 -6125 17350
rect -6155 17325 -6125 17330
rect -6075 17350 -6045 17355
rect -6075 17330 -6070 17350
rect -6070 17330 -6050 17350
rect -6050 17330 -6045 17350
rect -6075 17325 -6045 17330
rect -5995 17350 -5965 17355
rect -5995 17330 -5990 17350
rect -5990 17330 -5970 17350
rect -5970 17330 -5965 17350
rect -5995 17325 -5965 17330
rect -5915 17350 -5885 17355
rect -5915 17330 -5910 17350
rect -5910 17330 -5890 17350
rect -5890 17330 -5885 17350
rect -5915 17325 -5885 17330
rect -5835 17350 -5805 17355
rect -5835 17330 -5830 17350
rect -5830 17330 -5810 17350
rect -5810 17330 -5805 17350
rect -5835 17325 -5805 17330
rect -5755 17350 -5725 17355
rect -5755 17330 -5750 17350
rect -5750 17330 -5730 17350
rect -5730 17330 -5725 17350
rect -5755 17325 -5725 17330
rect -5435 17350 -5405 17355
rect -5435 17330 -5430 17350
rect -5430 17330 -5410 17350
rect -5410 17330 -5405 17350
rect -5435 17325 -5405 17330
rect -5275 17350 -5245 17355
rect -5275 17330 -5270 17350
rect -5270 17330 -5250 17350
rect -5250 17330 -5245 17350
rect -5275 17325 -5245 17330
rect -16555 17190 -16525 17195
rect -16555 17170 -16550 17190
rect -16550 17170 -16530 17190
rect -16530 17170 -16525 17190
rect -16555 17165 -16525 17170
rect -16475 17190 -16445 17195
rect -16475 17170 -16470 17190
rect -16470 17170 -16450 17190
rect -16450 17170 -16445 17190
rect -16475 17165 -16445 17170
rect -16395 17190 -16365 17195
rect -16395 17170 -16390 17190
rect -16390 17170 -16370 17190
rect -16370 17170 -16365 17190
rect -16395 17165 -16365 17170
rect -16315 17190 -16285 17195
rect -16315 17170 -16310 17190
rect -16310 17170 -16290 17190
rect -16290 17170 -16285 17190
rect -16315 17165 -16285 17170
rect -16235 17190 -16205 17195
rect -16235 17170 -16230 17190
rect -16230 17170 -16210 17190
rect -16210 17170 -16205 17190
rect -16235 17165 -16205 17170
rect -16155 17190 -16125 17195
rect -16155 17170 -16150 17190
rect -16150 17170 -16130 17190
rect -16130 17170 -16125 17190
rect -16155 17165 -16125 17170
rect -16075 17190 -16045 17195
rect -16075 17170 -16070 17190
rect -16070 17170 -16050 17190
rect -16050 17170 -16045 17190
rect -16075 17165 -16045 17170
rect -15995 17190 -15965 17195
rect -15995 17170 -15990 17190
rect -15990 17170 -15970 17190
rect -15970 17170 -15965 17190
rect -15995 17165 -15965 17170
rect -15915 17190 -15885 17195
rect -15915 17170 -15910 17190
rect -15910 17170 -15890 17190
rect -15890 17170 -15885 17190
rect -15915 17165 -15885 17170
rect -15835 17190 -15805 17195
rect -15835 17170 -15830 17190
rect -15830 17170 -15810 17190
rect -15810 17170 -15805 17190
rect -15835 17165 -15805 17170
rect -15755 17190 -15725 17195
rect -15755 17170 -15750 17190
rect -15750 17170 -15730 17190
rect -15730 17170 -15725 17190
rect -15755 17165 -15725 17170
rect -15675 17190 -15645 17195
rect -15675 17170 -15670 17190
rect -15670 17170 -15650 17190
rect -15650 17170 -15645 17190
rect -15675 17165 -15645 17170
rect -15595 17190 -15565 17195
rect -15595 17170 -15590 17190
rect -15590 17170 -15570 17190
rect -15570 17170 -15565 17190
rect -15595 17165 -15565 17170
rect -14955 17190 -14925 17195
rect -14955 17170 -14950 17190
rect -14950 17170 -14930 17190
rect -14930 17170 -14925 17190
rect -14955 17165 -14925 17170
rect -14875 17190 -14845 17195
rect -14875 17170 -14870 17190
rect -14870 17170 -14850 17190
rect -14850 17170 -14845 17190
rect -14875 17165 -14845 17170
rect -14795 17190 -14765 17195
rect -14795 17170 -14790 17190
rect -14790 17170 -14770 17190
rect -14770 17170 -14765 17190
rect -14795 17165 -14765 17170
rect -14715 17190 -14685 17195
rect -14715 17170 -14710 17190
rect -14710 17170 -14690 17190
rect -14690 17170 -14685 17190
rect -14715 17165 -14685 17170
rect -14635 17190 -14605 17195
rect -14635 17170 -14630 17190
rect -14630 17170 -14610 17190
rect -14610 17170 -14605 17190
rect -14635 17165 -14605 17170
rect -14555 17190 -14525 17195
rect -14555 17170 -14550 17190
rect -14550 17170 -14530 17190
rect -14530 17170 -14525 17190
rect -14555 17165 -14525 17170
rect -14475 17190 -14445 17195
rect -14475 17170 -14470 17190
rect -14470 17170 -14450 17190
rect -14450 17170 -14445 17190
rect -14475 17165 -14445 17170
rect -14395 17190 -14365 17195
rect -14395 17170 -14390 17190
rect -14390 17170 -14370 17190
rect -14370 17170 -14365 17190
rect -14395 17165 -14365 17170
rect -14315 17190 -14285 17195
rect -14315 17170 -14310 17190
rect -14310 17170 -14290 17190
rect -14290 17170 -14285 17190
rect -14315 17165 -14285 17170
rect -14235 17190 -14205 17195
rect -14235 17170 -14230 17190
rect -14230 17170 -14210 17190
rect -14210 17170 -14205 17190
rect -14235 17165 -14205 17170
rect -14155 17190 -14125 17195
rect -14155 17170 -14150 17190
rect -14150 17170 -14130 17190
rect -14130 17170 -14125 17190
rect -14155 17165 -14125 17170
rect -14075 17190 -14045 17195
rect -14075 17170 -14070 17190
rect -14070 17170 -14050 17190
rect -14050 17170 -14045 17190
rect -14075 17165 -14045 17170
rect -13995 17190 -13965 17195
rect -13995 17170 -13990 17190
rect -13990 17170 -13970 17190
rect -13970 17170 -13965 17190
rect -13995 17165 -13965 17170
rect -13915 17190 -13885 17195
rect -13915 17170 -13910 17190
rect -13910 17170 -13890 17190
rect -13890 17170 -13885 17190
rect -13915 17165 -13885 17170
rect -13835 17190 -13805 17195
rect -13835 17170 -13830 17190
rect -13830 17170 -13810 17190
rect -13810 17170 -13805 17190
rect -13835 17165 -13805 17170
rect -13755 17190 -13725 17195
rect -13755 17170 -13750 17190
rect -13750 17170 -13730 17190
rect -13730 17170 -13725 17190
rect -13755 17165 -13725 17170
rect -13675 17190 -13645 17195
rect -13675 17170 -13670 17190
rect -13670 17170 -13650 17190
rect -13650 17170 -13645 17190
rect -13675 17165 -13645 17170
rect -13595 17190 -13565 17195
rect -13595 17170 -13590 17190
rect -13590 17170 -13570 17190
rect -13570 17170 -13565 17190
rect -13595 17165 -13565 17170
rect -13515 17190 -13485 17195
rect -13515 17170 -13510 17190
rect -13510 17170 -13490 17190
rect -13490 17170 -13485 17190
rect -13515 17165 -13485 17170
rect -13435 17190 -13405 17195
rect -13435 17170 -13430 17190
rect -13430 17170 -13410 17190
rect -13410 17170 -13405 17190
rect -13435 17165 -13405 17170
rect -13355 17190 -13325 17195
rect -13355 17170 -13350 17190
rect -13350 17170 -13330 17190
rect -13330 17170 -13325 17190
rect -13355 17165 -13325 17170
rect -13275 17190 -13245 17195
rect -13275 17170 -13270 17190
rect -13270 17170 -13250 17190
rect -13250 17170 -13245 17190
rect -13275 17165 -13245 17170
rect -13195 17190 -13165 17195
rect -13195 17170 -13190 17190
rect -13190 17170 -13170 17190
rect -13170 17170 -13165 17190
rect -13195 17165 -13165 17170
rect -13115 17190 -13085 17195
rect -13115 17170 -13110 17190
rect -13110 17170 -13090 17190
rect -13090 17170 -13085 17190
rect -13115 17165 -13085 17170
rect -13035 17190 -13005 17195
rect -13035 17170 -13030 17190
rect -13030 17170 -13010 17190
rect -13010 17170 -13005 17190
rect -13035 17165 -13005 17170
rect -12955 17190 -12925 17195
rect -12955 17170 -12950 17190
rect -12950 17170 -12930 17190
rect -12930 17170 -12925 17190
rect -12955 17165 -12925 17170
rect -12875 17190 -12845 17195
rect -12875 17170 -12870 17190
rect -12870 17170 -12850 17190
rect -12850 17170 -12845 17190
rect -12875 17165 -12845 17170
rect -12795 17190 -12765 17195
rect -12795 17170 -12790 17190
rect -12790 17170 -12770 17190
rect -12770 17170 -12765 17190
rect -12795 17165 -12765 17170
rect -12715 17190 -12685 17195
rect -12715 17170 -12710 17190
rect -12710 17170 -12690 17190
rect -12690 17170 -12685 17190
rect -12715 17165 -12685 17170
rect -12635 17190 -12605 17195
rect -12635 17170 -12630 17190
rect -12630 17170 -12610 17190
rect -12610 17170 -12605 17190
rect -12635 17165 -12605 17170
rect -12555 17190 -12525 17195
rect -12555 17170 -12550 17190
rect -12550 17170 -12530 17190
rect -12530 17170 -12525 17190
rect -12555 17165 -12525 17170
rect -12475 17190 -12445 17195
rect -12475 17170 -12470 17190
rect -12470 17170 -12450 17190
rect -12450 17170 -12445 17190
rect -12475 17165 -12445 17170
rect -12395 17190 -12365 17195
rect -12395 17170 -12390 17190
rect -12390 17170 -12370 17190
rect -12370 17170 -12365 17190
rect -12395 17165 -12365 17170
rect -12315 17190 -12285 17195
rect -12315 17170 -12310 17190
rect -12310 17170 -12290 17190
rect -12290 17170 -12285 17190
rect -12315 17165 -12285 17170
rect -12235 17190 -12205 17195
rect -12235 17170 -12230 17190
rect -12230 17170 -12210 17190
rect -12210 17170 -12205 17190
rect -12235 17165 -12205 17170
rect -12155 17190 -12125 17195
rect -12155 17170 -12150 17190
rect -12150 17170 -12130 17190
rect -12130 17170 -12125 17190
rect -12155 17165 -12125 17170
rect -12075 17190 -12045 17195
rect -12075 17170 -12070 17190
rect -12070 17170 -12050 17190
rect -12050 17170 -12045 17190
rect -12075 17165 -12045 17170
rect -11995 17190 -11965 17195
rect -11995 17170 -11990 17190
rect -11990 17170 -11970 17190
rect -11970 17170 -11965 17190
rect -11995 17165 -11965 17170
rect -11915 17190 -11885 17195
rect -11915 17170 -11910 17190
rect -11910 17170 -11890 17190
rect -11890 17170 -11885 17190
rect -11915 17165 -11885 17170
rect -11835 17190 -11805 17195
rect -11835 17170 -11830 17190
rect -11830 17170 -11810 17190
rect -11810 17170 -11805 17190
rect -11835 17165 -11805 17170
rect -11755 17190 -11725 17195
rect -11755 17170 -11750 17190
rect -11750 17170 -11730 17190
rect -11730 17170 -11725 17190
rect -11755 17165 -11725 17170
rect -11675 17190 -11645 17195
rect -11675 17170 -11670 17190
rect -11670 17170 -11650 17190
rect -11650 17170 -11645 17190
rect -11675 17165 -11645 17170
rect -11595 17190 -11565 17195
rect -11595 17170 -11590 17190
rect -11590 17170 -11570 17190
rect -11570 17170 -11565 17190
rect -11595 17165 -11565 17170
rect -11515 17190 -11485 17195
rect -11515 17170 -11510 17190
rect -11510 17170 -11490 17190
rect -11490 17170 -11485 17190
rect -11515 17165 -11485 17170
rect -11435 17190 -11405 17195
rect -11435 17170 -11430 17190
rect -11430 17170 -11410 17190
rect -11410 17170 -11405 17190
rect -11435 17165 -11405 17170
rect -11355 17190 -11325 17195
rect -11355 17170 -11350 17190
rect -11350 17170 -11330 17190
rect -11330 17170 -11325 17190
rect -11355 17165 -11325 17170
rect -11275 17190 -11245 17195
rect -11275 17170 -11270 17190
rect -11270 17170 -11250 17190
rect -11250 17170 -11245 17190
rect -11275 17165 -11245 17170
rect -11195 17190 -11165 17195
rect -11195 17170 -11190 17190
rect -11190 17170 -11170 17190
rect -11170 17170 -11165 17190
rect -11195 17165 -11165 17170
rect -11115 17190 -11085 17195
rect -11115 17170 -11110 17190
rect -11110 17170 -11090 17190
rect -11090 17170 -11085 17190
rect -11115 17165 -11085 17170
rect -11035 17190 -11005 17195
rect -11035 17170 -11030 17190
rect -11030 17170 -11010 17190
rect -11010 17170 -11005 17190
rect -11035 17165 -11005 17170
rect -10955 17190 -10925 17195
rect -10955 17170 -10950 17190
rect -10950 17170 -10930 17190
rect -10930 17170 -10925 17190
rect -10955 17165 -10925 17170
rect -10875 17190 -10845 17195
rect -10875 17170 -10870 17190
rect -10870 17170 -10850 17190
rect -10850 17170 -10845 17190
rect -10875 17165 -10845 17170
rect -10795 17190 -10765 17195
rect -10795 17170 -10790 17190
rect -10790 17170 -10770 17190
rect -10770 17170 -10765 17190
rect -10795 17165 -10765 17170
rect -10715 17190 -10685 17195
rect -10715 17170 -10710 17190
rect -10710 17170 -10690 17190
rect -10690 17170 -10685 17190
rect -10715 17165 -10685 17170
rect -10635 17190 -10605 17195
rect -10635 17170 -10630 17190
rect -10630 17170 -10610 17190
rect -10610 17170 -10605 17190
rect -10635 17165 -10605 17170
rect -10555 17190 -10525 17195
rect -10555 17170 -10550 17190
rect -10550 17170 -10530 17190
rect -10530 17170 -10525 17190
rect -10555 17165 -10525 17170
rect -10475 17190 -10445 17195
rect -10475 17170 -10470 17190
rect -10470 17170 -10450 17190
rect -10450 17170 -10445 17190
rect -10475 17165 -10445 17170
rect -10395 17190 -10365 17195
rect -10395 17170 -10390 17190
rect -10390 17170 -10370 17190
rect -10370 17170 -10365 17190
rect -10395 17165 -10365 17170
rect -10315 17190 -10285 17195
rect -10315 17170 -10310 17190
rect -10310 17170 -10290 17190
rect -10290 17170 -10285 17190
rect -10315 17165 -10285 17170
rect -10235 17190 -10205 17195
rect -10235 17170 -10230 17190
rect -10230 17170 -10210 17190
rect -10210 17170 -10205 17190
rect -10235 17165 -10205 17170
rect -10155 17190 -10125 17195
rect -10155 17170 -10150 17190
rect -10150 17170 -10130 17190
rect -10130 17170 -10125 17190
rect -10155 17165 -10125 17170
rect -10075 17190 -10045 17195
rect -10075 17170 -10070 17190
rect -10070 17170 -10050 17190
rect -10050 17170 -10045 17190
rect -10075 17165 -10045 17170
rect -9995 17190 -9965 17195
rect -9995 17170 -9990 17190
rect -9990 17170 -9970 17190
rect -9970 17170 -9965 17190
rect -9995 17165 -9965 17170
rect -9915 17190 -9885 17195
rect -9915 17170 -9910 17190
rect -9910 17170 -9890 17190
rect -9890 17170 -9885 17190
rect -9915 17165 -9885 17170
rect -9835 17190 -9805 17195
rect -9835 17170 -9830 17190
rect -9830 17170 -9810 17190
rect -9810 17170 -9805 17190
rect -9835 17165 -9805 17170
rect -9755 17190 -9725 17195
rect -9755 17170 -9750 17190
rect -9750 17170 -9730 17190
rect -9730 17170 -9725 17190
rect -9755 17165 -9725 17170
rect -9675 17190 -9645 17195
rect -9675 17170 -9670 17190
rect -9670 17170 -9650 17190
rect -9650 17170 -9645 17190
rect -9675 17165 -9645 17170
rect -9595 17190 -9565 17195
rect -9595 17170 -9590 17190
rect -9590 17170 -9570 17190
rect -9570 17170 -9565 17190
rect -9595 17165 -9565 17170
rect -9515 17190 -9485 17195
rect -9515 17170 -9510 17190
rect -9510 17170 -9490 17190
rect -9490 17170 -9485 17190
rect -9515 17165 -9485 17170
rect -9435 17190 -9405 17195
rect -9435 17170 -9430 17190
rect -9430 17170 -9410 17190
rect -9410 17170 -9405 17190
rect -9435 17165 -9405 17170
rect -9355 17190 -9325 17195
rect -9355 17170 -9350 17190
rect -9350 17170 -9330 17190
rect -9330 17170 -9325 17190
rect -9355 17165 -9325 17170
rect -9275 17190 -9245 17195
rect -9275 17170 -9270 17190
rect -9270 17170 -9250 17190
rect -9250 17170 -9245 17190
rect -9275 17165 -9245 17170
rect -9195 17190 -9165 17195
rect -9195 17170 -9190 17190
rect -9190 17170 -9170 17190
rect -9170 17170 -9165 17190
rect -9195 17165 -9165 17170
rect -9115 17190 -9085 17195
rect -9115 17170 -9110 17190
rect -9110 17170 -9090 17190
rect -9090 17170 -9085 17190
rect -9115 17165 -9085 17170
rect -9035 17190 -9005 17195
rect -9035 17170 -9030 17190
rect -9030 17170 -9010 17190
rect -9010 17170 -9005 17190
rect -9035 17165 -9005 17170
rect -8955 17190 -8925 17195
rect -8955 17170 -8950 17190
rect -8950 17170 -8930 17190
rect -8930 17170 -8925 17190
rect -8955 17165 -8925 17170
rect -8875 17190 -8845 17195
rect -8875 17170 -8870 17190
rect -8870 17170 -8850 17190
rect -8850 17170 -8845 17190
rect -8875 17165 -8845 17170
rect -8795 17190 -8765 17195
rect -8795 17170 -8790 17190
rect -8790 17170 -8770 17190
rect -8770 17170 -8765 17190
rect -8795 17165 -8765 17170
rect -8715 17190 -8685 17195
rect -8715 17170 -8710 17190
rect -8710 17170 -8690 17190
rect -8690 17170 -8685 17190
rect -8715 17165 -8685 17170
rect -8635 17190 -8605 17195
rect -8635 17170 -8630 17190
rect -8630 17170 -8610 17190
rect -8610 17170 -8605 17190
rect -8635 17165 -8605 17170
rect -8555 17190 -8525 17195
rect -8555 17170 -8550 17190
rect -8550 17170 -8530 17190
rect -8530 17170 -8525 17190
rect -8555 17165 -8525 17170
rect -8475 17190 -8445 17195
rect -8475 17170 -8470 17190
rect -8470 17170 -8450 17190
rect -8450 17170 -8445 17190
rect -8475 17165 -8445 17170
rect -8395 17190 -8365 17195
rect -8395 17170 -8390 17190
rect -8390 17170 -8370 17190
rect -8370 17170 -8365 17190
rect -8395 17165 -8365 17170
rect -8315 17190 -8285 17195
rect -8315 17170 -8310 17190
rect -8310 17170 -8290 17190
rect -8290 17170 -8285 17190
rect -8315 17165 -8285 17170
rect -8235 17190 -8205 17195
rect -8235 17170 -8230 17190
rect -8230 17170 -8210 17190
rect -8210 17170 -8205 17190
rect -8235 17165 -8205 17170
rect -8155 17190 -8125 17195
rect -8155 17170 -8150 17190
rect -8150 17170 -8130 17190
rect -8130 17170 -8125 17190
rect -8155 17165 -8125 17170
rect -8075 17190 -8045 17195
rect -8075 17170 -8070 17190
rect -8070 17170 -8050 17190
rect -8050 17170 -8045 17190
rect -8075 17165 -8045 17170
rect -7995 17190 -7965 17195
rect -7995 17170 -7990 17190
rect -7990 17170 -7970 17190
rect -7970 17170 -7965 17190
rect -7995 17165 -7965 17170
rect -7915 17190 -7885 17195
rect -7915 17170 -7910 17190
rect -7910 17170 -7890 17190
rect -7890 17170 -7885 17190
rect -7915 17165 -7885 17170
rect -7835 17190 -7805 17195
rect -7835 17170 -7830 17190
rect -7830 17170 -7810 17190
rect -7810 17170 -7805 17190
rect -7835 17165 -7805 17170
rect -7755 17190 -7725 17195
rect -7755 17170 -7750 17190
rect -7750 17170 -7730 17190
rect -7730 17170 -7725 17190
rect -7755 17165 -7725 17170
rect -7675 17190 -7645 17195
rect -7675 17170 -7670 17190
rect -7670 17170 -7650 17190
rect -7650 17170 -7645 17190
rect -7675 17165 -7645 17170
rect -7595 17190 -7565 17195
rect -7595 17170 -7590 17190
rect -7590 17170 -7570 17190
rect -7570 17170 -7565 17190
rect -7595 17165 -7565 17170
rect -7515 17190 -7485 17195
rect -7515 17170 -7510 17190
rect -7510 17170 -7490 17190
rect -7490 17170 -7485 17190
rect -7515 17165 -7485 17170
rect -7435 17190 -7405 17195
rect -7435 17170 -7430 17190
rect -7430 17170 -7410 17190
rect -7410 17170 -7405 17190
rect -7435 17165 -7405 17170
rect -7355 17190 -7325 17195
rect -7355 17170 -7350 17190
rect -7350 17170 -7330 17190
rect -7330 17170 -7325 17190
rect -7355 17165 -7325 17170
rect -7275 17190 -7245 17195
rect -7275 17170 -7270 17190
rect -7270 17170 -7250 17190
rect -7250 17170 -7245 17190
rect -7275 17165 -7245 17170
rect -7195 17190 -7165 17195
rect -7195 17170 -7190 17190
rect -7190 17170 -7170 17190
rect -7170 17170 -7165 17190
rect -7195 17165 -7165 17170
rect -7115 17190 -7085 17195
rect -7115 17170 -7110 17190
rect -7110 17170 -7090 17190
rect -7090 17170 -7085 17190
rect -7115 17165 -7085 17170
rect -7035 17190 -7005 17195
rect -7035 17170 -7030 17190
rect -7030 17170 -7010 17190
rect -7010 17170 -7005 17190
rect -7035 17165 -7005 17170
rect -6955 17190 -6925 17195
rect -6955 17170 -6950 17190
rect -6950 17170 -6930 17190
rect -6930 17170 -6925 17190
rect -6955 17165 -6925 17170
rect -6875 17190 -6845 17195
rect -6875 17170 -6870 17190
rect -6870 17170 -6850 17190
rect -6850 17170 -6845 17190
rect -6875 17165 -6845 17170
rect -6795 17190 -6765 17195
rect -6795 17170 -6790 17190
rect -6790 17170 -6770 17190
rect -6770 17170 -6765 17190
rect -6795 17165 -6765 17170
rect -6715 17190 -6685 17195
rect -6715 17170 -6710 17190
rect -6710 17170 -6690 17190
rect -6690 17170 -6685 17190
rect -6715 17165 -6685 17170
rect -6635 17190 -6605 17195
rect -6635 17170 -6630 17190
rect -6630 17170 -6610 17190
rect -6610 17170 -6605 17190
rect -6635 17165 -6605 17170
rect -6555 17190 -6525 17195
rect -6555 17170 -6550 17190
rect -6550 17170 -6530 17190
rect -6530 17170 -6525 17190
rect -6555 17165 -6525 17170
rect -6475 17190 -6445 17195
rect -6475 17170 -6470 17190
rect -6470 17170 -6450 17190
rect -6450 17170 -6445 17190
rect -6475 17165 -6445 17170
rect -6395 17190 -6365 17195
rect -6395 17170 -6390 17190
rect -6390 17170 -6370 17190
rect -6370 17170 -6365 17190
rect -6395 17165 -6365 17170
rect -6315 17190 -6285 17195
rect -6315 17170 -6310 17190
rect -6310 17170 -6290 17190
rect -6290 17170 -6285 17190
rect -6315 17165 -6285 17170
rect -6235 17190 -6205 17195
rect -6235 17170 -6230 17190
rect -6230 17170 -6210 17190
rect -6210 17170 -6205 17190
rect -6235 17165 -6205 17170
rect -6155 17190 -6125 17195
rect -6155 17170 -6150 17190
rect -6150 17170 -6130 17190
rect -6130 17170 -6125 17190
rect -6155 17165 -6125 17170
rect -6075 17190 -6045 17195
rect -6075 17170 -6070 17190
rect -6070 17170 -6050 17190
rect -6050 17170 -6045 17190
rect -6075 17165 -6045 17170
rect -5995 17190 -5965 17195
rect -5995 17170 -5990 17190
rect -5990 17170 -5970 17190
rect -5970 17170 -5965 17190
rect -5995 17165 -5965 17170
rect -5915 17190 -5885 17195
rect -5915 17170 -5910 17190
rect -5910 17170 -5890 17190
rect -5890 17170 -5885 17190
rect -5915 17165 -5885 17170
rect -5835 17190 -5805 17195
rect -5835 17170 -5830 17190
rect -5830 17170 -5810 17190
rect -5810 17170 -5805 17190
rect -5835 17165 -5805 17170
rect -5755 17190 -5725 17195
rect -5755 17170 -5750 17190
rect -5750 17170 -5730 17190
rect -5730 17170 -5725 17190
rect -5755 17165 -5725 17170
rect -5435 17190 -5405 17195
rect -5435 17170 -5430 17190
rect -5430 17170 -5410 17190
rect -5410 17170 -5405 17190
rect -5435 17165 -5405 17170
rect -5275 17190 -5245 17195
rect -5275 17170 -5270 17190
rect -5270 17170 -5250 17190
rect -5250 17170 -5245 17190
rect -5275 17165 -5245 17170
rect -14955 16470 -14925 16475
rect -14955 16450 -14950 16470
rect -14950 16450 -14930 16470
rect -14930 16450 -14925 16470
rect -14955 16445 -14925 16450
rect -14875 16470 -14845 16475
rect -14875 16450 -14870 16470
rect -14870 16450 -14850 16470
rect -14850 16450 -14845 16470
rect -14875 16445 -14845 16450
rect -14795 16470 -14765 16475
rect -14795 16450 -14790 16470
rect -14790 16450 -14770 16470
rect -14770 16450 -14765 16470
rect -14795 16445 -14765 16450
rect -14715 16470 -14685 16475
rect -14715 16450 -14710 16470
rect -14710 16450 -14690 16470
rect -14690 16450 -14685 16470
rect -14715 16445 -14685 16450
rect -14635 16470 -14605 16475
rect -14635 16450 -14630 16470
rect -14630 16450 -14610 16470
rect -14610 16450 -14605 16470
rect -14635 16445 -14605 16450
rect -14555 16470 -14525 16475
rect -14555 16450 -14550 16470
rect -14550 16450 -14530 16470
rect -14530 16450 -14525 16470
rect -14555 16445 -14525 16450
rect -14475 16470 -14445 16475
rect -14475 16450 -14470 16470
rect -14470 16450 -14450 16470
rect -14450 16450 -14445 16470
rect -14475 16445 -14445 16450
rect -14395 16470 -14365 16475
rect -14395 16450 -14390 16470
rect -14390 16450 -14370 16470
rect -14370 16450 -14365 16470
rect -14395 16445 -14365 16450
rect -14315 16470 -14285 16475
rect -14315 16450 -14310 16470
rect -14310 16450 -14290 16470
rect -14290 16450 -14285 16470
rect -14315 16445 -14285 16450
rect -14235 16470 -14205 16475
rect -14235 16450 -14230 16470
rect -14230 16450 -14210 16470
rect -14210 16450 -14205 16470
rect -14235 16445 -14205 16450
rect -14155 16470 -14125 16475
rect -14155 16450 -14150 16470
rect -14150 16450 -14130 16470
rect -14130 16450 -14125 16470
rect -14155 16445 -14125 16450
rect -14075 16470 -14045 16475
rect -14075 16450 -14070 16470
rect -14070 16450 -14050 16470
rect -14050 16450 -14045 16470
rect -14075 16445 -14045 16450
rect -13995 16470 -13965 16475
rect -13995 16450 -13990 16470
rect -13990 16450 -13970 16470
rect -13970 16450 -13965 16470
rect -13995 16445 -13965 16450
rect -13915 16470 -13885 16475
rect -13915 16450 -13910 16470
rect -13910 16450 -13890 16470
rect -13890 16450 -13885 16470
rect -13915 16445 -13885 16450
rect -13835 16470 -13805 16475
rect -13835 16450 -13830 16470
rect -13830 16450 -13810 16470
rect -13810 16450 -13805 16470
rect -13835 16445 -13805 16450
rect -13755 16470 -13725 16475
rect -13755 16450 -13750 16470
rect -13750 16450 -13730 16470
rect -13730 16450 -13725 16470
rect -13755 16445 -13725 16450
rect -13675 16470 -13645 16475
rect -13675 16450 -13670 16470
rect -13670 16450 -13650 16470
rect -13650 16450 -13645 16470
rect -13675 16445 -13645 16450
rect -13595 16470 -13565 16475
rect -13595 16450 -13590 16470
rect -13590 16450 -13570 16470
rect -13570 16450 -13565 16470
rect -13595 16445 -13565 16450
rect -13515 16470 -13485 16475
rect -13515 16450 -13510 16470
rect -13510 16450 -13490 16470
rect -13490 16450 -13485 16470
rect -13515 16445 -13485 16450
rect -13435 16470 -13405 16475
rect -13435 16450 -13430 16470
rect -13430 16450 -13410 16470
rect -13410 16450 -13405 16470
rect -13435 16445 -13405 16450
rect -13355 16470 -13325 16475
rect -13355 16450 -13350 16470
rect -13350 16450 -13330 16470
rect -13330 16450 -13325 16470
rect -13355 16445 -13325 16450
rect -13275 16470 -13245 16475
rect -13275 16450 -13270 16470
rect -13270 16450 -13250 16470
rect -13250 16450 -13245 16470
rect -13275 16445 -13245 16450
rect -13195 16470 -13165 16475
rect -13195 16450 -13190 16470
rect -13190 16450 -13170 16470
rect -13170 16450 -13165 16470
rect -13195 16445 -13165 16450
rect -13115 16470 -13085 16475
rect -13115 16450 -13110 16470
rect -13110 16450 -13090 16470
rect -13090 16450 -13085 16470
rect -13115 16445 -13085 16450
rect -13035 16470 -13005 16475
rect -13035 16450 -13030 16470
rect -13030 16450 -13010 16470
rect -13010 16450 -13005 16470
rect -13035 16445 -13005 16450
rect -12955 16470 -12925 16475
rect -12955 16450 -12950 16470
rect -12950 16450 -12930 16470
rect -12930 16450 -12925 16470
rect -12955 16445 -12925 16450
rect -12875 16470 -12845 16475
rect -12875 16450 -12870 16470
rect -12870 16450 -12850 16470
rect -12850 16450 -12845 16470
rect -12875 16445 -12845 16450
rect -12795 16470 -12765 16475
rect -12795 16450 -12790 16470
rect -12790 16450 -12770 16470
rect -12770 16450 -12765 16470
rect -12795 16445 -12765 16450
rect -12715 16470 -12685 16475
rect -12715 16450 -12710 16470
rect -12710 16450 -12690 16470
rect -12690 16450 -12685 16470
rect -12715 16445 -12685 16450
rect -12635 16470 -12605 16475
rect -12635 16450 -12630 16470
rect -12630 16450 -12610 16470
rect -12610 16450 -12605 16470
rect -12635 16445 -12605 16450
rect -12555 16470 -12525 16475
rect -12555 16450 -12550 16470
rect -12550 16450 -12530 16470
rect -12530 16450 -12525 16470
rect -12555 16445 -12525 16450
rect -12475 16470 -12445 16475
rect -12475 16450 -12470 16470
rect -12470 16450 -12450 16470
rect -12450 16450 -12445 16470
rect -12475 16445 -12445 16450
rect -12395 16470 -12365 16475
rect -12395 16450 -12390 16470
rect -12390 16450 -12370 16470
rect -12370 16450 -12365 16470
rect -12395 16445 -12365 16450
rect -12315 16470 -12285 16475
rect -12315 16450 -12310 16470
rect -12310 16450 -12290 16470
rect -12290 16450 -12285 16470
rect -12315 16445 -12285 16450
rect -12235 16470 -12205 16475
rect -12235 16450 -12230 16470
rect -12230 16450 -12210 16470
rect -12210 16450 -12205 16470
rect -12235 16445 -12205 16450
rect -12155 16470 -12125 16475
rect -12155 16450 -12150 16470
rect -12150 16450 -12130 16470
rect -12130 16450 -12125 16470
rect -12155 16445 -12125 16450
rect -12075 16470 -12045 16475
rect -12075 16450 -12070 16470
rect -12070 16450 -12050 16470
rect -12050 16450 -12045 16470
rect -12075 16445 -12045 16450
rect -11995 16470 -11965 16475
rect -11995 16450 -11990 16470
rect -11990 16450 -11970 16470
rect -11970 16450 -11965 16470
rect -11995 16445 -11965 16450
rect -11915 16470 -11885 16475
rect -11915 16450 -11910 16470
rect -11910 16450 -11890 16470
rect -11890 16450 -11885 16470
rect -11915 16445 -11885 16450
rect -11835 16470 -11805 16475
rect -11835 16450 -11830 16470
rect -11830 16450 -11810 16470
rect -11810 16450 -11805 16470
rect -11835 16445 -11805 16450
rect -11755 16470 -11725 16475
rect -11755 16450 -11750 16470
rect -11750 16450 -11730 16470
rect -11730 16450 -11725 16470
rect -11755 16445 -11725 16450
rect -11675 16470 -11645 16475
rect -11675 16450 -11670 16470
rect -11670 16450 -11650 16470
rect -11650 16450 -11645 16470
rect -11675 16445 -11645 16450
rect -11595 16470 -11565 16475
rect -11595 16450 -11590 16470
rect -11590 16450 -11570 16470
rect -11570 16450 -11565 16470
rect -11595 16445 -11565 16450
rect -11515 16470 -11485 16475
rect -11515 16450 -11510 16470
rect -11510 16450 -11490 16470
rect -11490 16450 -11485 16470
rect -11515 16445 -11485 16450
rect -11435 16470 -11405 16475
rect -11435 16450 -11430 16470
rect -11430 16450 -11410 16470
rect -11410 16450 -11405 16470
rect -11435 16445 -11405 16450
rect -11355 16470 -11325 16475
rect -11355 16450 -11350 16470
rect -11350 16450 -11330 16470
rect -11330 16450 -11325 16470
rect -11355 16445 -11325 16450
rect -11275 16470 -11245 16475
rect -11275 16450 -11270 16470
rect -11270 16450 -11250 16470
rect -11250 16450 -11245 16470
rect -11275 16445 -11245 16450
rect -11195 16470 -11165 16475
rect -11195 16450 -11190 16470
rect -11190 16450 -11170 16470
rect -11170 16450 -11165 16470
rect -11195 16445 -11165 16450
rect -11115 16470 -11085 16475
rect -11115 16450 -11110 16470
rect -11110 16450 -11090 16470
rect -11090 16450 -11085 16470
rect -11115 16445 -11085 16450
rect -11035 16470 -11005 16475
rect -11035 16450 -11030 16470
rect -11030 16450 -11010 16470
rect -11010 16450 -11005 16470
rect -11035 16445 -11005 16450
rect -10955 16470 -10925 16475
rect -10955 16450 -10950 16470
rect -10950 16450 -10930 16470
rect -10930 16450 -10925 16470
rect -10955 16445 -10925 16450
rect -10875 16470 -10845 16475
rect -10875 16450 -10870 16470
rect -10870 16450 -10850 16470
rect -10850 16450 -10845 16470
rect -10875 16445 -10845 16450
rect -10795 16470 -10765 16475
rect -10795 16450 -10790 16470
rect -10790 16450 -10770 16470
rect -10770 16450 -10765 16470
rect -10795 16445 -10765 16450
rect -10715 16470 -10685 16475
rect -10715 16450 -10710 16470
rect -10710 16450 -10690 16470
rect -10690 16450 -10685 16470
rect -10715 16445 -10685 16450
rect -10635 16470 -10605 16475
rect -10635 16450 -10630 16470
rect -10630 16450 -10610 16470
rect -10610 16450 -10605 16470
rect -10635 16445 -10605 16450
rect -10555 16470 -10525 16475
rect -10555 16450 -10550 16470
rect -10550 16450 -10530 16470
rect -10530 16450 -10525 16470
rect -10555 16445 -10525 16450
rect -10475 16470 -10445 16475
rect -10475 16450 -10470 16470
rect -10470 16450 -10450 16470
rect -10450 16450 -10445 16470
rect -10475 16445 -10445 16450
rect -10395 16470 -10365 16475
rect -10395 16450 -10390 16470
rect -10390 16450 -10370 16470
rect -10370 16450 -10365 16470
rect -10395 16445 -10365 16450
rect -10315 16470 -10285 16475
rect -10315 16450 -10310 16470
rect -10310 16450 -10290 16470
rect -10290 16450 -10285 16470
rect -10315 16445 -10285 16450
rect -10235 16470 -10205 16475
rect -10235 16450 -10230 16470
rect -10230 16450 -10210 16470
rect -10210 16450 -10205 16470
rect -10235 16445 -10205 16450
rect -10155 16470 -10125 16475
rect -10155 16450 -10150 16470
rect -10150 16450 -10130 16470
rect -10130 16450 -10125 16470
rect -10155 16445 -10125 16450
rect -10075 16470 -10045 16475
rect -10075 16450 -10070 16470
rect -10070 16450 -10050 16470
rect -10050 16450 -10045 16470
rect -10075 16445 -10045 16450
rect -9995 16470 -9965 16475
rect -9995 16450 -9990 16470
rect -9990 16450 -9970 16470
rect -9970 16450 -9965 16470
rect -9995 16445 -9965 16450
rect -9915 16470 -9885 16475
rect -9915 16450 -9910 16470
rect -9910 16450 -9890 16470
rect -9890 16450 -9885 16470
rect -9915 16445 -9885 16450
rect -9835 16470 -9805 16475
rect -9835 16450 -9830 16470
rect -9830 16450 -9810 16470
rect -9810 16450 -9805 16470
rect -9835 16445 -9805 16450
rect -9755 16470 -9725 16475
rect -9755 16450 -9750 16470
rect -9750 16450 -9730 16470
rect -9730 16450 -9725 16470
rect -9755 16445 -9725 16450
rect -9675 16470 -9645 16475
rect -9675 16450 -9670 16470
rect -9670 16450 -9650 16470
rect -9650 16450 -9645 16470
rect -9675 16445 -9645 16450
rect -9595 16470 -9565 16475
rect -9595 16450 -9590 16470
rect -9590 16450 -9570 16470
rect -9570 16450 -9565 16470
rect -9595 16445 -9565 16450
rect -9515 16470 -9485 16475
rect -9515 16450 -9510 16470
rect -9510 16450 -9490 16470
rect -9490 16450 -9485 16470
rect -9515 16445 -9485 16450
rect -9435 16470 -9405 16475
rect -9435 16450 -9430 16470
rect -9430 16450 -9410 16470
rect -9410 16450 -9405 16470
rect -9435 16445 -9405 16450
rect -9355 16470 -9325 16475
rect -9355 16450 -9350 16470
rect -9350 16450 -9330 16470
rect -9330 16450 -9325 16470
rect -9355 16445 -9325 16450
rect -9275 16470 -9245 16475
rect -9275 16450 -9270 16470
rect -9270 16450 -9250 16470
rect -9250 16450 -9245 16470
rect -9275 16445 -9245 16450
rect -9195 16470 -9165 16475
rect -9195 16450 -9190 16470
rect -9190 16450 -9170 16470
rect -9170 16450 -9165 16470
rect -9195 16445 -9165 16450
rect -9115 16470 -9085 16475
rect -9115 16450 -9110 16470
rect -9110 16450 -9090 16470
rect -9090 16450 -9085 16470
rect -9115 16445 -9085 16450
rect -9035 16470 -9005 16475
rect -9035 16450 -9030 16470
rect -9030 16450 -9010 16470
rect -9010 16450 -9005 16470
rect -9035 16445 -9005 16450
rect -8955 16470 -8925 16475
rect -8955 16450 -8950 16470
rect -8950 16450 -8930 16470
rect -8930 16450 -8925 16470
rect -8955 16445 -8925 16450
rect -8875 16470 -8845 16475
rect -8875 16450 -8870 16470
rect -8870 16450 -8850 16470
rect -8850 16450 -8845 16470
rect -8875 16445 -8845 16450
rect -8795 16470 -8765 16475
rect -8795 16450 -8790 16470
rect -8790 16450 -8770 16470
rect -8770 16450 -8765 16470
rect -8795 16445 -8765 16450
rect -8715 16470 -8685 16475
rect -8715 16450 -8710 16470
rect -8710 16450 -8690 16470
rect -8690 16450 -8685 16470
rect -8715 16445 -8685 16450
rect -8635 16470 -8605 16475
rect -8635 16450 -8630 16470
rect -8630 16450 -8610 16470
rect -8610 16450 -8605 16470
rect -8635 16445 -8605 16450
rect -8555 16470 -8525 16475
rect -8555 16450 -8550 16470
rect -8550 16450 -8530 16470
rect -8530 16450 -8525 16470
rect -8555 16445 -8525 16450
rect -8475 16470 -8445 16475
rect -8475 16450 -8470 16470
rect -8470 16450 -8450 16470
rect -8450 16450 -8445 16470
rect -8475 16445 -8445 16450
rect -8395 16470 -8365 16475
rect -8395 16450 -8390 16470
rect -8390 16450 -8370 16470
rect -8370 16450 -8365 16470
rect -8395 16445 -8365 16450
rect -8315 16470 -8285 16475
rect -8315 16450 -8310 16470
rect -8310 16450 -8290 16470
rect -8290 16450 -8285 16470
rect -8315 16445 -8285 16450
rect -8235 16470 -8205 16475
rect -8235 16450 -8230 16470
rect -8230 16450 -8210 16470
rect -8210 16450 -8205 16470
rect -8235 16445 -8205 16450
rect -8155 16470 -8125 16475
rect -8155 16450 -8150 16470
rect -8150 16450 -8130 16470
rect -8130 16450 -8125 16470
rect -8155 16445 -8125 16450
rect -8075 16470 -8045 16475
rect -8075 16450 -8070 16470
rect -8070 16450 -8050 16470
rect -8050 16450 -8045 16470
rect -8075 16445 -8045 16450
rect -7995 16470 -7965 16475
rect -7995 16450 -7990 16470
rect -7990 16450 -7970 16470
rect -7970 16450 -7965 16470
rect -7995 16445 -7965 16450
rect -7915 16470 -7885 16475
rect -7915 16450 -7910 16470
rect -7910 16450 -7890 16470
rect -7890 16450 -7885 16470
rect -7915 16445 -7885 16450
rect -7835 16470 -7805 16475
rect -7835 16450 -7830 16470
rect -7830 16450 -7810 16470
rect -7810 16450 -7805 16470
rect -7835 16445 -7805 16450
rect -7755 16470 -7725 16475
rect -7755 16450 -7750 16470
rect -7750 16450 -7730 16470
rect -7730 16450 -7725 16470
rect -7755 16445 -7725 16450
rect -7675 16470 -7645 16475
rect -7675 16450 -7670 16470
rect -7670 16450 -7650 16470
rect -7650 16450 -7645 16470
rect -7675 16445 -7645 16450
rect -7595 16470 -7565 16475
rect -7595 16450 -7590 16470
rect -7590 16450 -7570 16470
rect -7570 16450 -7565 16470
rect -7595 16445 -7565 16450
rect -7515 16470 -7485 16475
rect -7515 16450 -7510 16470
rect -7510 16450 -7490 16470
rect -7490 16450 -7485 16470
rect -7515 16445 -7485 16450
rect -7435 16470 -7405 16475
rect -7435 16450 -7430 16470
rect -7430 16450 -7410 16470
rect -7410 16450 -7405 16470
rect -7435 16445 -7405 16450
rect -7355 16470 -7325 16475
rect -7355 16450 -7350 16470
rect -7350 16450 -7330 16470
rect -7330 16450 -7325 16470
rect -7355 16445 -7325 16450
rect -7275 16470 -7245 16475
rect -7275 16450 -7270 16470
rect -7270 16450 -7250 16470
rect -7250 16450 -7245 16470
rect -7275 16445 -7245 16450
rect -7195 16470 -7165 16475
rect -7195 16450 -7190 16470
rect -7190 16450 -7170 16470
rect -7170 16450 -7165 16470
rect -7195 16445 -7165 16450
rect -7115 16470 -7085 16475
rect -7115 16450 -7110 16470
rect -7110 16450 -7090 16470
rect -7090 16450 -7085 16470
rect -7115 16445 -7085 16450
rect -7035 16470 -7005 16475
rect -7035 16450 -7030 16470
rect -7030 16450 -7010 16470
rect -7010 16450 -7005 16470
rect -7035 16445 -7005 16450
rect -6955 16470 -6925 16475
rect -6955 16450 -6950 16470
rect -6950 16450 -6930 16470
rect -6930 16450 -6925 16470
rect -6955 16445 -6925 16450
rect -6875 16470 -6845 16475
rect -6875 16450 -6870 16470
rect -6870 16450 -6850 16470
rect -6850 16450 -6845 16470
rect -6875 16445 -6845 16450
rect -6795 16470 -6765 16475
rect -6795 16450 -6790 16470
rect -6790 16450 -6770 16470
rect -6770 16450 -6765 16470
rect -6795 16445 -6765 16450
rect -6715 16470 -6685 16475
rect -6715 16450 -6710 16470
rect -6710 16450 -6690 16470
rect -6690 16450 -6685 16470
rect -6715 16445 -6685 16450
rect -6635 16470 -6605 16475
rect -6635 16450 -6630 16470
rect -6630 16450 -6610 16470
rect -6610 16450 -6605 16470
rect -6635 16445 -6605 16450
rect -6555 16470 -6525 16475
rect -6555 16450 -6550 16470
rect -6550 16450 -6530 16470
rect -6530 16450 -6525 16470
rect -6555 16445 -6525 16450
rect -6475 16470 -6445 16475
rect -6475 16450 -6470 16470
rect -6470 16450 -6450 16470
rect -6450 16450 -6445 16470
rect -6475 16445 -6445 16450
rect -6395 16470 -6365 16475
rect -6395 16450 -6390 16470
rect -6390 16450 -6370 16470
rect -6370 16450 -6365 16470
rect -6395 16445 -6365 16450
rect -6315 16470 -6285 16475
rect -6315 16450 -6310 16470
rect -6310 16450 -6290 16470
rect -6290 16450 -6285 16470
rect -6315 16445 -6285 16450
rect -6235 16470 -6205 16475
rect -6235 16450 -6230 16470
rect -6230 16450 -6210 16470
rect -6210 16450 -6205 16470
rect -6235 16445 -6205 16450
rect -6155 16470 -6125 16475
rect -6155 16450 -6150 16470
rect -6150 16450 -6130 16470
rect -6130 16450 -6125 16470
rect -6155 16445 -6125 16450
rect -6075 16470 -6045 16475
rect -6075 16450 -6070 16470
rect -6070 16450 -6050 16470
rect -6050 16450 -6045 16470
rect -6075 16445 -6045 16450
rect -5995 16470 -5965 16475
rect -5995 16450 -5990 16470
rect -5990 16450 -5970 16470
rect -5970 16450 -5965 16470
rect -5995 16445 -5965 16450
rect -5915 16470 -5885 16475
rect -5915 16450 -5910 16470
rect -5910 16450 -5890 16470
rect -5890 16450 -5885 16470
rect -5915 16445 -5885 16450
rect -5835 16470 -5805 16475
rect -5835 16450 -5830 16470
rect -5830 16450 -5810 16470
rect -5810 16450 -5805 16470
rect -5835 16445 -5805 16450
rect -5755 16470 -5725 16475
rect -5755 16450 -5750 16470
rect -5750 16450 -5730 16470
rect -5730 16450 -5725 16470
rect -5755 16445 -5725 16450
rect -5595 16470 -5565 16475
rect -5595 16450 -5590 16470
rect -5590 16450 -5570 16470
rect -5570 16450 -5565 16470
rect -5595 16445 -5565 16450
rect -5435 16470 -5405 16475
rect -5435 16450 -5430 16470
rect -5430 16450 -5410 16470
rect -5410 16450 -5405 16470
rect -5435 16445 -5405 16450
rect -5355 16470 -5325 16475
rect -5355 16450 -5350 16470
rect -5350 16450 -5330 16470
rect -5330 16450 -5325 16470
rect -5355 16445 -5325 16450
rect -5275 16470 -5245 16475
rect -5275 16450 -5270 16470
rect -5270 16450 -5250 16470
rect -5250 16450 -5245 16470
rect -5275 16445 -5245 16450
rect -5195 16470 -5165 16475
rect -5195 16450 -5190 16470
rect -5190 16450 -5170 16470
rect -5170 16450 -5165 16470
rect -5195 16445 -5165 16450
rect -5115 16470 -5085 16475
rect -5115 16450 -5110 16470
rect -5110 16450 -5090 16470
rect -5090 16450 -5085 16470
rect -5115 16445 -5085 16450
rect -5035 16470 -5005 16475
rect -5035 16450 -5030 16470
rect -5030 16450 -5010 16470
rect -5010 16450 -5005 16470
rect -5035 16445 -5005 16450
rect -4955 16470 -4925 16475
rect -4955 16450 -4950 16470
rect -4950 16450 -4930 16470
rect -4930 16450 -4925 16470
rect -4955 16445 -4925 16450
rect -4875 16470 -4845 16475
rect -4875 16450 -4870 16470
rect -4870 16450 -4850 16470
rect -4850 16450 -4845 16470
rect -4875 16445 -4845 16450
rect -4795 16470 -4765 16475
rect -4795 16450 -4790 16470
rect -4790 16450 -4770 16470
rect -4770 16450 -4765 16470
rect -4795 16445 -4765 16450
rect -4715 16470 -4685 16475
rect -4715 16450 -4710 16470
rect -4710 16450 -4690 16470
rect -4690 16450 -4685 16470
rect -4715 16445 -4685 16450
rect -4635 16470 -4605 16475
rect -4635 16450 -4630 16470
rect -4630 16450 -4610 16470
rect -4610 16450 -4605 16470
rect -4635 16445 -4605 16450
rect -4555 16470 -4525 16475
rect -4555 16450 -4550 16470
rect -4550 16450 -4530 16470
rect -4530 16450 -4525 16470
rect -4555 16445 -4525 16450
rect -4475 16470 -4445 16475
rect -4475 16450 -4470 16470
rect -4470 16450 -4450 16470
rect -4450 16450 -4445 16470
rect -4475 16445 -4445 16450
rect -4395 16470 -4365 16475
rect -4395 16450 -4390 16470
rect -4390 16450 -4370 16470
rect -4370 16450 -4365 16470
rect -4395 16445 -4365 16450
rect -4315 16470 -4285 16475
rect -4315 16450 -4310 16470
rect -4310 16450 -4290 16470
rect -4290 16450 -4285 16470
rect -4315 16445 -4285 16450
rect -4235 16470 -4205 16475
rect -4235 16450 -4230 16470
rect -4230 16450 -4210 16470
rect -4210 16450 -4205 16470
rect -4235 16445 -4205 16450
rect -4155 16470 -4125 16475
rect -4155 16450 -4150 16470
rect -4150 16450 -4130 16470
rect -4130 16450 -4125 16470
rect -4155 16445 -4125 16450
rect -4075 16470 -4045 16475
rect -4075 16450 -4070 16470
rect -4070 16450 -4050 16470
rect -4050 16450 -4045 16470
rect -4075 16445 -4045 16450
rect -3995 16470 -3965 16475
rect -3995 16450 -3990 16470
rect -3990 16450 -3970 16470
rect -3970 16450 -3965 16470
rect -3995 16445 -3965 16450
rect -3915 16470 -3885 16475
rect -3915 16450 -3910 16470
rect -3910 16450 -3890 16470
rect -3890 16450 -3885 16470
rect -3915 16445 -3885 16450
rect -3835 16470 -3805 16475
rect -3835 16450 -3830 16470
rect -3830 16450 -3810 16470
rect -3810 16450 -3805 16470
rect -3835 16445 -3805 16450
rect -3755 16470 -3725 16475
rect -3755 16450 -3750 16470
rect -3750 16450 -3730 16470
rect -3730 16450 -3725 16470
rect -3755 16445 -3725 16450
rect -3675 16470 -3645 16475
rect -3675 16450 -3670 16470
rect -3670 16450 -3650 16470
rect -3650 16450 -3645 16470
rect -3675 16445 -3645 16450
rect -3595 16470 -3565 16475
rect -3595 16450 -3590 16470
rect -3590 16450 -3570 16470
rect -3570 16450 -3565 16470
rect -3595 16445 -3565 16450
rect -3515 16470 -3485 16475
rect -3515 16450 -3510 16470
rect -3510 16450 -3490 16470
rect -3490 16450 -3485 16470
rect -3515 16445 -3485 16450
rect -3435 16470 -3405 16475
rect -3435 16450 -3430 16470
rect -3430 16450 -3410 16470
rect -3410 16450 -3405 16470
rect -3435 16445 -3405 16450
rect -3355 16470 -3325 16475
rect -3355 16450 -3350 16470
rect -3350 16450 -3330 16470
rect -3330 16450 -3325 16470
rect -3355 16445 -3325 16450
rect -3275 16470 -3245 16475
rect -3275 16450 -3270 16470
rect -3270 16450 -3250 16470
rect -3250 16450 -3245 16470
rect -3275 16445 -3245 16450
rect -3195 16470 -3165 16475
rect -3195 16450 -3190 16470
rect -3190 16450 -3170 16470
rect -3170 16450 -3165 16470
rect -3195 16445 -3165 16450
rect -3115 16470 -3085 16475
rect -3115 16450 -3110 16470
rect -3110 16450 -3090 16470
rect -3090 16450 -3085 16470
rect -3115 16445 -3085 16450
rect -3035 16470 -3005 16475
rect -3035 16450 -3030 16470
rect -3030 16450 -3010 16470
rect -3010 16450 -3005 16470
rect -3035 16445 -3005 16450
rect -2955 16470 -2925 16475
rect -2955 16450 -2950 16470
rect -2950 16450 -2930 16470
rect -2930 16450 -2925 16470
rect -2955 16445 -2925 16450
rect -2875 16470 -2845 16475
rect -2875 16450 -2870 16470
rect -2870 16450 -2850 16470
rect -2850 16450 -2845 16470
rect -2875 16445 -2845 16450
rect -2795 16470 -2765 16475
rect -2795 16450 -2790 16470
rect -2790 16450 -2770 16470
rect -2770 16450 -2765 16470
rect -2795 16445 -2765 16450
rect -2715 16470 -2685 16475
rect -2715 16450 -2710 16470
rect -2710 16450 -2690 16470
rect -2690 16450 -2685 16470
rect -2715 16445 -2685 16450
rect -2635 16470 -2605 16475
rect -2635 16450 -2630 16470
rect -2630 16450 -2610 16470
rect -2610 16450 -2605 16470
rect -2635 16445 -2605 16450
rect -2555 16470 -2525 16475
rect -2555 16450 -2550 16470
rect -2550 16450 -2530 16470
rect -2530 16450 -2525 16470
rect -2555 16445 -2525 16450
rect -2475 16470 -2445 16475
rect -2475 16450 -2470 16470
rect -2470 16450 -2450 16470
rect -2450 16450 -2445 16470
rect -2475 16445 -2445 16450
rect -2395 16470 -2365 16475
rect -2395 16450 -2390 16470
rect -2390 16450 -2370 16470
rect -2370 16450 -2365 16470
rect -2395 16445 -2365 16450
rect -2315 16470 -2285 16475
rect -2315 16450 -2310 16470
rect -2310 16450 -2290 16470
rect -2290 16450 -2285 16470
rect -2315 16445 -2285 16450
rect -2235 16470 -2205 16475
rect -2235 16450 -2230 16470
rect -2230 16450 -2210 16470
rect -2210 16450 -2205 16470
rect -2235 16445 -2205 16450
rect -2155 16470 -2125 16475
rect -2155 16450 -2150 16470
rect -2150 16450 -2130 16470
rect -2130 16450 -2125 16470
rect -2155 16445 -2125 16450
rect -2075 16470 -2045 16475
rect -2075 16450 -2070 16470
rect -2070 16450 -2050 16470
rect -2050 16450 -2045 16470
rect -2075 16445 -2045 16450
rect -1995 16470 -1965 16475
rect -1995 16450 -1990 16470
rect -1990 16450 -1970 16470
rect -1970 16450 -1965 16470
rect -1995 16445 -1965 16450
rect -1835 16470 -1805 16475
rect -1835 16450 -1830 16470
rect -1830 16450 -1810 16470
rect -1810 16450 -1805 16470
rect -1835 16445 -1805 16450
rect -1755 16470 -1725 16475
rect -1755 16450 -1750 16470
rect -1750 16450 -1730 16470
rect -1730 16450 -1725 16470
rect -1755 16445 -1725 16450
rect -1675 16470 -1645 16475
rect -1675 16450 -1670 16470
rect -1670 16450 -1650 16470
rect -1650 16450 -1645 16470
rect -1675 16445 -1645 16450
rect -1595 16470 -1565 16475
rect -1595 16450 -1590 16470
rect -1590 16450 -1570 16470
rect -1570 16450 -1565 16470
rect -1595 16445 -1565 16450
rect -1515 16470 -1485 16475
rect -1515 16450 -1510 16470
rect -1510 16450 -1490 16470
rect -1490 16450 -1485 16470
rect -1515 16445 -1485 16450
rect -1435 16470 -1405 16475
rect -1435 16450 -1430 16470
rect -1430 16450 -1410 16470
rect -1410 16450 -1405 16470
rect -1435 16445 -1405 16450
rect -1355 16470 -1325 16475
rect -1355 16450 -1350 16470
rect -1350 16450 -1330 16470
rect -1330 16450 -1325 16470
rect -1355 16445 -1325 16450
rect -1195 16470 -1165 16475
rect -1195 16450 -1190 16470
rect -1190 16450 -1170 16470
rect -1170 16450 -1165 16470
rect -1195 16445 -1165 16450
rect -1035 16470 -1005 16475
rect -1035 16450 -1030 16470
rect -1030 16450 -1010 16470
rect -1010 16450 -1005 16470
rect -1035 16445 -1005 16450
rect -875 16470 -845 16475
rect -875 16450 -870 16470
rect -870 16450 -850 16470
rect -850 16450 -845 16470
rect -875 16445 -845 16450
rect -715 16470 -685 16475
rect -715 16450 -710 16470
rect -710 16450 -690 16470
rect -690 16450 -685 16470
rect -715 16445 -685 16450
rect -555 16470 -525 16475
rect -555 16450 -550 16470
rect -550 16450 -530 16470
rect -530 16450 -525 16470
rect -555 16445 -525 16450
rect -14955 16310 -14925 16315
rect -14955 16290 -14950 16310
rect -14950 16290 -14930 16310
rect -14930 16290 -14925 16310
rect -14955 16285 -14925 16290
rect -14875 16310 -14845 16315
rect -14875 16290 -14870 16310
rect -14870 16290 -14850 16310
rect -14850 16290 -14845 16310
rect -14875 16285 -14845 16290
rect -14795 16310 -14765 16315
rect -14795 16290 -14790 16310
rect -14790 16290 -14770 16310
rect -14770 16290 -14765 16310
rect -14795 16285 -14765 16290
rect -14715 16310 -14685 16315
rect -14715 16290 -14710 16310
rect -14710 16290 -14690 16310
rect -14690 16290 -14685 16310
rect -14715 16285 -14685 16290
rect -14635 16310 -14605 16315
rect -14635 16290 -14630 16310
rect -14630 16290 -14610 16310
rect -14610 16290 -14605 16310
rect -14635 16285 -14605 16290
rect -14555 16310 -14525 16315
rect -14555 16290 -14550 16310
rect -14550 16290 -14530 16310
rect -14530 16290 -14525 16310
rect -14555 16285 -14525 16290
rect -14475 16310 -14445 16315
rect -14475 16290 -14470 16310
rect -14470 16290 -14450 16310
rect -14450 16290 -14445 16310
rect -14475 16285 -14445 16290
rect -14395 16310 -14365 16315
rect -14395 16290 -14390 16310
rect -14390 16290 -14370 16310
rect -14370 16290 -14365 16310
rect -14395 16285 -14365 16290
rect -14315 16310 -14285 16315
rect -14315 16290 -14310 16310
rect -14310 16290 -14290 16310
rect -14290 16290 -14285 16310
rect -14315 16285 -14285 16290
rect -14235 16310 -14205 16315
rect -14235 16290 -14230 16310
rect -14230 16290 -14210 16310
rect -14210 16290 -14205 16310
rect -14235 16285 -14205 16290
rect -14155 16310 -14125 16315
rect -14155 16290 -14150 16310
rect -14150 16290 -14130 16310
rect -14130 16290 -14125 16310
rect -14155 16285 -14125 16290
rect -14075 16310 -14045 16315
rect -14075 16290 -14070 16310
rect -14070 16290 -14050 16310
rect -14050 16290 -14045 16310
rect -14075 16285 -14045 16290
rect -13995 16310 -13965 16315
rect -13995 16290 -13990 16310
rect -13990 16290 -13970 16310
rect -13970 16290 -13965 16310
rect -13995 16285 -13965 16290
rect -13915 16310 -13885 16315
rect -13915 16290 -13910 16310
rect -13910 16290 -13890 16310
rect -13890 16290 -13885 16310
rect -13915 16285 -13885 16290
rect -13835 16310 -13805 16315
rect -13835 16290 -13830 16310
rect -13830 16290 -13810 16310
rect -13810 16290 -13805 16310
rect -13835 16285 -13805 16290
rect -13755 16310 -13725 16315
rect -13755 16290 -13750 16310
rect -13750 16290 -13730 16310
rect -13730 16290 -13725 16310
rect -13755 16285 -13725 16290
rect -13675 16310 -13645 16315
rect -13675 16290 -13670 16310
rect -13670 16290 -13650 16310
rect -13650 16290 -13645 16310
rect -13675 16285 -13645 16290
rect -13595 16310 -13565 16315
rect -13595 16290 -13590 16310
rect -13590 16290 -13570 16310
rect -13570 16290 -13565 16310
rect -13595 16285 -13565 16290
rect -13515 16310 -13485 16315
rect -13515 16290 -13510 16310
rect -13510 16290 -13490 16310
rect -13490 16290 -13485 16310
rect -13515 16285 -13485 16290
rect -13435 16310 -13405 16315
rect -13435 16290 -13430 16310
rect -13430 16290 -13410 16310
rect -13410 16290 -13405 16310
rect -13435 16285 -13405 16290
rect -13355 16310 -13325 16315
rect -13355 16290 -13350 16310
rect -13350 16290 -13330 16310
rect -13330 16290 -13325 16310
rect -13355 16285 -13325 16290
rect -13275 16310 -13245 16315
rect -13275 16290 -13270 16310
rect -13270 16290 -13250 16310
rect -13250 16290 -13245 16310
rect -13275 16285 -13245 16290
rect -13195 16310 -13165 16315
rect -13195 16290 -13190 16310
rect -13190 16290 -13170 16310
rect -13170 16290 -13165 16310
rect -13195 16285 -13165 16290
rect -13115 16310 -13085 16315
rect -13115 16290 -13110 16310
rect -13110 16290 -13090 16310
rect -13090 16290 -13085 16310
rect -13115 16285 -13085 16290
rect -13035 16310 -13005 16315
rect -13035 16290 -13030 16310
rect -13030 16290 -13010 16310
rect -13010 16290 -13005 16310
rect -13035 16285 -13005 16290
rect -12955 16310 -12925 16315
rect -12955 16290 -12950 16310
rect -12950 16290 -12930 16310
rect -12930 16290 -12925 16310
rect -12955 16285 -12925 16290
rect -12875 16310 -12845 16315
rect -12875 16290 -12870 16310
rect -12870 16290 -12850 16310
rect -12850 16290 -12845 16310
rect -12875 16285 -12845 16290
rect -12795 16310 -12765 16315
rect -12795 16290 -12790 16310
rect -12790 16290 -12770 16310
rect -12770 16290 -12765 16310
rect -12795 16285 -12765 16290
rect -12715 16310 -12685 16315
rect -12715 16290 -12710 16310
rect -12710 16290 -12690 16310
rect -12690 16290 -12685 16310
rect -12715 16285 -12685 16290
rect -12635 16310 -12605 16315
rect -12635 16290 -12630 16310
rect -12630 16290 -12610 16310
rect -12610 16290 -12605 16310
rect -12635 16285 -12605 16290
rect -12555 16310 -12525 16315
rect -12555 16290 -12550 16310
rect -12550 16290 -12530 16310
rect -12530 16290 -12525 16310
rect -12555 16285 -12525 16290
rect -12475 16310 -12445 16315
rect -12475 16290 -12470 16310
rect -12470 16290 -12450 16310
rect -12450 16290 -12445 16310
rect -12475 16285 -12445 16290
rect -12395 16310 -12365 16315
rect -12395 16290 -12390 16310
rect -12390 16290 -12370 16310
rect -12370 16290 -12365 16310
rect -12395 16285 -12365 16290
rect -12315 16310 -12285 16315
rect -12315 16290 -12310 16310
rect -12310 16290 -12290 16310
rect -12290 16290 -12285 16310
rect -12315 16285 -12285 16290
rect -12235 16310 -12205 16315
rect -12235 16290 -12230 16310
rect -12230 16290 -12210 16310
rect -12210 16290 -12205 16310
rect -12235 16285 -12205 16290
rect -12155 16310 -12125 16315
rect -12155 16290 -12150 16310
rect -12150 16290 -12130 16310
rect -12130 16290 -12125 16310
rect -12155 16285 -12125 16290
rect -12075 16310 -12045 16315
rect -12075 16290 -12070 16310
rect -12070 16290 -12050 16310
rect -12050 16290 -12045 16310
rect -12075 16285 -12045 16290
rect -11995 16310 -11965 16315
rect -11995 16290 -11990 16310
rect -11990 16290 -11970 16310
rect -11970 16290 -11965 16310
rect -11995 16285 -11965 16290
rect -11915 16310 -11885 16315
rect -11915 16290 -11910 16310
rect -11910 16290 -11890 16310
rect -11890 16290 -11885 16310
rect -11915 16285 -11885 16290
rect -11835 16310 -11805 16315
rect -11835 16290 -11830 16310
rect -11830 16290 -11810 16310
rect -11810 16290 -11805 16310
rect -11835 16285 -11805 16290
rect -11755 16310 -11725 16315
rect -11755 16290 -11750 16310
rect -11750 16290 -11730 16310
rect -11730 16290 -11725 16310
rect -11755 16285 -11725 16290
rect -11675 16310 -11645 16315
rect -11675 16290 -11670 16310
rect -11670 16290 -11650 16310
rect -11650 16290 -11645 16310
rect -11675 16285 -11645 16290
rect -11595 16310 -11565 16315
rect -11595 16290 -11590 16310
rect -11590 16290 -11570 16310
rect -11570 16290 -11565 16310
rect -11595 16285 -11565 16290
rect -11515 16310 -11485 16315
rect -11515 16290 -11510 16310
rect -11510 16290 -11490 16310
rect -11490 16290 -11485 16310
rect -11515 16285 -11485 16290
rect -11435 16310 -11405 16315
rect -11435 16290 -11430 16310
rect -11430 16290 -11410 16310
rect -11410 16290 -11405 16310
rect -11435 16285 -11405 16290
rect -11355 16310 -11325 16315
rect -11355 16290 -11350 16310
rect -11350 16290 -11330 16310
rect -11330 16290 -11325 16310
rect -11355 16285 -11325 16290
rect -11275 16310 -11245 16315
rect -11275 16290 -11270 16310
rect -11270 16290 -11250 16310
rect -11250 16290 -11245 16310
rect -11275 16285 -11245 16290
rect -11195 16310 -11165 16315
rect -11195 16290 -11190 16310
rect -11190 16290 -11170 16310
rect -11170 16290 -11165 16310
rect -11195 16285 -11165 16290
rect -11115 16310 -11085 16315
rect -11115 16290 -11110 16310
rect -11110 16290 -11090 16310
rect -11090 16290 -11085 16310
rect -11115 16285 -11085 16290
rect -11035 16310 -11005 16315
rect -11035 16290 -11030 16310
rect -11030 16290 -11010 16310
rect -11010 16290 -11005 16310
rect -11035 16285 -11005 16290
rect -10955 16310 -10925 16315
rect -10955 16290 -10950 16310
rect -10950 16290 -10930 16310
rect -10930 16290 -10925 16310
rect -10955 16285 -10925 16290
rect -10875 16310 -10845 16315
rect -10875 16290 -10870 16310
rect -10870 16290 -10850 16310
rect -10850 16290 -10845 16310
rect -10875 16285 -10845 16290
rect -10795 16310 -10765 16315
rect -10795 16290 -10790 16310
rect -10790 16290 -10770 16310
rect -10770 16290 -10765 16310
rect -10795 16285 -10765 16290
rect -10715 16310 -10685 16315
rect -10715 16290 -10710 16310
rect -10710 16290 -10690 16310
rect -10690 16290 -10685 16310
rect -10715 16285 -10685 16290
rect -10635 16310 -10605 16315
rect -10635 16290 -10630 16310
rect -10630 16290 -10610 16310
rect -10610 16290 -10605 16310
rect -10635 16285 -10605 16290
rect -10555 16310 -10525 16315
rect -10555 16290 -10550 16310
rect -10550 16290 -10530 16310
rect -10530 16290 -10525 16310
rect -10555 16285 -10525 16290
rect -10475 16310 -10445 16315
rect -10475 16290 -10470 16310
rect -10470 16290 -10450 16310
rect -10450 16290 -10445 16310
rect -10475 16285 -10445 16290
rect -10395 16310 -10365 16315
rect -10395 16290 -10390 16310
rect -10390 16290 -10370 16310
rect -10370 16290 -10365 16310
rect -10395 16285 -10365 16290
rect -10315 16310 -10285 16315
rect -10315 16290 -10310 16310
rect -10310 16290 -10290 16310
rect -10290 16290 -10285 16310
rect -10315 16285 -10285 16290
rect -10235 16310 -10205 16315
rect -10235 16290 -10230 16310
rect -10230 16290 -10210 16310
rect -10210 16290 -10205 16310
rect -10235 16285 -10205 16290
rect -10155 16310 -10125 16315
rect -10155 16290 -10150 16310
rect -10150 16290 -10130 16310
rect -10130 16290 -10125 16310
rect -10155 16285 -10125 16290
rect -10075 16310 -10045 16315
rect -10075 16290 -10070 16310
rect -10070 16290 -10050 16310
rect -10050 16290 -10045 16310
rect -10075 16285 -10045 16290
rect -9995 16310 -9965 16315
rect -9995 16290 -9990 16310
rect -9990 16290 -9970 16310
rect -9970 16290 -9965 16310
rect -9995 16285 -9965 16290
rect -9915 16310 -9885 16315
rect -9915 16290 -9910 16310
rect -9910 16290 -9890 16310
rect -9890 16290 -9885 16310
rect -9915 16285 -9885 16290
rect -9835 16310 -9805 16315
rect -9835 16290 -9830 16310
rect -9830 16290 -9810 16310
rect -9810 16290 -9805 16310
rect -9835 16285 -9805 16290
rect -9755 16310 -9725 16315
rect -9755 16290 -9750 16310
rect -9750 16290 -9730 16310
rect -9730 16290 -9725 16310
rect -9755 16285 -9725 16290
rect -9675 16310 -9645 16315
rect -9675 16290 -9670 16310
rect -9670 16290 -9650 16310
rect -9650 16290 -9645 16310
rect -9675 16285 -9645 16290
rect -9595 16310 -9565 16315
rect -9595 16290 -9590 16310
rect -9590 16290 -9570 16310
rect -9570 16290 -9565 16310
rect -9595 16285 -9565 16290
rect -9515 16310 -9485 16315
rect -9515 16290 -9510 16310
rect -9510 16290 -9490 16310
rect -9490 16290 -9485 16310
rect -9515 16285 -9485 16290
rect -9435 16310 -9405 16315
rect -9435 16290 -9430 16310
rect -9430 16290 -9410 16310
rect -9410 16290 -9405 16310
rect -9435 16285 -9405 16290
rect -9355 16310 -9325 16315
rect -9355 16290 -9350 16310
rect -9350 16290 -9330 16310
rect -9330 16290 -9325 16310
rect -9355 16285 -9325 16290
rect -9275 16310 -9245 16315
rect -9275 16290 -9270 16310
rect -9270 16290 -9250 16310
rect -9250 16290 -9245 16310
rect -9275 16285 -9245 16290
rect -9195 16310 -9165 16315
rect -9195 16290 -9190 16310
rect -9190 16290 -9170 16310
rect -9170 16290 -9165 16310
rect -9195 16285 -9165 16290
rect -9115 16310 -9085 16315
rect -9115 16290 -9110 16310
rect -9110 16290 -9090 16310
rect -9090 16290 -9085 16310
rect -9115 16285 -9085 16290
rect -9035 16310 -9005 16315
rect -9035 16290 -9030 16310
rect -9030 16290 -9010 16310
rect -9010 16290 -9005 16310
rect -9035 16285 -9005 16290
rect -8955 16310 -8925 16315
rect -8955 16290 -8950 16310
rect -8950 16290 -8930 16310
rect -8930 16290 -8925 16310
rect -8955 16285 -8925 16290
rect -8875 16310 -8845 16315
rect -8875 16290 -8870 16310
rect -8870 16290 -8850 16310
rect -8850 16290 -8845 16310
rect -8875 16285 -8845 16290
rect -8795 16310 -8765 16315
rect -8795 16290 -8790 16310
rect -8790 16290 -8770 16310
rect -8770 16290 -8765 16310
rect -8795 16285 -8765 16290
rect -8715 16310 -8685 16315
rect -8715 16290 -8710 16310
rect -8710 16290 -8690 16310
rect -8690 16290 -8685 16310
rect -8715 16285 -8685 16290
rect -8635 16310 -8605 16315
rect -8635 16290 -8630 16310
rect -8630 16290 -8610 16310
rect -8610 16290 -8605 16310
rect -8635 16285 -8605 16290
rect -8555 16310 -8525 16315
rect -8555 16290 -8550 16310
rect -8550 16290 -8530 16310
rect -8530 16290 -8525 16310
rect -8555 16285 -8525 16290
rect -8475 16310 -8445 16315
rect -8475 16290 -8470 16310
rect -8470 16290 -8450 16310
rect -8450 16290 -8445 16310
rect -8475 16285 -8445 16290
rect -8395 16310 -8365 16315
rect -8395 16290 -8390 16310
rect -8390 16290 -8370 16310
rect -8370 16290 -8365 16310
rect -8395 16285 -8365 16290
rect -8315 16310 -8285 16315
rect -8315 16290 -8310 16310
rect -8310 16290 -8290 16310
rect -8290 16290 -8285 16310
rect -8315 16285 -8285 16290
rect -8235 16310 -8205 16315
rect -8235 16290 -8230 16310
rect -8230 16290 -8210 16310
rect -8210 16290 -8205 16310
rect -8235 16285 -8205 16290
rect -8155 16310 -8125 16315
rect -8155 16290 -8150 16310
rect -8150 16290 -8130 16310
rect -8130 16290 -8125 16310
rect -8155 16285 -8125 16290
rect -8075 16310 -8045 16315
rect -8075 16290 -8070 16310
rect -8070 16290 -8050 16310
rect -8050 16290 -8045 16310
rect -8075 16285 -8045 16290
rect -7995 16310 -7965 16315
rect -7995 16290 -7990 16310
rect -7990 16290 -7970 16310
rect -7970 16290 -7965 16310
rect -7995 16285 -7965 16290
rect -7915 16310 -7885 16315
rect -7915 16290 -7910 16310
rect -7910 16290 -7890 16310
rect -7890 16290 -7885 16310
rect -7915 16285 -7885 16290
rect -7835 16310 -7805 16315
rect -7835 16290 -7830 16310
rect -7830 16290 -7810 16310
rect -7810 16290 -7805 16310
rect -7835 16285 -7805 16290
rect -7755 16310 -7725 16315
rect -7755 16290 -7750 16310
rect -7750 16290 -7730 16310
rect -7730 16290 -7725 16310
rect -7755 16285 -7725 16290
rect -7675 16310 -7645 16315
rect -7675 16290 -7670 16310
rect -7670 16290 -7650 16310
rect -7650 16290 -7645 16310
rect -7675 16285 -7645 16290
rect -7595 16310 -7565 16315
rect -7595 16290 -7590 16310
rect -7590 16290 -7570 16310
rect -7570 16290 -7565 16310
rect -7595 16285 -7565 16290
rect -7515 16310 -7485 16315
rect -7515 16290 -7510 16310
rect -7510 16290 -7490 16310
rect -7490 16290 -7485 16310
rect -7515 16285 -7485 16290
rect -7435 16310 -7405 16315
rect -7435 16290 -7430 16310
rect -7430 16290 -7410 16310
rect -7410 16290 -7405 16310
rect -7435 16285 -7405 16290
rect -7355 16310 -7325 16315
rect -7355 16290 -7350 16310
rect -7350 16290 -7330 16310
rect -7330 16290 -7325 16310
rect -7355 16285 -7325 16290
rect -7275 16310 -7245 16315
rect -7275 16290 -7270 16310
rect -7270 16290 -7250 16310
rect -7250 16290 -7245 16310
rect -7275 16285 -7245 16290
rect -7195 16310 -7165 16315
rect -7195 16290 -7190 16310
rect -7190 16290 -7170 16310
rect -7170 16290 -7165 16310
rect -7195 16285 -7165 16290
rect -7115 16310 -7085 16315
rect -7115 16290 -7110 16310
rect -7110 16290 -7090 16310
rect -7090 16290 -7085 16310
rect -7115 16285 -7085 16290
rect -7035 16310 -7005 16315
rect -7035 16290 -7030 16310
rect -7030 16290 -7010 16310
rect -7010 16290 -7005 16310
rect -7035 16285 -7005 16290
rect -6955 16310 -6925 16315
rect -6955 16290 -6950 16310
rect -6950 16290 -6930 16310
rect -6930 16290 -6925 16310
rect -6955 16285 -6925 16290
rect -6875 16310 -6845 16315
rect -6875 16290 -6870 16310
rect -6870 16290 -6850 16310
rect -6850 16290 -6845 16310
rect -6875 16285 -6845 16290
rect -6795 16310 -6765 16315
rect -6795 16290 -6790 16310
rect -6790 16290 -6770 16310
rect -6770 16290 -6765 16310
rect -6795 16285 -6765 16290
rect -6715 16310 -6685 16315
rect -6715 16290 -6710 16310
rect -6710 16290 -6690 16310
rect -6690 16290 -6685 16310
rect -6715 16285 -6685 16290
rect -6635 16310 -6605 16315
rect -6635 16290 -6630 16310
rect -6630 16290 -6610 16310
rect -6610 16290 -6605 16310
rect -6635 16285 -6605 16290
rect -6555 16310 -6525 16315
rect -6555 16290 -6550 16310
rect -6550 16290 -6530 16310
rect -6530 16290 -6525 16310
rect -6555 16285 -6525 16290
rect -6475 16310 -6445 16315
rect -6475 16290 -6470 16310
rect -6470 16290 -6450 16310
rect -6450 16290 -6445 16310
rect -6475 16285 -6445 16290
rect -6395 16310 -6365 16315
rect -6395 16290 -6390 16310
rect -6390 16290 -6370 16310
rect -6370 16290 -6365 16310
rect -6395 16285 -6365 16290
rect -6315 16310 -6285 16315
rect -6315 16290 -6310 16310
rect -6310 16290 -6290 16310
rect -6290 16290 -6285 16310
rect -6315 16285 -6285 16290
rect -6235 16310 -6205 16315
rect -6235 16290 -6230 16310
rect -6230 16290 -6210 16310
rect -6210 16290 -6205 16310
rect -6235 16285 -6205 16290
rect -6155 16310 -6125 16315
rect -6155 16290 -6150 16310
rect -6150 16290 -6130 16310
rect -6130 16290 -6125 16310
rect -6155 16285 -6125 16290
rect -6075 16310 -6045 16315
rect -6075 16290 -6070 16310
rect -6070 16290 -6050 16310
rect -6050 16290 -6045 16310
rect -6075 16285 -6045 16290
rect -5995 16310 -5965 16315
rect -5995 16290 -5990 16310
rect -5990 16290 -5970 16310
rect -5970 16290 -5965 16310
rect -5995 16285 -5965 16290
rect -5915 16310 -5885 16315
rect -5915 16290 -5910 16310
rect -5910 16290 -5890 16310
rect -5890 16290 -5885 16310
rect -5915 16285 -5885 16290
rect -5835 16310 -5805 16315
rect -5835 16290 -5830 16310
rect -5830 16290 -5810 16310
rect -5810 16290 -5805 16310
rect -5835 16285 -5805 16290
rect -5755 16310 -5725 16315
rect -5755 16290 -5750 16310
rect -5750 16290 -5730 16310
rect -5730 16290 -5725 16310
rect -5755 16285 -5725 16290
rect -5595 16310 -5565 16315
rect -5595 16290 -5590 16310
rect -5590 16290 -5570 16310
rect -5570 16290 -5565 16310
rect -5595 16285 -5565 16290
rect -5435 16310 -5405 16315
rect -5435 16290 -5430 16310
rect -5430 16290 -5410 16310
rect -5410 16290 -5405 16310
rect -5435 16285 -5405 16290
rect -5355 16310 -5325 16315
rect -5355 16290 -5350 16310
rect -5350 16290 -5330 16310
rect -5330 16290 -5325 16310
rect -5355 16285 -5325 16290
rect -5275 16310 -5245 16315
rect -5275 16290 -5270 16310
rect -5270 16290 -5250 16310
rect -5250 16290 -5245 16310
rect -5275 16285 -5245 16290
rect -5195 16310 -5165 16315
rect -5195 16290 -5190 16310
rect -5190 16290 -5170 16310
rect -5170 16290 -5165 16310
rect -5195 16285 -5165 16290
rect -5115 16310 -5085 16315
rect -5115 16290 -5110 16310
rect -5110 16290 -5090 16310
rect -5090 16290 -5085 16310
rect -5115 16285 -5085 16290
rect -5035 16310 -5005 16315
rect -5035 16290 -5030 16310
rect -5030 16290 -5010 16310
rect -5010 16290 -5005 16310
rect -5035 16285 -5005 16290
rect -4955 16310 -4925 16315
rect -4955 16290 -4950 16310
rect -4950 16290 -4930 16310
rect -4930 16290 -4925 16310
rect -4955 16285 -4925 16290
rect -4875 16310 -4845 16315
rect -4875 16290 -4870 16310
rect -4870 16290 -4850 16310
rect -4850 16290 -4845 16310
rect -4875 16285 -4845 16290
rect -4795 16310 -4765 16315
rect -4795 16290 -4790 16310
rect -4790 16290 -4770 16310
rect -4770 16290 -4765 16310
rect -4795 16285 -4765 16290
rect -4715 16310 -4685 16315
rect -4715 16290 -4710 16310
rect -4710 16290 -4690 16310
rect -4690 16290 -4685 16310
rect -4715 16285 -4685 16290
rect -4635 16310 -4605 16315
rect -4635 16290 -4630 16310
rect -4630 16290 -4610 16310
rect -4610 16290 -4605 16310
rect -4635 16285 -4605 16290
rect -4555 16310 -4525 16315
rect -4555 16290 -4550 16310
rect -4550 16290 -4530 16310
rect -4530 16290 -4525 16310
rect -4555 16285 -4525 16290
rect -4475 16310 -4445 16315
rect -4475 16290 -4470 16310
rect -4470 16290 -4450 16310
rect -4450 16290 -4445 16310
rect -4475 16285 -4445 16290
rect -4395 16310 -4365 16315
rect -4395 16290 -4390 16310
rect -4390 16290 -4370 16310
rect -4370 16290 -4365 16310
rect -4395 16285 -4365 16290
rect -4315 16310 -4285 16315
rect -4315 16290 -4310 16310
rect -4310 16290 -4290 16310
rect -4290 16290 -4285 16310
rect -4315 16285 -4285 16290
rect -4235 16310 -4205 16315
rect -4235 16290 -4230 16310
rect -4230 16290 -4210 16310
rect -4210 16290 -4205 16310
rect -4235 16285 -4205 16290
rect -4155 16310 -4125 16315
rect -4155 16290 -4150 16310
rect -4150 16290 -4130 16310
rect -4130 16290 -4125 16310
rect -4155 16285 -4125 16290
rect -4075 16310 -4045 16315
rect -4075 16290 -4070 16310
rect -4070 16290 -4050 16310
rect -4050 16290 -4045 16310
rect -4075 16285 -4045 16290
rect -3995 16310 -3965 16315
rect -3995 16290 -3990 16310
rect -3990 16290 -3970 16310
rect -3970 16290 -3965 16310
rect -3995 16285 -3965 16290
rect -3915 16310 -3885 16315
rect -3915 16290 -3910 16310
rect -3910 16290 -3890 16310
rect -3890 16290 -3885 16310
rect -3915 16285 -3885 16290
rect -3835 16310 -3805 16315
rect -3835 16290 -3830 16310
rect -3830 16290 -3810 16310
rect -3810 16290 -3805 16310
rect -3835 16285 -3805 16290
rect -3755 16310 -3725 16315
rect -3755 16290 -3750 16310
rect -3750 16290 -3730 16310
rect -3730 16290 -3725 16310
rect -3755 16285 -3725 16290
rect -3675 16310 -3645 16315
rect -3675 16290 -3670 16310
rect -3670 16290 -3650 16310
rect -3650 16290 -3645 16310
rect -3675 16285 -3645 16290
rect -3595 16310 -3565 16315
rect -3595 16290 -3590 16310
rect -3590 16290 -3570 16310
rect -3570 16290 -3565 16310
rect -3595 16285 -3565 16290
rect -3515 16310 -3485 16315
rect -3515 16290 -3510 16310
rect -3510 16290 -3490 16310
rect -3490 16290 -3485 16310
rect -3515 16285 -3485 16290
rect -3435 16310 -3405 16315
rect -3435 16290 -3430 16310
rect -3430 16290 -3410 16310
rect -3410 16290 -3405 16310
rect -3435 16285 -3405 16290
rect -3355 16310 -3325 16315
rect -3355 16290 -3350 16310
rect -3350 16290 -3330 16310
rect -3330 16290 -3325 16310
rect -3355 16285 -3325 16290
rect -3275 16310 -3245 16315
rect -3275 16290 -3270 16310
rect -3270 16290 -3250 16310
rect -3250 16290 -3245 16310
rect -3275 16285 -3245 16290
rect -3195 16310 -3165 16315
rect -3195 16290 -3190 16310
rect -3190 16290 -3170 16310
rect -3170 16290 -3165 16310
rect -3195 16285 -3165 16290
rect -3115 16310 -3085 16315
rect -3115 16290 -3110 16310
rect -3110 16290 -3090 16310
rect -3090 16290 -3085 16310
rect -3115 16285 -3085 16290
rect -3035 16310 -3005 16315
rect -3035 16290 -3030 16310
rect -3030 16290 -3010 16310
rect -3010 16290 -3005 16310
rect -3035 16285 -3005 16290
rect -2955 16310 -2925 16315
rect -2955 16290 -2950 16310
rect -2950 16290 -2930 16310
rect -2930 16290 -2925 16310
rect -2955 16285 -2925 16290
rect -2875 16310 -2845 16315
rect -2875 16290 -2870 16310
rect -2870 16290 -2850 16310
rect -2850 16290 -2845 16310
rect -2875 16285 -2845 16290
rect -2795 16310 -2765 16315
rect -2795 16290 -2790 16310
rect -2790 16290 -2770 16310
rect -2770 16290 -2765 16310
rect -2795 16285 -2765 16290
rect -2715 16310 -2685 16315
rect -2715 16290 -2710 16310
rect -2710 16290 -2690 16310
rect -2690 16290 -2685 16310
rect -2715 16285 -2685 16290
rect -2635 16310 -2605 16315
rect -2635 16290 -2630 16310
rect -2630 16290 -2610 16310
rect -2610 16290 -2605 16310
rect -2635 16285 -2605 16290
rect -2555 16310 -2525 16315
rect -2555 16290 -2550 16310
rect -2550 16290 -2530 16310
rect -2530 16290 -2525 16310
rect -2555 16285 -2525 16290
rect -2475 16310 -2445 16315
rect -2475 16290 -2470 16310
rect -2470 16290 -2450 16310
rect -2450 16290 -2445 16310
rect -2475 16285 -2445 16290
rect -2395 16310 -2365 16315
rect -2395 16290 -2390 16310
rect -2390 16290 -2370 16310
rect -2370 16290 -2365 16310
rect -2395 16285 -2365 16290
rect -2315 16310 -2285 16315
rect -2315 16290 -2310 16310
rect -2310 16290 -2290 16310
rect -2290 16290 -2285 16310
rect -2315 16285 -2285 16290
rect -2235 16310 -2205 16315
rect -2235 16290 -2230 16310
rect -2230 16290 -2210 16310
rect -2210 16290 -2205 16310
rect -2235 16285 -2205 16290
rect -2155 16310 -2125 16315
rect -2155 16290 -2150 16310
rect -2150 16290 -2130 16310
rect -2130 16290 -2125 16310
rect -2155 16285 -2125 16290
rect -2075 16310 -2045 16315
rect -2075 16290 -2070 16310
rect -2070 16290 -2050 16310
rect -2050 16290 -2045 16310
rect -2075 16285 -2045 16290
rect -1995 16310 -1965 16315
rect -1995 16290 -1990 16310
rect -1990 16290 -1970 16310
rect -1970 16290 -1965 16310
rect -1995 16285 -1965 16290
rect -1835 16310 -1805 16315
rect -1835 16290 -1830 16310
rect -1830 16290 -1810 16310
rect -1810 16290 -1805 16310
rect -1835 16285 -1805 16290
rect -1755 16310 -1725 16315
rect -1755 16290 -1750 16310
rect -1750 16290 -1730 16310
rect -1730 16290 -1725 16310
rect -1755 16285 -1725 16290
rect -1675 16310 -1645 16315
rect -1675 16290 -1670 16310
rect -1670 16290 -1650 16310
rect -1650 16290 -1645 16310
rect -1675 16285 -1645 16290
rect -1595 16310 -1565 16315
rect -1595 16290 -1590 16310
rect -1590 16290 -1570 16310
rect -1570 16290 -1565 16310
rect -1595 16285 -1565 16290
rect -1515 16310 -1485 16315
rect -1515 16290 -1510 16310
rect -1510 16290 -1490 16310
rect -1490 16290 -1485 16310
rect -1515 16285 -1485 16290
rect -1435 16310 -1405 16315
rect -1435 16290 -1430 16310
rect -1430 16290 -1410 16310
rect -1410 16290 -1405 16310
rect -1435 16285 -1405 16290
rect -1355 16310 -1325 16315
rect -1355 16290 -1350 16310
rect -1350 16290 -1330 16310
rect -1330 16290 -1325 16310
rect -1355 16285 -1325 16290
rect -1195 16310 -1165 16315
rect -1195 16290 -1190 16310
rect -1190 16290 -1170 16310
rect -1170 16290 -1165 16310
rect -1195 16285 -1165 16290
rect -1035 16310 -1005 16315
rect -1035 16290 -1030 16310
rect -1030 16290 -1010 16310
rect -1010 16290 -1005 16310
rect -1035 16285 -1005 16290
rect -875 16310 -845 16315
rect -875 16290 -870 16310
rect -870 16290 -850 16310
rect -850 16290 -845 16310
rect -875 16285 -845 16290
rect -715 16310 -685 16315
rect -715 16290 -710 16310
rect -710 16290 -690 16310
rect -690 16290 -685 16310
rect -715 16285 -685 16290
rect -555 16310 -525 16315
rect -555 16290 -550 16310
rect -550 16290 -530 16310
rect -530 16290 -525 16310
rect -555 16285 -525 16290
rect -14955 16150 -14925 16155
rect -14955 16130 -14950 16150
rect -14950 16130 -14930 16150
rect -14930 16130 -14925 16150
rect -14955 16125 -14925 16130
rect -14875 16150 -14845 16155
rect -14875 16130 -14870 16150
rect -14870 16130 -14850 16150
rect -14850 16130 -14845 16150
rect -14875 16125 -14845 16130
rect -14795 16150 -14765 16155
rect -14795 16130 -14790 16150
rect -14790 16130 -14770 16150
rect -14770 16130 -14765 16150
rect -14795 16125 -14765 16130
rect -14715 16150 -14685 16155
rect -14715 16130 -14710 16150
rect -14710 16130 -14690 16150
rect -14690 16130 -14685 16150
rect -14715 16125 -14685 16130
rect -14635 16150 -14605 16155
rect -14635 16130 -14630 16150
rect -14630 16130 -14610 16150
rect -14610 16130 -14605 16150
rect -14635 16125 -14605 16130
rect -14555 16150 -14525 16155
rect -14555 16130 -14550 16150
rect -14550 16130 -14530 16150
rect -14530 16130 -14525 16150
rect -14555 16125 -14525 16130
rect -14475 16150 -14445 16155
rect -14475 16130 -14470 16150
rect -14470 16130 -14450 16150
rect -14450 16130 -14445 16150
rect -14475 16125 -14445 16130
rect -14395 16150 -14365 16155
rect -14395 16130 -14390 16150
rect -14390 16130 -14370 16150
rect -14370 16130 -14365 16150
rect -14395 16125 -14365 16130
rect -14315 16150 -14285 16155
rect -14315 16130 -14310 16150
rect -14310 16130 -14290 16150
rect -14290 16130 -14285 16150
rect -14315 16125 -14285 16130
rect -14235 16150 -14205 16155
rect -14235 16130 -14230 16150
rect -14230 16130 -14210 16150
rect -14210 16130 -14205 16150
rect -14235 16125 -14205 16130
rect -14155 16150 -14125 16155
rect -14155 16130 -14150 16150
rect -14150 16130 -14130 16150
rect -14130 16130 -14125 16150
rect -14155 16125 -14125 16130
rect -14075 16150 -14045 16155
rect -14075 16130 -14070 16150
rect -14070 16130 -14050 16150
rect -14050 16130 -14045 16150
rect -14075 16125 -14045 16130
rect -13995 16150 -13965 16155
rect -13995 16130 -13990 16150
rect -13990 16130 -13970 16150
rect -13970 16130 -13965 16150
rect -13995 16125 -13965 16130
rect -13915 16150 -13885 16155
rect -13915 16130 -13910 16150
rect -13910 16130 -13890 16150
rect -13890 16130 -13885 16150
rect -13915 16125 -13885 16130
rect -13835 16150 -13805 16155
rect -13835 16130 -13830 16150
rect -13830 16130 -13810 16150
rect -13810 16130 -13805 16150
rect -13835 16125 -13805 16130
rect -13755 16150 -13725 16155
rect -13755 16130 -13750 16150
rect -13750 16130 -13730 16150
rect -13730 16130 -13725 16150
rect -13755 16125 -13725 16130
rect -13675 16150 -13645 16155
rect -13675 16130 -13670 16150
rect -13670 16130 -13650 16150
rect -13650 16130 -13645 16150
rect -13675 16125 -13645 16130
rect -13595 16150 -13565 16155
rect -13595 16130 -13590 16150
rect -13590 16130 -13570 16150
rect -13570 16130 -13565 16150
rect -13595 16125 -13565 16130
rect -13515 16150 -13485 16155
rect -13515 16130 -13510 16150
rect -13510 16130 -13490 16150
rect -13490 16130 -13485 16150
rect -13515 16125 -13485 16130
rect -13435 16150 -13405 16155
rect -13435 16130 -13430 16150
rect -13430 16130 -13410 16150
rect -13410 16130 -13405 16150
rect -13435 16125 -13405 16130
rect -13355 16150 -13325 16155
rect -13355 16130 -13350 16150
rect -13350 16130 -13330 16150
rect -13330 16130 -13325 16150
rect -13355 16125 -13325 16130
rect -13275 16150 -13245 16155
rect -13275 16130 -13270 16150
rect -13270 16130 -13250 16150
rect -13250 16130 -13245 16150
rect -13275 16125 -13245 16130
rect -13195 16150 -13165 16155
rect -13195 16130 -13190 16150
rect -13190 16130 -13170 16150
rect -13170 16130 -13165 16150
rect -13195 16125 -13165 16130
rect -13115 16150 -13085 16155
rect -13115 16130 -13110 16150
rect -13110 16130 -13090 16150
rect -13090 16130 -13085 16150
rect -13115 16125 -13085 16130
rect -13035 16150 -13005 16155
rect -13035 16130 -13030 16150
rect -13030 16130 -13010 16150
rect -13010 16130 -13005 16150
rect -13035 16125 -13005 16130
rect -12955 16150 -12925 16155
rect -12955 16130 -12950 16150
rect -12950 16130 -12930 16150
rect -12930 16130 -12925 16150
rect -12955 16125 -12925 16130
rect -12875 16150 -12845 16155
rect -12875 16130 -12870 16150
rect -12870 16130 -12850 16150
rect -12850 16130 -12845 16150
rect -12875 16125 -12845 16130
rect -12795 16150 -12765 16155
rect -12795 16130 -12790 16150
rect -12790 16130 -12770 16150
rect -12770 16130 -12765 16150
rect -12795 16125 -12765 16130
rect -12715 16150 -12685 16155
rect -12715 16130 -12710 16150
rect -12710 16130 -12690 16150
rect -12690 16130 -12685 16150
rect -12715 16125 -12685 16130
rect -12635 16150 -12605 16155
rect -12635 16130 -12630 16150
rect -12630 16130 -12610 16150
rect -12610 16130 -12605 16150
rect -12635 16125 -12605 16130
rect -12555 16150 -12525 16155
rect -12555 16130 -12550 16150
rect -12550 16130 -12530 16150
rect -12530 16130 -12525 16150
rect -12555 16125 -12525 16130
rect -12475 16150 -12445 16155
rect -12475 16130 -12470 16150
rect -12470 16130 -12450 16150
rect -12450 16130 -12445 16150
rect -12475 16125 -12445 16130
rect -12395 16150 -12365 16155
rect -12395 16130 -12390 16150
rect -12390 16130 -12370 16150
rect -12370 16130 -12365 16150
rect -12395 16125 -12365 16130
rect -12315 16150 -12285 16155
rect -12315 16130 -12310 16150
rect -12310 16130 -12290 16150
rect -12290 16130 -12285 16150
rect -12315 16125 -12285 16130
rect -12235 16150 -12205 16155
rect -12235 16130 -12230 16150
rect -12230 16130 -12210 16150
rect -12210 16130 -12205 16150
rect -12235 16125 -12205 16130
rect -12155 16150 -12125 16155
rect -12155 16130 -12150 16150
rect -12150 16130 -12130 16150
rect -12130 16130 -12125 16150
rect -12155 16125 -12125 16130
rect -12075 16150 -12045 16155
rect -12075 16130 -12070 16150
rect -12070 16130 -12050 16150
rect -12050 16130 -12045 16150
rect -12075 16125 -12045 16130
rect -11995 16150 -11965 16155
rect -11995 16130 -11990 16150
rect -11990 16130 -11970 16150
rect -11970 16130 -11965 16150
rect -11995 16125 -11965 16130
rect -11915 16150 -11885 16155
rect -11915 16130 -11910 16150
rect -11910 16130 -11890 16150
rect -11890 16130 -11885 16150
rect -11915 16125 -11885 16130
rect -11835 16150 -11805 16155
rect -11835 16130 -11830 16150
rect -11830 16130 -11810 16150
rect -11810 16130 -11805 16150
rect -11835 16125 -11805 16130
rect -11755 16150 -11725 16155
rect -11755 16130 -11750 16150
rect -11750 16130 -11730 16150
rect -11730 16130 -11725 16150
rect -11755 16125 -11725 16130
rect -11675 16150 -11645 16155
rect -11675 16130 -11670 16150
rect -11670 16130 -11650 16150
rect -11650 16130 -11645 16150
rect -11675 16125 -11645 16130
rect -11595 16150 -11565 16155
rect -11595 16130 -11590 16150
rect -11590 16130 -11570 16150
rect -11570 16130 -11565 16150
rect -11595 16125 -11565 16130
rect -11515 16150 -11485 16155
rect -11515 16130 -11510 16150
rect -11510 16130 -11490 16150
rect -11490 16130 -11485 16150
rect -11515 16125 -11485 16130
rect -11435 16150 -11405 16155
rect -11435 16130 -11430 16150
rect -11430 16130 -11410 16150
rect -11410 16130 -11405 16150
rect -11435 16125 -11405 16130
rect -11355 16150 -11325 16155
rect -11355 16130 -11350 16150
rect -11350 16130 -11330 16150
rect -11330 16130 -11325 16150
rect -11355 16125 -11325 16130
rect -11275 16150 -11245 16155
rect -11275 16130 -11270 16150
rect -11270 16130 -11250 16150
rect -11250 16130 -11245 16150
rect -11275 16125 -11245 16130
rect -11195 16150 -11165 16155
rect -11195 16130 -11190 16150
rect -11190 16130 -11170 16150
rect -11170 16130 -11165 16150
rect -11195 16125 -11165 16130
rect -11115 16150 -11085 16155
rect -11115 16130 -11110 16150
rect -11110 16130 -11090 16150
rect -11090 16130 -11085 16150
rect -11115 16125 -11085 16130
rect -11035 16150 -11005 16155
rect -11035 16130 -11030 16150
rect -11030 16130 -11010 16150
rect -11010 16130 -11005 16150
rect -11035 16125 -11005 16130
rect -10955 16150 -10925 16155
rect -10955 16130 -10950 16150
rect -10950 16130 -10930 16150
rect -10930 16130 -10925 16150
rect -10955 16125 -10925 16130
rect -10875 16150 -10845 16155
rect -10875 16130 -10870 16150
rect -10870 16130 -10850 16150
rect -10850 16130 -10845 16150
rect -10875 16125 -10845 16130
rect -10795 16150 -10765 16155
rect -10795 16130 -10790 16150
rect -10790 16130 -10770 16150
rect -10770 16130 -10765 16150
rect -10795 16125 -10765 16130
rect -10715 16150 -10685 16155
rect -10715 16130 -10710 16150
rect -10710 16130 -10690 16150
rect -10690 16130 -10685 16150
rect -10715 16125 -10685 16130
rect -10635 16150 -10605 16155
rect -10635 16130 -10630 16150
rect -10630 16130 -10610 16150
rect -10610 16130 -10605 16150
rect -10635 16125 -10605 16130
rect -10555 16150 -10525 16155
rect -10555 16130 -10550 16150
rect -10550 16130 -10530 16150
rect -10530 16130 -10525 16150
rect -10555 16125 -10525 16130
rect -10475 16150 -10445 16155
rect -10475 16130 -10470 16150
rect -10470 16130 -10450 16150
rect -10450 16130 -10445 16150
rect -10475 16125 -10445 16130
rect -10395 16150 -10365 16155
rect -10395 16130 -10390 16150
rect -10390 16130 -10370 16150
rect -10370 16130 -10365 16150
rect -10395 16125 -10365 16130
rect -10315 16150 -10285 16155
rect -10315 16130 -10310 16150
rect -10310 16130 -10290 16150
rect -10290 16130 -10285 16150
rect -10315 16125 -10285 16130
rect -10235 16150 -10205 16155
rect -10235 16130 -10230 16150
rect -10230 16130 -10210 16150
rect -10210 16130 -10205 16150
rect -10235 16125 -10205 16130
rect -10155 16150 -10125 16155
rect -10155 16130 -10150 16150
rect -10150 16130 -10130 16150
rect -10130 16130 -10125 16150
rect -10155 16125 -10125 16130
rect -10075 16150 -10045 16155
rect -10075 16130 -10070 16150
rect -10070 16130 -10050 16150
rect -10050 16130 -10045 16150
rect -10075 16125 -10045 16130
rect -9995 16150 -9965 16155
rect -9995 16130 -9990 16150
rect -9990 16130 -9970 16150
rect -9970 16130 -9965 16150
rect -9995 16125 -9965 16130
rect -9915 16150 -9885 16155
rect -9915 16130 -9910 16150
rect -9910 16130 -9890 16150
rect -9890 16130 -9885 16150
rect -9915 16125 -9885 16130
rect -9835 16150 -9805 16155
rect -9835 16130 -9830 16150
rect -9830 16130 -9810 16150
rect -9810 16130 -9805 16150
rect -9835 16125 -9805 16130
rect -9755 16150 -9725 16155
rect -9755 16130 -9750 16150
rect -9750 16130 -9730 16150
rect -9730 16130 -9725 16150
rect -9755 16125 -9725 16130
rect -9675 16150 -9645 16155
rect -9675 16130 -9670 16150
rect -9670 16130 -9650 16150
rect -9650 16130 -9645 16150
rect -9675 16125 -9645 16130
rect -9595 16150 -9565 16155
rect -9595 16130 -9590 16150
rect -9590 16130 -9570 16150
rect -9570 16130 -9565 16150
rect -9595 16125 -9565 16130
rect -9515 16150 -9485 16155
rect -9515 16130 -9510 16150
rect -9510 16130 -9490 16150
rect -9490 16130 -9485 16150
rect -9515 16125 -9485 16130
rect -9435 16150 -9405 16155
rect -9435 16130 -9430 16150
rect -9430 16130 -9410 16150
rect -9410 16130 -9405 16150
rect -9435 16125 -9405 16130
rect -9355 16150 -9325 16155
rect -9355 16130 -9350 16150
rect -9350 16130 -9330 16150
rect -9330 16130 -9325 16150
rect -9355 16125 -9325 16130
rect -9275 16150 -9245 16155
rect -9275 16130 -9270 16150
rect -9270 16130 -9250 16150
rect -9250 16130 -9245 16150
rect -9275 16125 -9245 16130
rect -9195 16150 -9165 16155
rect -9195 16130 -9190 16150
rect -9190 16130 -9170 16150
rect -9170 16130 -9165 16150
rect -9195 16125 -9165 16130
rect -9115 16150 -9085 16155
rect -9115 16130 -9110 16150
rect -9110 16130 -9090 16150
rect -9090 16130 -9085 16150
rect -9115 16125 -9085 16130
rect -9035 16150 -9005 16155
rect -9035 16130 -9030 16150
rect -9030 16130 -9010 16150
rect -9010 16130 -9005 16150
rect -9035 16125 -9005 16130
rect -8955 16150 -8925 16155
rect -8955 16130 -8950 16150
rect -8950 16130 -8930 16150
rect -8930 16130 -8925 16150
rect -8955 16125 -8925 16130
rect -8875 16150 -8845 16155
rect -8875 16130 -8870 16150
rect -8870 16130 -8850 16150
rect -8850 16130 -8845 16150
rect -8875 16125 -8845 16130
rect -8795 16150 -8765 16155
rect -8795 16130 -8790 16150
rect -8790 16130 -8770 16150
rect -8770 16130 -8765 16150
rect -8795 16125 -8765 16130
rect -8715 16150 -8685 16155
rect -8715 16130 -8710 16150
rect -8710 16130 -8690 16150
rect -8690 16130 -8685 16150
rect -8715 16125 -8685 16130
rect -8635 16150 -8605 16155
rect -8635 16130 -8630 16150
rect -8630 16130 -8610 16150
rect -8610 16130 -8605 16150
rect -8635 16125 -8605 16130
rect -8555 16150 -8525 16155
rect -8555 16130 -8550 16150
rect -8550 16130 -8530 16150
rect -8530 16130 -8525 16150
rect -8555 16125 -8525 16130
rect -8475 16150 -8445 16155
rect -8475 16130 -8470 16150
rect -8470 16130 -8450 16150
rect -8450 16130 -8445 16150
rect -8475 16125 -8445 16130
rect -8395 16150 -8365 16155
rect -8395 16130 -8390 16150
rect -8390 16130 -8370 16150
rect -8370 16130 -8365 16150
rect -8395 16125 -8365 16130
rect -8315 16150 -8285 16155
rect -8315 16130 -8310 16150
rect -8310 16130 -8290 16150
rect -8290 16130 -8285 16150
rect -8315 16125 -8285 16130
rect -8235 16150 -8205 16155
rect -8235 16130 -8230 16150
rect -8230 16130 -8210 16150
rect -8210 16130 -8205 16150
rect -8235 16125 -8205 16130
rect -8155 16150 -8125 16155
rect -8155 16130 -8150 16150
rect -8150 16130 -8130 16150
rect -8130 16130 -8125 16150
rect -8155 16125 -8125 16130
rect -8075 16150 -8045 16155
rect -8075 16130 -8070 16150
rect -8070 16130 -8050 16150
rect -8050 16130 -8045 16150
rect -8075 16125 -8045 16130
rect -7995 16150 -7965 16155
rect -7995 16130 -7990 16150
rect -7990 16130 -7970 16150
rect -7970 16130 -7965 16150
rect -7995 16125 -7965 16130
rect -7915 16150 -7885 16155
rect -7915 16130 -7910 16150
rect -7910 16130 -7890 16150
rect -7890 16130 -7885 16150
rect -7915 16125 -7885 16130
rect -7835 16150 -7805 16155
rect -7835 16130 -7830 16150
rect -7830 16130 -7810 16150
rect -7810 16130 -7805 16150
rect -7835 16125 -7805 16130
rect -7755 16150 -7725 16155
rect -7755 16130 -7750 16150
rect -7750 16130 -7730 16150
rect -7730 16130 -7725 16150
rect -7755 16125 -7725 16130
rect -7675 16150 -7645 16155
rect -7675 16130 -7670 16150
rect -7670 16130 -7650 16150
rect -7650 16130 -7645 16150
rect -7675 16125 -7645 16130
rect -7595 16150 -7565 16155
rect -7595 16130 -7590 16150
rect -7590 16130 -7570 16150
rect -7570 16130 -7565 16150
rect -7595 16125 -7565 16130
rect -7515 16150 -7485 16155
rect -7515 16130 -7510 16150
rect -7510 16130 -7490 16150
rect -7490 16130 -7485 16150
rect -7515 16125 -7485 16130
rect -7435 16150 -7405 16155
rect -7435 16130 -7430 16150
rect -7430 16130 -7410 16150
rect -7410 16130 -7405 16150
rect -7435 16125 -7405 16130
rect -7355 16150 -7325 16155
rect -7355 16130 -7350 16150
rect -7350 16130 -7330 16150
rect -7330 16130 -7325 16150
rect -7355 16125 -7325 16130
rect -7275 16150 -7245 16155
rect -7275 16130 -7270 16150
rect -7270 16130 -7250 16150
rect -7250 16130 -7245 16150
rect -7275 16125 -7245 16130
rect -7195 16150 -7165 16155
rect -7195 16130 -7190 16150
rect -7190 16130 -7170 16150
rect -7170 16130 -7165 16150
rect -7195 16125 -7165 16130
rect -7115 16150 -7085 16155
rect -7115 16130 -7110 16150
rect -7110 16130 -7090 16150
rect -7090 16130 -7085 16150
rect -7115 16125 -7085 16130
rect -7035 16150 -7005 16155
rect -7035 16130 -7030 16150
rect -7030 16130 -7010 16150
rect -7010 16130 -7005 16150
rect -7035 16125 -7005 16130
rect -6955 16150 -6925 16155
rect -6955 16130 -6950 16150
rect -6950 16130 -6930 16150
rect -6930 16130 -6925 16150
rect -6955 16125 -6925 16130
rect -6875 16150 -6845 16155
rect -6875 16130 -6870 16150
rect -6870 16130 -6850 16150
rect -6850 16130 -6845 16150
rect -6875 16125 -6845 16130
rect -6795 16150 -6765 16155
rect -6795 16130 -6790 16150
rect -6790 16130 -6770 16150
rect -6770 16130 -6765 16150
rect -6795 16125 -6765 16130
rect -6715 16150 -6685 16155
rect -6715 16130 -6710 16150
rect -6710 16130 -6690 16150
rect -6690 16130 -6685 16150
rect -6715 16125 -6685 16130
rect -6635 16150 -6605 16155
rect -6635 16130 -6630 16150
rect -6630 16130 -6610 16150
rect -6610 16130 -6605 16150
rect -6635 16125 -6605 16130
rect -6555 16150 -6525 16155
rect -6555 16130 -6550 16150
rect -6550 16130 -6530 16150
rect -6530 16130 -6525 16150
rect -6555 16125 -6525 16130
rect -6475 16150 -6445 16155
rect -6475 16130 -6470 16150
rect -6470 16130 -6450 16150
rect -6450 16130 -6445 16150
rect -6475 16125 -6445 16130
rect -6395 16150 -6365 16155
rect -6395 16130 -6390 16150
rect -6390 16130 -6370 16150
rect -6370 16130 -6365 16150
rect -6395 16125 -6365 16130
rect -6315 16150 -6285 16155
rect -6315 16130 -6310 16150
rect -6310 16130 -6290 16150
rect -6290 16130 -6285 16150
rect -6315 16125 -6285 16130
rect -6235 16150 -6205 16155
rect -6235 16130 -6230 16150
rect -6230 16130 -6210 16150
rect -6210 16130 -6205 16150
rect -6235 16125 -6205 16130
rect -6155 16150 -6125 16155
rect -6155 16130 -6150 16150
rect -6150 16130 -6130 16150
rect -6130 16130 -6125 16150
rect -6155 16125 -6125 16130
rect -6075 16150 -6045 16155
rect -6075 16130 -6070 16150
rect -6070 16130 -6050 16150
rect -6050 16130 -6045 16150
rect -6075 16125 -6045 16130
rect -5995 16150 -5965 16155
rect -5995 16130 -5990 16150
rect -5990 16130 -5970 16150
rect -5970 16130 -5965 16150
rect -5995 16125 -5965 16130
rect -5915 16150 -5885 16155
rect -5915 16130 -5910 16150
rect -5910 16130 -5890 16150
rect -5890 16130 -5885 16150
rect -5915 16125 -5885 16130
rect -5835 16150 -5805 16155
rect -5835 16130 -5830 16150
rect -5830 16130 -5810 16150
rect -5810 16130 -5805 16150
rect -5835 16125 -5805 16130
rect -5755 16150 -5725 16155
rect -5755 16130 -5750 16150
rect -5750 16130 -5730 16150
rect -5730 16130 -5725 16150
rect -5755 16125 -5725 16130
rect -5675 16150 -5645 16155
rect -5675 16130 -5670 16150
rect -5670 16130 -5650 16150
rect -5650 16130 -5645 16150
rect -5675 16125 -5645 16130
rect -5595 16150 -5565 16155
rect -5595 16130 -5590 16150
rect -5590 16130 -5570 16150
rect -5570 16130 -5565 16150
rect -5595 16125 -5565 16130
rect -5435 16150 -5405 16155
rect -5435 16130 -5430 16150
rect -5430 16130 -5410 16150
rect -5410 16130 -5405 16150
rect -5435 16125 -5405 16130
rect -5355 16150 -5325 16155
rect -5355 16130 -5350 16150
rect -5350 16130 -5330 16150
rect -5330 16130 -5325 16150
rect -5355 16125 -5325 16130
rect -5275 16150 -5245 16155
rect -5275 16130 -5270 16150
rect -5270 16130 -5250 16150
rect -5250 16130 -5245 16150
rect -5275 16125 -5245 16130
rect -5195 16150 -5165 16155
rect -5195 16130 -5190 16150
rect -5190 16130 -5170 16150
rect -5170 16130 -5165 16150
rect -5195 16125 -5165 16130
rect -5115 16150 -5085 16155
rect -5115 16130 -5110 16150
rect -5110 16130 -5090 16150
rect -5090 16130 -5085 16150
rect -5115 16125 -5085 16130
rect -5035 16150 -5005 16155
rect -5035 16130 -5030 16150
rect -5030 16130 -5010 16150
rect -5010 16130 -5005 16150
rect -5035 16125 -5005 16130
rect -4955 16150 -4925 16155
rect -4955 16130 -4950 16150
rect -4950 16130 -4930 16150
rect -4930 16130 -4925 16150
rect -4955 16125 -4925 16130
rect -4875 16150 -4845 16155
rect -4875 16130 -4870 16150
rect -4870 16130 -4850 16150
rect -4850 16130 -4845 16150
rect -4875 16125 -4845 16130
rect -4795 16150 -4765 16155
rect -4795 16130 -4790 16150
rect -4790 16130 -4770 16150
rect -4770 16130 -4765 16150
rect -4795 16125 -4765 16130
rect -4715 16150 -4685 16155
rect -4715 16130 -4710 16150
rect -4710 16130 -4690 16150
rect -4690 16130 -4685 16150
rect -4715 16125 -4685 16130
rect -4635 16150 -4605 16155
rect -4635 16130 -4630 16150
rect -4630 16130 -4610 16150
rect -4610 16130 -4605 16150
rect -4635 16125 -4605 16130
rect -4555 16150 -4525 16155
rect -4555 16130 -4550 16150
rect -4550 16130 -4530 16150
rect -4530 16130 -4525 16150
rect -4555 16125 -4525 16130
rect -4475 16150 -4445 16155
rect -4475 16130 -4470 16150
rect -4470 16130 -4450 16150
rect -4450 16130 -4445 16150
rect -4475 16125 -4445 16130
rect -4395 16150 -4365 16155
rect -4395 16130 -4390 16150
rect -4390 16130 -4370 16150
rect -4370 16130 -4365 16150
rect -4395 16125 -4365 16130
rect -4315 16150 -4285 16155
rect -4315 16130 -4310 16150
rect -4310 16130 -4290 16150
rect -4290 16130 -4285 16150
rect -4315 16125 -4285 16130
rect -4235 16150 -4205 16155
rect -4235 16130 -4230 16150
rect -4230 16130 -4210 16150
rect -4210 16130 -4205 16150
rect -4235 16125 -4205 16130
rect -4155 16150 -4125 16155
rect -4155 16130 -4150 16150
rect -4150 16130 -4130 16150
rect -4130 16130 -4125 16150
rect -4155 16125 -4125 16130
rect -4075 16150 -4045 16155
rect -4075 16130 -4070 16150
rect -4070 16130 -4050 16150
rect -4050 16130 -4045 16150
rect -4075 16125 -4045 16130
rect -3995 16150 -3965 16155
rect -3995 16130 -3990 16150
rect -3990 16130 -3970 16150
rect -3970 16130 -3965 16150
rect -3995 16125 -3965 16130
rect -3915 16150 -3885 16155
rect -3915 16130 -3910 16150
rect -3910 16130 -3890 16150
rect -3890 16130 -3885 16150
rect -3915 16125 -3885 16130
rect -3835 16150 -3805 16155
rect -3835 16130 -3830 16150
rect -3830 16130 -3810 16150
rect -3810 16130 -3805 16150
rect -3835 16125 -3805 16130
rect -3755 16150 -3725 16155
rect -3755 16130 -3750 16150
rect -3750 16130 -3730 16150
rect -3730 16130 -3725 16150
rect -3755 16125 -3725 16130
rect -3675 16150 -3645 16155
rect -3675 16130 -3670 16150
rect -3670 16130 -3650 16150
rect -3650 16130 -3645 16150
rect -3675 16125 -3645 16130
rect -3595 16150 -3565 16155
rect -3595 16130 -3590 16150
rect -3590 16130 -3570 16150
rect -3570 16130 -3565 16150
rect -3595 16125 -3565 16130
rect -3515 16150 -3485 16155
rect -3515 16130 -3510 16150
rect -3510 16130 -3490 16150
rect -3490 16130 -3485 16150
rect -3515 16125 -3485 16130
rect -3435 16150 -3405 16155
rect -3435 16130 -3430 16150
rect -3430 16130 -3410 16150
rect -3410 16130 -3405 16150
rect -3435 16125 -3405 16130
rect -3355 16150 -3325 16155
rect -3355 16130 -3350 16150
rect -3350 16130 -3330 16150
rect -3330 16130 -3325 16150
rect -3355 16125 -3325 16130
rect -3275 16150 -3245 16155
rect -3275 16130 -3270 16150
rect -3270 16130 -3250 16150
rect -3250 16130 -3245 16150
rect -3275 16125 -3245 16130
rect -3195 16150 -3165 16155
rect -3195 16130 -3190 16150
rect -3190 16130 -3170 16150
rect -3170 16130 -3165 16150
rect -3195 16125 -3165 16130
rect -3115 16150 -3085 16155
rect -3115 16130 -3110 16150
rect -3110 16130 -3090 16150
rect -3090 16130 -3085 16150
rect -3115 16125 -3085 16130
rect -3035 16150 -3005 16155
rect -3035 16130 -3030 16150
rect -3030 16130 -3010 16150
rect -3010 16130 -3005 16150
rect -3035 16125 -3005 16130
rect -2955 16150 -2925 16155
rect -2955 16130 -2950 16150
rect -2950 16130 -2930 16150
rect -2930 16130 -2925 16150
rect -2955 16125 -2925 16130
rect -2875 16150 -2845 16155
rect -2875 16130 -2870 16150
rect -2870 16130 -2850 16150
rect -2850 16130 -2845 16150
rect -2875 16125 -2845 16130
rect -2795 16150 -2765 16155
rect -2795 16130 -2790 16150
rect -2790 16130 -2770 16150
rect -2770 16130 -2765 16150
rect -2795 16125 -2765 16130
rect -2715 16150 -2685 16155
rect -2715 16130 -2710 16150
rect -2710 16130 -2690 16150
rect -2690 16130 -2685 16150
rect -2715 16125 -2685 16130
rect -2635 16150 -2605 16155
rect -2635 16130 -2630 16150
rect -2630 16130 -2610 16150
rect -2610 16130 -2605 16150
rect -2635 16125 -2605 16130
rect -2555 16150 -2525 16155
rect -2555 16130 -2550 16150
rect -2550 16130 -2530 16150
rect -2530 16130 -2525 16150
rect -2555 16125 -2525 16130
rect -2475 16150 -2445 16155
rect -2475 16130 -2470 16150
rect -2470 16130 -2450 16150
rect -2450 16130 -2445 16150
rect -2475 16125 -2445 16130
rect -2395 16150 -2365 16155
rect -2395 16130 -2390 16150
rect -2390 16130 -2370 16150
rect -2370 16130 -2365 16150
rect -2395 16125 -2365 16130
rect -2315 16150 -2285 16155
rect -2315 16130 -2310 16150
rect -2310 16130 -2290 16150
rect -2290 16130 -2285 16150
rect -2315 16125 -2285 16130
rect -2235 16150 -2205 16155
rect -2235 16130 -2230 16150
rect -2230 16130 -2210 16150
rect -2210 16130 -2205 16150
rect -2235 16125 -2205 16130
rect -2155 16150 -2125 16155
rect -2155 16130 -2150 16150
rect -2150 16130 -2130 16150
rect -2130 16130 -2125 16150
rect -2155 16125 -2125 16130
rect -2075 16150 -2045 16155
rect -2075 16130 -2070 16150
rect -2070 16130 -2050 16150
rect -2050 16130 -2045 16150
rect -2075 16125 -2045 16130
rect -1995 16150 -1965 16155
rect -1995 16130 -1990 16150
rect -1990 16130 -1970 16150
rect -1970 16130 -1965 16150
rect -1995 16125 -1965 16130
rect -1835 16150 -1805 16155
rect -1835 16130 -1830 16150
rect -1830 16130 -1810 16150
rect -1810 16130 -1805 16150
rect -1835 16125 -1805 16130
rect -1755 16150 -1725 16155
rect -1755 16130 -1750 16150
rect -1750 16130 -1730 16150
rect -1730 16130 -1725 16150
rect -1755 16125 -1725 16130
rect -1675 16150 -1645 16155
rect -1675 16130 -1670 16150
rect -1670 16130 -1650 16150
rect -1650 16130 -1645 16150
rect -1675 16125 -1645 16130
rect -1595 16150 -1565 16155
rect -1595 16130 -1590 16150
rect -1590 16130 -1570 16150
rect -1570 16130 -1565 16150
rect -1595 16125 -1565 16130
rect -1515 16150 -1485 16155
rect -1515 16130 -1510 16150
rect -1510 16130 -1490 16150
rect -1490 16130 -1485 16150
rect -1515 16125 -1485 16130
rect -1435 16150 -1405 16155
rect -1435 16130 -1430 16150
rect -1430 16130 -1410 16150
rect -1410 16130 -1405 16150
rect -1435 16125 -1405 16130
rect -1355 16150 -1325 16155
rect -1355 16130 -1350 16150
rect -1350 16130 -1330 16150
rect -1330 16130 -1325 16150
rect -1355 16125 -1325 16130
rect -1195 16150 -1165 16155
rect -1195 16130 -1190 16150
rect -1190 16130 -1170 16150
rect -1170 16130 -1165 16150
rect -1195 16125 -1165 16130
rect -1035 16150 -1005 16155
rect -1035 16130 -1030 16150
rect -1030 16130 -1010 16150
rect -1010 16130 -1005 16150
rect -1035 16125 -1005 16130
rect -875 16150 -845 16155
rect -875 16130 -870 16150
rect -870 16130 -850 16150
rect -850 16130 -845 16150
rect -875 16125 -845 16130
rect -715 16150 -685 16155
rect -715 16130 -710 16150
rect -710 16130 -690 16150
rect -690 16130 -685 16150
rect -715 16125 -685 16130
rect -555 16150 -525 16155
rect -555 16130 -550 16150
rect -550 16130 -530 16150
rect -530 16130 -525 16150
rect -555 16125 -525 16130
rect -14955 15990 -14925 15995
rect -14955 15970 -14950 15990
rect -14950 15970 -14930 15990
rect -14930 15970 -14925 15990
rect -14955 15965 -14925 15970
rect -14875 15990 -14845 15995
rect -14875 15970 -14870 15990
rect -14870 15970 -14850 15990
rect -14850 15970 -14845 15990
rect -14875 15965 -14845 15970
rect -14795 15990 -14765 15995
rect -14795 15970 -14790 15990
rect -14790 15970 -14770 15990
rect -14770 15970 -14765 15990
rect -14795 15965 -14765 15970
rect -14715 15990 -14685 15995
rect -14715 15970 -14710 15990
rect -14710 15970 -14690 15990
rect -14690 15970 -14685 15990
rect -14715 15965 -14685 15970
rect -14635 15990 -14605 15995
rect -14635 15970 -14630 15990
rect -14630 15970 -14610 15990
rect -14610 15970 -14605 15990
rect -14635 15965 -14605 15970
rect -14555 15990 -14525 15995
rect -14555 15970 -14550 15990
rect -14550 15970 -14530 15990
rect -14530 15970 -14525 15990
rect -14555 15965 -14525 15970
rect -14475 15990 -14445 15995
rect -14475 15970 -14470 15990
rect -14470 15970 -14450 15990
rect -14450 15970 -14445 15990
rect -14475 15965 -14445 15970
rect -14395 15990 -14365 15995
rect -14395 15970 -14390 15990
rect -14390 15970 -14370 15990
rect -14370 15970 -14365 15990
rect -14395 15965 -14365 15970
rect -14315 15990 -14285 15995
rect -14315 15970 -14310 15990
rect -14310 15970 -14290 15990
rect -14290 15970 -14285 15990
rect -14315 15965 -14285 15970
rect -14235 15990 -14205 15995
rect -14235 15970 -14230 15990
rect -14230 15970 -14210 15990
rect -14210 15970 -14205 15990
rect -14235 15965 -14205 15970
rect -14155 15990 -14125 15995
rect -14155 15970 -14150 15990
rect -14150 15970 -14130 15990
rect -14130 15970 -14125 15990
rect -14155 15965 -14125 15970
rect -14075 15990 -14045 15995
rect -14075 15970 -14070 15990
rect -14070 15970 -14050 15990
rect -14050 15970 -14045 15990
rect -14075 15965 -14045 15970
rect -13995 15990 -13965 15995
rect -13995 15970 -13990 15990
rect -13990 15970 -13970 15990
rect -13970 15970 -13965 15990
rect -13995 15965 -13965 15970
rect -13915 15990 -13885 15995
rect -13915 15970 -13910 15990
rect -13910 15970 -13890 15990
rect -13890 15970 -13885 15990
rect -13915 15965 -13885 15970
rect -13835 15990 -13805 15995
rect -13835 15970 -13830 15990
rect -13830 15970 -13810 15990
rect -13810 15970 -13805 15990
rect -13835 15965 -13805 15970
rect -13755 15990 -13725 15995
rect -13755 15970 -13750 15990
rect -13750 15970 -13730 15990
rect -13730 15970 -13725 15990
rect -13755 15965 -13725 15970
rect -13675 15990 -13645 15995
rect -13675 15970 -13670 15990
rect -13670 15970 -13650 15990
rect -13650 15970 -13645 15990
rect -13675 15965 -13645 15970
rect -13595 15990 -13565 15995
rect -13595 15970 -13590 15990
rect -13590 15970 -13570 15990
rect -13570 15970 -13565 15990
rect -13595 15965 -13565 15970
rect -13515 15990 -13485 15995
rect -13515 15970 -13510 15990
rect -13510 15970 -13490 15990
rect -13490 15970 -13485 15990
rect -13515 15965 -13485 15970
rect -13435 15990 -13405 15995
rect -13435 15970 -13430 15990
rect -13430 15970 -13410 15990
rect -13410 15970 -13405 15990
rect -13435 15965 -13405 15970
rect -13355 15990 -13325 15995
rect -13355 15970 -13350 15990
rect -13350 15970 -13330 15990
rect -13330 15970 -13325 15990
rect -13355 15965 -13325 15970
rect -13275 15990 -13245 15995
rect -13275 15970 -13270 15990
rect -13270 15970 -13250 15990
rect -13250 15970 -13245 15990
rect -13275 15965 -13245 15970
rect -13195 15990 -13165 15995
rect -13195 15970 -13190 15990
rect -13190 15970 -13170 15990
rect -13170 15970 -13165 15990
rect -13195 15965 -13165 15970
rect -13115 15990 -13085 15995
rect -13115 15970 -13110 15990
rect -13110 15970 -13090 15990
rect -13090 15970 -13085 15990
rect -13115 15965 -13085 15970
rect -13035 15990 -13005 15995
rect -13035 15970 -13030 15990
rect -13030 15970 -13010 15990
rect -13010 15970 -13005 15990
rect -13035 15965 -13005 15970
rect -12955 15990 -12925 15995
rect -12955 15970 -12950 15990
rect -12950 15970 -12930 15990
rect -12930 15970 -12925 15990
rect -12955 15965 -12925 15970
rect -12875 15990 -12845 15995
rect -12875 15970 -12870 15990
rect -12870 15970 -12850 15990
rect -12850 15970 -12845 15990
rect -12875 15965 -12845 15970
rect -12795 15990 -12765 15995
rect -12795 15970 -12790 15990
rect -12790 15970 -12770 15990
rect -12770 15970 -12765 15990
rect -12795 15965 -12765 15970
rect -12715 15990 -12685 15995
rect -12715 15970 -12710 15990
rect -12710 15970 -12690 15990
rect -12690 15970 -12685 15990
rect -12715 15965 -12685 15970
rect -12635 15990 -12605 15995
rect -12635 15970 -12630 15990
rect -12630 15970 -12610 15990
rect -12610 15970 -12605 15990
rect -12635 15965 -12605 15970
rect -12555 15990 -12525 15995
rect -12555 15970 -12550 15990
rect -12550 15970 -12530 15990
rect -12530 15970 -12525 15990
rect -12555 15965 -12525 15970
rect -12475 15990 -12445 15995
rect -12475 15970 -12470 15990
rect -12470 15970 -12450 15990
rect -12450 15970 -12445 15990
rect -12475 15965 -12445 15970
rect -12395 15990 -12365 15995
rect -12395 15970 -12390 15990
rect -12390 15970 -12370 15990
rect -12370 15970 -12365 15990
rect -12395 15965 -12365 15970
rect -12315 15990 -12285 15995
rect -12315 15970 -12310 15990
rect -12310 15970 -12290 15990
rect -12290 15970 -12285 15990
rect -12315 15965 -12285 15970
rect -12235 15990 -12205 15995
rect -12235 15970 -12230 15990
rect -12230 15970 -12210 15990
rect -12210 15970 -12205 15990
rect -12235 15965 -12205 15970
rect -12155 15990 -12125 15995
rect -12155 15970 -12150 15990
rect -12150 15970 -12130 15990
rect -12130 15970 -12125 15990
rect -12155 15965 -12125 15970
rect -12075 15990 -12045 15995
rect -12075 15970 -12070 15990
rect -12070 15970 -12050 15990
rect -12050 15970 -12045 15990
rect -12075 15965 -12045 15970
rect -11995 15990 -11965 15995
rect -11995 15970 -11990 15990
rect -11990 15970 -11970 15990
rect -11970 15970 -11965 15990
rect -11995 15965 -11965 15970
rect -11915 15990 -11885 15995
rect -11915 15970 -11910 15990
rect -11910 15970 -11890 15990
rect -11890 15970 -11885 15990
rect -11915 15965 -11885 15970
rect -11835 15990 -11805 15995
rect -11835 15970 -11830 15990
rect -11830 15970 -11810 15990
rect -11810 15970 -11805 15990
rect -11835 15965 -11805 15970
rect -11755 15990 -11725 15995
rect -11755 15970 -11750 15990
rect -11750 15970 -11730 15990
rect -11730 15970 -11725 15990
rect -11755 15965 -11725 15970
rect -11675 15990 -11645 15995
rect -11675 15970 -11670 15990
rect -11670 15970 -11650 15990
rect -11650 15970 -11645 15990
rect -11675 15965 -11645 15970
rect -11595 15990 -11565 15995
rect -11595 15970 -11590 15990
rect -11590 15970 -11570 15990
rect -11570 15970 -11565 15990
rect -11595 15965 -11565 15970
rect -11515 15990 -11485 15995
rect -11515 15970 -11510 15990
rect -11510 15970 -11490 15990
rect -11490 15970 -11485 15990
rect -11515 15965 -11485 15970
rect -11435 15990 -11405 15995
rect -11435 15970 -11430 15990
rect -11430 15970 -11410 15990
rect -11410 15970 -11405 15990
rect -11435 15965 -11405 15970
rect -11355 15990 -11325 15995
rect -11355 15970 -11350 15990
rect -11350 15970 -11330 15990
rect -11330 15970 -11325 15990
rect -11355 15965 -11325 15970
rect -11275 15990 -11245 15995
rect -11275 15970 -11270 15990
rect -11270 15970 -11250 15990
rect -11250 15970 -11245 15990
rect -11275 15965 -11245 15970
rect -11195 15990 -11165 15995
rect -11195 15970 -11190 15990
rect -11190 15970 -11170 15990
rect -11170 15970 -11165 15990
rect -11195 15965 -11165 15970
rect -11115 15990 -11085 15995
rect -11115 15970 -11110 15990
rect -11110 15970 -11090 15990
rect -11090 15970 -11085 15990
rect -11115 15965 -11085 15970
rect -11035 15990 -11005 15995
rect -11035 15970 -11030 15990
rect -11030 15970 -11010 15990
rect -11010 15970 -11005 15990
rect -11035 15965 -11005 15970
rect -10955 15990 -10925 15995
rect -10955 15970 -10950 15990
rect -10950 15970 -10930 15990
rect -10930 15970 -10925 15990
rect -10955 15965 -10925 15970
rect -10875 15990 -10845 15995
rect -10875 15970 -10870 15990
rect -10870 15970 -10850 15990
rect -10850 15970 -10845 15990
rect -10875 15965 -10845 15970
rect -10795 15990 -10765 15995
rect -10795 15970 -10790 15990
rect -10790 15970 -10770 15990
rect -10770 15970 -10765 15990
rect -10795 15965 -10765 15970
rect -10715 15990 -10685 15995
rect -10715 15970 -10710 15990
rect -10710 15970 -10690 15990
rect -10690 15970 -10685 15990
rect -10715 15965 -10685 15970
rect -10635 15990 -10605 15995
rect -10635 15970 -10630 15990
rect -10630 15970 -10610 15990
rect -10610 15970 -10605 15990
rect -10635 15965 -10605 15970
rect -10555 15990 -10525 15995
rect -10555 15970 -10550 15990
rect -10550 15970 -10530 15990
rect -10530 15970 -10525 15990
rect -10555 15965 -10525 15970
rect -10475 15990 -10445 15995
rect -10475 15970 -10470 15990
rect -10470 15970 -10450 15990
rect -10450 15970 -10445 15990
rect -10475 15965 -10445 15970
rect -10395 15990 -10365 15995
rect -10395 15970 -10390 15990
rect -10390 15970 -10370 15990
rect -10370 15970 -10365 15990
rect -10395 15965 -10365 15970
rect -10315 15990 -10285 15995
rect -10315 15970 -10310 15990
rect -10310 15970 -10290 15990
rect -10290 15970 -10285 15990
rect -10315 15965 -10285 15970
rect -10235 15990 -10205 15995
rect -10235 15970 -10230 15990
rect -10230 15970 -10210 15990
rect -10210 15970 -10205 15990
rect -10235 15965 -10205 15970
rect -10155 15990 -10125 15995
rect -10155 15970 -10150 15990
rect -10150 15970 -10130 15990
rect -10130 15970 -10125 15990
rect -10155 15965 -10125 15970
rect -10075 15990 -10045 15995
rect -10075 15970 -10070 15990
rect -10070 15970 -10050 15990
rect -10050 15970 -10045 15990
rect -10075 15965 -10045 15970
rect -9995 15990 -9965 15995
rect -9995 15970 -9990 15990
rect -9990 15970 -9970 15990
rect -9970 15970 -9965 15990
rect -9995 15965 -9965 15970
rect -9915 15990 -9885 15995
rect -9915 15970 -9910 15990
rect -9910 15970 -9890 15990
rect -9890 15970 -9885 15990
rect -9915 15965 -9885 15970
rect -9835 15990 -9805 15995
rect -9835 15970 -9830 15990
rect -9830 15970 -9810 15990
rect -9810 15970 -9805 15990
rect -9835 15965 -9805 15970
rect -9755 15990 -9725 15995
rect -9755 15970 -9750 15990
rect -9750 15970 -9730 15990
rect -9730 15970 -9725 15990
rect -9755 15965 -9725 15970
rect -9675 15990 -9645 15995
rect -9675 15970 -9670 15990
rect -9670 15970 -9650 15990
rect -9650 15970 -9645 15990
rect -9675 15965 -9645 15970
rect -9595 15990 -9565 15995
rect -9595 15970 -9590 15990
rect -9590 15970 -9570 15990
rect -9570 15970 -9565 15990
rect -9595 15965 -9565 15970
rect -9515 15990 -9485 15995
rect -9515 15970 -9510 15990
rect -9510 15970 -9490 15990
rect -9490 15970 -9485 15990
rect -9515 15965 -9485 15970
rect -9435 15990 -9405 15995
rect -9435 15970 -9430 15990
rect -9430 15970 -9410 15990
rect -9410 15970 -9405 15990
rect -9435 15965 -9405 15970
rect -9355 15990 -9325 15995
rect -9355 15970 -9350 15990
rect -9350 15970 -9330 15990
rect -9330 15970 -9325 15990
rect -9355 15965 -9325 15970
rect -9275 15990 -9245 15995
rect -9275 15970 -9270 15990
rect -9270 15970 -9250 15990
rect -9250 15970 -9245 15990
rect -9275 15965 -9245 15970
rect -9195 15990 -9165 15995
rect -9195 15970 -9190 15990
rect -9190 15970 -9170 15990
rect -9170 15970 -9165 15990
rect -9195 15965 -9165 15970
rect -9115 15990 -9085 15995
rect -9115 15970 -9110 15990
rect -9110 15970 -9090 15990
rect -9090 15970 -9085 15990
rect -9115 15965 -9085 15970
rect -9035 15990 -9005 15995
rect -9035 15970 -9030 15990
rect -9030 15970 -9010 15990
rect -9010 15970 -9005 15990
rect -9035 15965 -9005 15970
rect -8955 15990 -8925 15995
rect -8955 15970 -8950 15990
rect -8950 15970 -8930 15990
rect -8930 15970 -8925 15990
rect -8955 15965 -8925 15970
rect -8875 15990 -8845 15995
rect -8875 15970 -8870 15990
rect -8870 15970 -8850 15990
rect -8850 15970 -8845 15990
rect -8875 15965 -8845 15970
rect -8795 15990 -8765 15995
rect -8795 15970 -8790 15990
rect -8790 15970 -8770 15990
rect -8770 15970 -8765 15990
rect -8795 15965 -8765 15970
rect -8715 15990 -8685 15995
rect -8715 15970 -8710 15990
rect -8710 15970 -8690 15990
rect -8690 15970 -8685 15990
rect -8715 15965 -8685 15970
rect -8635 15990 -8605 15995
rect -8635 15970 -8630 15990
rect -8630 15970 -8610 15990
rect -8610 15970 -8605 15990
rect -8635 15965 -8605 15970
rect -8555 15990 -8525 15995
rect -8555 15970 -8550 15990
rect -8550 15970 -8530 15990
rect -8530 15970 -8525 15990
rect -8555 15965 -8525 15970
rect -8475 15990 -8445 15995
rect -8475 15970 -8470 15990
rect -8470 15970 -8450 15990
rect -8450 15970 -8445 15990
rect -8475 15965 -8445 15970
rect -8395 15990 -8365 15995
rect -8395 15970 -8390 15990
rect -8390 15970 -8370 15990
rect -8370 15970 -8365 15990
rect -8395 15965 -8365 15970
rect -8315 15990 -8285 15995
rect -8315 15970 -8310 15990
rect -8310 15970 -8290 15990
rect -8290 15970 -8285 15990
rect -8315 15965 -8285 15970
rect -8235 15990 -8205 15995
rect -8235 15970 -8230 15990
rect -8230 15970 -8210 15990
rect -8210 15970 -8205 15990
rect -8235 15965 -8205 15970
rect -8155 15990 -8125 15995
rect -8155 15970 -8150 15990
rect -8150 15970 -8130 15990
rect -8130 15970 -8125 15990
rect -8155 15965 -8125 15970
rect -8075 15990 -8045 15995
rect -8075 15970 -8070 15990
rect -8070 15970 -8050 15990
rect -8050 15970 -8045 15990
rect -8075 15965 -8045 15970
rect -7995 15990 -7965 15995
rect -7995 15970 -7990 15990
rect -7990 15970 -7970 15990
rect -7970 15970 -7965 15990
rect -7995 15965 -7965 15970
rect -7915 15990 -7885 15995
rect -7915 15970 -7910 15990
rect -7910 15970 -7890 15990
rect -7890 15970 -7885 15990
rect -7915 15965 -7885 15970
rect -7835 15990 -7805 15995
rect -7835 15970 -7830 15990
rect -7830 15970 -7810 15990
rect -7810 15970 -7805 15990
rect -7835 15965 -7805 15970
rect -7755 15990 -7725 15995
rect -7755 15970 -7750 15990
rect -7750 15970 -7730 15990
rect -7730 15970 -7725 15990
rect -7755 15965 -7725 15970
rect -7675 15990 -7645 15995
rect -7675 15970 -7670 15990
rect -7670 15970 -7650 15990
rect -7650 15970 -7645 15990
rect -7675 15965 -7645 15970
rect -7595 15990 -7565 15995
rect -7595 15970 -7590 15990
rect -7590 15970 -7570 15990
rect -7570 15970 -7565 15990
rect -7595 15965 -7565 15970
rect -7515 15990 -7485 15995
rect -7515 15970 -7510 15990
rect -7510 15970 -7490 15990
rect -7490 15970 -7485 15990
rect -7515 15965 -7485 15970
rect -7435 15990 -7405 15995
rect -7435 15970 -7430 15990
rect -7430 15970 -7410 15990
rect -7410 15970 -7405 15990
rect -7435 15965 -7405 15970
rect -7355 15990 -7325 15995
rect -7355 15970 -7350 15990
rect -7350 15970 -7330 15990
rect -7330 15970 -7325 15990
rect -7355 15965 -7325 15970
rect -7275 15990 -7245 15995
rect -7275 15970 -7270 15990
rect -7270 15970 -7250 15990
rect -7250 15970 -7245 15990
rect -7275 15965 -7245 15970
rect -7195 15990 -7165 15995
rect -7195 15970 -7190 15990
rect -7190 15970 -7170 15990
rect -7170 15970 -7165 15990
rect -7195 15965 -7165 15970
rect -7115 15990 -7085 15995
rect -7115 15970 -7110 15990
rect -7110 15970 -7090 15990
rect -7090 15970 -7085 15990
rect -7115 15965 -7085 15970
rect -7035 15990 -7005 15995
rect -7035 15970 -7030 15990
rect -7030 15970 -7010 15990
rect -7010 15970 -7005 15990
rect -7035 15965 -7005 15970
rect -6955 15990 -6925 15995
rect -6955 15970 -6950 15990
rect -6950 15970 -6930 15990
rect -6930 15970 -6925 15990
rect -6955 15965 -6925 15970
rect -6875 15990 -6845 15995
rect -6875 15970 -6870 15990
rect -6870 15970 -6850 15990
rect -6850 15970 -6845 15990
rect -6875 15965 -6845 15970
rect -6795 15990 -6765 15995
rect -6795 15970 -6790 15990
rect -6790 15970 -6770 15990
rect -6770 15970 -6765 15990
rect -6795 15965 -6765 15970
rect -6715 15990 -6685 15995
rect -6715 15970 -6710 15990
rect -6710 15970 -6690 15990
rect -6690 15970 -6685 15990
rect -6715 15965 -6685 15970
rect -6635 15990 -6605 15995
rect -6635 15970 -6630 15990
rect -6630 15970 -6610 15990
rect -6610 15970 -6605 15990
rect -6635 15965 -6605 15970
rect -6555 15990 -6525 15995
rect -6555 15970 -6550 15990
rect -6550 15970 -6530 15990
rect -6530 15970 -6525 15990
rect -6555 15965 -6525 15970
rect -6475 15990 -6445 15995
rect -6475 15970 -6470 15990
rect -6470 15970 -6450 15990
rect -6450 15970 -6445 15990
rect -6475 15965 -6445 15970
rect -6395 15990 -6365 15995
rect -6395 15970 -6390 15990
rect -6390 15970 -6370 15990
rect -6370 15970 -6365 15990
rect -6395 15965 -6365 15970
rect -6315 15990 -6285 15995
rect -6315 15970 -6310 15990
rect -6310 15970 -6290 15990
rect -6290 15970 -6285 15990
rect -6315 15965 -6285 15970
rect -6235 15990 -6205 15995
rect -6235 15970 -6230 15990
rect -6230 15970 -6210 15990
rect -6210 15970 -6205 15990
rect -6235 15965 -6205 15970
rect -6155 15990 -6125 15995
rect -6155 15970 -6150 15990
rect -6150 15970 -6130 15990
rect -6130 15970 -6125 15990
rect -6155 15965 -6125 15970
rect -6075 15990 -6045 15995
rect -6075 15970 -6070 15990
rect -6070 15970 -6050 15990
rect -6050 15970 -6045 15990
rect -6075 15965 -6045 15970
rect -5995 15990 -5965 15995
rect -5995 15970 -5990 15990
rect -5990 15970 -5970 15990
rect -5970 15970 -5965 15990
rect -5995 15965 -5965 15970
rect -5915 15990 -5885 15995
rect -5915 15970 -5910 15990
rect -5910 15970 -5890 15990
rect -5890 15970 -5885 15990
rect -5915 15965 -5885 15970
rect -5835 15990 -5805 15995
rect -5835 15970 -5830 15990
rect -5830 15970 -5810 15990
rect -5810 15970 -5805 15990
rect -5835 15965 -5805 15970
rect -5755 15990 -5725 15995
rect -5755 15970 -5750 15990
rect -5750 15970 -5730 15990
rect -5730 15970 -5725 15990
rect -5755 15965 -5725 15970
rect -5675 15990 -5645 15995
rect -5675 15970 -5670 15990
rect -5670 15970 -5650 15990
rect -5650 15970 -5645 15990
rect -5675 15965 -5645 15970
rect -5595 15990 -5565 15995
rect -5595 15970 -5590 15990
rect -5590 15970 -5570 15990
rect -5570 15970 -5565 15990
rect -5595 15965 -5565 15970
rect -5435 15990 -5405 15995
rect -5435 15970 -5430 15990
rect -5430 15970 -5410 15990
rect -5410 15970 -5405 15990
rect -5435 15965 -5405 15970
rect -5355 15990 -5325 15995
rect -5355 15970 -5350 15990
rect -5350 15970 -5330 15990
rect -5330 15970 -5325 15990
rect -5355 15965 -5325 15970
rect -5275 15990 -5245 15995
rect -5275 15970 -5270 15990
rect -5270 15970 -5250 15990
rect -5250 15970 -5245 15990
rect -5275 15965 -5245 15970
rect -5195 15990 -5165 15995
rect -5195 15970 -5190 15990
rect -5190 15970 -5170 15990
rect -5170 15970 -5165 15990
rect -5195 15965 -5165 15970
rect -5115 15990 -5085 15995
rect -5115 15970 -5110 15990
rect -5110 15970 -5090 15990
rect -5090 15970 -5085 15990
rect -5115 15965 -5085 15970
rect -5035 15990 -5005 15995
rect -5035 15970 -5030 15990
rect -5030 15970 -5010 15990
rect -5010 15970 -5005 15990
rect -5035 15965 -5005 15970
rect -4955 15990 -4925 15995
rect -4955 15970 -4950 15990
rect -4950 15970 -4930 15990
rect -4930 15970 -4925 15990
rect -4955 15965 -4925 15970
rect -4875 15990 -4845 15995
rect -4875 15970 -4870 15990
rect -4870 15970 -4850 15990
rect -4850 15970 -4845 15990
rect -4875 15965 -4845 15970
rect -4795 15990 -4765 15995
rect -4795 15970 -4790 15990
rect -4790 15970 -4770 15990
rect -4770 15970 -4765 15990
rect -4795 15965 -4765 15970
rect -4715 15990 -4685 15995
rect -4715 15970 -4710 15990
rect -4710 15970 -4690 15990
rect -4690 15970 -4685 15990
rect -4715 15965 -4685 15970
rect -4635 15990 -4605 15995
rect -4635 15970 -4630 15990
rect -4630 15970 -4610 15990
rect -4610 15970 -4605 15990
rect -4635 15965 -4605 15970
rect -4555 15990 -4525 15995
rect -4555 15970 -4550 15990
rect -4550 15970 -4530 15990
rect -4530 15970 -4525 15990
rect -4555 15965 -4525 15970
rect -4475 15990 -4445 15995
rect -4475 15970 -4470 15990
rect -4470 15970 -4450 15990
rect -4450 15970 -4445 15990
rect -4475 15965 -4445 15970
rect -4395 15990 -4365 15995
rect -4395 15970 -4390 15990
rect -4390 15970 -4370 15990
rect -4370 15970 -4365 15990
rect -4395 15965 -4365 15970
rect -4315 15990 -4285 15995
rect -4315 15970 -4310 15990
rect -4310 15970 -4290 15990
rect -4290 15970 -4285 15990
rect -4315 15965 -4285 15970
rect -4235 15990 -4205 15995
rect -4235 15970 -4230 15990
rect -4230 15970 -4210 15990
rect -4210 15970 -4205 15990
rect -4235 15965 -4205 15970
rect -4155 15990 -4125 15995
rect -4155 15970 -4150 15990
rect -4150 15970 -4130 15990
rect -4130 15970 -4125 15990
rect -4155 15965 -4125 15970
rect -4075 15990 -4045 15995
rect -4075 15970 -4070 15990
rect -4070 15970 -4050 15990
rect -4050 15970 -4045 15990
rect -4075 15965 -4045 15970
rect -3995 15990 -3965 15995
rect -3995 15970 -3990 15990
rect -3990 15970 -3970 15990
rect -3970 15970 -3965 15990
rect -3995 15965 -3965 15970
rect -3915 15990 -3885 15995
rect -3915 15970 -3910 15990
rect -3910 15970 -3890 15990
rect -3890 15970 -3885 15990
rect -3915 15965 -3885 15970
rect -3835 15990 -3805 15995
rect -3835 15970 -3830 15990
rect -3830 15970 -3810 15990
rect -3810 15970 -3805 15990
rect -3835 15965 -3805 15970
rect -3755 15990 -3725 15995
rect -3755 15970 -3750 15990
rect -3750 15970 -3730 15990
rect -3730 15970 -3725 15990
rect -3755 15965 -3725 15970
rect -3675 15990 -3645 15995
rect -3675 15970 -3670 15990
rect -3670 15970 -3650 15990
rect -3650 15970 -3645 15990
rect -3675 15965 -3645 15970
rect -3595 15990 -3565 15995
rect -3595 15970 -3590 15990
rect -3590 15970 -3570 15990
rect -3570 15970 -3565 15990
rect -3595 15965 -3565 15970
rect -3515 15990 -3485 15995
rect -3515 15970 -3510 15990
rect -3510 15970 -3490 15990
rect -3490 15970 -3485 15990
rect -3515 15965 -3485 15970
rect -3435 15990 -3405 15995
rect -3435 15970 -3430 15990
rect -3430 15970 -3410 15990
rect -3410 15970 -3405 15990
rect -3435 15965 -3405 15970
rect -3355 15990 -3325 15995
rect -3355 15970 -3350 15990
rect -3350 15970 -3330 15990
rect -3330 15970 -3325 15990
rect -3355 15965 -3325 15970
rect -3275 15990 -3245 15995
rect -3275 15970 -3270 15990
rect -3270 15970 -3250 15990
rect -3250 15970 -3245 15990
rect -3275 15965 -3245 15970
rect -3195 15990 -3165 15995
rect -3195 15970 -3190 15990
rect -3190 15970 -3170 15990
rect -3170 15970 -3165 15990
rect -3195 15965 -3165 15970
rect -3115 15990 -3085 15995
rect -3115 15970 -3110 15990
rect -3110 15970 -3090 15990
rect -3090 15970 -3085 15990
rect -3115 15965 -3085 15970
rect -3035 15990 -3005 15995
rect -3035 15970 -3030 15990
rect -3030 15970 -3010 15990
rect -3010 15970 -3005 15990
rect -3035 15965 -3005 15970
rect -2955 15990 -2925 15995
rect -2955 15970 -2950 15990
rect -2950 15970 -2930 15990
rect -2930 15970 -2925 15990
rect -2955 15965 -2925 15970
rect -2875 15990 -2845 15995
rect -2875 15970 -2870 15990
rect -2870 15970 -2850 15990
rect -2850 15970 -2845 15990
rect -2875 15965 -2845 15970
rect -2795 15990 -2765 15995
rect -2795 15970 -2790 15990
rect -2790 15970 -2770 15990
rect -2770 15970 -2765 15990
rect -2795 15965 -2765 15970
rect -2715 15990 -2685 15995
rect -2715 15970 -2710 15990
rect -2710 15970 -2690 15990
rect -2690 15970 -2685 15990
rect -2715 15965 -2685 15970
rect -2635 15990 -2605 15995
rect -2635 15970 -2630 15990
rect -2630 15970 -2610 15990
rect -2610 15970 -2605 15990
rect -2635 15965 -2605 15970
rect -2555 15990 -2525 15995
rect -2555 15970 -2550 15990
rect -2550 15970 -2530 15990
rect -2530 15970 -2525 15990
rect -2555 15965 -2525 15970
rect -2475 15990 -2445 15995
rect -2475 15970 -2470 15990
rect -2470 15970 -2450 15990
rect -2450 15970 -2445 15990
rect -2475 15965 -2445 15970
rect -2395 15990 -2365 15995
rect -2395 15970 -2390 15990
rect -2390 15970 -2370 15990
rect -2370 15970 -2365 15990
rect -2395 15965 -2365 15970
rect -2315 15990 -2285 15995
rect -2315 15970 -2310 15990
rect -2310 15970 -2290 15990
rect -2290 15970 -2285 15990
rect -2315 15965 -2285 15970
rect -2235 15990 -2205 15995
rect -2235 15970 -2230 15990
rect -2230 15970 -2210 15990
rect -2210 15970 -2205 15990
rect -2235 15965 -2205 15970
rect -2155 15990 -2125 15995
rect -2155 15970 -2150 15990
rect -2150 15970 -2130 15990
rect -2130 15970 -2125 15990
rect -2155 15965 -2125 15970
rect -2075 15990 -2045 15995
rect -2075 15970 -2070 15990
rect -2070 15970 -2050 15990
rect -2050 15970 -2045 15990
rect -2075 15965 -2045 15970
rect -1995 15990 -1965 15995
rect -1995 15970 -1990 15990
rect -1990 15970 -1970 15990
rect -1970 15970 -1965 15990
rect -1995 15965 -1965 15970
rect -1835 15990 -1805 15995
rect -1835 15970 -1830 15990
rect -1830 15970 -1810 15990
rect -1810 15970 -1805 15990
rect -1835 15965 -1805 15970
rect -1755 15990 -1725 15995
rect -1755 15970 -1750 15990
rect -1750 15970 -1730 15990
rect -1730 15970 -1725 15990
rect -1755 15965 -1725 15970
rect -1675 15990 -1645 15995
rect -1675 15970 -1670 15990
rect -1670 15970 -1650 15990
rect -1650 15970 -1645 15990
rect -1675 15965 -1645 15970
rect -1595 15990 -1565 15995
rect -1595 15970 -1590 15990
rect -1590 15970 -1570 15990
rect -1570 15970 -1565 15990
rect -1595 15965 -1565 15970
rect -1515 15990 -1485 15995
rect -1515 15970 -1510 15990
rect -1510 15970 -1490 15990
rect -1490 15970 -1485 15990
rect -1515 15965 -1485 15970
rect -1435 15990 -1405 15995
rect -1435 15970 -1430 15990
rect -1430 15970 -1410 15990
rect -1410 15970 -1405 15990
rect -1435 15965 -1405 15970
rect -1355 15990 -1325 15995
rect -1355 15970 -1350 15990
rect -1350 15970 -1330 15990
rect -1330 15970 -1325 15990
rect -1355 15965 -1325 15970
rect -1195 15990 -1165 15995
rect -1195 15970 -1190 15990
rect -1190 15970 -1170 15990
rect -1170 15970 -1165 15990
rect -1195 15965 -1165 15970
rect -1035 15990 -1005 15995
rect -1035 15970 -1030 15990
rect -1030 15970 -1010 15990
rect -1010 15970 -1005 15990
rect -1035 15965 -1005 15970
rect -875 15990 -845 15995
rect -875 15970 -870 15990
rect -870 15970 -850 15990
rect -850 15970 -845 15990
rect -875 15965 -845 15970
rect -715 15990 -685 15995
rect -715 15970 -710 15990
rect -710 15970 -690 15990
rect -690 15970 -685 15990
rect -715 15965 -685 15970
rect -555 15990 -525 15995
rect -555 15970 -550 15990
rect -550 15970 -530 15990
rect -530 15970 -525 15990
rect -555 15965 -525 15970
<< metal2 >>
rect -15520 21435 -520 21440
rect -15520 21405 -15515 21435
rect -15485 21405 -15355 21435
rect -15325 21405 -15195 21435
rect -15165 21405 -15035 21435
rect -15005 21405 -14955 21435
rect -14925 21405 -14875 21435
rect -14845 21405 -14795 21435
rect -14765 21405 -14715 21435
rect -14685 21405 -14635 21435
rect -14605 21405 -14555 21435
rect -14525 21405 -14475 21435
rect -14445 21405 -14395 21435
rect -14365 21405 -14315 21435
rect -14285 21405 -14235 21435
rect -14205 21405 -14155 21435
rect -14125 21405 -14075 21435
rect -14045 21405 -13995 21435
rect -13965 21405 -13915 21435
rect -13885 21405 -13835 21435
rect -13805 21405 -13755 21435
rect -13725 21405 -13675 21435
rect -13645 21405 -13595 21435
rect -13565 21405 -13515 21435
rect -13485 21405 -13435 21435
rect -13405 21405 -13355 21435
rect -13325 21405 -13275 21435
rect -13245 21405 -13195 21435
rect -13165 21405 -13115 21435
rect -13085 21405 -13035 21435
rect -13005 21405 -12955 21435
rect -12925 21405 -12875 21435
rect -12845 21405 -12795 21435
rect -12765 21405 -12715 21435
rect -12685 21405 -12635 21435
rect -12605 21405 -12555 21435
rect -12525 21405 -12475 21435
rect -12445 21405 -12395 21435
rect -12365 21405 -12315 21435
rect -12285 21405 -12235 21435
rect -12205 21405 -12155 21435
rect -12125 21405 -12075 21435
rect -12045 21405 -11995 21435
rect -11965 21405 -11915 21435
rect -11885 21405 -11835 21435
rect -11805 21405 -11755 21435
rect -11725 21405 -11675 21435
rect -11645 21405 -11595 21435
rect -11565 21405 -11515 21435
rect -11485 21405 -11435 21435
rect -11405 21405 -11355 21435
rect -11325 21405 -11275 21435
rect -11245 21405 -11195 21435
rect -11165 21405 -11115 21435
rect -11085 21405 -11035 21435
rect -11005 21405 -10955 21435
rect -10925 21405 -10875 21435
rect -10845 21405 -10795 21435
rect -10765 21405 -10715 21435
rect -10685 21405 -10635 21435
rect -10605 21405 -10555 21435
rect -10525 21405 -10475 21435
rect -10445 21405 -10395 21435
rect -10365 21405 -10315 21435
rect -10285 21405 -10235 21435
rect -10205 21405 -10155 21435
rect -10125 21405 -10075 21435
rect -10045 21405 -9995 21435
rect -9965 21405 -9915 21435
rect -9885 21405 -9835 21435
rect -9805 21405 -9755 21435
rect -9725 21405 -9675 21435
rect -9645 21405 -9595 21435
rect -9565 21405 -9515 21435
rect -9485 21405 -9435 21435
rect -9405 21405 -9355 21435
rect -9325 21405 -9275 21435
rect -9245 21405 -9195 21435
rect -9165 21405 -9115 21435
rect -9085 21405 -9035 21435
rect -9005 21405 -8955 21435
rect -8925 21405 -8875 21435
rect -8845 21405 -8795 21435
rect -8765 21405 -8715 21435
rect -8685 21405 -8635 21435
rect -8605 21405 -8555 21435
rect -8525 21405 -8475 21435
rect -8445 21405 -8395 21435
rect -8365 21405 -8315 21435
rect -8285 21405 -8235 21435
rect -8205 21405 -8155 21435
rect -8125 21405 -8075 21435
rect -8045 21405 -7995 21435
rect -7965 21405 -7915 21435
rect -7885 21405 -7835 21435
rect -7805 21405 -7755 21435
rect -7725 21405 -7675 21435
rect -7645 21405 -7595 21435
rect -7565 21405 -7515 21435
rect -7485 21405 -7435 21435
rect -7405 21405 -7355 21435
rect -7325 21405 -7275 21435
rect -7245 21405 -7195 21435
rect -7165 21405 -7115 21435
rect -7085 21405 -7035 21435
rect -7005 21405 -6955 21435
rect -6925 21405 -6875 21435
rect -6845 21405 -6795 21435
rect -6765 21405 -6715 21435
rect -6685 21405 -6635 21435
rect -6605 21405 -6555 21435
rect -6525 21405 -6475 21435
rect -6445 21405 -6395 21435
rect -6365 21405 -6315 21435
rect -6285 21405 -6235 21435
rect -6205 21405 -6155 21435
rect -6125 21405 -6075 21435
rect -6045 21405 -5915 21435
rect -5885 21405 -5755 21435
rect -5725 21405 -5675 21435
rect -5645 21405 -5595 21435
rect -5565 21405 -5515 21435
rect -5485 21405 -5435 21435
rect -5405 21405 -5355 21435
rect -5325 21405 -5275 21435
rect -5245 21405 -5195 21435
rect -5165 21405 -5115 21435
rect -5085 21405 -5035 21435
rect -5005 21405 -4955 21435
rect -4925 21405 -4875 21435
rect -4845 21405 -4795 21435
rect -4765 21405 -4715 21435
rect -4685 21405 -4635 21435
rect -4605 21405 -4555 21435
rect -4525 21405 -4475 21435
rect -4445 21405 -4395 21435
rect -4365 21405 -4315 21435
rect -4285 21405 -4235 21435
rect -4205 21405 -4155 21435
rect -4125 21405 -4075 21435
rect -4045 21405 -3995 21435
rect -3965 21405 -3915 21435
rect -3885 21405 -3835 21435
rect -3805 21405 -3755 21435
rect -3725 21405 -3675 21435
rect -3645 21405 -3595 21435
rect -3565 21405 -3515 21435
rect -3485 21405 -3435 21435
rect -3405 21405 -3355 21435
rect -3325 21405 -3275 21435
rect -3245 21405 -3195 21435
rect -3165 21405 -3115 21435
rect -3085 21405 -3035 21435
rect -3005 21405 -2955 21435
rect -2925 21405 -2875 21435
rect -2845 21405 -2795 21435
rect -2765 21405 -2715 21435
rect -2685 21405 -2635 21435
rect -2605 21405 -2555 21435
rect -2525 21405 -2475 21435
rect -2445 21405 -2395 21435
rect -2365 21405 -2315 21435
rect -2285 21405 -2235 21435
rect -2205 21405 -2155 21435
rect -2125 21405 -2075 21435
rect -2045 21405 -1995 21435
rect -1965 21405 -1835 21435
rect -1805 21405 -1755 21435
rect -1725 21405 -1675 21435
rect -1645 21405 -1595 21435
rect -1565 21405 -1515 21435
rect -1485 21405 -1355 21435
rect -1325 21405 -1275 21435
rect -1245 21405 -1195 21435
rect -1165 21405 -1115 21435
rect -1085 21405 -1035 21435
rect -1005 21405 -875 21435
rect -845 21405 -715 21435
rect -685 21405 -555 21435
rect -525 21405 -520 21435
rect -15520 21400 -520 21405
rect -15520 21355 -15160 21360
rect -15520 21325 -15515 21355
rect -15485 21325 -15355 21355
rect -15325 21325 -15195 21355
rect -15165 21325 -15160 21355
rect -15520 21320 -15160 21325
rect -15120 21355 -1400 21360
rect -15120 21325 -15115 21355
rect -15085 21325 -5995 21355
rect -5965 21325 -1435 21355
rect -1405 21325 -1400 21355
rect -15120 21320 -1400 21325
rect -1360 21320 -1320 21360
rect -1280 21320 -1240 21360
rect -1200 21320 -1160 21360
rect -1120 21320 -1080 21360
rect -1040 21320 -1000 21360
rect -880 21320 -840 21360
rect -720 21320 -680 21360
rect -560 21320 -520 21360
rect -15520 21275 -520 21280
rect -15520 21245 -15515 21275
rect -15485 21245 -15355 21275
rect -15325 21245 -15195 21275
rect -15165 21245 -15035 21275
rect -15005 21245 -14955 21275
rect -14925 21245 -14875 21275
rect -14845 21245 -14795 21275
rect -14765 21245 -14715 21275
rect -14685 21245 -14635 21275
rect -14605 21245 -14555 21275
rect -14525 21245 -14475 21275
rect -14445 21245 -14395 21275
rect -14365 21245 -14315 21275
rect -14285 21245 -14235 21275
rect -14205 21245 -14155 21275
rect -14125 21245 -14075 21275
rect -14045 21245 -13995 21275
rect -13965 21245 -13915 21275
rect -13885 21245 -13835 21275
rect -13805 21245 -13755 21275
rect -13725 21245 -13675 21275
rect -13645 21245 -13595 21275
rect -13565 21245 -13515 21275
rect -13485 21245 -13435 21275
rect -13405 21245 -13355 21275
rect -13325 21245 -13275 21275
rect -13245 21245 -13195 21275
rect -13165 21245 -13115 21275
rect -13085 21245 -13035 21275
rect -13005 21245 -12955 21275
rect -12925 21245 -12875 21275
rect -12845 21245 -12795 21275
rect -12765 21245 -12715 21275
rect -12685 21245 -12635 21275
rect -12605 21245 -12555 21275
rect -12525 21245 -12475 21275
rect -12445 21245 -12395 21275
rect -12365 21245 -12315 21275
rect -12285 21245 -12235 21275
rect -12205 21245 -12155 21275
rect -12125 21245 -12075 21275
rect -12045 21245 -11995 21275
rect -11965 21245 -11915 21275
rect -11885 21245 -11835 21275
rect -11805 21245 -11755 21275
rect -11725 21245 -11675 21275
rect -11645 21245 -11595 21275
rect -11565 21245 -11515 21275
rect -11485 21245 -11435 21275
rect -11405 21245 -11355 21275
rect -11325 21245 -11275 21275
rect -11245 21245 -11195 21275
rect -11165 21245 -11115 21275
rect -11085 21245 -11035 21275
rect -11005 21245 -10955 21275
rect -10925 21245 -10875 21275
rect -10845 21245 -10795 21275
rect -10765 21245 -10715 21275
rect -10685 21245 -10635 21275
rect -10605 21245 -10555 21275
rect -10525 21245 -10475 21275
rect -10445 21245 -10395 21275
rect -10365 21245 -10315 21275
rect -10285 21245 -10235 21275
rect -10205 21245 -10155 21275
rect -10125 21245 -10075 21275
rect -10045 21245 -9995 21275
rect -9965 21245 -9915 21275
rect -9885 21245 -9835 21275
rect -9805 21245 -9755 21275
rect -9725 21245 -9675 21275
rect -9645 21245 -9595 21275
rect -9565 21245 -9515 21275
rect -9485 21245 -9435 21275
rect -9405 21245 -9355 21275
rect -9325 21245 -9275 21275
rect -9245 21245 -9195 21275
rect -9165 21245 -9115 21275
rect -9085 21245 -9035 21275
rect -9005 21245 -8955 21275
rect -8925 21245 -8875 21275
rect -8845 21245 -8795 21275
rect -8765 21245 -8715 21275
rect -8685 21245 -8635 21275
rect -8605 21245 -8555 21275
rect -8525 21245 -8475 21275
rect -8445 21245 -8395 21275
rect -8365 21245 -8315 21275
rect -8285 21245 -8235 21275
rect -8205 21245 -8155 21275
rect -8125 21245 -8075 21275
rect -8045 21245 -7995 21275
rect -7965 21245 -7915 21275
rect -7885 21245 -7835 21275
rect -7805 21245 -7755 21275
rect -7725 21245 -7675 21275
rect -7645 21245 -7595 21275
rect -7565 21245 -7515 21275
rect -7485 21245 -7435 21275
rect -7405 21245 -7355 21275
rect -7325 21245 -7275 21275
rect -7245 21245 -7195 21275
rect -7165 21245 -7115 21275
rect -7085 21245 -7035 21275
rect -7005 21245 -6955 21275
rect -6925 21245 -6875 21275
rect -6845 21245 -6795 21275
rect -6765 21245 -6715 21275
rect -6685 21245 -6635 21275
rect -6605 21245 -6555 21275
rect -6525 21245 -6475 21275
rect -6445 21245 -6395 21275
rect -6365 21245 -6315 21275
rect -6285 21245 -6235 21275
rect -6205 21245 -6155 21275
rect -6125 21245 -6075 21275
rect -6045 21245 -5915 21275
rect -5885 21245 -5755 21275
rect -5725 21245 -5675 21275
rect -5645 21245 -5595 21275
rect -5565 21245 -5515 21275
rect -5485 21245 -5435 21275
rect -5405 21245 -5355 21275
rect -5325 21245 -5275 21275
rect -5245 21245 -5195 21275
rect -5165 21245 -5115 21275
rect -5085 21245 -5035 21275
rect -5005 21245 -4955 21275
rect -4925 21245 -4875 21275
rect -4845 21245 -4795 21275
rect -4765 21245 -4715 21275
rect -4685 21245 -4635 21275
rect -4605 21245 -4555 21275
rect -4525 21245 -4475 21275
rect -4445 21245 -4395 21275
rect -4365 21245 -4315 21275
rect -4285 21245 -4235 21275
rect -4205 21245 -4155 21275
rect -4125 21245 -4075 21275
rect -4045 21245 -3995 21275
rect -3965 21245 -3915 21275
rect -3885 21245 -3835 21275
rect -3805 21245 -3755 21275
rect -3725 21245 -3675 21275
rect -3645 21245 -3595 21275
rect -3565 21245 -3515 21275
rect -3485 21245 -3435 21275
rect -3405 21245 -3355 21275
rect -3325 21245 -3275 21275
rect -3245 21245 -3195 21275
rect -3165 21245 -3115 21275
rect -3085 21245 -3035 21275
rect -3005 21245 -2955 21275
rect -2925 21245 -2875 21275
rect -2845 21245 -2795 21275
rect -2765 21245 -2715 21275
rect -2685 21245 -2635 21275
rect -2605 21245 -2555 21275
rect -2525 21245 -2475 21275
rect -2445 21245 -2395 21275
rect -2365 21245 -2315 21275
rect -2285 21245 -2235 21275
rect -2205 21245 -2155 21275
rect -2125 21245 -2075 21275
rect -2045 21245 -1995 21275
rect -1965 21245 -1835 21275
rect -1805 21245 -1755 21275
rect -1725 21245 -1675 21275
rect -1645 21245 -1595 21275
rect -1565 21245 -1515 21275
rect -1485 21245 -1355 21275
rect -1325 21245 -1275 21275
rect -1245 21245 -1195 21275
rect -1165 21245 -1115 21275
rect -1085 21245 -1035 21275
rect -1005 21245 -875 21275
rect -845 21245 -715 21275
rect -685 21245 -555 21275
rect -525 21245 -520 21275
rect -15520 21240 -520 21245
rect -15520 21195 -15320 21200
rect -15520 21165 -15515 21195
rect -15485 21165 -15355 21195
rect -15325 21165 -15320 21195
rect -15520 21160 -15320 21165
rect -15280 21195 -1560 21200
rect -15280 21165 -15275 21195
rect -15245 21165 -5835 21195
rect -5805 21165 -1595 21195
rect -1565 21165 -1560 21195
rect -15280 21160 -1560 21165
rect -1520 21160 -1480 21200
rect -1360 21160 -1320 21200
rect -1280 21160 -1240 21200
rect -1200 21160 -1160 21200
rect -1120 21160 -1080 21200
rect -1040 21160 -1000 21200
rect -880 21160 -840 21200
rect -720 21160 -680 21200
rect -560 21160 -520 21200
rect -15520 21115 -520 21120
rect -15520 21085 -15515 21115
rect -15485 21085 -15355 21115
rect -15325 21085 -15195 21115
rect -15165 21085 -15035 21115
rect -15005 21085 -14955 21115
rect -14925 21085 -14875 21115
rect -14845 21085 -14795 21115
rect -14765 21085 -14715 21115
rect -14685 21085 -14635 21115
rect -14605 21085 -14555 21115
rect -14525 21085 -14475 21115
rect -14445 21085 -14395 21115
rect -14365 21085 -14315 21115
rect -14285 21085 -14235 21115
rect -14205 21085 -14155 21115
rect -14125 21085 -14075 21115
rect -14045 21085 -13995 21115
rect -13965 21085 -13915 21115
rect -13885 21085 -13835 21115
rect -13805 21085 -13755 21115
rect -13725 21085 -13675 21115
rect -13645 21085 -13595 21115
rect -13565 21085 -13515 21115
rect -13485 21085 -13435 21115
rect -13405 21085 -13355 21115
rect -13325 21085 -13275 21115
rect -13245 21085 -13195 21115
rect -13165 21085 -13115 21115
rect -13085 21085 -13035 21115
rect -13005 21085 -12955 21115
rect -12925 21085 -12875 21115
rect -12845 21085 -12795 21115
rect -12765 21085 -12715 21115
rect -12685 21085 -12635 21115
rect -12605 21085 -12555 21115
rect -12525 21085 -12475 21115
rect -12445 21085 -12395 21115
rect -12365 21085 -12315 21115
rect -12285 21085 -12235 21115
rect -12205 21085 -12155 21115
rect -12125 21085 -12075 21115
rect -12045 21085 -11995 21115
rect -11965 21085 -11915 21115
rect -11885 21085 -11835 21115
rect -11805 21085 -11755 21115
rect -11725 21085 -11675 21115
rect -11645 21085 -11595 21115
rect -11565 21085 -11515 21115
rect -11485 21085 -11435 21115
rect -11405 21085 -11355 21115
rect -11325 21085 -11275 21115
rect -11245 21085 -11195 21115
rect -11165 21085 -11115 21115
rect -11085 21085 -11035 21115
rect -11005 21085 -10955 21115
rect -10925 21085 -10875 21115
rect -10845 21085 -10795 21115
rect -10765 21085 -10715 21115
rect -10685 21085 -10635 21115
rect -10605 21085 -10555 21115
rect -10525 21085 -10475 21115
rect -10445 21085 -10395 21115
rect -10365 21085 -10315 21115
rect -10285 21085 -10235 21115
rect -10205 21085 -10155 21115
rect -10125 21085 -10075 21115
rect -10045 21085 -9995 21115
rect -9965 21085 -9915 21115
rect -9885 21085 -9835 21115
rect -9805 21085 -9755 21115
rect -9725 21085 -9675 21115
rect -9645 21085 -9595 21115
rect -9565 21085 -9515 21115
rect -9485 21085 -9435 21115
rect -9405 21085 -9355 21115
rect -9325 21085 -9275 21115
rect -9245 21085 -9195 21115
rect -9165 21085 -9115 21115
rect -9085 21085 -9035 21115
rect -9005 21085 -8955 21115
rect -8925 21085 -8875 21115
rect -8845 21085 -8795 21115
rect -8765 21085 -8715 21115
rect -8685 21085 -8635 21115
rect -8605 21085 -8555 21115
rect -8525 21085 -8475 21115
rect -8445 21085 -8395 21115
rect -8365 21085 -8315 21115
rect -8285 21085 -8235 21115
rect -8205 21085 -8155 21115
rect -8125 21085 -8075 21115
rect -8045 21085 -7995 21115
rect -7965 21085 -7915 21115
rect -7885 21085 -7835 21115
rect -7805 21085 -7755 21115
rect -7725 21085 -7675 21115
rect -7645 21085 -7595 21115
rect -7565 21085 -7515 21115
rect -7485 21085 -7435 21115
rect -7405 21085 -7355 21115
rect -7325 21085 -7275 21115
rect -7245 21085 -7195 21115
rect -7165 21085 -7115 21115
rect -7085 21085 -7035 21115
rect -7005 21085 -6955 21115
rect -6925 21085 -6875 21115
rect -6845 21085 -6795 21115
rect -6765 21085 -6715 21115
rect -6685 21085 -6635 21115
rect -6605 21085 -6555 21115
rect -6525 21085 -6475 21115
rect -6445 21085 -6395 21115
rect -6365 21085 -6315 21115
rect -6285 21085 -6235 21115
rect -6205 21085 -6155 21115
rect -6125 21085 -6075 21115
rect -6045 21085 -5915 21115
rect -5885 21085 -5755 21115
rect -5725 21085 -5675 21115
rect -5645 21085 -5595 21115
rect -5565 21085 -5515 21115
rect -5485 21085 -5435 21115
rect -5405 21085 -5355 21115
rect -5325 21085 -5275 21115
rect -5245 21085 -5195 21115
rect -5165 21085 -5115 21115
rect -5085 21085 -5035 21115
rect -5005 21085 -4955 21115
rect -4925 21085 -4875 21115
rect -4845 21085 -4795 21115
rect -4765 21085 -4715 21115
rect -4685 21085 -4635 21115
rect -4605 21085 -4555 21115
rect -4525 21085 -4475 21115
rect -4445 21085 -4395 21115
rect -4365 21085 -4315 21115
rect -4285 21085 -4235 21115
rect -4205 21085 -4155 21115
rect -4125 21085 -4075 21115
rect -4045 21085 -3995 21115
rect -3965 21085 -3915 21115
rect -3885 21085 -3835 21115
rect -3805 21085 -3755 21115
rect -3725 21085 -3675 21115
rect -3645 21085 -3595 21115
rect -3565 21085 -3515 21115
rect -3485 21085 -3435 21115
rect -3405 21085 -3355 21115
rect -3325 21085 -3275 21115
rect -3245 21085 -3195 21115
rect -3165 21085 -3115 21115
rect -3085 21085 -3035 21115
rect -3005 21085 -2955 21115
rect -2925 21085 -2875 21115
rect -2845 21085 -2795 21115
rect -2765 21085 -2715 21115
rect -2685 21085 -2635 21115
rect -2605 21085 -2555 21115
rect -2525 21085 -2475 21115
rect -2445 21085 -2395 21115
rect -2365 21085 -2315 21115
rect -2285 21085 -2235 21115
rect -2205 21085 -2155 21115
rect -2125 21085 -2075 21115
rect -2045 21085 -1995 21115
rect -1965 21085 -1835 21115
rect -1805 21085 -1755 21115
rect -1725 21085 -1675 21115
rect -1645 21085 -1515 21115
rect -1485 21085 -1355 21115
rect -1325 21085 -1275 21115
rect -1245 21085 -1195 21115
rect -1165 21085 -1115 21115
rect -1085 21085 -1035 21115
rect -1005 21085 -875 21115
rect -845 21085 -715 21115
rect -685 21085 -555 21115
rect -525 21085 -520 21115
rect -15520 21080 -520 21085
rect -15520 21035 -15160 21040
rect -15520 21005 -15515 21035
rect -15485 21005 -15355 21035
rect -15325 21005 -15195 21035
rect -15165 21005 -15160 21035
rect -15520 21000 -15160 21005
rect -15120 21035 -600 21040
rect -15120 21005 -15115 21035
rect -15085 21005 -635 21035
rect -605 21005 -600 21035
rect -15120 21000 -600 21005
rect -560 21000 -520 21040
rect -15520 20955 -520 20960
rect -15520 20925 -15515 20955
rect -15485 20925 -15355 20955
rect -15325 20925 -15195 20955
rect -15165 20925 -15035 20955
rect -15005 20925 -14955 20955
rect -14925 20925 -14875 20955
rect -14845 20925 -14795 20955
rect -14765 20925 -14715 20955
rect -14685 20925 -14635 20955
rect -14605 20925 -14555 20955
rect -14525 20925 -14475 20955
rect -14445 20925 -14395 20955
rect -14365 20925 -14315 20955
rect -14285 20925 -14235 20955
rect -14205 20925 -14155 20955
rect -14125 20925 -14075 20955
rect -14045 20925 -13995 20955
rect -13965 20925 -13915 20955
rect -13885 20925 -13835 20955
rect -13805 20925 -13755 20955
rect -13725 20925 -13675 20955
rect -13645 20925 -13595 20955
rect -13565 20925 -13515 20955
rect -13485 20925 -13435 20955
rect -13405 20925 -13355 20955
rect -13325 20925 -13275 20955
rect -13245 20925 -13195 20955
rect -13165 20925 -13115 20955
rect -13085 20925 -13035 20955
rect -13005 20925 -12955 20955
rect -12925 20925 -12875 20955
rect -12845 20925 -12795 20955
rect -12765 20925 -12715 20955
rect -12685 20925 -12635 20955
rect -12605 20925 -12555 20955
rect -12525 20925 -12475 20955
rect -12445 20925 -12395 20955
rect -12365 20925 -12315 20955
rect -12285 20925 -12235 20955
rect -12205 20925 -12155 20955
rect -12125 20925 -12075 20955
rect -12045 20925 -11995 20955
rect -11965 20925 -11915 20955
rect -11885 20925 -11835 20955
rect -11805 20925 -11755 20955
rect -11725 20925 -11675 20955
rect -11645 20925 -11595 20955
rect -11565 20925 -11515 20955
rect -11485 20925 -11435 20955
rect -11405 20925 -11355 20955
rect -11325 20925 -11275 20955
rect -11245 20925 -11195 20955
rect -11165 20925 -11115 20955
rect -11085 20925 -11035 20955
rect -11005 20925 -10955 20955
rect -10925 20925 -10875 20955
rect -10845 20925 -10795 20955
rect -10765 20925 -10715 20955
rect -10685 20925 -10635 20955
rect -10605 20925 -10555 20955
rect -10525 20925 -10475 20955
rect -10445 20925 -10395 20955
rect -10365 20925 -10315 20955
rect -10285 20925 -10235 20955
rect -10205 20925 -10155 20955
rect -10125 20925 -10075 20955
rect -10045 20925 -9995 20955
rect -9965 20925 -9915 20955
rect -9885 20925 -9835 20955
rect -9805 20925 -9755 20955
rect -9725 20925 -9675 20955
rect -9645 20925 -9595 20955
rect -9565 20925 -9515 20955
rect -9485 20925 -9435 20955
rect -9405 20925 -9355 20955
rect -9325 20925 -9275 20955
rect -9245 20925 -9195 20955
rect -9165 20925 -9115 20955
rect -9085 20925 -9035 20955
rect -9005 20925 -8955 20955
rect -8925 20925 -8875 20955
rect -8845 20925 -8795 20955
rect -8765 20925 -8715 20955
rect -8685 20925 -8635 20955
rect -8605 20925 -8555 20955
rect -8525 20925 -8475 20955
rect -8445 20925 -8395 20955
rect -8365 20925 -8315 20955
rect -8285 20925 -8235 20955
rect -8205 20925 -8155 20955
rect -8125 20925 -8075 20955
rect -8045 20925 -7995 20955
rect -7965 20925 -7915 20955
rect -7885 20925 -7835 20955
rect -7805 20925 -7755 20955
rect -7725 20925 -7675 20955
rect -7645 20925 -7595 20955
rect -7565 20925 -7515 20955
rect -7485 20925 -7435 20955
rect -7405 20925 -7355 20955
rect -7325 20925 -7275 20955
rect -7245 20925 -7195 20955
rect -7165 20925 -7115 20955
rect -7085 20925 -7035 20955
rect -7005 20925 -6955 20955
rect -6925 20925 -6875 20955
rect -6845 20925 -6795 20955
rect -6765 20925 -6715 20955
rect -6685 20925 -6635 20955
rect -6605 20925 -6555 20955
rect -6525 20925 -6475 20955
rect -6445 20925 -6395 20955
rect -6365 20925 -6315 20955
rect -6285 20925 -6235 20955
rect -6205 20925 -6155 20955
rect -6125 20925 -6075 20955
rect -6045 20925 -5915 20955
rect -5885 20925 -5755 20955
rect -5725 20925 -5675 20955
rect -5645 20925 -5595 20955
rect -5565 20925 -5515 20955
rect -5485 20925 -5435 20955
rect -5405 20925 -5355 20955
rect -5325 20925 -5275 20955
rect -5245 20925 -5195 20955
rect -5165 20925 -5115 20955
rect -5085 20925 -5035 20955
rect -5005 20925 -4955 20955
rect -4925 20925 -4875 20955
rect -4845 20925 -4795 20955
rect -4765 20925 -4715 20955
rect -4685 20925 -4635 20955
rect -4605 20925 -4555 20955
rect -4525 20925 -4475 20955
rect -4445 20925 -4395 20955
rect -4365 20925 -4315 20955
rect -4285 20925 -4235 20955
rect -4205 20925 -4155 20955
rect -4125 20925 -4075 20955
rect -4045 20925 -3995 20955
rect -3965 20925 -3915 20955
rect -3885 20925 -3835 20955
rect -3805 20925 -3755 20955
rect -3725 20925 -3675 20955
rect -3645 20925 -3595 20955
rect -3565 20925 -3515 20955
rect -3485 20925 -3435 20955
rect -3405 20925 -3355 20955
rect -3325 20925 -3275 20955
rect -3245 20925 -3195 20955
rect -3165 20925 -3115 20955
rect -3085 20925 -3035 20955
rect -3005 20925 -2955 20955
rect -2925 20925 -2875 20955
rect -2845 20925 -2795 20955
rect -2765 20925 -2715 20955
rect -2685 20925 -2635 20955
rect -2605 20925 -2555 20955
rect -2525 20925 -2475 20955
rect -2445 20925 -2395 20955
rect -2365 20925 -2315 20955
rect -2285 20925 -2235 20955
rect -2205 20925 -2155 20955
rect -2125 20925 -2075 20955
rect -2045 20925 -1995 20955
rect -1965 20925 -1835 20955
rect -1805 20925 -1755 20955
rect -1725 20925 -1675 20955
rect -1645 20925 -1515 20955
rect -1485 20925 -1355 20955
rect -1325 20925 -1275 20955
rect -1245 20925 -1195 20955
rect -1165 20925 -1115 20955
rect -1085 20925 -1035 20955
rect -1005 20925 -875 20955
rect -845 20925 -715 20955
rect -685 20925 -555 20955
rect -525 20925 -520 20955
rect -15520 20920 -520 20925
rect -15520 20875 -15000 20880
rect -15520 20845 -15515 20875
rect -15485 20845 -15355 20875
rect -15325 20845 -15195 20875
rect -15165 20845 -15035 20875
rect -15005 20845 -15000 20875
rect -15520 20840 -15000 20845
rect -6080 20875 -5720 20880
rect -6080 20845 -6075 20875
rect -6045 20845 -5915 20875
rect -5885 20845 -5755 20875
rect -5725 20845 -5720 20875
rect -6080 20840 -5720 20845
rect -1680 20875 -520 20880
rect -1680 20845 -1675 20875
rect -1645 20845 -1515 20875
rect -1485 20845 -1355 20875
rect -1325 20845 -1195 20875
rect -1165 20845 -1035 20875
rect -1005 20845 -875 20875
rect -845 20845 -715 20875
rect -685 20845 -555 20875
rect -525 20845 -520 20875
rect -1680 20840 -520 20845
rect -15520 20795 -15000 20800
rect -15520 20765 -15515 20795
rect -15485 20765 -15355 20795
rect -15325 20765 -15195 20795
rect -15165 20765 -15035 20795
rect -15005 20765 -15000 20795
rect -15520 20760 -15000 20765
rect -6080 20795 -5720 20800
rect -6080 20765 -6075 20795
rect -6045 20765 -5915 20795
rect -5885 20765 -5755 20795
rect -5725 20765 -5720 20795
rect -6080 20760 -5720 20765
rect -1680 20795 -520 20800
rect -1680 20765 -1675 20795
rect -1645 20765 -1515 20795
rect -1485 20765 -1355 20795
rect -1325 20765 -1195 20795
rect -1165 20765 -1035 20795
rect -1005 20765 -875 20795
rect -845 20765 -715 20795
rect -685 20765 -555 20795
rect -525 20765 -520 20795
rect -1680 20760 -520 20765
rect -16560 20675 -480 20680
rect -16560 20645 -16555 20675
rect -16525 20645 -16475 20675
rect -16445 20645 -16395 20675
rect -16365 20645 -16315 20675
rect -16285 20645 -16235 20675
rect -16205 20645 -16155 20675
rect -16125 20645 -16075 20675
rect -16045 20645 -15995 20675
rect -15965 20645 -15915 20675
rect -15885 20645 -15835 20675
rect -15805 20645 -15755 20675
rect -15725 20645 -15675 20675
rect -15645 20645 -15595 20675
rect -15565 20645 -14955 20675
rect -14925 20645 -14875 20675
rect -14845 20645 -14795 20675
rect -14765 20645 -14715 20675
rect -14685 20645 -14635 20675
rect -14605 20645 -14555 20675
rect -14525 20645 -14475 20675
rect -14445 20645 -14395 20675
rect -14365 20645 -14315 20675
rect -14285 20645 -14235 20675
rect -14205 20645 -14155 20675
rect -14125 20645 -14075 20675
rect -14045 20645 -13995 20675
rect -13965 20645 -13915 20675
rect -13885 20645 -13835 20675
rect -13805 20645 -13755 20675
rect -13725 20645 -13675 20675
rect -13645 20645 -13595 20675
rect -13565 20645 -13515 20675
rect -13485 20645 -13435 20675
rect -13405 20645 -13355 20675
rect -13325 20645 -13275 20675
rect -13245 20645 -13195 20675
rect -13165 20645 -13115 20675
rect -13085 20645 -13035 20675
rect -13005 20645 -12955 20675
rect -12925 20645 -12875 20675
rect -12845 20645 -12795 20675
rect -12765 20645 -12715 20675
rect -12685 20645 -12635 20675
rect -12605 20645 -12555 20675
rect -12525 20645 -12475 20675
rect -12445 20645 -12395 20675
rect -12365 20645 -12315 20675
rect -12285 20645 -12235 20675
rect -12205 20645 -12155 20675
rect -12125 20645 -12075 20675
rect -12045 20645 -11995 20675
rect -11965 20645 -11915 20675
rect -11885 20645 -11835 20675
rect -11805 20645 -11755 20675
rect -11725 20645 -11675 20675
rect -11645 20645 -11595 20675
rect -11565 20645 -11515 20675
rect -11485 20645 -11435 20675
rect -11405 20645 -11355 20675
rect -11325 20645 -11275 20675
rect -11245 20645 -11195 20675
rect -11165 20645 -11115 20675
rect -11085 20645 -11035 20675
rect -11005 20645 -10955 20675
rect -10925 20645 -10875 20675
rect -10845 20645 -10795 20675
rect -10765 20645 -10715 20675
rect -10685 20645 -10635 20675
rect -10605 20645 -10555 20675
rect -10525 20645 -10475 20675
rect -10445 20645 -10395 20675
rect -10365 20645 -10315 20675
rect -10285 20645 -10235 20675
rect -10205 20645 -10155 20675
rect -10125 20645 -10075 20675
rect -10045 20645 -9995 20675
rect -9965 20645 -9915 20675
rect -9885 20645 -9835 20675
rect -9805 20645 -9755 20675
rect -9725 20645 -9675 20675
rect -9645 20645 -9595 20675
rect -9565 20645 -9515 20675
rect -9485 20645 -9435 20675
rect -9405 20645 -9355 20675
rect -9325 20645 -9275 20675
rect -9245 20645 -9195 20675
rect -9165 20645 -9115 20675
rect -9085 20645 -9035 20675
rect -9005 20645 -8955 20675
rect -8925 20645 -8875 20675
rect -8845 20645 -8795 20675
rect -8765 20645 -8715 20675
rect -8685 20645 -8635 20675
rect -8605 20645 -8555 20675
rect -8525 20645 -8475 20675
rect -8445 20645 -8395 20675
rect -8365 20645 -8315 20675
rect -8285 20645 -8235 20675
rect -8205 20645 -8155 20675
rect -8125 20645 -8075 20675
rect -8045 20645 -7995 20675
rect -7965 20645 -7915 20675
rect -7885 20645 -7835 20675
rect -7805 20645 -7755 20675
rect -7725 20645 -7675 20675
rect -7645 20645 -7595 20675
rect -7565 20645 -7515 20675
rect -7485 20645 -7435 20675
rect -7405 20645 -7355 20675
rect -7325 20645 -7275 20675
rect -7245 20645 -7195 20675
rect -7165 20645 -7115 20675
rect -7085 20645 -7035 20675
rect -7005 20645 -6955 20675
rect -6925 20645 -6875 20675
rect -6845 20645 -6795 20675
rect -6765 20645 -6715 20675
rect -6685 20645 -6635 20675
rect -6605 20645 -6555 20675
rect -6525 20645 -6475 20675
rect -6445 20645 -6395 20675
rect -6365 20645 -6315 20675
rect -6285 20645 -6235 20675
rect -6205 20645 -6155 20675
rect -6125 20645 -5675 20675
rect -5645 20645 -5595 20675
rect -5565 20645 -5515 20675
rect -5485 20645 -5435 20675
rect -5405 20645 -5355 20675
rect -5325 20645 -5275 20675
rect -5245 20645 -5195 20675
rect -5165 20645 -5115 20675
rect -5085 20645 -5035 20675
rect -5005 20645 -4955 20675
rect -4925 20645 -4875 20675
rect -4845 20645 -4795 20675
rect -4765 20645 -4715 20675
rect -4685 20645 -4635 20675
rect -4605 20645 -4555 20675
rect -4525 20645 -4475 20675
rect -4445 20645 -4395 20675
rect -4365 20645 -4315 20675
rect -4285 20645 -4235 20675
rect -4205 20645 -4155 20675
rect -4125 20645 -4075 20675
rect -4045 20645 -3995 20675
rect -3965 20645 -3915 20675
rect -3885 20645 -3835 20675
rect -3805 20645 -3755 20675
rect -3725 20645 -3675 20675
rect -3645 20645 -3595 20675
rect -3565 20645 -3515 20675
rect -3485 20645 -3435 20675
rect -3405 20645 -3355 20675
rect -3325 20645 -3275 20675
rect -3245 20645 -3195 20675
rect -3165 20645 -3115 20675
rect -3085 20645 -3035 20675
rect -3005 20645 -2955 20675
rect -2925 20645 -2875 20675
rect -2845 20645 -2795 20675
rect -2765 20645 -2715 20675
rect -2685 20645 -2635 20675
rect -2605 20645 -2555 20675
rect -2525 20645 -2475 20675
rect -2445 20645 -2395 20675
rect -2365 20645 -2315 20675
rect -2285 20645 -2235 20675
rect -2205 20645 -2155 20675
rect -2125 20645 -2075 20675
rect -2045 20645 -1995 20675
rect -1965 20645 -1915 20675
rect -1885 20645 -1835 20675
rect -1805 20645 -1755 20675
rect -1725 20645 -480 20675
rect -16560 20640 -480 20645
rect 20480 20675 21600 20680
rect 20480 20645 20525 20675
rect 20555 20645 20605 20675
rect 20635 20645 20685 20675
rect 20715 20645 20765 20675
rect 20795 20645 20845 20675
rect 20875 20645 20925 20675
rect 20955 20645 21005 20675
rect 21035 20645 21085 20675
rect 21115 20645 21165 20675
rect 21195 20645 21245 20675
rect 21275 20645 21325 20675
rect 21355 20645 21405 20675
rect 21435 20645 21485 20675
rect 21515 20645 21565 20675
rect 21595 20645 21600 20675
rect 20480 20640 21600 20645
rect -16640 20560 21680 20600
rect -16560 20515 -480 20520
rect -16560 20485 -16555 20515
rect -16525 20485 -16475 20515
rect -16445 20485 -16395 20515
rect -16365 20485 -16315 20515
rect -16285 20485 -16235 20515
rect -16205 20485 -16155 20515
rect -16125 20485 -16075 20515
rect -16045 20485 -15995 20515
rect -15965 20485 -15915 20515
rect -15885 20485 -15835 20515
rect -15805 20485 -15755 20515
rect -15725 20485 -15675 20515
rect -15645 20485 -15595 20515
rect -15565 20485 -14955 20515
rect -14925 20485 -14875 20515
rect -14845 20485 -14795 20515
rect -14765 20485 -14715 20515
rect -14685 20485 -14635 20515
rect -14605 20485 -14555 20515
rect -14525 20485 -14475 20515
rect -14445 20485 -14395 20515
rect -14365 20485 -14315 20515
rect -14285 20485 -14235 20515
rect -14205 20485 -14155 20515
rect -14125 20485 -14075 20515
rect -14045 20485 -13995 20515
rect -13965 20485 -13915 20515
rect -13885 20485 -13835 20515
rect -13805 20485 -13755 20515
rect -13725 20485 -13675 20515
rect -13645 20485 -13595 20515
rect -13565 20485 -13515 20515
rect -13485 20485 -13435 20515
rect -13405 20485 -13355 20515
rect -13325 20485 -13275 20515
rect -13245 20485 -13195 20515
rect -13165 20485 -13115 20515
rect -13085 20485 -13035 20515
rect -13005 20485 -12955 20515
rect -12925 20485 -12875 20515
rect -12845 20485 -12795 20515
rect -12765 20485 -12715 20515
rect -12685 20485 -12635 20515
rect -12605 20485 -12555 20515
rect -12525 20485 -12475 20515
rect -12445 20485 -12395 20515
rect -12365 20485 -12315 20515
rect -12285 20485 -12235 20515
rect -12205 20485 -12155 20515
rect -12125 20485 -12075 20515
rect -12045 20485 -11995 20515
rect -11965 20485 -11915 20515
rect -11885 20485 -11835 20515
rect -11805 20485 -11755 20515
rect -11725 20485 -11675 20515
rect -11645 20485 -11595 20515
rect -11565 20485 -11515 20515
rect -11485 20485 -11435 20515
rect -11405 20485 -11355 20515
rect -11325 20485 -11275 20515
rect -11245 20485 -11195 20515
rect -11165 20485 -11115 20515
rect -11085 20485 -11035 20515
rect -11005 20485 -10955 20515
rect -10925 20485 -10875 20515
rect -10845 20485 -10795 20515
rect -10765 20485 -10715 20515
rect -10685 20485 -10635 20515
rect -10605 20485 -10555 20515
rect -10525 20485 -10475 20515
rect -10445 20485 -10395 20515
rect -10365 20485 -10315 20515
rect -10285 20485 -10235 20515
rect -10205 20485 -10155 20515
rect -10125 20485 -10075 20515
rect -10045 20485 -9995 20515
rect -9965 20485 -9915 20515
rect -9885 20485 -9835 20515
rect -9805 20485 -9755 20515
rect -9725 20485 -9675 20515
rect -9645 20485 -9595 20515
rect -9565 20485 -9515 20515
rect -9485 20485 -9435 20515
rect -9405 20485 -9355 20515
rect -9325 20485 -9275 20515
rect -9245 20485 -9195 20515
rect -9165 20485 -9115 20515
rect -9085 20485 -9035 20515
rect -9005 20485 -8955 20515
rect -8925 20485 -8875 20515
rect -8845 20485 -8795 20515
rect -8765 20485 -8715 20515
rect -8685 20485 -8635 20515
rect -8605 20485 -8555 20515
rect -8525 20485 -8475 20515
rect -8445 20485 -8395 20515
rect -8365 20485 -8315 20515
rect -8285 20485 -8235 20515
rect -8205 20485 -8155 20515
rect -8125 20485 -8075 20515
rect -8045 20485 -7995 20515
rect -7965 20485 -7915 20515
rect -7885 20485 -7835 20515
rect -7805 20485 -7755 20515
rect -7725 20485 -7675 20515
rect -7645 20485 -7595 20515
rect -7565 20485 -7515 20515
rect -7485 20485 -7435 20515
rect -7405 20485 -7355 20515
rect -7325 20485 -7275 20515
rect -7245 20485 -7195 20515
rect -7165 20485 -7115 20515
rect -7085 20485 -7035 20515
rect -7005 20485 -6955 20515
rect -6925 20485 -6875 20515
rect -6845 20485 -6795 20515
rect -6765 20485 -6715 20515
rect -6685 20485 -6635 20515
rect -6605 20485 -6555 20515
rect -6525 20485 -6475 20515
rect -6445 20485 -6395 20515
rect -6365 20485 -6315 20515
rect -6285 20485 -6235 20515
rect -6205 20485 -6155 20515
rect -6125 20485 -5675 20515
rect -5645 20485 -5595 20515
rect -5565 20485 -5515 20515
rect -5485 20485 -5435 20515
rect -5405 20485 -5355 20515
rect -5325 20485 -5275 20515
rect -5245 20485 -5195 20515
rect -5165 20485 -5115 20515
rect -5085 20485 -5035 20515
rect -5005 20485 -4955 20515
rect -4925 20485 -4875 20515
rect -4845 20485 -4795 20515
rect -4765 20485 -4715 20515
rect -4685 20485 -4635 20515
rect -4605 20485 -4555 20515
rect -4525 20485 -4475 20515
rect -4445 20485 -4395 20515
rect -4365 20485 -4315 20515
rect -4285 20485 -4235 20515
rect -4205 20485 -4155 20515
rect -4125 20485 -4075 20515
rect -4045 20485 -3995 20515
rect -3965 20485 -3915 20515
rect -3885 20485 -3835 20515
rect -3805 20485 -3755 20515
rect -3725 20485 -3675 20515
rect -3645 20485 -3595 20515
rect -3565 20485 -3515 20515
rect -3485 20485 -3435 20515
rect -3405 20485 -3355 20515
rect -3325 20485 -3275 20515
rect -3245 20485 -3195 20515
rect -3165 20485 -3115 20515
rect -3085 20485 -3035 20515
rect -3005 20485 -2955 20515
rect -2925 20485 -2875 20515
rect -2845 20485 -2795 20515
rect -2765 20485 -2715 20515
rect -2685 20485 -2635 20515
rect -2605 20485 -2555 20515
rect -2525 20485 -2475 20515
rect -2445 20485 -2395 20515
rect -2365 20485 -2315 20515
rect -2285 20485 -2235 20515
rect -2205 20485 -2155 20515
rect -2125 20485 -2075 20515
rect -2045 20485 -1995 20515
rect -1965 20485 -1915 20515
rect -1885 20485 -1835 20515
rect -1805 20485 -1755 20515
rect -1725 20485 -480 20515
rect -16560 20480 -480 20485
rect 20480 20515 21600 20520
rect 20480 20485 20525 20515
rect 20555 20485 20605 20515
rect 20635 20485 20685 20515
rect 20715 20485 20765 20515
rect 20795 20485 20845 20515
rect 20875 20485 20925 20515
rect 20955 20485 21005 20515
rect 21035 20485 21085 20515
rect 21115 20485 21165 20515
rect 21195 20485 21245 20515
rect 21275 20485 21325 20515
rect 21355 20485 21405 20515
rect 21435 20485 21485 20515
rect 21515 20485 21565 20515
rect 21595 20485 21600 20515
rect 20480 20480 21600 20485
rect -6080 20435 -5720 20440
rect -6080 20405 -6075 20435
rect -6045 20405 -5915 20435
rect -5885 20405 -5755 20435
rect -5725 20405 -5720 20435
rect -6080 20400 -5720 20405
rect -1680 20435 -520 20440
rect -1680 20405 -1675 20435
rect -1645 20405 -1515 20435
rect -1485 20405 -1355 20435
rect -1325 20405 -1195 20435
rect -1165 20405 -1035 20435
rect -1005 20405 -875 20435
rect -845 20405 -715 20435
rect -685 20405 -555 20435
rect -525 20405 -520 20435
rect -1680 20400 -520 20405
rect -15520 20395 -15000 20400
rect -15520 20365 -15515 20395
rect -15485 20365 -15355 20395
rect -15325 20365 -15195 20395
rect -15165 20365 -15035 20395
rect -15005 20365 -15000 20395
rect -15520 20360 -15000 20365
rect -6080 20355 -5720 20360
rect -6080 20325 -6075 20355
rect -6045 20325 -5915 20355
rect -5885 20325 -5755 20355
rect -5725 20325 -5720 20355
rect -6080 20320 -5720 20325
rect -5280 20355 -520 20360
rect -5280 20325 -5275 20355
rect -5245 20325 -5115 20355
rect -5085 20325 -5035 20355
rect -5005 20325 -4955 20355
rect -4925 20325 -4875 20355
rect -4845 20325 -4795 20355
rect -4765 20325 -4715 20355
rect -4685 20325 -4635 20355
rect -4605 20325 -4555 20355
rect -4525 20325 -4475 20355
rect -4445 20325 -4395 20355
rect -4365 20325 -4315 20355
rect -4285 20325 -4235 20355
rect -4205 20325 -4155 20355
rect -4125 20325 -4075 20355
rect -4045 20325 -3995 20355
rect -3965 20325 -3915 20355
rect -3885 20325 -3835 20355
rect -3805 20325 -3755 20355
rect -3725 20325 -3675 20355
rect -3645 20325 -3595 20355
rect -3565 20325 -3515 20355
rect -3485 20325 -3435 20355
rect -3405 20325 -3355 20355
rect -3325 20325 -3275 20355
rect -3245 20325 -3195 20355
rect -3165 20325 -3115 20355
rect -3085 20325 -3035 20355
rect -3005 20325 -2955 20355
rect -2925 20325 -2875 20355
rect -2845 20325 -2795 20355
rect -2765 20325 -2715 20355
rect -2685 20325 -2635 20355
rect -2605 20325 -2555 20355
rect -2525 20325 -2475 20355
rect -2445 20325 -2395 20355
rect -2365 20325 -2315 20355
rect -2285 20325 -2235 20355
rect -2205 20325 -2155 20355
rect -2125 20325 -2075 20355
rect -2045 20325 -1995 20355
rect -1965 20325 -1835 20355
rect -1805 20325 -1755 20355
rect -1725 20325 -1675 20355
rect -1645 20325 -1515 20355
rect -1485 20325 -1355 20355
rect -1325 20325 -1195 20355
rect -1165 20325 -1035 20355
rect -1005 20325 -875 20355
rect -845 20325 -715 20355
rect -685 20325 -555 20355
rect -525 20325 -520 20355
rect -5280 20320 -520 20325
rect -15520 20315 -15000 20320
rect -15520 20285 -15515 20315
rect -15485 20285 -15355 20315
rect -15325 20285 -15195 20315
rect -15165 20285 -15035 20315
rect -15005 20285 -15000 20315
rect -15520 20280 -15000 20285
rect -5200 20275 -600 20280
rect -5200 20245 -5195 20275
rect -5165 20245 -635 20275
rect -605 20245 -600 20275
rect -5200 20240 -600 20245
rect -15520 20235 -15000 20240
rect -15520 20205 -15515 20235
rect -15485 20205 -15355 20235
rect -15325 20205 -15195 20235
rect -15165 20205 -15035 20235
rect -15005 20205 -15000 20235
rect -15520 20200 -15000 20205
rect -6080 20195 -5720 20200
rect -6080 20165 -6075 20195
rect -6045 20165 -5915 20195
rect -5885 20165 -5755 20195
rect -5725 20165 -5720 20195
rect -6080 20160 -5720 20165
rect -5280 20195 -520 20200
rect -5280 20165 -5275 20195
rect -5245 20165 -5115 20195
rect -5085 20165 -5035 20195
rect -5005 20165 -4955 20195
rect -4925 20165 -4875 20195
rect -4845 20165 -4795 20195
rect -4765 20165 -4715 20195
rect -4685 20165 -4635 20195
rect -4605 20165 -4555 20195
rect -4525 20165 -4475 20195
rect -4445 20165 -4395 20195
rect -4365 20165 -4315 20195
rect -4285 20165 -4235 20195
rect -4205 20165 -4155 20195
rect -4125 20165 -4075 20195
rect -4045 20165 -3995 20195
rect -3965 20165 -3915 20195
rect -3885 20165 -3835 20195
rect -3805 20165 -3755 20195
rect -3725 20165 -3675 20195
rect -3645 20165 -3595 20195
rect -3565 20165 -3515 20195
rect -3485 20165 -3435 20195
rect -3405 20165 -3355 20195
rect -3325 20165 -3275 20195
rect -3245 20165 -3195 20195
rect -3165 20165 -3115 20195
rect -3085 20165 -3035 20195
rect -3005 20165 -2955 20195
rect -2925 20165 -2875 20195
rect -2845 20165 -2795 20195
rect -2765 20165 -2715 20195
rect -2685 20165 -2635 20195
rect -2605 20165 -2555 20195
rect -2525 20165 -2475 20195
rect -2445 20165 -2395 20195
rect -2365 20165 -2315 20195
rect -2285 20165 -2235 20195
rect -2205 20165 -2155 20195
rect -2125 20165 -2075 20195
rect -2045 20165 -1995 20195
rect -1965 20165 -1835 20195
rect -1805 20165 -1755 20195
rect -1725 20165 -1675 20195
rect -1645 20165 -1515 20195
rect -1485 20165 -1355 20195
rect -1325 20165 -1195 20195
rect -1165 20165 -1035 20195
rect -1005 20165 -875 20195
rect -845 20165 -715 20195
rect -685 20165 -555 20195
rect -525 20165 -520 20195
rect -5280 20160 -520 20165
rect -15520 20155 -15000 20160
rect -15520 20125 -15515 20155
rect -15485 20125 -15355 20155
rect -15325 20125 -15195 20155
rect -15165 20125 -15035 20155
rect -15005 20125 -15000 20155
rect -15520 20120 -15000 20125
rect -1680 20115 -1320 20120
rect -1680 20085 -1675 20115
rect -1645 20085 -1515 20115
rect -1485 20085 -1355 20115
rect -1325 20085 -1320 20115
rect -1680 20080 -1320 20085
rect -1280 20115 -480 20120
rect -1280 20085 -1275 20115
rect -1245 20085 -955 20115
rect -925 20085 -480 20115
rect -1280 20080 -480 20085
rect -15520 20075 -15000 20080
rect -15520 20045 -15515 20075
rect -15485 20045 -15355 20075
rect -15325 20045 -15195 20075
rect -15165 20045 -15035 20075
rect -15005 20045 -15000 20075
rect -15520 20040 -15000 20045
rect -1680 20035 -520 20040
rect -1680 20005 -1675 20035
rect -1645 20005 -1515 20035
rect -1485 20005 -1355 20035
rect -1325 20005 -1195 20035
rect -1165 20005 -1035 20035
rect -1005 20005 -875 20035
rect -845 20005 -715 20035
rect -685 20005 -555 20035
rect -525 20005 -520 20035
rect -1680 20000 -520 20005
rect 20480 20035 21600 20040
rect 20480 20005 20525 20035
rect 20555 20005 20605 20035
rect 20635 20005 20685 20035
rect 20715 20005 20765 20035
rect 20795 20005 20845 20035
rect 20875 20005 20925 20035
rect 20955 20005 21005 20035
rect 21035 20005 21085 20035
rect 21115 20005 21165 20035
rect 21195 20005 21245 20035
rect 21275 20005 21325 20035
rect 21355 20005 21405 20035
rect 21435 20005 21485 20035
rect 21515 20005 21565 20035
rect 21595 20005 21600 20035
rect 20480 20000 21600 20005
rect -15520 19995 -15000 20000
rect -15520 19965 -15515 19995
rect -15485 19965 -15355 19995
rect -15325 19965 -15195 19995
rect -15165 19965 -15035 19995
rect -15005 19965 -15000 19995
rect -15520 19960 -15000 19965
rect -1680 19955 -1160 19960
rect -1680 19925 -1675 19955
rect -1645 19925 -1515 19955
rect -1485 19925 -1355 19955
rect -1325 19925 -1195 19955
rect -1165 19925 -1160 19955
rect -1680 19920 -1160 19925
rect -1120 19955 21680 19960
rect -1120 19925 -1115 19955
rect -1085 19925 -795 19955
rect -765 19925 21680 19955
rect -1120 19920 21680 19925
rect -15520 19915 -15000 19920
rect -15520 19885 -15515 19915
rect -15485 19885 -15355 19915
rect -15325 19885 -15195 19915
rect -15165 19885 -15035 19915
rect -15005 19885 -15000 19915
rect -15520 19880 -15000 19885
rect -1680 19875 -520 19880
rect -1680 19845 -1675 19875
rect -1645 19845 -1515 19875
rect -1485 19845 -1355 19875
rect -1325 19845 -1195 19875
rect -1165 19845 -1035 19875
rect -1005 19845 -875 19875
rect -845 19845 -715 19875
rect -685 19845 -555 19875
rect -525 19845 -520 19875
rect -1680 19840 -520 19845
rect 20480 19875 21600 19880
rect 20480 19845 20525 19875
rect 20555 19845 20605 19875
rect 20635 19845 20685 19875
rect 20715 19845 20765 19875
rect 20795 19845 20845 19875
rect 20875 19845 20925 19875
rect 20955 19845 21005 19875
rect 21035 19845 21085 19875
rect 21115 19845 21165 19875
rect 21195 19845 21245 19875
rect 21275 19845 21325 19875
rect 21355 19845 21405 19875
rect 21435 19845 21485 19875
rect 21515 19845 21565 19875
rect 21595 19845 21600 19875
rect 20480 19840 21600 19845
rect -15520 19835 -15000 19840
rect -15520 19805 -15515 19835
rect -15485 19805 -15355 19835
rect -15325 19805 -15195 19835
rect -15165 19805 -15035 19835
rect -15005 19805 -15000 19835
rect -15520 19800 -15000 19805
rect -1680 19795 -520 19800
rect -1680 19765 -1675 19795
rect -1645 19765 -1515 19795
rect -1485 19765 -1355 19795
rect -1325 19765 -1195 19795
rect -1165 19765 -1035 19795
rect -1005 19765 -875 19795
rect -845 19765 -715 19795
rect -685 19765 -555 19795
rect -525 19765 -520 19795
rect -1680 19760 -520 19765
rect -15520 19755 -15000 19760
rect -15520 19725 -15515 19755
rect -15485 19725 -15355 19755
rect -15325 19725 -15195 19755
rect -15165 19725 -15035 19755
rect -15005 19725 -15000 19755
rect -15520 19720 -15000 19725
rect -1680 19715 -520 19720
rect -1680 19685 -1675 19715
rect -1645 19685 -1515 19715
rect -1485 19685 -1355 19715
rect -1325 19685 -1195 19715
rect -1165 19685 -1035 19715
rect -1005 19685 -875 19715
rect -845 19685 -715 19715
rect -685 19685 -555 19715
rect -525 19685 -520 19715
rect -1680 19680 -520 19685
rect -15520 19675 -15000 19680
rect -15520 19645 -15515 19675
rect -15485 19645 -15355 19675
rect -15325 19645 -15195 19675
rect -15165 19645 -15035 19675
rect -15005 19645 -15000 19675
rect -15520 19640 -15000 19645
rect -1680 19635 -520 19640
rect -1680 19605 -1675 19635
rect -1645 19605 -1515 19635
rect -1485 19605 -1355 19635
rect -1325 19605 -1195 19635
rect -1165 19605 -1035 19635
rect -1005 19605 -875 19635
rect -845 19605 -715 19635
rect -685 19605 -555 19635
rect -525 19605 -520 19635
rect -1680 19600 -520 19605
rect -15520 19595 -15000 19600
rect -15520 19565 -15515 19595
rect -15485 19565 -15355 19595
rect -15325 19565 -15195 19595
rect -15165 19565 -15035 19595
rect -15005 19565 -15000 19595
rect -15520 19560 -15000 19565
rect -1680 19555 -520 19560
rect -1680 19525 -1675 19555
rect -1645 19525 -1515 19555
rect -1485 19525 -1355 19555
rect -1325 19525 -1195 19555
rect -1165 19525 -1035 19555
rect -1005 19525 -875 19555
rect -845 19525 -715 19555
rect -685 19525 -555 19555
rect -525 19525 -520 19555
rect -1680 19520 -520 19525
rect -15520 19515 -15000 19520
rect -15520 19485 -15515 19515
rect -15485 19485 -15355 19515
rect -15325 19485 -15195 19515
rect -15165 19485 -15035 19515
rect -15005 19485 -15000 19515
rect -15520 19480 -15000 19485
rect -1680 19475 -520 19480
rect -1680 19445 -1675 19475
rect -1645 19445 -1515 19475
rect -1485 19445 -1355 19475
rect -1325 19445 -1195 19475
rect -1165 19445 -1035 19475
rect -1005 19445 -875 19475
rect -845 19445 -715 19475
rect -685 19445 -555 19475
rect -525 19445 -520 19475
rect -1680 19440 -520 19445
rect -15520 19435 -15000 19440
rect -15520 19405 -15515 19435
rect -15485 19405 -15355 19435
rect -15325 19405 -15195 19435
rect -15165 19405 -15035 19435
rect -15005 19405 -15000 19435
rect -15520 19400 -15000 19405
rect -1680 19395 -520 19400
rect -1680 19365 -1675 19395
rect -1645 19365 -1515 19395
rect -1485 19365 -1355 19395
rect -1325 19365 -1195 19395
rect -1165 19365 -1035 19395
rect -1005 19365 -875 19395
rect -845 19365 -715 19395
rect -685 19365 -555 19395
rect -525 19365 -520 19395
rect -1680 19360 -520 19365
rect -15520 19355 -15000 19360
rect -15520 19325 -15515 19355
rect -15485 19325 -15355 19355
rect -15325 19325 -15195 19355
rect -15165 19325 -15035 19355
rect -15005 19325 -15000 19355
rect -15520 19320 -15000 19325
rect -1680 19315 -520 19320
rect -1680 19285 -1675 19315
rect -1645 19285 -1515 19315
rect -1485 19285 -1355 19315
rect -1325 19285 -1195 19315
rect -1165 19285 -1035 19315
rect -1005 19285 -875 19315
rect -845 19285 -715 19315
rect -685 19285 -555 19315
rect -525 19285 -520 19315
rect -1680 19280 -520 19285
rect -15520 19275 -15000 19280
rect -15520 19245 -15515 19275
rect -15485 19245 -15355 19275
rect -15325 19245 -15195 19275
rect -15165 19245 -15035 19275
rect -15005 19245 -15000 19275
rect -15520 19240 -15000 19245
rect -1680 19235 -520 19240
rect -1680 19205 -1675 19235
rect -1645 19205 -1515 19235
rect -1485 19205 -1355 19235
rect -1325 19205 -1195 19235
rect -1165 19205 -1035 19235
rect -1005 19205 -875 19235
rect -845 19205 -715 19235
rect -685 19205 -555 19235
rect -525 19205 -520 19235
rect -1680 19200 -520 19205
rect -15520 19195 -15000 19200
rect -15520 19165 -15515 19195
rect -15485 19165 -15355 19195
rect -15325 19165 -15195 19195
rect -15165 19165 -15035 19195
rect -15005 19165 -15000 19195
rect -15520 19160 -15000 19165
rect -1680 19155 -520 19160
rect -1680 19125 -1675 19155
rect -1645 19125 -1515 19155
rect -1485 19125 -1355 19155
rect -1325 19125 -1195 19155
rect -1165 19125 -1035 19155
rect -1005 19125 -875 19155
rect -845 19125 -715 19155
rect -685 19125 -555 19155
rect -525 19125 -520 19155
rect -1680 19120 -520 19125
rect -15520 19115 -15000 19120
rect -15520 19085 -15515 19115
rect -15485 19085 -15355 19115
rect -15325 19085 -15195 19115
rect -15165 19085 -15035 19115
rect -15005 19085 -15000 19115
rect -15520 19080 -15000 19085
rect -1680 19075 -520 19080
rect -1680 19045 -1675 19075
rect -1645 19045 -1515 19075
rect -1485 19045 -1355 19075
rect -1325 19045 -1195 19075
rect -1165 19045 -1035 19075
rect -1005 19045 -875 19075
rect -845 19045 -715 19075
rect -685 19045 -555 19075
rect -525 19045 -520 19075
rect -1680 19040 -520 19045
rect -15520 19035 -15000 19040
rect -15520 19005 -15515 19035
rect -15485 19005 -15355 19035
rect -15325 19005 -15195 19035
rect -15165 19005 -15035 19035
rect -15005 19005 -15000 19035
rect -15520 19000 -15000 19005
rect -1680 18995 -520 19000
rect -1680 18965 -1675 18995
rect -1645 18965 -1515 18995
rect -1485 18965 -1355 18995
rect -1325 18965 -1195 18995
rect -1165 18965 -1035 18995
rect -1005 18965 -875 18995
rect -845 18965 -715 18995
rect -685 18965 -555 18995
rect -525 18965 -520 18995
rect -1680 18960 -520 18965
rect -15520 18955 -15000 18960
rect -15520 18925 -15515 18955
rect -15485 18925 -15355 18955
rect -15325 18925 -15195 18955
rect -15165 18925 -15035 18955
rect -15005 18925 -15000 18955
rect -15520 18920 -15000 18925
rect -1680 18915 -520 18920
rect -1680 18885 -1675 18915
rect -1645 18885 -1515 18915
rect -1485 18885 -1355 18915
rect -1325 18885 -1195 18915
rect -1165 18885 -1035 18915
rect -1005 18885 -875 18915
rect -845 18885 -715 18915
rect -685 18885 -555 18915
rect -525 18885 -520 18915
rect -1680 18880 -520 18885
rect -16560 18875 -15000 18880
rect -16560 18845 -16555 18875
rect -16525 18845 -16475 18875
rect -16445 18845 -16395 18875
rect -16365 18845 -16315 18875
rect -16285 18845 -16235 18875
rect -16205 18845 -16155 18875
rect -16125 18845 -16075 18875
rect -16045 18845 -15995 18875
rect -15965 18845 -15915 18875
rect -15885 18845 -15835 18875
rect -15805 18845 -15755 18875
rect -15725 18845 -15675 18875
rect -15645 18845 -15595 18875
rect -15565 18845 -15515 18875
rect -15485 18845 -15355 18875
rect -15325 18845 -15195 18875
rect -15165 18845 -15035 18875
rect -15005 18845 -15000 18875
rect -16560 18840 -15000 18845
rect -1680 18835 -680 18840
rect -1680 18805 -1675 18835
rect -1645 18805 -1515 18835
rect -1485 18805 -1355 18835
rect -1325 18805 -1195 18835
rect -1165 18805 -1035 18835
rect -1005 18805 -875 18835
rect -845 18805 -715 18835
rect -685 18805 -680 18835
rect -1680 18800 -680 18805
rect -640 18835 20480 18840
rect -640 18805 -635 18835
rect -605 18805 20480 18835
rect -640 18800 20480 18805
rect -16640 18795 -15240 18800
rect -16640 18765 -15435 18795
rect -15405 18765 -15275 18795
rect -15245 18765 -15240 18795
rect -16640 18760 -15240 18765
rect -1680 18755 -520 18760
rect -1680 18725 -1675 18755
rect -1645 18725 -1515 18755
rect -1485 18725 -1355 18755
rect -1325 18725 -1195 18755
rect -1165 18725 -1035 18755
rect -1005 18725 -875 18755
rect -845 18725 -715 18755
rect -685 18725 -555 18755
rect -525 18725 -520 18755
rect -1680 18720 -520 18725
rect -16560 18715 -15000 18720
rect -16560 18685 -16555 18715
rect -16525 18685 -16475 18715
rect -16445 18685 -16395 18715
rect -16365 18685 -16315 18715
rect -16285 18685 -16235 18715
rect -16205 18685 -16155 18715
rect -16125 18685 -16075 18715
rect -16045 18685 -15995 18715
rect -15965 18685 -15915 18715
rect -15885 18685 -15835 18715
rect -15805 18685 -15755 18715
rect -15725 18685 -15675 18715
rect -15645 18685 -15595 18715
rect -15565 18685 -15515 18715
rect -15485 18685 -15355 18715
rect -15325 18685 -15195 18715
rect -15165 18685 -15035 18715
rect -15005 18685 -15000 18715
rect -16560 18680 -15000 18685
rect -1680 18675 -520 18680
rect -1680 18645 -1675 18675
rect -1645 18645 -1515 18675
rect -1485 18645 -1355 18675
rect -1325 18645 -1195 18675
rect -1165 18645 -1035 18675
rect -1005 18645 -875 18675
rect -845 18645 -715 18675
rect -685 18645 -555 18675
rect -525 18645 -520 18675
rect -1680 18640 -520 18645
rect -16640 18635 -15080 18640
rect -16640 18605 -15435 18635
rect -15405 18605 -15115 18635
rect -15085 18605 -15080 18635
rect -16640 18600 -15080 18605
rect -1680 18595 -520 18600
rect -1680 18565 -1675 18595
rect -1645 18565 -1515 18595
rect -1485 18565 -1355 18595
rect -1325 18565 -1195 18595
rect -1165 18565 -1035 18595
rect -1005 18565 -875 18595
rect -845 18565 -715 18595
rect -685 18565 -555 18595
rect -525 18565 -520 18595
rect -1680 18560 -520 18565
rect -16560 18555 -15000 18560
rect -16560 18525 -16555 18555
rect -16525 18525 -16475 18555
rect -16445 18525 -16395 18555
rect -16365 18525 -16315 18555
rect -16285 18525 -16235 18555
rect -16205 18525 -16155 18555
rect -16125 18525 -16075 18555
rect -16045 18525 -15995 18555
rect -15965 18525 -15915 18555
rect -15885 18525 -15835 18555
rect -15805 18525 -15755 18555
rect -15725 18525 -15675 18555
rect -15645 18525 -15595 18555
rect -15565 18525 -15515 18555
rect -15485 18525 -15355 18555
rect -15325 18525 -15195 18555
rect -15165 18525 -15035 18555
rect -15005 18525 -15000 18555
rect -16560 18520 -15000 18525
rect -1680 18515 -520 18520
rect -1680 18485 -1675 18515
rect -1645 18485 -1515 18515
rect -1485 18485 -1355 18515
rect -1325 18485 -1195 18515
rect -1165 18485 -1035 18515
rect -1005 18485 -875 18515
rect -845 18485 -715 18515
rect -685 18485 -555 18515
rect -525 18485 -520 18515
rect -1680 18480 -520 18485
rect -15520 18475 -15000 18480
rect -15520 18445 -15515 18475
rect -15485 18445 -15355 18475
rect -15325 18445 -15195 18475
rect -15165 18445 -15035 18475
rect -15005 18445 -15000 18475
rect -15520 18440 -15000 18445
rect -1680 18435 -520 18440
rect -1680 18405 -1675 18435
rect -1645 18405 -1515 18435
rect -1485 18405 -1355 18435
rect -1325 18405 -1195 18435
rect -1165 18405 -1035 18435
rect -1005 18405 -875 18435
rect -845 18405 -715 18435
rect -685 18405 -555 18435
rect -525 18405 -520 18435
rect -1680 18400 -520 18405
rect -15520 18395 -15000 18400
rect -15520 18365 -15515 18395
rect -15485 18365 -15355 18395
rect -15325 18365 -15195 18395
rect -15165 18365 -15035 18395
rect -15005 18365 -15000 18395
rect -15520 18360 -15000 18365
rect -1680 18355 -520 18360
rect -1680 18325 -1675 18355
rect -1645 18325 -1515 18355
rect -1485 18325 -1355 18355
rect -1325 18325 -1195 18355
rect -1165 18325 -1035 18355
rect -1005 18325 -875 18355
rect -845 18325 -715 18355
rect -685 18325 -555 18355
rect -525 18325 -520 18355
rect -1680 18320 -520 18325
rect -15520 18315 -15000 18320
rect -15520 18285 -15515 18315
rect -15485 18285 -15355 18315
rect -15325 18285 -15195 18315
rect -15165 18285 -15035 18315
rect -15005 18285 -15000 18315
rect -15520 18280 -15000 18285
rect -1680 18275 -520 18280
rect -1680 18245 -1675 18275
rect -1645 18245 -1515 18275
rect -1485 18245 -1355 18275
rect -1325 18245 -1195 18275
rect -1165 18245 -1035 18275
rect -1005 18245 -875 18275
rect -845 18245 -715 18275
rect -685 18245 -555 18275
rect -525 18245 -520 18275
rect -1680 18240 -520 18245
rect -15520 18235 -15000 18240
rect -15520 18205 -15515 18235
rect -15485 18205 -15355 18235
rect -15325 18205 -15195 18235
rect -15165 18205 -15035 18235
rect -15005 18205 -15000 18235
rect -15520 18200 -15000 18205
rect -1680 18195 -520 18200
rect -1680 18165 -1675 18195
rect -1645 18165 -1515 18195
rect -1485 18165 -1355 18195
rect -1325 18165 -1195 18195
rect -1165 18165 -1035 18195
rect -1005 18165 -875 18195
rect -845 18165 -715 18195
rect -685 18165 -555 18195
rect -525 18165 -520 18195
rect -1680 18160 -520 18165
rect -15520 18155 -15000 18160
rect -15520 18125 -15515 18155
rect -15485 18125 -15355 18155
rect -15325 18125 -15195 18155
rect -15165 18125 -15035 18155
rect -15005 18125 -15000 18155
rect -15520 18120 -15000 18125
rect -1680 18115 -1480 18120
rect -1680 18085 -1675 18115
rect -1645 18085 -1515 18115
rect -1485 18085 -1480 18115
rect -1680 18080 -1480 18085
rect -1440 18115 -480 18120
rect -1440 18085 -1435 18115
rect -1405 18085 -955 18115
rect -925 18085 -480 18115
rect -1440 18080 -480 18085
rect -15520 18075 -15000 18080
rect -15520 18045 -15515 18075
rect -15485 18045 -15355 18075
rect -15325 18045 -15195 18075
rect -15165 18045 -15035 18075
rect -15005 18045 -15000 18075
rect -15520 18040 -15000 18045
rect -1680 18035 -520 18040
rect -1680 18005 -1675 18035
rect -1645 18005 -1515 18035
rect -1485 18005 -1355 18035
rect -1325 18005 -1195 18035
rect -1165 18005 -1035 18035
rect -1005 18005 -875 18035
rect -845 18005 -715 18035
rect -685 18005 -555 18035
rect -525 18005 -520 18035
rect -1680 18000 -520 18005
rect 20480 18035 21600 18040
rect 20480 18005 20525 18035
rect 20555 18005 20605 18035
rect 20635 18005 20685 18035
rect 20715 18005 20765 18035
rect 20795 18005 20845 18035
rect 20875 18005 20925 18035
rect 20955 18005 21005 18035
rect 21035 18005 21085 18035
rect 21115 18005 21165 18035
rect 21195 18005 21245 18035
rect 21275 18005 21325 18035
rect 21355 18005 21405 18035
rect 21435 18005 21485 18035
rect 21515 18005 21565 18035
rect 21595 18005 21600 18035
rect 20480 18000 21600 18005
rect -15520 17995 -15000 18000
rect -15520 17965 -15515 17995
rect -15485 17965 -15355 17995
rect -15325 17965 -15195 17995
rect -15165 17965 -15035 17995
rect -15005 17965 -15000 17995
rect -15520 17960 -15000 17965
rect -1600 17955 21680 17960
rect -1600 17925 -1595 17955
rect -1565 17925 -795 17955
rect -765 17925 21680 17955
rect -1600 17920 21680 17925
rect -15520 17915 -15000 17920
rect -15520 17885 -15515 17915
rect -15485 17885 -15355 17915
rect -15325 17885 -15195 17915
rect -15165 17885 -15035 17915
rect -15005 17885 -15000 17915
rect -15520 17880 -15000 17885
rect -1680 17875 -520 17880
rect -1680 17845 -1675 17875
rect -1645 17845 -1515 17875
rect -1485 17845 -1355 17875
rect -1325 17845 -1195 17875
rect -1165 17845 -1035 17875
rect -1005 17845 -875 17875
rect -845 17845 -715 17875
rect -685 17845 -555 17875
rect -525 17845 -520 17875
rect -1680 17840 -520 17845
rect 20480 17875 21600 17880
rect 20480 17845 20525 17875
rect 20555 17845 20605 17875
rect 20635 17845 20685 17875
rect 20715 17845 20765 17875
rect 20795 17845 20845 17875
rect 20875 17845 20925 17875
rect 20955 17845 21005 17875
rect 21035 17845 21085 17875
rect 21115 17845 21165 17875
rect 21195 17845 21245 17875
rect 21275 17845 21325 17875
rect 21355 17845 21405 17875
rect 21435 17845 21485 17875
rect 21515 17845 21565 17875
rect 21595 17845 21600 17875
rect 20480 17840 21600 17845
rect -15520 17835 -15000 17840
rect -15520 17805 -15515 17835
rect -15485 17805 -15355 17835
rect -15325 17805 -15195 17835
rect -15165 17805 -15035 17835
rect -15005 17805 -15000 17835
rect -15520 17800 -15000 17805
rect -1680 17795 -520 17800
rect -1680 17765 -1675 17795
rect -1645 17765 -1515 17795
rect -1485 17765 -1355 17795
rect -1325 17765 -1195 17795
rect -1165 17765 -1035 17795
rect -1005 17765 -875 17795
rect -845 17765 -715 17795
rect -685 17765 -555 17795
rect -525 17765 -520 17795
rect -1680 17760 -520 17765
rect -15520 17755 -15000 17760
rect -15520 17725 -15515 17755
rect -15485 17725 -15355 17755
rect -15325 17725 -15195 17755
rect -15165 17725 -15035 17755
rect -15005 17725 -15000 17755
rect -15520 17720 -15000 17725
rect -1680 17715 -520 17720
rect -1680 17685 -1675 17715
rect -1645 17685 -1515 17715
rect -1485 17685 -1355 17715
rect -1325 17685 -1195 17715
rect -1165 17685 -1035 17715
rect -1005 17685 -875 17715
rect -845 17685 -715 17715
rect -685 17685 -555 17715
rect -525 17685 -520 17715
rect -1680 17680 -520 17685
rect -15520 17675 -15000 17680
rect -15520 17645 -15515 17675
rect -15485 17645 -15355 17675
rect -15325 17645 -15195 17675
rect -15165 17645 -15035 17675
rect -15005 17645 -15000 17675
rect -15520 17640 -15000 17645
rect -1680 17635 -520 17640
rect -1680 17605 -1675 17635
rect -1645 17605 -1515 17635
rect -1485 17605 -1355 17635
rect -1325 17605 -1195 17635
rect -1165 17605 -1035 17635
rect -1005 17605 -875 17635
rect -845 17605 -715 17635
rect -685 17605 -555 17635
rect -525 17605 -520 17635
rect -1680 17600 -520 17605
rect -15520 17595 -15000 17600
rect -15520 17565 -15515 17595
rect -15485 17565 -15355 17595
rect -15325 17565 -15195 17595
rect -15165 17565 -15035 17595
rect -15005 17565 -15000 17595
rect -15520 17560 -15000 17565
rect -1680 17555 -520 17560
rect -1680 17525 -1675 17555
rect -1645 17525 -1515 17555
rect -1485 17525 -1355 17555
rect -1325 17525 -1195 17555
rect -1165 17525 -1035 17555
rect -1005 17525 -875 17555
rect -845 17525 -715 17555
rect -685 17525 -555 17555
rect -525 17525 -520 17555
rect -1680 17520 -520 17525
rect -15520 17515 -15000 17520
rect -15520 17485 -15515 17515
rect -15485 17485 -15355 17515
rect -15325 17485 -15195 17515
rect -15165 17485 -15035 17515
rect -15005 17485 -15000 17515
rect -15520 17480 -15000 17485
rect -1680 17475 -520 17480
rect -1680 17445 -1675 17475
rect -1645 17445 -1515 17475
rect -1485 17445 -1355 17475
rect -1325 17445 -1195 17475
rect -1165 17445 -1035 17475
rect -1005 17445 -875 17475
rect -845 17445 -715 17475
rect -685 17445 -555 17475
rect -525 17445 -520 17475
rect -1680 17440 -520 17445
rect -15520 17435 -15000 17440
rect -15520 17405 -15515 17435
rect -15485 17405 -15355 17435
rect -15325 17405 -15195 17435
rect -15165 17405 -15035 17435
rect -15005 17405 -15000 17435
rect -15520 17400 -15000 17405
rect -1680 17395 -520 17400
rect -1680 17365 -1675 17395
rect -1645 17365 -1515 17395
rect -1485 17365 -1355 17395
rect -1325 17365 -1195 17395
rect -1165 17365 -1035 17395
rect -1005 17365 -875 17395
rect -845 17365 -715 17395
rect -685 17365 -555 17395
rect -525 17365 -520 17395
rect -1680 17360 -520 17365
rect -16560 17355 -5240 17360
rect -16560 17325 -16555 17355
rect -16525 17325 -16475 17355
rect -16445 17325 -16395 17355
rect -16365 17325 -16315 17355
rect -16285 17325 -16235 17355
rect -16205 17325 -16155 17355
rect -16125 17325 -16075 17355
rect -16045 17325 -15995 17355
rect -15965 17325 -15915 17355
rect -15885 17325 -15835 17355
rect -15805 17325 -15755 17355
rect -15725 17325 -15675 17355
rect -15645 17325 -15595 17355
rect -15565 17325 -15515 17355
rect -15485 17325 -15355 17355
rect -15325 17325 -15195 17355
rect -15165 17325 -15035 17355
rect -15005 17325 -14955 17355
rect -14925 17325 -14875 17355
rect -14845 17325 -14795 17355
rect -14765 17325 -14715 17355
rect -14685 17325 -14635 17355
rect -14605 17325 -14555 17355
rect -14525 17325 -14475 17355
rect -14445 17325 -14395 17355
rect -14365 17325 -14315 17355
rect -14285 17325 -14235 17355
rect -14205 17325 -14155 17355
rect -14125 17325 -14075 17355
rect -14045 17325 -13995 17355
rect -13965 17325 -13915 17355
rect -13885 17325 -13835 17355
rect -13805 17325 -13755 17355
rect -13725 17325 -13675 17355
rect -13645 17325 -13595 17355
rect -13565 17325 -13515 17355
rect -13485 17325 -13435 17355
rect -13405 17325 -13355 17355
rect -13325 17325 -13275 17355
rect -13245 17325 -13195 17355
rect -13165 17325 -13115 17355
rect -13085 17325 -13035 17355
rect -13005 17325 -12955 17355
rect -12925 17325 -12875 17355
rect -12845 17325 -12795 17355
rect -12765 17325 -12715 17355
rect -12685 17325 -12635 17355
rect -12605 17325 -12555 17355
rect -12525 17325 -12475 17355
rect -12445 17325 -12395 17355
rect -12365 17325 -12315 17355
rect -12285 17325 -12235 17355
rect -12205 17325 -12155 17355
rect -12125 17325 -12075 17355
rect -12045 17325 -11995 17355
rect -11965 17325 -11915 17355
rect -11885 17325 -11835 17355
rect -11805 17325 -11755 17355
rect -11725 17325 -11675 17355
rect -11645 17325 -11595 17355
rect -11565 17325 -11515 17355
rect -11485 17325 -11435 17355
rect -11405 17325 -11355 17355
rect -11325 17325 -11275 17355
rect -11245 17325 -11195 17355
rect -11165 17325 -11115 17355
rect -11085 17325 -11035 17355
rect -11005 17325 -10955 17355
rect -10925 17325 -10875 17355
rect -10845 17325 -10795 17355
rect -10765 17325 -10715 17355
rect -10685 17325 -10635 17355
rect -10605 17325 -10555 17355
rect -10525 17325 -10475 17355
rect -10445 17325 -10395 17355
rect -10365 17325 -10315 17355
rect -10285 17325 -10235 17355
rect -10205 17325 -10155 17355
rect -10125 17325 -10075 17355
rect -10045 17325 -9995 17355
rect -9965 17325 -9915 17355
rect -9885 17325 -9835 17355
rect -9805 17325 -9755 17355
rect -9725 17325 -9675 17355
rect -9645 17325 -9595 17355
rect -9565 17325 -9515 17355
rect -9485 17325 -9435 17355
rect -9405 17325 -9355 17355
rect -9325 17325 -9275 17355
rect -9245 17325 -9195 17355
rect -9165 17325 -9115 17355
rect -9085 17325 -9035 17355
rect -9005 17325 -8955 17355
rect -8925 17325 -8875 17355
rect -8845 17325 -8795 17355
rect -8765 17325 -8715 17355
rect -8685 17325 -8635 17355
rect -8605 17325 -8555 17355
rect -8525 17325 -8475 17355
rect -8445 17325 -8395 17355
rect -8365 17325 -8315 17355
rect -8285 17325 -8235 17355
rect -8205 17325 -8155 17355
rect -8125 17325 -8075 17355
rect -8045 17325 -7995 17355
rect -7965 17325 -7915 17355
rect -7885 17325 -7835 17355
rect -7805 17325 -7755 17355
rect -7725 17325 -7675 17355
rect -7645 17325 -7595 17355
rect -7565 17325 -7515 17355
rect -7485 17325 -7435 17355
rect -7405 17325 -7355 17355
rect -7325 17325 -7275 17355
rect -7245 17325 -7195 17355
rect -7165 17325 -7115 17355
rect -7085 17325 -7035 17355
rect -7005 17325 -6955 17355
rect -6925 17325 -6875 17355
rect -6845 17325 -6795 17355
rect -6765 17325 -6715 17355
rect -6685 17325 -6635 17355
rect -6605 17325 -6555 17355
rect -6525 17325 -6475 17355
rect -6445 17325 -6395 17355
rect -6365 17325 -6315 17355
rect -6285 17325 -6235 17355
rect -6205 17325 -6155 17355
rect -6125 17325 -6075 17355
rect -6045 17325 -5995 17355
rect -5965 17325 -5915 17355
rect -5885 17325 -5835 17355
rect -5805 17325 -5755 17355
rect -5725 17325 -5595 17355
rect -5565 17325 -5435 17355
rect -5405 17325 -5275 17355
rect -5245 17325 -5240 17355
rect -16560 17320 -5240 17325
rect -1680 17315 -520 17320
rect -1680 17285 -1675 17315
rect -1645 17285 -1515 17315
rect -1485 17285 -1355 17315
rect -1325 17285 -1195 17315
rect -1165 17285 -1035 17315
rect -1005 17285 -875 17315
rect -845 17285 -715 17315
rect -685 17285 -555 17315
rect -525 17285 -520 17315
rect -1680 17280 -520 17285
rect -16640 17275 -5320 17280
rect -16640 17245 -5355 17275
rect -5325 17245 -5320 17275
rect -16640 17240 -5320 17245
rect -5280 17240 -5240 17280
rect -1680 17235 -520 17240
rect -1680 17205 -1675 17235
rect -1645 17205 -1515 17235
rect -1485 17205 -1355 17235
rect -1325 17205 -1195 17235
rect -1165 17205 -1035 17235
rect -1005 17205 -875 17235
rect -845 17205 -715 17235
rect -685 17205 -555 17235
rect -525 17205 -520 17235
rect -1680 17200 -520 17205
rect -16560 17195 -5240 17200
rect -16560 17165 -16555 17195
rect -16525 17165 -16475 17195
rect -16445 17165 -16395 17195
rect -16365 17165 -16315 17195
rect -16285 17165 -16235 17195
rect -16205 17165 -16155 17195
rect -16125 17165 -16075 17195
rect -16045 17165 -15995 17195
rect -15965 17165 -15915 17195
rect -15885 17165 -15835 17195
rect -15805 17165 -15755 17195
rect -15725 17165 -15675 17195
rect -15645 17165 -15595 17195
rect -15565 17165 -15515 17195
rect -15485 17165 -15355 17195
rect -15325 17165 -15195 17195
rect -15165 17165 -15035 17195
rect -15005 17165 -14955 17195
rect -14925 17165 -14875 17195
rect -14845 17165 -14795 17195
rect -14765 17165 -14715 17195
rect -14685 17165 -14635 17195
rect -14605 17165 -14555 17195
rect -14525 17165 -14475 17195
rect -14445 17165 -14395 17195
rect -14365 17165 -14315 17195
rect -14285 17165 -14235 17195
rect -14205 17165 -14155 17195
rect -14125 17165 -14075 17195
rect -14045 17165 -13995 17195
rect -13965 17165 -13915 17195
rect -13885 17165 -13835 17195
rect -13805 17165 -13755 17195
rect -13725 17165 -13675 17195
rect -13645 17165 -13595 17195
rect -13565 17165 -13515 17195
rect -13485 17165 -13435 17195
rect -13405 17165 -13355 17195
rect -13325 17165 -13275 17195
rect -13245 17165 -13195 17195
rect -13165 17165 -13115 17195
rect -13085 17165 -13035 17195
rect -13005 17165 -12955 17195
rect -12925 17165 -12875 17195
rect -12845 17165 -12795 17195
rect -12765 17165 -12715 17195
rect -12685 17165 -12635 17195
rect -12605 17165 -12555 17195
rect -12525 17165 -12475 17195
rect -12445 17165 -12395 17195
rect -12365 17165 -12315 17195
rect -12285 17165 -12235 17195
rect -12205 17165 -12155 17195
rect -12125 17165 -12075 17195
rect -12045 17165 -11995 17195
rect -11965 17165 -11915 17195
rect -11885 17165 -11835 17195
rect -11805 17165 -11755 17195
rect -11725 17165 -11675 17195
rect -11645 17165 -11595 17195
rect -11565 17165 -11515 17195
rect -11485 17165 -11435 17195
rect -11405 17165 -11355 17195
rect -11325 17165 -11275 17195
rect -11245 17165 -11195 17195
rect -11165 17165 -11115 17195
rect -11085 17165 -11035 17195
rect -11005 17165 -10955 17195
rect -10925 17165 -10875 17195
rect -10845 17165 -10795 17195
rect -10765 17165 -10715 17195
rect -10685 17165 -10635 17195
rect -10605 17165 -10555 17195
rect -10525 17165 -10475 17195
rect -10445 17165 -10395 17195
rect -10365 17165 -10315 17195
rect -10285 17165 -10235 17195
rect -10205 17165 -10155 17195
rect -10125 17165 -10075 17195
rect -10045 17165 -9995 17195
rect -9965 17165 -9915 17195
rect -9885 17165 -9835 17195
rect -9805 17165 -9755 17195
rect -9725 17165 -9675 17195
rect -9645 17165 -9595 17195
rect -9565 17165 -9515 17195
rect -9485 17165 -9435 17195
rect -9405 17165 -9355 17195
rect -9325 17165 -9275 17195
rect -9245 17165 -9195 17195
rect -9165 17165 -9115 17195
rect -9085 17165 -9035 17195
rect -9005 17165 -8955 17195
rect -8925 17165 -8875 17195
rect -8845 17165 -8795 17195
rect -8765 17165 -8715 17195
rect -8685 17165 -8635 17195
rect -8605 17165 -8555 17195
rect -8525 17165 -8475 17195
rect -8445 17165 -8395 17195
rect -8365 17165 -8315 17195
rect -8285 17165 -8235 17195
rect -8205 17165 -8155 17195
rect -8125 17165 -8075 17195
rect -8045 17165 -7995 17195
rect -7965 17165 -7915 17195
rect -7885 17165 -7835 17195
rect -7805 17165 -7755 17195
rect -7725 17165 -7675 17195
rect -7645 17165 -7595 17195
rect -7565 17165 -7515 17195
rect -7485 17165 -7435 17195
rect -7405 17165 -7355 17195
rect -7325 17165 -7275 17195
rect -7245 17165 -7195 17195
rect -7165 17165 -7115 17195
rect -7085 17165 -7035 17195
rect -7005 17165 -6955 17195
rect -6925 17165 -6875 17195
rect -6845 17165 -6795 17195
rect -6765 17165 -6715 17195
rect -6685 17165 -6635 17195
rect -6605 17165 -6555 17195
rect -6525 17165 -6475 17195
rect -6445 17165 -6395 17195
rect -6365 17165 -6315 17195
rect -6285 17165 -6235 17195
rect -6205 17165 -6155 17195
rect -6125 17165 -6075 17195
rect -6045 17165 -5995 17195
rect -5965 17165 -5915 17195
rect -5885 17165 -5835 17195
rect -5805 17165 -5755 17195
rect -5725 17165 -5595 17195
rect -5565 17165 -5435 17195
rect -5405 17165 -5275 17195
rect -5245 17165 -5240 17195
rect -16560 17160 -5240 17165
rect -1680 17155 -520 17160
rect -1680 17125 -1675 17155
rect -1645 17125 -1515 17155
rect -1485 17125 -1355 17155
rect -1325 17125 -1195 17155
rect -1165 17125 -1035 17155
rect -1005 17125 -875 17155
rect -845 17125 -715 17155
rect -685 17125 -555 17155
rect -525 17125 -520 17155
rect -1680 17120 -520 17125
rect -15520 17115 -15000 17120
rect -15520 17085 -15515 17115
rect -15485 17085 -15355 17115
rect -15325 17085 -15195 17115
rect -15165 17085 -15035 17115
rect -15005 17085 -15000 17115
rect -15520 17080 -15000 17085
rect -1680 17075 -520 17080
rect -1680 17045 -1675 17075
rect -1645 17045 -1515 17075
rect -1485 17045 -1355 17075
rect -1325 17045 -1195 17075
rect -1165 17045 -1035 17075
rect -1005 17045 -875 17075
rect -845 17045 -715 17075
rect -685 17045 -555 17075
rect -525 17045 -520 17075
rect -1680 17040 -520 17045
rect -15520 17035 -15000 17040
rect -15520 17005 -15515 17035
rect -15485 17005 -15355 17035
rect -15325 17005 -15195 17035
rect -15165 17005 -15035 17035
rect -15005 17005 -15000 17035
rect -15520 17000 -15000 17005
rect -1680 16995 -520 17000
rect -1680 16965 -1675 16995
rect -1645 16965 -1515 16995
rect -1485 16965 -1355 16995
rect -1325 16965 -1195 16995
rect -1165 16965 -1035 16995
rect -1005 16965 -875 16995
rect -845 16965 -715 16995
rect -685 16965 -555 16995
rect -525 16965 -520 16995
rect -1680 16960 -520 16965
rect -15520 16955 -15000 16960
rect -15520 16925 -15515 16955
rect -15485 16925 -15355 16955
rect -15325 16925 -15195 16955
rect -15165 16925 -15035 16955
rect -15005 16925 -15000 16955
rect -15520 16920 -15000 16925
rect -1680 16915 -520 16920
rect -1680 16885 -1675 16915
rect -1645 16885 -1515 16915
rect -1485 16885 -1355 16915
rect -1325 16885 -1195 16915
rect -1165 16885 -1035 16915
rect -1005 16885 -875 16915
rect -845 16885 -715 16915
rect -685 16885 -555 16915
rect -525 16885 -520 16915
rect -1680 16880 -520 16885
rect -15520 16875 -15000 16880
rect -15520 16845 -15515 16875
rect -15485 16845 -15355 16875
rect -15325 16845 -15195 16875
rect -15165 16845 -15035 16875
rect -15005 16845 -15000 16875
rect -15520 16840 -15000 16845
rect -1680 16835 -520 16840
rect -1680 16805 -1675 16835
rect -1645 16805 -1515 16835
rect -1485 16805 -1355 16835
rect -1325 16805 -1195 16835
rect -1165 16805 -1035 16835
rect -1005 16805 -875 16835
rect -845 16805 -715 16835
rect -685 16805 -555 16835
rect -525 16805 -520 16835
rect -1680 16800 -520 16805
rect -15520 16795 -15000 16800
rect -15520 16765 -15515 16795
rect -15485 16765 -15355 16795
rect -15325 16765 -15195 16795
rect -15165 16765 -15035 16795
rect -15005 16765 -15000 16795
rect -15520 16760 -15000 16765
rect -1680 16755 -520 16760
rect -1680 16725 -1675 16755
rect -1645 16725 -1515 16755
rect -1485 16725 -1355 16755
rect -1325 16725 -1195 16755
rect -1165 16725 -1035 16755
rect -1005 16725 -875 16755
rect -845 16725 -715 16755
rect -685 16725 -555 16755
rect -525 16725 -520 16755
rect -1680 16720 -520 16725
rect -15520 16715 -15000 16720
rect -15520 16685 -15515 16715
rect -15485 16685 -15355 16715
rect -15325 16685 -15195 16715
rect -15165 16685 -15035 16715
rect -15005 16685 -15000 16715
rect -15520 16680 -15000 16685
rect -15520 16635 -15000 16640
rect -15520 16605 -15515 16635
rect -15485 16605 -15355 16635
rect -15325 16605 -15195 16635
rect -15165 16605 -15035 16635
rect -15005 16605 -15000 16635
rect -15520 16600 -15000 16605
rect -1680 16635 -520 16640
rect -1680 16605 -1675 16635
rect -1645 16605 -1515 16635
rect -1485 16605 -1355 16635
rect -1325 16605 -1195 16635
rect -1165 16605 -1035 16635
rect -1005 16605 -875 16635
rect -845 16605 -715 16635
rect -685 16605 -555 16635
rect -525 16605 -520 16635
rect -1680 16600 -520 16605
rect -15520 16555 -15000 16560
rect -15520 16525 -15515 16555
rect -15485 16525 -15355 16555
rect -15325 16525 -15195 16555
rect -15165 16525 -15035 16555
rect -15005 16525 -15000 16555
rect -15520 16520 -15000 16525
rect -1680 16555 -520 16560
rect -1680 16525 -1675 16555
rect -1645 16525 -1515 16555
rect -1485 16525 -1355 16555
rect -1325 16525 -1195 16555
rect -1165 16525 -1035 16555
rect -1005 16525 -875 16555
rect -845 16525 -715 16555
rect -685 16525 -555 16555
rect -525 16525 -520 16555
rect -1680 16520 -520 16525
rect -15520 16475 -520 16480
rect -15520 16445 -15515 16475
rect -15485 16445 -15355 16475
rect -15325 16445 -15195 16475
rect -15165 16445 -15035 16475
rect -15005 16445 -14955 16475
rect -14925 16445 -14875 16475
rect -14845 16445 -14795 16475
rect -14765 16445 -14715 16475
rect -14685 16445 -14635 16475
rect -14605 16445 -14555 16475
rect -14525 16445 -14475 16475
rect -14445 16445 -14395 16475
rect -14365 16445 -14315 16475
rect -14285 16445 -14235 16475
rect -14205 16445 -14155 16475
rect -14125 16445 -14075 16475
rect -14045 16445 -13995 16475
rect -13965 16445 -13915 16475
rect -13885 16445 -13835 16475
rect -13805 16445 -13755 16475
rect -13725 16445 -13675 16475
rect -13645 16445 -13595 16475
rect -13565 16445 -13515 16475
rect -13485 16445 -13435 16475
rect -13405 16445 -13355 16475
rect -13325 16445 -13275 16475
rect -13245 16445 -13195 16475
rect -13165 16445 -13115 16475
rect -13085 16445 -13035 16475
rect -13005 16445 -12955 16475
rect -12925 16445 -12875 16475
rect -12845 16445 -12795 16475
rect -12765 16445 -12715 16475
rect -12685 16445 -12635 16475
rect -12605 16445 -12555 16475
rect -12525 16445 -12475 16475
rect -12445 16445 -12395 16475
rect -12365 16445 -12315 16475
rect -12285 16445 -12235 16475
rect -12205 16445 -12155 16475
rect -12125 16445 -12075 16475
rect -12045 16445 -11995 16475
rect -11965 16445 -11915 16475
rect -11885 16445 -11835 16475
rect -11805 16445 -11755 16475
rect -11725 16445 -11675 16475
rect -11645 16445 -11595 16475
rect -11565 16445 -11515 16475
rect -11485 16445 -11435 16475
rect -11405 16445 -11355 16475
rect -11325 16445 -11275 16475
rect -11245 16445 -11195 16475
rect -11165 16445 -11115 16475
rect -11085 16445 -11035 16475
rect -11005 16445 -10955 16475
rect -10925 16445 -10875 16475
rect -10845 16445 -10795 16475
rect -10765 16445 -10715 16475
rect -10685 16445 -10635 16475
rect -10605 16445 -10555 16475
rect -10525 16445 -10475 16475
rect -10445 16445 -10395 16475
rect -10365 16445 -10315 16475
rect -10285 16445 -10235 16475
rect -10205 16445 -10155 16475
rect -10125 16445 -10075 16475
rect -10045 16445 -9995 16475
rect -9965 16445 -9915 16475
rect -9885 16445 -9835 16475
rect -9805 16445 -9755 16475
rect -9725 16445 -9675 16475
rect -9645 16445 -9595 16475
rect -9565 16445 -9515 16475
rect -9485 16445 -9435 16475
rect -9405 16445 -9355 16475
rect -9325 16445 -9275 16475
rect -9245 16445 -9195 16475
rect -9165 16445 -9115 16475
rect -9085 16445 -9035 16475
rect -9005 16445 -8955 16475
rect -8925 16445 -8875 16475
rect -8845 16445 -8795 16475
rect -8765 16445 -8715 16475
rect -8685 16445 -8635 16475
rect -8605 16445 -8555 16475
rect -8525 16445 -8475 16475
rect -8445 16445 -8395 16475
rect -8365 16445 -8315 16475
rect -8285 16445 -8235 16475
rect -8205 16445 -8155 16475
rect -8125 16445 -8075 16475
rect -8045 16445 -7995 16475
rect -7965 16445 -7915 16475
rect -7885 16445 -7835 16475
rect -7805 16445 -7755 16475
rect -7725 16445 -7675 16475
rect -7645 16445 -7595 16475
rect -7565 16445 -7515 16475
rect -7485 16445 -7435 16475
rect -7405 16445 -7355 16475
rect -7325 16445 -7275 16475
rect -7245 16445 -7195 16475
rect -7165 16445 -7115 16475
rect -7085 16445 -7035 16475
rect -7005 16445 -6955 16475
rect -6925 16445 -6875 16475
rect -6845 16445 -6795 16475
rect -6765 16445 -6715 16475
rect -6685 16445 -6635 16475
rect -6605 16445 -6555 16475
rect -6525 16445 -6475 16475
rect -6445 16445 -6395 16475
rect -6365 16445 -6315 16475
rect -6285 16445 -6235 16475
rect -6205 16445 -6155 16475
rect -6125 16445 -6075 16475
rect -6045 16445 -5995 16475
rect -5965 16445 -5915 16475
rect -5885 16445 -5835 16475
rect -5805 16445 -5755 16475
rect -5725 16445 -5595 16475
rect -5565 16445 -5435 16475
rect -5405 16445 -5355 16475
rect -5325 16445 -5275 16475
rect -5245 16445 -5195 16475
rect -5165 16445 -5115 16475
rect -5085 16445 -5035 16475
rect -5005 16445 -4955 16475
rect -4925 16445 -4875 16475
rect -4845 16445 -4795 16475
rect -4765 16445 -4715 16475
rect -4685 16445 -4635 16475
rect -4605 16445 -4555 16475
rect -4525 16445 -4475 16475
rect -4445 16445 -4395 16475
rect -4365 16445 -4315 16475
rect -4285 16445 -4235 16475
rect -4205 16445 -4155 16475
rect -4125 16445 -4075 16475
rect -4045 16445 -3995 16475
rect -3965 16445 -3915 16475
rect -3885 16445 -3835 16475
rect -3805 16445 -3755 16475
rect -3725 16445 -3675 16475
rect -3645 16445 -3595 16475
rect -3565 16445 -3515 16475
rect -3485 16445 -3435 16475
rect -3405 16445 -3355 16475
rect -3325 16445 -3275 16475
rect -3245 16445 -3195 16475
rect -3165 16445 -3115 16475
rect -3085 16445 -3035 16475
rect -3005 16445 -2955 16475
rect -2925 16445 -2875 16475
rect -2845 16445 -2795 16475
rect -2765 16445 -2715 16475
rect -2685 16445 -2635 16475
rect -2605 16445 -2555 16475
rect -2525 16445 -2475 16475
rect -2445 16445 -2395 16475
rect -2365 16445 -2315 16475
rect -2285 16445 -2235 16475
rect -2205 16445 -2155 16475
rect -2125 16445 -2075 16475
rect -2045 16445 -1995 16475
rect -1965 16445 -1835 16475
rect -1805 16445 -1755 16475
rect -1725 16445 -1675 16475
rect -1645 16445 -1595 16475
rect -1565 16445 -1515 16475
rect -1485 16445 -1435 16475
rect -1405 16445 -1355 16475
rect -1325 16445 -1195 16475
rect -1165 16445 -1035 16475
rect -1005 16445 -875 16475
rect -845 16445 -715 16475
rect -685 16445 -555 16475
rect -525 16445 -520 16475
rect -15520 16440 -520 16445
rect -15520 16395 -15320 16400
rect -15520 16365 -15515 16395
rect -15485 16365 -15355 16395
rect -15325 16365 -15320 16395
rect -15520 16360 -15320 16365
rect -15280 16395 -600 16400
rect -15280 16365 -15275 16395
rect -15245 16365 -635 16395
rect -605 16365 -600 16395
rect -15280 16360 -600 16365
rect -560 16360 -520 16400
rect -15520 16315 -520 16320
rect -15520 16285 -15515 16315
rect -15485 16285 -15355 16315
rect -15325 16285 -15195 16315
rect -15165 16285 -15035 16315
rect -15005 16285 -14955 16315
rect -14925 16285 -14875 16315
rect -14845 16285 -14795 16315
rect -14765 16285 -14715 16315
rect -14685 16285 -14635 16315
rect -14605 16285 -14555 16315
rect -14525 16285 -14475 16315
rect -14445 16285 -14395 16315
rect -14365 16285 -14315 16315
rect -14285 16285 -14235 16315
rect -14205 16285 -14155 16315
rect -14125 16285 -14075 16315
rect -14045 16285 -13995 16315
rect -13965 16285 -13915 16315
rect -13885 16285 -13835 16315
rect -13805 16285 -13755 16315
rect -13725 16285 -13675 16315
rect -13645 16285 -13595 16315
rect -13565 16285 -13515 16315
rect -13485 16285 -13435 16315
rect -13405 16285 -13355 16315
rect -13325 16285 -13275 16315
rect -13245 16285 -13195 16315
rect -13165 16285 -13115 16315
rect -13085 16285 -13035 16315
rect -13005 16285 -12955 16315
rect -12925 16285 -12875 16315
rect -12845 16285 -12795 16315
rect -12765 16285 -12715 16315
rect -12685 16285 -12635 16315
rect -12605 16285 -12555 16315
rect -12525 16285 -12475 16315
rect -12445 16285 -12395 16315
rect -12365 16285 -12315 16315
rect -12285 16285 -12235 16315
rect -12205 16285 -12155 16315
rect -12125 16285 -12075 16315
rect -12045 16285 -11995 16315
rect -11965 16285 -11915 16315
rect -11885 16285 -11835 16315
rect -11805 16285 -11755 16315
rect -11725 16285 -11675 16315
rect -11645 16285 -11595 16315
rect -11565 16285 -11515 16315
rect -11485 16285 -11435 16315
rect -11405 16285 -11355 16315
rect -11325 16285 -11275 16315
rect -11245 16285 -11195 16315
rect -11165 16285 -11115 16315
rect -11085 16285 -11035 16315
rect -11005 16285 -10955 16315
rect -10925 16285 -10875 16315
rect -10845 16285 -10795 16315
rect -10765 16285 -10715 16315
rect -10685 16285 -10635 16315
rect -10605 16285 -10555 16315
rect -10525 16285 -10475 16315
rect -10445 16285 -10395 16315
rect -10365 16285 -10315 16315
rect -10285 16285 -10235 16315
rect -10205 16285 -10155 16315
rect -10125 16285 -10075 16315
rect -10045 16285 -9995 16315
rect -9965 16285 -9915 16315
rect -9885 16285 -9835 16315
rect -9805 16285 -9755 16315
rect -9725 16285 -9675 16315
rect -9645 16285 -9595 16315
rect -9565 16285 -9515 16315
rect -9485 16285 -9435 16315
rect -9405 16285 -9355 16315
rect -9325 16285 -9275 16315
rect -9245 16285 -9195 16315
rect -9165 16285 -9115 16315
rect -9085 16285 -9035 16315
rect -9005 16285 -8955 16315
rect -8925 16285 -8875 16315
rect -8845 16285 -8795 16315
rect -8765 16285 -8715 16315
rect -8685 16285 -8635 16315
rect -8605 16285 -8555 16315
rect -8525 16285 -8475 16315
rect -8445 16285 -8395 16315
rect -8365 16285 -8315 16315
rect -8285 16285 -8235 16315
rect -8205 16285 -8155 16315
rect -8125 16285 -8075 16315
rect -8045 16285 -7995 16315
rect -7965 16285 -7915 16315
rect -7885 16285 -7835 16315
rect -7805 16285 -7755 16315
rect -7725 16285 -7675 16315
rect -7645 16285 -7595 16315
rect -7565 16285 -7515 16315
rect -7485 16285 -7435 16315
rect -7405 16285 -7355 16315
rect -7325 16285 -7275 16315
rect -7245 16285 -7195 16315
rect -7165 16285 -7115 16315
rect -7085 16285 -7035 16315
rect -7005 16285 -6955 16315
rect -6925 16285 -6875 16315
rect -6845 16285 -6795 16315
rect -6765 16285 -6715 16315
rect -6685 16285 -6635 16315
rect -6605 16285 -6555 16315
rect -6525 16285 -6475 16315
rect -6445 16285 -6395 16315
rect -6365 16285 -6315 16315
rect -6285 16285 -6235 16315
rect -6205 16285 -6155 16315
rect -6125 16285 -6075 16315
rect -6045 16285 -5995 16315
rect -5965 16285 -5915 16315
rect -5885 16285 -5835 16315
rect -5805 16285 -5755 16315
rect -5725 16285 -5595 16315
rect -5565 16285 -5435 16315
rect -5405 16285 -5355 16315
rect -5325 16285 -5275 16315
rect -5245 16285 -5195 16315
rect -5165 16285 -5115 16315
rect -5085 16285 -5035 16315
rect -5005 16285 -4955 16315
rect -4925 16285 -4875 16315
rect -4845 16285 -4795 16315
rect -4765 16285 -4715 16315
rect -4685 16285 -4635 16315
rect -4605 16285 -4555 16315
rect -4525 16285 -4475 16315
rect -4445 16285 -4395 16315
rect -4365 16285 -4315 16315
rect -4285 16285 -4235 16315
rect -4205 16285 -4155 16315
rect -4125 16285 -4075 16315
rect -4045 16285 -3995 16315
rect -3965 16285 -3915 16315
rect -3885 16285 -3835 16315
rect -3805 16285 -3755 16315
rect -3725 16285 -3675 16315
rect -3645 16285 -3595 16315
rect -3565 16285 -3515 16315
rect -3485 16285 -3435 16315
rect -3405 16285 -3355 16315
rect -3325 16285 -3275 16315
rect -3245 16285 -3195 16315
rect -3165 16285 -3115 16315
rect -3085 16285 -3035 16315
rect -3005 16285 -2955 16315
rect -2925 16285 -2875 16315
rect -2845 16285 -2795 16315
rect -2765 16285 -2715 16315
rect -2685 16285 -2635 16315
rect -2605 16285 -2555 16315
rect -2525 16285 -2475 16315
rect -2445 16285 -2395 16315
rect -2365 16285 -2315 16315
rect -2285 16285 -2235 16315
rect -2205 16285 -2155 16315
rect -2125 16285 -2075 16315
rect -2045 16285 -1995 16315
rect -1965 16285 -1835 16315
rect -1805 16285 -1755 16315
rect -1725 16285 -1675 16315
rect -1645 16285 -1595 16315
rect -1565 16285 -1515 16315
rect -1485 16285 -1435 16315
rect -1405 16285 -1355 16315
rect -1325 16285 -1195 16315
rect -1165 16285 -1035 16315
rect -1005 16285 -875 16315
rect -845 16285 -715 16315
rect -685 16285 -555 16315
rect -525 16285 -520 16315
rect -15520 16280 -520 16285
rect -15520 16235 -15160 16240
rect -15520 16205 -15515 16235
rect -15485 16205 -15355 16235
rect -15325 16205 -15160 16235
rect -15520 16200 -15160 16205
rect -15120 16235 -1240 16240
rect -15120 16205 -15115 16235
rect -15085 16205 -5675 16235
rect -5645 16205 -1275 16235
rect -1245 16205 -1240 16235
rect -15120 16200 -1240 16205
rect -1200 16200 -1160 16240
rect -1040 16200 -1000 16240
rect -880 16200 -840 16240
rect -720 16200 -680 16240
rect -560 16200 -520 16240
rect -15520 16155 -520 16160
rect -15520 16125 -15515 16155
rect -15485 16125 -15355 16155
rect -15325 16125 -15195 16155
rect -15165 16125 -15035 16155
rect -15005 16125 -14955 16155
rect -14925 16125 -14875 16155
rect -14845 16125 -14795 16155
rect -14765 16125 -14715 16155
rect -14685 16125 -14635 16155
rect -14605 16125 -14555 16155
rect -14525 16125 -14475 16155
rect -14445 16125 -14395 16155
rect -14365 16125 -14315 16155
rect -14285 16125 -14235 16155
rect -14205 16125 -14155 16155
rect -14125 16125 -14075 16155
rect -14045 16125 -13995 16155
rect -13965 16125 -13915 16155
rect -13885 16125 -13835 16155
rect -13805 16125 -13755 16155
rect -13725 16125 -13675 16155
rect -13645 16125 -13595 16155
rect -13565 16125 -13515 16155
rect -13485 16125 -13435 16155
rect -13405 16125 -13355 16155
rect -13325 16125 -13275 16155
rect -13245 16125 -13195 16155
rect -13165 16125 -13115 16155
rect -13085 16125 -13035 16155
rect -13005 16125 -12955 16155
rect -12925 16125 -12875 16155
rect -12845 16125 -12795 16155
rect -12765 16125 -12715 16155
rect -12685 16125 -12635 16155
rect -12605 16125 -12555 16155
rect -12525 16125 -12475 16155
rect -12445 16125 -12395 16155
rect -12365 16125 -12315 16155
rect -12285 16125 -12235 16155
rect -12205 16125 -12155 16155
rect -12125 16125 -12075 16155
rect -12045 16125 -11995 16155
rect -11965 16125 -11915 16155
rect -11885 16125 -11835 16155
rect -11805 16125 -11755 16155
rect -11725 16125 -11675 16155
rect -11645 16125 -11595 16155
rect -11565 16125 -11515 16155
rect -11485 16125 -11435 16155
rect -11405 16125 -11355 16155
rect -11325 16125 -11275 16155
rect -11245 16125 -11195 16155
rect -11165 16125 -11115 16155
rect -11085 16125 -11035 16155
rect -11005 16125 -10955 16155
rect -10925 16125 -10875 16155
rect -10845 16125 -10795 16155
rect -10765 16125 -10715 16155
rect -10685 16125 -10635 16155
rect -10605 16125 -10555 16155
rect -10525 16125 -10475 16155
rect -10445 16125 -10395 16155
rect -10365 16125 -10315 16155
rect -10285 16125 -10235 16155
rect -10205 16125 -10155 16155
rect -10125 16125 -10075 16155
rect -10045 16125 -9995 16155
rect -9965 16125 -9915 16155
rect -9885 16125 -9835 16155
rect -9805 16125 -9755 16155
rect -9725 16125 -9675 16155
rect -9645 16125 -9595 16155
rect -9565 16125 -9515 16155
rect -9485 16125 -9435 16155
rect -9405 16125 -9355 16155
rect -9325 16125 -9275 16155
rect -9245 16125 -9195 16155
rect -9165 16125 -9115 16155
rect -9085 16125 -9035 16155
rect -9005 16125 -8955 16155
rect -8925 16125 -8875 16155
rect -8845 16125 -8795 16155
rect -8765 16125 -8715 16155
rect -8685 16125 -8635 16155
rect -8605 16125 -8555 16155
rect -8525 16125 -8475 16155
rect -8445 16125 -8395 16155
rect -8365 16125 -8315 16155
rect -8285 16125 -8235 16155
rect -8205 16125 -8155 16155
rect -8125 16125 -8075 16155
rect -8045 16125 -7995 16155
rect -7965 16125 -7915 16155
rect -7885 16125 -7835 16155
rect -7805 16125 -7755 16155
rect -7725 16125 -7675 16155
rect -7645 16125 -7595 16155
rect -7565 16125 -7515 16155
rect -7485 16125 -7435 16155
rect -7405 16125 -7355 16155
rect -7325 16125 -7275 16155
rect -7245 16125 -7195 16155
rect -7165 16125 -7115 16155
rect -7085 16125 -7035 16155
rect -7005 16125 -6955 16155
rect -6925 16125 -6875 16155
rect -6845 16125 -6795 16155
rect -6765 16125 -6715 16155
rect -6685 16125 -6635 16155
rect -6605 16125 -6555 16155
rect -6525 16125 -6475 16155
rect -6445 16125 -6395 16155
rect -6365 16125 -6315 16155
rect -6285 16125 -6235 16155
rect -6205 16125 -6155 16155
rect -6125 16125 -6075 16155
rect -6045 16125 -5995 16155
rect -5965 16125 -5915 16155
rect -5885 16125 -5835 16155
rect -5805 16125 -5755 16155
rect -5725 16125 -5675 16155
rect -5645 16125 -5595 16155
rect -5565 16125 -5435 16155
rect -5405 16125 -5355 16155
rect -5325 16125 -5275 16155
rect -5245 16125 -5195 16155
rect -5165 16125 -5115 16155
rect -5085 16125 -5035 16155
rect -5005 16125 -4955 16155
rect -4925 16125 -4875 16155
rect -4845 16125 -4795 16155
rect -4765 16125 -4715 16155
rect -4685 16125 -4635 16155
rect -4605 16125 -4555 16155
rect -4525 16125 -4475 16155
rect -4445 16125 -4395 16155
rect -4365 16125 -4315 16155
rect -4285 16125 -4235 16155
rect -4205 16125 -4155 16155
rect -4125 16125 -4075 16155
rect -4045 16125 -3995 16155
rect -3965 16125 -3915 16155
rect -3885 16125 -3835 16155
rect -3805 16125 -3755 16155
rect -3725 16125 -3675 16155
rect -3645 16125 -3595 16155
rect -3565 16125 -3515 16155
rect -3485 16125 -3435 16155
rect -3405 16125 -3355 16155
rect -3325 16125 -3275 16155
rect -3245 16125 -3195 16155
rect -3165 16125 -3115 16155
rect -3085 16125 -3035 16155
rect -3005 16125 -2955 16155
rect -2925 16125 -2875 16155
rect -2845 16125 -2795 16155
rect -2765 16125 -2715 16155
rect -2685 16125 -2635 16155
rect -2605 16125 -2555 16155
rect -2525 16125 -2475 16155
rect -2445 16125 -2395 16155
rect -2365 16125 -2315 16155
rect -2285 16125 -2235 16155
rect -2205 16125 -2155 16155
rect -2125 16125 -2075 16155
rect -2045 16125 -1995 16155
rect -1965 16125 -1835 16155
rect -1805 16125 -1755 16155
rect -1725 16125 -1675 16155
rect -1645 16125 -1595 16155
rect -1565 16125 -1515 16155
rect -1485 16125 -1435 16155
rect -1405 16125 -1355 16155
rect -1325 16125 -1195 16155
rect -1165 16125 -1035 16155
rect -1005 16125 -875 16155
rect -845 16125 -715 16155
rect -685 16125 -555 16155
rect -525 16125 -520 16155
rect -15520 16120 -520 16125
rect -15520 16075 -15320 16080
rect -15520 16045 -15515 16075
rect -15485 16045 -15355 16075
rect -15325 16045 -15320 16075
rect -15520 16040 -15320 16045
rect -15280 16075 -1080 16080
rect -15280 16045 -15275 16075
rect -15245 16045 -5515 16075
rect -5485 16045 -1115 16075
rect -1085 16045 -1080 16075
rect -15280 16040 -1080 16045
rect -1040 16040 -1000 16080
rect -880 16040 -840 16080
rect -720 16040 -680 16080
rect -560 16040 -520 16080
rect -15520 15995 -520 16000
rect -15520 15965 -15515 15995
rect -15485 15965 -15355 15995
rect -15325 15965 -15195 15995
rect -15165 15965 -15035 15995
rect -15005 15965 -14955 15995
rect -14925 15965 -14875 15995
rect -14845 15965 -14795 15995
rect -14765 15965 -14715 15995
rect -14685 15965 -14635 15995
rect -14605 15965 -14555 15995
rect -14525 15965 -14475 15995
rect -14445 15965 -14395 15995
rect -14365 15965 -14315 15995
rect -14285 15965 -14235 15995
rect -14205 15965 -14155 15995
rect -14125 15965 -14075 15995
rect -14045 15965 -13995 15995
rect -13965 15965 -13915 15995
rect -13885 15965 -13835 15995
rect -13805 15965 -13755 15995
rect -13725 15965 -13675 15995
rect -13645 15965 -13595 15995
rect -13565 15965 -13515 15995
rect -13485 15965 -13435 15995
rect -13405 15965 -13355 15995
rect -13325 15965 -13275 15995
rect -13245 15965 -13195 15995
rect -13165 15965 -13115 15995
rect -13085 15965 -13035 15995
rect -13005 15965 -12955 15995
rect -12925 15965 -12875 15995
rect -12845 15965 -12795 15995
rect -12765 15965 -12715 15995
rect -12685 15965 -12635 15995
rect -12605 15965 -12555 15995
rect -12525 15965 -12475 15995
rect -12445 15965 -12395 15995
rect -12365 15965 -12315 15995
rect -12285 15965 -12235 15995
rect -12205 15965 -12155 15995
rect -12125 15965 -12075 15995
rect -12045 15965 -11995 15995
rect -11965 15965 -11915 15995
rect -11885 15965 -11835 15995
rect -11805 15965 -11755 15995
rect -11725 15965 -11675 15995
rect -11645 15965 -11595 15995
rect -11565 15965 -11515 15995
rect -11485 15965 -11435 15995
rect -11405 15965 -11355 15995
rect -11325 15965 -11275 15995
rect -11245 15965 -11195 15995
rect -11165 15965 -11115 15995
rect -11085 15965 -11035 15995
rect -11005 15965 -10955 15995
rect -10925 15965 -10875 15995
rect -10845 15965 -10795 15995
rect -10765 15965 -10715 15995
rect -10685 15965 -10635 15995
rect -10605 15965 -10555 15995
rect -10525 15965 -10475 15995
rect -10445 15965 -10395 15995
rect -10365 15965 -10315 15995
rect -10285 15965 -10235 15995
rect -10205 15965 -10155 15995
rect -10125 15965 -10075 15995
rect -10045 15965 -9995 15995
rect -9965 15965 -9915 15995
rect -9885 15965 -9835 15995
rect -9805 15965 -9755 15995
rect -9725 15965 -9675 15995
rect -9645 15965 -9595 15995
rect -9565 15965 -9515 15995
rect -9485 15965 -9435 15995
rect -9405 15965 -9355 15995
rect -9325 15965 -9275 15995
rect -9245 15965 -9195 15995
rect -9165 15965 -9115 15995
rect -9085 15965 -9035 15995
rect -9005 15965 -8955 15995
rect -8925 15965 -8875 15995
rect -8845 15965 -8795 15995
rect -8765 15965 -8715 15995
rect -8685 15965 -8635 15995
rect -8605 15965 -8555 15995
rect -8525 15965 -8475 15995
rect -8445 15965 -8395 15995
rect -8365 15965 -8315 15995
rect -8285 15965 -8235 15995
rect -8205 15965 -8155 15995
rect -8125 15965 -8075 15995
rect -8045 15965 -7995 15995
rect -7965 15965 -7915 15995
rect -7885 15965 -7835 15995
rect -7805 15965 -7755 15995
rect -7725 15965 -7675 15995
rect -7645 15965 -7595 15995
rect -7565 15965 -7515 15995
rect -7485 15965 -7435 15995
rect -7405 15965 -7355 15995
rect -7325 15965 -7275 15995
rect -7245 15965 -7195 15995
rect -7165 15965 -7115 15995
rect -7085 15965 -7035 15995
rect -7005 15965 -6955 15995
rect -6925 15965 -6875 15995
rect -6845 15965 -6795 15995
rect -6765 15965 -6715 15995
rect -6685 15965 -6635 15995
rect -6605 15965 -6555 15995
rect -6525 15965 -6475 15995
rect -6445 15965 -6395 15995
rect -6365 15965 -6315 15995
rect -6285 15965 -6235 15995
rect -6205 15965 -6155 15995
rect -6125 15965 -6075 15995
rect -6045 15965 -5995 15995
rect -5965 15965 -5915 15995
rect -5885 15965 -5835 15995
rect -5805 15965 -5755 15995
rect -5725 15965 -5675 15995
rect -5645 15965 -5595 15995
rect -5565 15965 -5435 15995
rect -5405 15965 -5355 15995
rect -5325 15965 -5275 15995
rect -5245 15965 -5195 15995
rect -5165 15965 -5115 15995
rect -5085 15965 -5035 15995
rect -5005 15965 -4955 15995
rect -4925 15965 -4875 15995
rect -4845 15965 -4795 15995
rect -4765 15965 -4715 15995
rect -4685 15965 -4635 15995
rect -4605 15965 -4555 15995
rect -4525 15965 -4475 15995
rect -4445 15965 -4395 15995
rect -4365 15965 -4315 15995
rect -4285 15965 -4235 15995
rect -4205 15965 -4155 15995
rect -4125 15965 -4075 15995
rect -4045 15965 -3995 15995
rect -3965 15965 -3915 15995
rect -3885 15965 -3835 15995
rect -3805 15965 -3755 15995
rect -3725 15965 -3675 15995
rect -3645 15965 -3595 15995
rect -3565 15965 -3515 15995
rect -3485 15965 -3435 15995
rect -3405 15965 -3355 15995
rect -3325 15965 -3275 15995
rect -3245 15965 -3195 15995
rect -3165 15965 -3115 15995
rect -3085 15965 -3035 15995
rect -3005 15965 -2955 15995
rect -2925 15965 -2875 15995
rect -2845 15965 -2795 15995
rect -2765 15965 -2715 15995
rect -2685 15965 -2635 15995
rect -2605 15965 -2555 15995
rect -2525 15965 -2475 15995
rect -2445 15965 -2395 15995
rect -2365 15965 -2315 15995
rect -2285 15965 -2235 15995
rect -2205 15965 -2155 15995
rect -2125 15965 -2075 15995
rect -2045 15965 -1995 15995
rect -1965 15965 -1835 15995
rect -1805 15965 -1755 15995
rect -1725 15965 -1675 15995
rect -1645 15965 -1595 15995
rect -1565 15965 -1515 15995
rect -1485 15965 -1435 15995
rect -1405 15965 -1355 15995
rect -1325 15965 -1195 15995
rect -1165 15965 -1035 15995
rect -1005 15965 -875 15995
rect -845 15965 -715 15995
rect -685 15965 -555 15995
rect -525 15965 -520 15995
rect -15520 15960 -520 15965
<< via2 >>
rect -15515 21405 -15485 21435
rect -15355 21405 -15325 21435
rect -15195 21405 -15165 21435
rect -15035 21405 -15005 21435
rect -14955 21405 -14925 21435
rect -14875 21405 -14845 21435
rect -14795 21405 -14765 21435
rect -14715 21405 -14685 21435
rect -14635 21405 -14605 21435
rect -14555 21405 -14525 21435
rect -14475 21405 -14445 21435
rect -14395 21405 -14365 21435
rect -14315 21405 -14285 21435
rect -14235 21405 -14205 21435
rect -14155 21405 -14125 21435
rect -14075 21405 -14045 21435
rect -13995 21405 -13965 21435
rect -13915 21405 -13885 21435
rect -13835 21405 -13805 21435
rect -13755 21405 -13725 21435
rect -13675 21405 -13645 21435
rect -13595 21405 -13565 21435
rect -13515 21405 -13485 21435
rect -13435 21405 -13405 21435
rect -13355 21405 -13325 21435
rect -13275 21405 -13245 21435
rect -13195 21405 -13165 21435
rect -13115 21405 -13085 21435
rect -13035 21405 -13005 21435
rect -12955 21405 -12925 21435
rect -12875 21405 -12845 21435
rect -12795 21405 -12765 21435
rect -12715 21405 -12685 21435
rect -12635 21405 -12605 21435
rect -12555 21405 -12525 21435
rect -12475 21405 -12445 21435
rect -12395 21405 -12365 21435
rect -12315 21405 -12285 21435
rect -12235 21405 -12205 21435
rect -12155 21405 -12125 21435
rect -12075 21405 -12045 21435
rect -11995 21405 -11965 21435
rect -11915 21405 -11885 21435
rect -11835 21405 -11805 21435
rect -11755 21405 -11725 21435
rect -11675 21405 -11645 21435
rect -11595 21405 -11565 21435
rect -11515 21405 -11485 21435
rect -11435 21405 -11405 21435
rect -11355 21405 -11325 21435
rect -11275 21405 -11245 21435
rect -11195 21405 -11165 21435
rect -11115 21405 -11085 21435
rect -11035 21405 -11005 21435
rect -10955 21405 -10925 21435
rect -10875 21405 -10845 21435
rect -10795 21405 -10765 21435
rect -10715 21405 -10685 21435
rect -10635 21405 -10605 21435
rect -10555 21405 -10525 21435
rect -10475 21405 -10445 21435
rect -10395 21405 -10365 21435
rect -10315 21405 -10285 21435
rect -10235 21405 -10205 21435
rect -10155 21405 -10125 21435
rect -10075 21405 -10045 21435
rect -9995 21405 -9965 21435
rect -9915 21405 -9885 21435
rect -9835 21405 -9805 21435
rect -9755 21405 -9725 21435
rect -9675 21405 -9645 21435
rect -9595 21405 -9565 21435
rect -9515 21405 -9485 21435
rect -9435 21405 -9405 21435
rect -9355 21405 -9325 21435
rect -9275 21405 -9245 21435
rect -9195 21405 -9165 21435
rect -9115 21405 -9085 21435
rect -9035 21405 -9005 21435
rect -8955 21405 -8925 21435
rect -8875 21405 -8845 21435
rect -8795 21405 -8765 21435
rect -8715 21405 -8685 21435
rect -8635 21405 -8605 21435
rect -8555 21405 -8525 21435
rect -8475 21405 -8445 21435
rect -8395 21405 -8365 21435
rect -8315 21405 -8285 21435
rect -8235 21405 -8205 21435
rect -8155 21405 -8125 21435
rect -8075 21405 -8045 21435
rect -7995 21405 -7965 21435
rect -7915 21405 -7885 21435
rect -7835 21405 -7805 21435
rect -7755 21405 -7725 21435
rect -7675 21405 -7645 21435
rect -7595 21405 -7565 21435
rect -7515 21405 -7485 21435
rect -7435 21405 -7405 21435
rect -7355 21405 -7325 21435
rect -7275 21405 -7245 21435
rect -7195 21405 -7165 21435
rect -7115 21405 -7085 21435
rect -7035 21405 -7005 21435
rect -6955 21405 -6925 21435
rect -6875 21405 -6845 21435
rect -6795 21405 -6765 21435
rect -6715 21405 -6685 21435
rect -6635 21405 -6605 21435
rect -6555 21405 -6525 21435
rect -6475 21405 -6445 21435
rect -6395 21405 -6365 21435
rect -6315 21405 -6285 21435
rect -6235 21405 -6205 21435
rect -6155 21405 -6125 21435
rect -6075 21405 -6045 21435
rect -5915 21405 -5885 21435
rect -5755 21405 -5725 21435
rect -5675 21405 -5645 21435
rect -5595 21405 -5565 21435
rect -5515 21405 -5485 21435
rect -5435 21405 -5405 21435
rect -5355 21405 -5325 21435
rect -5275 21405 -5245 21435
rect -5195 21405 -5165 21435
rect -5115 21405 -5085 21435
rect -5035 21405 -5005 21435
rect -4955 21405 -4925 21435
rect -4875 21405 -4845 21435
rect -4795 21405 -4765 21435
rect -4715 21405 -4685 21435
rect -4635 21405 -4605 21435
rect -4555 21405 -4525 21435
rect -4475 21405 -4445 21435
rect -4395 21405 -4365 21435
rect -4315 21405 -4285 21435
rect -4235 21405 -4205 21435
rect -4155 21405 -4125 21435
rect -4075 21405 -4045 21435
rect -3995 21405 -3965 21435
rect -3915 21405 -3885 21435
rect -3835 21405 -3805 21435
rect -3755 21405 -3725 21435
rect -3675 21405 -3645 21435
rect -3595 21405 -3565 21435
rect -3515 21405 -3485 21435
rect -3435 21405 -3405 21435
rect -3355 21405 -3325 21435
rect -3275 21405 -3245 21435
rect -3195 21405 -3165 21435
rect -3115 21405 -3085 21435
rect -3035 21405 -3005 21435
rect -2955 21405 -2925 21435
rect -2875 21405 -2845 21435
rect -2795 21405 -2765 21435
rect -2715 21405 -2685 21435
rect -2635 21405 -2605 21435
rect -2555 21405 -2525 21435
rect -2475 21405 -2445 21435
rect -2395 21405 -2365 21435
rect -2315 21405 -2285 21435
rect -2235 21405 -2205 21435
rect -2155 21405 -2125 21435
rect -2075 21405 -2045 21435
rect -1995 21405 -1965 21435
rect -1835 21405 -1805 21435
rect -1755 21405 -1725 21435
rect -1675 21405 -1645 21435
rect -1595 21405 -1565 21435
rect -1515 21405 -1485 21435
rect -1355 21405 -1325 21435
rect -1275 21405 -1245 21435
rect -1195 21405 -1165 21435
rect -1115 21405 -1085 21435
rect -1035 21405 -1005 21435
rect -875 21405 -845 21435
rect -715 21405 -685 21435
rect -555 21405 -525 21435
rect -15515 21325 -15485 21355
rect -15355 21325 -15325 21355
rect -15195 21325 -15165 21355
rect -15115 21325 -15085 21355
rect -5995 21325 -5965 21355
rect -1435 21325 -1405 21355
rect -15515 21245 -15485 21275
rect -15355 21245 -15325 21275
rect -15195 21245 -15165 21275
rect -15035 21245 -15005 21275
rect -14955 21245 -14925 21275
rect -14875 21245 -14845 21275
rect -14795 21245 -14765 21275
rect -14715 21245 -14685 21275
rect -14635 21245 -14605 21275
rect -14555 21245 -14525 21275
rect -14475 21245 -14445 21275
rect -14395 21245 -14365 21275
rect -14315 21245 -14285 21275
rect -14235 21245 -14205 21275
rect -14155 21245 -14125 21275
rect -14075 21245 -14045 21275
rect -13995 21245 -13965 21275
rect -13915 21245 -13885 21275
rect -13835 21245 -13805 21275
rect -13755 21245 -13725 21275
rect -13675 21245 -13645 21275
rect -13595 21245 -13565 21275
rect -13515 21245 -13485 21275
rect -13435 21245 -13405 21275
rect -13355 21245 -13325 21275
rect -13275 21245 -13245 21275
rect -13195 21245 -13165 21275
rect -13115 21245 -13085 21275
rect -13035 21245 -13005 21275
rect -12955 21245 -12925 21275
rect -12875 21245 -12845 21275
rect -12795 21245 -12765 21275
rect -12715 21245 -12685 21275
rect -12635 21245 -12605 21275
rect -12555 21245 -12525 21275
rect -12475 21245 -12445 21275
rect -12395 21245 -12365 21275
rect -12315 21245 -12285 21275
rect -12235 21245 -12205 21275
rect -12155 21245 -12125 21275
rect -12075 21245 -12045 21275
rect -11995 21245 -11965 21275
rect -11915 21245 -11885 21275
rect -11835 21245 -11805 21275
rect -11755 21245 -11725 21275
rect -11675 21245 -11645 21275
rect -11595 21245 -11565 21275
rect -11515 21245 -11485 21275
rect -11435 21245 -11405 21275
rect -11355 21245 -11325 21275
rect -11275 21245 -11245 21275
rect -11195 21245 -11165 21275
rect -11115 21245 -11085 21275
rect -11035 21245 -11005 21275
rect -10955 21245 -10925 21275
rect -10875 21245 -10845 21275
rect -10795 21245 -10765 21275
rect -10715 21245 -10685 21275
rect -10635 21245 -10605 21275
rect -10555 21245 -10525 21275
rect -10475 21245 -10445 21275
rect -10395 21245 -10365 21275
rect -10315 21245 -10285 21275
rect -10235 21245 -10205 21275
rect -10155 21245 -10125 21275
rect -10075 21245 -10045 21275
rect -9995 21245 -9965 21275
rect -9915 21245 -9885 21275
rect -9835 21245 -9805 21275
rect -9755 21245 -9725 21275
rect -9675 21245 -9645 21275
rect -9595 21245 -9565 21275
rect -9515 21245 -9485 21275
rect -9435 21245 -9405 21275
rect -9355 21245 -9325 21275
rect -9275 21245 -9245 21275
rect -9195 21245 -9165 21275
rect -9115 21245 -9085 21275
rect -9035 21245 -9005 21275
rect -8955 21245 -8925 21275
rect -8875 21245 -8845 21275
rect -8795 21245 -8765 21275
rect -8715 21245 -8685 21275
rect -8635 21245 -8605 21275
rect -8555 21245 -8525 21275
rect -8475 21245 -8445 21275
rect -8395 21245 -8365 21275
rect -8315 21245 -8285 21275
rect -8235 21245 -8205 21275
rect -8155 21245 -8125 21275
rect -8075 21245 -8045 21275
rect -7995 21245 -7965 21275
rect -7915 21245 -7885 21275
rect -7835 21245 -7805 21275
rect -7755 21245 -7725 21275
rect -7675 21245 -7645 21275
rect -7595 21245 -7565 21275
rect -7515 21245 -7485 21275
rect -7435 21245 -7405 21275
rect -7355 21245 -7325 21275
rect -7275 21245 -7245 21275
rect -7195 21245 -7165 21275
rect -7115 21245 -7085 21275
rect -7035 21245 -7005 21275
rect -6955 21245 -6925 21275
rect -6875 21245 -6845 21275
rect -6795 21245 -6765 21275
rect -6715 21245 -6685 21275
rect -6635 21245 -6605 21275
rect -6555 21245 -6525 21275
rect -6475 21245 -6445 21275
rect -6395 21245 -6365 21275
rect -6315 21245 -6285 21275
rect -6235 21245 -6205 21275
rect -6155 21245 -6125 21275
rect -6075 21245 -6045 21275
rect -5915 21245 -5885 21275
rect -5755 21245 -5725 21275
rect -5675 21245 -5645 21275
rect -5595 21245 -5565 21275
rect -5515 21245 -5485 21275
rect -5435 21245 -5405 21275
rect -5355 21245 -5325 21275
rect -5275 21245 -5245 21275
rect -5195 21245 -5165 21275
rect -5115 21245 -5085 21275
rect -5035 21245 -5005 21275
rect -4955 21245 -4925 21275
rect -4875 21245 -4845 21275
rect -4795 21245 -4765 21275
rect -4715 21245 -4685 21275
rect -4635 21245 -4605 21275
rect -4555 21245 -4525 21275
rect -4475 21245 -4445 21275
rect -4395 21245 -4365 21275
rect -4315 21245 -4285 21275
rect -4235 21245 -4205 21275
rect -4155 21245 -4125 21275
rect -4075 21245 -4045 21275
rect -3995 21245 -3965 21275
rect -3915 21245 -3885 21275
rect -3835 21245 -3805 21275
rect -3755 21245 -3725 21275
rect -3675 21245 -3645 21275
rect -3595 21245 -3565 21275
rect -3515 21245 -3485 21275
rect -3435 21245 -3405 21275
rect -3355 21245 -3325 21275
rect -3275 21245 -3245 21275
rect -3195 21245 -3165 21275
rect -3115 21245 -3085 21275
rect -3035 21245 -3005 21275
rect -2955 21245 -2925 21275
rect -2875 21245 -2845 21275
rect -2795 21245 -2765 21275
rect -2715 21245 -2685 21275
rect -2635 21245 -2605 21275
rect -2555 21245 -2525 21275
rect -2475 21245 -2445 21275
rect -2395 21245 -2365 21275
rect -2315 21245 -2285 21275
rect -2235 21245 -2205 21275
rect -2155 21245 -2125 21275
rect -2075 21245 -2045 21275
rect -1995 21245 -1965 21275
rect -1835 21245 -1805 21275
rect -1755 21245 -1725 21275
rect -1675 21245 -1645 21275
rect -1595 21245 -1565 21275
rect -1515 21245 -1485 21275
rect -1355 21245 -1325 21275
rect -1275 21245 -1245 21275
rect -1195 21245 -1165 21275
rect -1115 21245 -1085 21275
rect -1035 21245 -1005 21275
rect -875 21245 -845 21275
rect -715 21245 -685 21275
rect -555 21245 -525 21275
rect -15515 21165 -15485 21195
rect -15355 21165 -15325 21195
rect -15275 21165 -15245 21195
rect -5835 21165 -5805 21195
rect -1595 21165 -1565 21195
rect -15515 21085 -15485 21115
rect -15355 21085 -15325 21115
rect -15195 21085 -15165 21115
rect -15035 21085 -15005 21115
rect -14955 21085 -14925 21115
rect -14875 21085 -14845 21115
rect -14795 21085 -14765 21115
rect -14715 21085 -14685 21115
rect -14635 21085 -14605 21115
rect -14555 21085 -14525 21115
rect -14475 21085 -14445 21115
rect -14395 21085 -14365 21115
rect -14315 21085 -14285 21115
rect -14235 21085 -14205 21115
rect -14155 21085 -14125 21115
rect -14075 21085 -14045 21115
rect -13995 21085 -13965 21115
rect -13915 21085 -13885 21115
rect -13835 21085 -13805 21115
rect -13755 21085 -13725 21115
rect -13675 21085 -13645 21115
rect -13595 21085 -13565 21115
rect -13515 21085 -13485 21115
rect -13435 21085 -13405 21115
rect -13355 21085 -13325 21115
rect -13275 21085 -13245 21115
rect -13195 21085 -13165 21115
rect -13115 21085 -13085 21115
rect -13035 21085 -13005 21115
rect -12955 21085 -12925 21115
rect -12875 21085 -12845 21115
rect -12795 21085 -12765 21115
rect -12715 21085 -12685 21115
rect -12635 21085 -12605 21115
rect -12555 21085 -12525 21115
rect -12475 21085 -12445 21115
rect -12395 21085 -12365 21115
rect -12315 21085 -12285 21115
rect -12235 21085 -12205 21115
rect -12155 21085 -12125 21115
rect -12075 21085 -12045 21115
rect -11995 21085 -11965 21115
rect -11915 21085 -11885 21115
rect -11835 21085 -11805 21115
rect -11755 21085 -11725 21115
rect -11675 21085 -11645 21115
rect -11595 21085 -11565 21115
rect -11515 21085 -11485 21115
rect -11435 21085 -11405 21115
rect -11355 21085 -11325 21115
rect -11275 21085 -11245 21115
rect -11195 21085 -11165 21115
rect -11115 21085 -11085 21115
rect -11035 21085 -11005 21115
rect -10955 21085 -10925 21115
rect -10875 21085 -10845 21115
rect -10795 21085 -10765 21115
rect -10715 21085 -10685 21115
rect -10635 21085 -10605 21115
rect -10555 21085 -10525 21115
rect -10475 21085 -10445 21115
rect -10395 21085 -10365 21115
rect -10315 21085 -10285 21115
rect -10235 21085 -10205 21115
rect -10155 21085 -10125 21115
rect -10075 21085 -10045 21115
rect -9995 21085 -9965 21115
rect -9915 21085 -9885 21115
rect -9835 21085 -9805 21115
rect -9755 21085 -9725 21115
rect -9675 21085 -9645 21115
rect -9595 21085 -9565 21115
rect -9515 21085 -9485 21115
rect -9435 21085 -9405 21115
rect -9355 21085 -9325 21115
rect -9275 21085 -9245 21115
rect -9195 21085 -9165 21115
rect -9115 21085 -9085 21115
rect -9035 21085 -9005 21115
rect -8955 21085 -8925 21115
rect -8875 21085 -8845 21115
rect -8795 21085 -8765 21115
rect -8715 21085 -8685 21115
rect -8635 21085 -8605 21115
rect -8555 21085 -8525 21115
rect -8475 21085 -8445 21115
rect -8395 21085 -8365 21115
rect -8315 21085 -8285 21115
rect -8235 21085 -8205 21115
rect -8155 21085 -8125 21115
rect -8075 21085 -8045 21115
rect -7995 21085 -7965 21115
rect -7915 21085 -7885 21115
rect -7835 21085 -7805 21115
rect -7755 21085 -7725 21115
rect -7675 21085 -7645 21115
rect -7595 21085 -7565 21115
rect -7515 21085 -7485 21115
rect -7435 21085 -7405 21115
rect -7355 21085 -7325 21115
rect -7275 21085 -7245 21115
rect -7195 21085 -7165 21115
rect -7115 21085 -7085 21115
rect -7035 21085 -7005 21115
rect -6955 21085 -6925 21115
rect -6875 21085 -6845 21115
rect -6795 21085 -6765 21115
rect -6715 21085 -6685 21115
rect -6635 21085 -6605 21115
rect -6555 21085 -6525 21115
rect -6475 21085 -6445 21115
rect -6395 21085 -6365 21115
rect -6315 21085 -6285 21115
rect -6235 21085 -6205 21115
rect -6155 21085 -6125 21115
rect -6075 21085 -6045 21115
rect -5915 21085 -5885 21115
rect -5755 21085 -5725 21115
rect -5675 21085 -5645 21115
rect -5595 21085 -5565 21115
rect -5515 21085 -5485 21115
rect -5435 21085 -5405 21115
rect -5355 21085 -5325 21115
rect -5275 21085 -5245 21115
rect -5195 21085 -5165 21115
rect -5115 21085 -5085 21115
rect -5035 21085 -5005 21115
rect -4955 21085 -4925 21115
rect -4875 21085 -4845 21115
rect -4795 21085 -4765 21115
rect -4715 21085 -4685 21115
rect -4635 21085 -4605 21115
rect -4555 21085 -4525 21115
rect -4475 21085 -4445 21115
rect -4395 21085 -4365 21115
rect -4315 21085 -4285 21115
rect -4235 21085 -4205 21115
rect -4155 21085 -4125 21115
rect -4075 21085 -4045 21115
rect -3995 21085 -3965 21115
rect -3915 21085 -3885 21115
rect -3835 21085 -3805 21115
rect -3755 21085 -3725 21115
rect -3675 21085 -3645 21115
rect -3595 21085 -3565 21115
rect -3515 21085 -3485 21115
rect -3435 21085 -3405 21115
rect -3355 21085 -3325 21115
rect -3275 21085 -3245 21115
rect -3195 21085 -3165 21115
rect -3115 21085 -3085 21115
rect -3035 21085 -3005 21115
rect -2955 21085 -2925 21115
rect -2875 21085 -2845 21115
rect -2795 21085 -2765 21115
rect -2715 21085 -2685 21115
rect -2635 21085 -2605 21115
rect -2555 21085 -2525 21115
rect -2475 21085 -2445 21115
rect -2395 21085 -2365 21115
rect -2315 21085 -2285 21115
rect -2235 21085 -2205 21115
rect -2155 21085 -2125 21115
rect -2075 21085 -2045 21115
rect -1995 21085 -1965 21115
rect -1835 21085 -1805 21115
rect -1755 21085 -1725 21115
rect -1675 21085 -1645 21115
rect -1515 21085 -1485 21115
rect -1355 21085 -1325 21115
rect -1275 21085 -1245 21115
rect -1195 21085 -1165 21115
rect -1115 21085 -1085 21115
rect -1035 21085 -1005 21115
rect -875 21085 -845 21115
rect -715 21085 -685 21115
rect -555 21085 -525 21115
rect -15515 21005 -15485 21035
rect -15355 21005 -15325 21035
rect -15195 21005 -15165 21035
rect -15115 21005 -15085 21035
rect -635 21005 -605 21035
rect -15515 20925 -15485 20955
rect -15355 20925 -15325 20955
rect -15195 20925 -15165 20955
rect -15035 20925 -15005 20955
rect -14955 20925 -14925 20955
rect -14875 20925 -14845 20955
rect -14795 20925 -14765 20955
rect -14715 20925 -14685 20955
rect -14635 20925 -14605 20955
rect -14555 20925 -14525 20955
rect -14475 20925 -14445 20955
rect -14395 20925 -14365 20955
rect -14315 20925 -14285 20955
rect -14235 20925 -14205 20955
rect -14155 20925 -14125 20955
rect -14075 20925 -14045 20955
rect -13995 20925 -13965 20955
rect -13915 20925 -13885 20955
rect -13835 20925 -13805 20955
rect -13755 20925 -13725 20955
rect -13675 20925 -13645 20955
rect -13595 20925 -13565 20955
rect -13515 20925 -13485 20955
rect -13435 20925 -13405 20955
rect -13355 20925 -13325 20955
rect -13275 20925 -13245 20955
rect -13195 20925 -13165 20955
rect -13115 20925 -13085 20955
rect -13035 20925 -13005 20955
rect -12955 20925 -12925 20955
rect -12875 20925 -12845 20955
rect -12795 20925 -12765 20955
rect -12715 20925 -12685 20955
rect -12635 20925 -12605 20955
rect -12555 20925 -12525 20955
rect -12475 20925 -12445 20955
rect -12395 20925 -12365 20955
rect -12315 20925 -12285 20955
rect -12235 20925 -12205 20955
rect -12155 20925 -12125 20955
rect -12075 20925 -12045 20955
rect -11995 20925 -11965 20955
rect -11915 20925 -11885 20955
rect -11835 20925 -11805 20955
rect -11755 20925 -11725 20955
rect -11675 20925 -11645 20955
rect -11595 20925 -11565 20955
rect -11515 20925 -11485 20955
rect -11435 20925 -11405 20955
rect -11355 20925 -11325 20955
rect -11275 20925 -11245 20955
rect -11195 20925 -11165 20955
rect -11115 20925 -11085 20955
rect -11035 20925 -11005 20955
rect -10955 20925 -10925 20955
rect -10875 20925 -10845 20955
rect -10795 20925 -10765 20955
rect -10715 20925 -10685 20955
rect -10635 20925 -10605 20955
rect -10555 20925 -10525 20955
rect -10475 20925 -10445 20955
rect -10395 20925 -10365 20955
rect -10315 20925 -10285 20955
rect -10235 20925 -10205 20955
rect -10155 20925 -10125 20955
rect -10075 20925 -10045 20955
rect -9995 20925 -9965 20955
rect -9915 20925 -9885 20955
rect -9835 20925 -9805 20955
rect -9755 20925 -9725 20955
rect -9675 20925 -9645 20955
rect -9595 20925 -9565 20955
rect -9515 20925 -9485 20955
rect -9435 20925 -9405 20955
rect -9355 20925 -9325 20955
rect -9275 20925 -9245 20955
rect -9195 20925 -9165 20955
rect -9115 20925 -9085 20955
rect -9035 20925 -9005 20955
rect -8955 20925 -8925 20955
rect -8875 20925 -8845 20955
rect -8795 20925 -8765 20955
rect -8715 20925 -8685 20955
rect -8635 20925 -8605 20955
rect -8555 20925 -8525 20955
rect -8475 20925 -8445 20955
rect -8395 20925 -8365 20955
rect -8315 20925 -8285 20955
rect -8235 20925 -8205 20955
rect -8155 20925 -8125 20955
rect -8075 20925 -8045 20955
rect -7995 20925 -7965 20955
rect -7915 20925 -7885 20955
rect -7835 20925 -7805 20955
rect -7755 20925 -7725 20955
rect -7675 20925 -7645 20955
rect -7595 20925 -7565 20955
rect -7515 20925 -7485 20955
rect -7435 20925 -7405 20955
rect -7355 20925 -7325 20955
rect -7275 20925 -7245 20955
rect -7195 20925 -7165 20955
rect -7115 20925 -7085 20955
rect -7035 20925 -7005 20955
rect -6955 20925 -6925 20955
rect -6875 20925 -6845 20955
rect -6795 20925 -6765 20955
rect -6715 20925 -6685 20955
rect -6635 20925 -6605 20955
rect -6555 20925 -6525 20955
rect -6475 20925 -6445 20955
rect -6395 20925 -6365 20955
rect -6315 20925 -6285 20955
rect -6235 20925 -6205 20955
rect -6155 20925 -6125 20955
rect -6075 20925 -6045 20955
rect -5915 20925 -5885 20955
rect -5755 20925 -5725 20955
rect -5675 20925 -5645 20955
rect -5595 20925 -5565 20955
rect -5515 20925 -5485 20955
rect -5435 20925 -5405 20955
rect -5355 20925 -5325 20955
rect -5275 20925 -5245 20955
rect -5195 20925 -5165 20955
rect -5115 20925 -5085 20955
rect -5035 20925 -5005 20955
rect -4955 20925 -4925 20955
rect -4875 20925 -4845 20955
rect -4795 20925 -4765 20955
rect -4715 20925 -4685 20955
rect -4635 20925 -4605 20955
rect -4555 20925 -4525 20955
rect -4475 20925 -4445 20955
rect -4395 20925 -4365 20955
rect -4315 20925 -4285 20955
rect -4235 20925 -4205 20955
rect -4155 20925 -4125 20955
rect -4075 20925 -4045 20955
rect -3995 20925 -3965 20955
rect -3915 20925 -3885 20955
rect -3835 20925 -3805 20955
rect -3755 20925 -3725 20955
rect -3675 20925 -3645 20955
rect -3595 20925 -3565 20955
rect -3515 20925 -3485 20955
rect -3435 20925 -3405 20955
rect -3355 20925 -3325 20955
rect -3275 20925 -3245 20955
rect -3195 20925 -3165 20955
rect -3115 20925 -3085 20955
rect -3035 20925 -3005 20955
rect -2955 20925 -2925 20955
rect -2875 20925 -2845 20955
rect -2795 20925 -2765 20955
rect -2715 20925 -2685 20955
rect -2635 20925 -2605 20955
rect -2555 20925 -2525 20955
rect -2475 20925 -2445 20955
rect -2395 20925 -2365 20955
rect -2315 20925 -2285 20955
rect -2235 20925 -2205 20955
rect -2155 20925 -2125 20955
rect -2075 20925 -2045 20955
rect -1995 20925 -1965 20955
rect -1835 20925 -1805 20955
rect -1755 20925 -1725 20955
rect -1675 20925 -1645 20955
rect -1515 20925 -1485 20955
rect -1355 20925 -1325 20955
rect -1275 20925 -1245 20955
rect -1195 20925 -1165 20955
rect -1115 20925 -1085 20955
rect -1035 20925 -1005 20955
rect -875 20925 -845 20955
rect -715 20925 -685 20955
rect -555 20925 -525 20955
rect -15515 20845 -15485 20875
rect -15355 20845 -15325 20875
rect -15195 20845 -15165 20875
rect -15035 20845 -15005 20875
rect -6075 20845 -6045 20875
rect -5915 20845 -5885 20875
rect -5755 20845 -5725 20875
rect -1675 20845 -1645 20875
rect -1515 20845 -1485 20875
rect -1355 20845 -1325 20875
rect -1195 20845 -1165 20875
rect -1035 20845 -1005 20875
rect -875 20845 -845 20875
rect -715 20845 -685 20875
rect -555 20845 -525 20875
rect -15515 20765 -15485 20795
rect -15355 20765 -15325 20795
rect -15195 20765 -15165 20795
rect -15035 20765 -15005 20795
rect -6075 20765 -6045 20795
rect -5915 20765 -5885 20795
rect -5755 20765 -5725 20795
rect -1675 20765 -1645 20795
rect -1515 20765 -1485 20795
rect -1355 20765 -1325 20795
rect -1195 20765 -1165 20795
rect -1035 20765 -1005 20795
rect -875 20765 -845 20795
rect -715 20765 -685 20795
rect -555 20765 -525 20795
rect -16555 20645 -16525 20675
rect -16475 20645 -16445 20675
rect -16395 20645 -16365 20675
rect -16315 20645 -16285 20675
rect -16235 20645 -16205 20675
rect -16155 20645 -16125 20675
rect -16075 20645 -16045 20675
rect -15995 20645 -15965 20675
rect -15915 20645 -15885 20675
rect -15835 20645 -15805 20675
rect -15755 20645 -15725 20675
rect -15675 20645 -15645 20675
rect -15595 20645 -15565 20675
rect -14955 20645 -14925 20675
rect -14875 20645 -14845 20675
rect -14795 20645 -14765 20675
rect -14715 20645 -14685 20675
rect -14635 20645 -14605 20675
rect -14555 20645 -14525 20675
rect -14475 20645 -14445 20675
rect -14395 20645 -14365 20675
rect -14315 20645 -14285 20675
rect -14235 20645 -14205 20675
rect -14155 20645 -14125 20675
rect -14075 20645 -14045 20675
rect -13995 20645 -13965 20675
rect -13915 20645 -13885 20675
rect -13835 20645 -13805 20675
rect -13755 20645 -13725 20675
rect -13675 20645 -13645 20675
rect -13595 20645 -13565 20675
rect -13515 20645 -13485 20675
rect -13435 20645 -13405 20675
rect -13355 20645 -13325 20675
rect -13275 20645 -13245 20675
rect -13195 20645 -13165 20675
rect -13115 20645 -13085 20675
rect -13035 20645 -13005 20675
rect -12955 20645 -12925 20675
rect -12875 20645 -12845 20675
rect -12795 20645 -12765 20675
rect -12715 20645 -12685 20675
rect -12635 20645 -12605 20675
rect -12555 20645 -12525 20675
rect -12475 20645 -12445 20675
rect -12395 20645 -12365 20675
rect -12315 20645 -12285 20675
rect -12235 20645 -12205 20675
rect -12155 20645 -12125 20675
rect -12075 20645 -12045 20675
rect -11995 20645 -11965 20675
rect -11915 20645 -11885 20675
rect -11835 20645 -11805 20675
rect -11755 20645 -11725 20675
rect -11675 20645 -11645 20675
rect -11595 20645 -11565 20675
rect -11515 20645 -11485 20675
rect -11435 20645 -11405 20675
rect -11355 20645 -11325 20675
rect -11275 20645 -11245 20675
rect -11195 20645 -11165 20675
rect -11115 20645 -11085 20675
rect -11035 20645 -11005 20675
rect -10955 20645 -10925 20675
rect -10875 20645 -10845 20675
rect -10795 20645 -10765 20675
rect -10715 20645 -10685 20675
rect -10635 20645 -10605 20675
rect -10555 20645 -10525 20675
rect -10475 20645 -10445 20675
rect -10395 20645 -10365 20675
rect -10315 20645 -10285 20675
rect -10235 20645 -10205 20675
rect -10155 20645 -10125 20675
rect -10075 20645 -10045 20675
rect -9995 20645 -9965 20675
rect -9915 20645 -9885 20675
rect -9835 20645 -9805 20675
rect -9755 20645 -9725 20675
rect -9675 20645 -9645 20675
rect -9595 20645 -9565 20675
rect -9515 20645 -9485 20675
rect -9435 20645 -9405 20675
rect -9355 20645 -9325 20675
rect -9275 20645 -9245 20675
rect -9195 20645 -9165 20675
rect -9115 20645 -9085 20675
rect -9035 20645 -9005 20675
rect -8955 20645 -8925 20675
rect -8875 20645 -8845 20675
rect -8795 20645 -8765 20675
rect -8715 20645 -8685 20675
rect -8635 20645 -8605 20675
rect -8555 20645 -8525 20675
rect -8475 20645 -8445 20675
rect -8395 20645 -8365 20675
rect -8315 20645 -8285 20675
rect -8235 20645 -8205 20675
rect -8155 20645 -8125 20675
rect -8075 20645 -8045 20675
rect -7995 20645 -7965 20675
rect -7915 20645 -7885 20675
rect -7835 20645 -7805 20675
rect -7755 20645 -7725 20675
rect -7675 20645 -7645 20675
rect -7595 20645 -7565 20675
rect -7515 20645 -7485 20675
rect -7435 20645 -7405 20675
rect -7355 20645 -7325 20675
rect -7275 20645 -7245 20675
rect -7195 20645 -7165 20675
rect -7115 20645 -7085 20675
rect -7035 20645 -7005 20675
rect -6955 20645 -6925 20675
rect -6875 20645 -6845 20675
rect -6795 20645 -6765 20675
rect -6715 20645 -6685 20675
rect -6635 20645 -6605 20675
rect -6555 20645 -6525 20675
rect -6475 20645 -6445 20675
rect -6395 20645 -6365 20675
rect -6315 20645 -6285 20675
rect -6235 20645 -6205 20675
rect -6155 20645 -6125 20675
rect -5675 20645 -5645 20675
rect -5595 20645 -5565 20675
rect -5515 20645 -5485 20675
rect -5435 20645 -5405 20675
rect -5355 20645 -5325 20675
rect -5275 20645 -5245 20675
rect -5195 20645 -5165 20675
rect -5115 20645 -5085 20675
rect -5035 20645 -5005 20675
rect -4955 20645 -4925 20675
rect -4875 20645 -4845 20675
rect -4795 20645 -4765 20675
rect -4715 20645 -4685 20675
rect -4635 20645 -4605 20675
rect -4555 20645 -4525 20675
rect -4475 20645 -4445 20675
rect -4395 20645 -4365 20675
rect -4315 20645 -4285 20675
rect -4235 20645 -4205 20675
rect -4155 20645 -4125 20675
rect -4075 20645 -4045 20675
rect -3995 20645 -3965 20675
rect -3915 20645 -3885 20675
rect -3835 20645 -3805 20675
rect -3755 20645 -3725 20675
rect -3675 20645 -3645 20675
rect -3595 20645 -3565 20675
rect -3515 20645 -3485 20675
rect -3435 20645 -3405 20675
rect -3355 20645 -3325 20675
rect -3275 20645 -3245 20675
rect -3195 20645 -3165 20675
rect -3115 20645 -3085 20675
rect -3035 20645 -3005 20675
rect -2955 20645 -2925 20675
rect -2875 20645 -2845 20675
rect -2795 20645 -2765 20675
rect -2715 20645 -2685 20675
rect -2635 20645 -2605 20675
rect -2555 20645 -2525 20675
rect -2475 20645 -2445 20675
rect -2395 20645 -2365 20675
rect -2315 20645 -2285 20675
rect -2235 20645 -2205 20675
rect -2155 20645 -2125 20675
rect -2075 20645 -2045 20675
rect -1995 20645 -1965 20675
rect -1915 20645 -1885 20675
rect -1835 20645 -1805 20675
rect -1755 20645 -1725 20675
rect 20525 20645 20555 20675
rect 20605 20645 20635 20675
rect 20685 20645 20715 20675
rect 20765 20645 20795 20675
rect 20845 20645 20875 20675
rect 20925 20645 20955 20675
rect 21005 20645 21035 20675
rect 21085 20645 21115 20675
rect 21165 20645 21195 20675
rect 21245 20645 21275 20675
rect 21325 20645 21355 20675
rect 21405 20645 21435 20675
rect 21485 20645 21515 20675
rect 21565 20645 21595 20675
rect -16555 20485 -16525 20515
rect -16475 20485 -16445 20515
rect -16395 20485 -16365 20515
rect -16315 20485 -16285 20515
rect -16235 20485 -16205 20515
rect -16155 20485 -16125 20515
rect -16075 20485 -16045 20515
rect -15995 20485 -15965 20515
rect -15915 20485 -15885 20515
rect -15835 20485 -15805 20515
rect -15755 20485 -15725 20515
rect -15675 20485 -15645 20515
rect -15595 20485 -15565 20515
rect -14955 20485 -14925 20515
rect -14875 20485 -14845 20515
rect -14795 20485 -14765 20515
rect -14715 20485 -14685 20515
rect -14635 20485 -14605 20515
rect -14555 20485 -14525 20515
rect -14475 20485 -14445 20515
rect -14395 20485 -14365 20515
rect -14315 20485 -14285 20515
rect -14235 20485 -14205 20515
rect -14155 20485 -14125 20515
rect -14075 20485 -14045 20515
rect -13995 20485 -13965 20515
rect -13915 20485 -13885 20515
rect -13835 20485 -13805 20515
rect -13755 20485 -13725 20515
rect -13675 20485 -13645 20515
rect -13595 20485 -13565 20515
rect -13515 20485 -13485 20515
rect -13435 20485 -13405 20515
rect -13355 20485 -13325 20515
rect -13275 20485 -13245 20515
rect -13195 20485 -13165 20515
rect -13115 20485 -13085 20515
rect -13035 20485 -13005 20515
rect -12955 20485 -12925 20515
rect -12875 20485 -12845 20515
rect -12795 20485 -12765 20515
rect -12715 20485 -12685 20515
rect -12635 20485 -12605 20515
rect -12555 20485 -12525 20515
rect -12475 20485 -12445 20515
rect -12395 20485 -12365 20515
rect -12315 20485 -12285 20515
rect -12235 20485 -12205 20515
rect -12155 20485 -12125 20515
rect -12075 20485 -12045 20515
rect -11995 20485 -11965 20515
rect -11915 20485 -11885 20515
rect -11835 20485 -11805 20515
rect -11755 20485 -11725 20515
rect -11675 20485 -11645 20515
rect -11595 20485 -11565 20515
rect -11515 20485 -11485 20515
rect -11435 20485 -11405 20515
rect -11355 20485 -11325 20515
rect -11275 20485 -11245 20515
rect -11195 20485 -11165 20515
rect -11115 20485 -11085 20515
rect -11035 20485 -11005 20515
rect -10955 20485 -10925 20515
rect -10875 20485 -10845 20515
rect -10795 20485 -10765 20515
rect -10715 20485 -10685 20515
rect -10635 20485 -10605 20515
rect -10555 20485 -10525 20515
rect -10475 20485 -10445 20515
rect -10395 20485 -10365 20515
rect -10315 20485 -10285 20515
rect -10235 20485 -10205 20515
rect -10155 20485 -10125 20515
rect -10075 20485 -10045 20515
rect -9995 20485 -9965 20515
rect -9915 20485 -9885 20515
rect -9835 20485 -9805 20515
rect -9755 20485 -9725 20515
rect -9675 20485 -9645 20515
rect -9595 20485 -9565 20515
rect -9515 20485 -9485 20515
rect -9435 20485 -9405 20515
rect -9355 20485 -9325 20515
rect -9275 20485 -9245 20515
rect -9195 20485 -9165 20515
rect -9115 20485 -9085 20515
rect -9035 20485 -9005 20515
rect -8955 20485 -8925 20515
rect -8875 20485 -8845 20515
rect -8795 20485 -8765 20515
rect -8715 20485 -8685 20515
rect -8635 20485 -8605 20515
rect -8555 20485 -8525 20515
rect -8475 20485 -8445 20515
rect -8395 20485 -8365 20515
rect -8315 20485 -8285 20515
rect -8235 20485 -8205 20515
rect -8155 20485 -8125 20515
rect -8075 20485 -8045 20515
rect -7995 20485 -7965 20515
rect -7915 20485 -7885 20515
rect -7835 20485 -7805 20515
rect -7755 20485 -7725 20515
rect -7675 20485 -7645 20515
rect -7595 20485 -7565 20515
rect -7515 20485 -7485 20515
rect -7435 20485 -7405 20515
rect -7355 20485 -7325 20515
rect -7275 20485 -7245 20515
rect -7195 20485 -7165 20515
rect -7115 20485 -7085 20515
rect -7035 20485 -7005 20515
rect -6955 20485 -6925 20515
rect -6875 20485 -6845 20515
rect -6795 20485 -6765 20515
rect -6715 20485 -6685 20515
rect -6635 20485 -6605 20515
rect -6555 20485 -6525 20515
rect -6475 20485 -6445 20515
rect -6395 20485 -6365 20515
rect -6315 20485 -6285 20515
rect -6235 20485 -6205 20515
rect -6155 20485 -6125 20515
rect -5675 20485 -5645 20515
rect -5595 20485 -5565 20515
rect -5515 20485 -5485 20515
rect -5435 20485 -5405 20515
rect -5355 20485 -5325 20515
rect -5275 20485 -5245 20515
rect -5195 20485 -5165 20515
rect -5115 20485 -5085 20515
rect -5035 20485 -5005 20515
rect -4955 20485 -4925 20515
rect -4875 20485 -4845 20515
rect -4795 20485 -4765 20515
rect -4715 20485 -4685 20515
rect -4635 20485 -4605 20515
rect -4555 20485 -4525 20515
rect -4475 20485 -4445 20515
rect -4395 20485 -4365 20515
rect -4315 20485 -4285 20515
rect -4235 20485 -4205 20515
rect -4155 20485 -4125 20515
rect -4075 20485 -4045 20515
rect -3995 20485 -3965 20515
rect -3915 20485 -3885 20515
rect -3835 20485 -3805 20515
rect -3755 20485 -3725 20515
rect -3675 20485 -3645 20515
rect -3595 20485 -3565 20515
rect -3515 20485 -3485 20515
rect -3435 20485 -3405 20515
rect -3355 20485 -3325 20515
rect -3275 20485 -3245 20515
rect -3195 20485 -3165 20515
rect -3115 20485 -3085 20515
rect -3035 20485 -3005 20515
rect -2955 20485 -2925 20515
rect -2875 20485 -2845 20515
rect -2795 20485 -2765 20515
rect -2715 20485 -2685 20515
rect -2635 20485 -2605 20515
rect -2555 20485 -2525 20515
rect -2475 20485 -2445 20515
rect -2395 20485 -2365 20515
rect -2315 20485 -2285 20515
rect -2235 20485 -2205 20515
rect -2155 20485 -2125 20515
rect -2075 20485 -2045 20515
rect -1995 20485 -1965 20515
rect -1915 20485 -1885 20515
rect -1835 20485 -1805 20515
rect -1755 20485 -1725 20515
rect 20525 20485 20555 20515
rect 20605 20485 20635 20515
rect 20685 20485 20715 20515
rect 20765 20485 20795 20515
rect 20845 20485 20875 20515
rect 20925 20485 20955 20515
rect 21005 20485 21035 20515
rect 21085 20485 21115 20515
rect 21165 20485 21195 20515
rect 21245 20485 21275 20515
rect 21325 20485 21355 20515
rect 21405 20485 21435 20515
rect 21485 20485 21515 20515
rect 21565 20485 21595 20515
rect -6075 20405 -6045 20435
rect -5915 20405 -5885 20435
rect -5755 20405 -5725 20435
rect -1675 20405 -1645 20435
rect -1515 20405 -1485 20435
rect -1355 20405 -1325 20435
rect -1195 20405 -1165 20435
rect -1035 20405 -1005 20435
rect -875 20405 -845 20435
rect -715 20405 -685 20435
rect -555 20405 -525 20435
rect -15515 20365 -15485 20395
rect -15355 20365 -15325 20395
rect -15195 20365 -15165 20395
rect -15035 20365 -15005 20395
rect -6075 20325 -6045 20355
rect -5915 20325 -5885 20355
rect -5755 20325 -5725 20355
rect -5275 20325 -5245 20355
rect -5115 20325 -5085 20355
rect -5035 20325 -5005 20355
rect -4955 20325 -4925 20355
rect -4875 20325 -4845 20355
rect -4795 20325 -4765 20355
rect -4715 20325 -4685 20355
rect -4635 20325 -4605 20355
rect -4555 20325 -4525 20355
rect -4475 20325 -4445 20355
rect -4395 20325 -4365 20355
rect -4315 20325 -4285 20355
rect -4235 20325 -4205 20355
rect -4155 20325 -4125 20355
rect -4075 20325 -4045 20355
rect -3995 20325 -3965 20355
rect -3915 20325 -3885 20355
rect -3835 20325 -3805 20355
rect -3755 20325 -3725 20355
rect -3675 20325 -3645 20355
rect -3595 20325 -3565 20355
rect -3515 20325 -3485 20355
rect -3435 20325 -3405 20355
rect -3355 20325 -3325 20355
rect -3275 20325 -3245 20355
rect -3195 20325 -3165 20355
rect -3115 20325 -3085 20355
rect -3035 20325 -3005 20355
rect -2955 20325 -2925 20355
rect -2875 20325 -2845 20355
rect -2795 20325 -2765 20355
rect -2715 20325 -2685 20355
rect -2635 20325 -2605 20355
rect -2555 20325 -2525 20355
rect -2475 20325 -2445 20355
rect -2395 20325 -2365 20355
rect -2315 20325 -2285 20355
rect -2235 20325 -2205 20355
rect -2155 20325 -2125 20355
rect -2075 20325 -2045 20355
rect -1995 20325 -1965 20355
rect -1835 20325 -1805 20355
rect -1755 20325 -1725 20355
rect -1675 20325 -1645 20355
rect -1515 20325 -1485 20355
rect -1355 20325 -1325 20355
rect -1195 20325 -1165 20355
rect -1035 20325 -1005 20355
rect -875 20325 -845 20355
rect -715 20325 -685 20355
rect -555 20325 -525 20355
rect -15515 20285 -15485 20315
rect -15355 20285 -15325 20315
rect -15195 20285 -15165 20315
rect -15035 20285 -15005 20315
rect -5195 20245 -5165 20275
rect -635 20245 -605 20275
rect -15515 20205 -15485 20235
rect -15355 20205 -15325 20235
rect -15195 20205 -15165 20235
rect -15035 20205 -15005 20235
rect -6075 20165 -6045 20195
rect -5915 20165 -5885 20195
rect -5755 20165 -5725 20195
rect -5275 20165 -5245 20195
rect -5115 20165 -5085 20195
rect -5035 20165 -5005 20195
rect -4955 20165 -4925 20195
rect -4875 20165 -4845 20195
rect -4795 20165 -4765 20195
rect -4715 20165 -4685 20195
rect -4635 20165 -4605 20195
rect -4555 20165 -4525 20195
rect -4475 20165 -4445 20195
rect -4395 20165 -4365 20195
rect -4315 20165 -4285 20195
rect -4235 20165 -4205 20195
rect -4155 20165 -4125 20195
rect -4075 20165 -4045 20195
rect -3995 20165 -3965 20195
rect -3915 20165 -3885 20195
rect -3835 20165 -3805 20195
rect -3755 20165 -3725 20195
rect -3675 20165 -3645 20195
rect -3595 20165 -3565 20195
rect -3515 20165 -3485 20195
rect -3435 20165 -3405 20195
rect -3355 20165 -3325 20195
rect -3275 20165 -3245 20195
rect -3195 20165 -3165 20195
rect -3115 20165 -3085 20195
rect -3035 20165 -3005 20195
rect -2955 20165 -2925 20195
rect -2875 20165 -2845 20195
rect -2795 20165 -2765 20195
rect -2715 20165 -2685 20195
rect -2635 20165 -2605 20195
rect -2555 20165 -2525 20195
rect -2475 20165 -2445 20195
rect -2395 20165 -2365 20195
rect -2315 20165 -2285 20195
rect -2235 20165 -2205 20195
rect -2155 20165 -2125 20195
rect -2075 20165 -2045 20195
rect -1995 20165 -1965 20195
rect -1835 20165 -1805 20195
rect -1755 20165 -1725 20195
rect -1675 20165 -1645 20195
rect -1515 20165 -1485 20195
rect -1355 20165 -1325 20195
rect -1195 20165 -1165 20195
rect -1035 20165 -1005 20195
rect -875 20165 -845 20195
rect -715 20165 -685 20195
rect -555 20165 -525 20195
rect -15515 20125 -15485 20155
rect -15355 20125 -15325 20155
rect -15195 20125 -15165 20155
rect -15035 20125 -15005 20155
rect -1675 20085 -1645 20115
rect -1515 20085 -1485 20115
rect -1355 20085 -1325 20115
rect -1275 20085 -1245 20115
rect -955 20085 -925 20115
rect -15515 20045 -15485 20075
rect -15355 20045 -15325 20075
rect -15195 20045 -15165 20075
rect -15035 20045 -15005 20075
rect -1675 20005 -1645 20035
rect -1515 20005 -1485 20035
rect -1355 20005 -1325 20035
rect -1195 20005 -1165 20035
rect -1035 20005 -1005 20035
rect -875 20005 -845 20035
rect -715 20005 -685 20035
rect -555 20005 -525 20035
rect 20525 20005 20555 20035
rect 20605 20005 20635 20035
rect 20685 20005 20715 20035
rect 20765 20005 20795 20035
rect 20845 20005 20875 20035
rect 20925 20005 20955 20035
rect 21005 20005 21035 20035
rect 21085 20005 21115 20035
rect 21165 20005 21195 20035
rect 21245 20005 21275 20035
rect 21325 20005 21355 20035
rect 21405 20005 21435 20035
rect 21485 20005 21515 20035
rect 21565 20005 21595 20035
rect -15515 19965 -15485 19995
rect -15355 19965 -15325 19995
rect -15195 19965 -15165 19995
rect -15035 19965 -15005 19995
rect -1675 19925 -1645 19955
rect -1515 19925 -1485 19955
rect -1355 19925 -1325 19955
rect -1195 19925 -1165 19955
rect -1115 19925 -1085 19955
rect -795 19925 -765 19955
rect -15515 19885 -15485 19915
rect -15355 19885 -15325 19915
rect -15195 19885 -15165 19915
rect -15035 19885 -15005 19915
rect -1675 19845 -1645 19875
rect -1515 19845 -1485 19875
rect -1355 19845 -1325 19875
rect -1195 19845 -1165 19875
rect -1035 19845 -1005 19875
rect -875 19845 -845 19875
rect -715 19845 -685 19875
rect -555 19845 -525 19875
rect 20525 19845 20555 19875
rect 20605 19845 20635 19875
rect 20685 19845 20715 19875
rect 20765 19845 20795 19875
rect 20845 19845 20875 19875
rect 20925 19845 20955 19875
rect 21005 19845 21035 19875
rect 21085 19845 21115 19875
rect 21165 19845 21195 19875
rect 21245 19845 21275 19875
rect 21325 19845 21355 19875
rect 21405 19845 21435 19875
rect 21485 19845 21515 19875
rect 21565 19845 21595 19875
rect -15515 19805 -15485 19835
rect -15355 19805 -15325 19835
rect -15195 19805 -15165 19835
rect -15035 19805 -15005 19835
rect -1675 19765 -1645 19795
rect -1515 19765 -1485 19795
rect -1355 19765 -1325 19795
rect -1195 19765 -1165 19795
rect -1035 19765 -1005 19795
rect -875 19765 -845 19795
rect -715 19765 -685 19795
rect -555 19765 -525 19795
rect -15515 19725 -15485 19755
rect -15355 19725 -15325 19755
rect -15195 19725 -15165 19755
rect -15035 19725 -15005 19755
rect -1675 19685 -1645 19715
rect -1515 19685 -1485 19715
rect -1355 19685 -1325 19715
rect -1195 19685 -1165 19715
rect -1035 19685 -1005 19715
rect -875 19685 -845 19715
rect -715 19685 -685 19715
rect -555 19685 -525 19715
rect -15515 19645 -15485 19675
rect -15355 19645 -15325 19675
rect -15195 19645 -15165 19675
rect -15035 19645 -15005 19675
rect -1675 19605 -1645 19635
rect -1515 19605 -1485 19635
rect -1355 19605 -1325 19635
rect -1195 19605 -1165 19635
rect -1035 19605 -1005 19635
rect -875 19605 -845 19635
rect -715 19605 -685 19635
rect -555 19605 -525 19635
rect -15515 19565 -15485 19595
rect -15355 19565 -15325 19595
rect -15195 19565 -15165 19595
rect -15035 19565 -15005 19595
rect -1675 19525 -1645 19555
rect -1515 19525 -1485 19555
rect -1355 19525 -1325 19555
rect -1195 19525 -1165 19555
rect -1035 19525 -1005 19555
rect -875 19525 -845 19555
rect -715 19525 -685 19555
rect -555 19525 -525 19555
rect -15515 19485 -15485 19515
rect -15355 19485 -15325 19515
rect -15195 19485 -15165 19515
rect -15035 19485 -15005 19515
rect -1675 19445 -1645 19475
rect -1515 19445 -1485 19475
rect -1355 19445 -1325 19475
rect -1195 19445 -1165 19475
rect -1035 19445 -1005 19475
rect -875 19445 -845 19475
rect -715 19445 -685 19475
rect -555 19445 -525 19475
rect -15515 19405 -15485 19435
rect -15355 19405 -15325 19435
rect -15195 19405 -15165 19435
rect -15035 19405 -15005 19435
rect -1675 19365 -1645 19395
rect -1515 19365 -1485 19395
rect -1355 19365 -1325 19395
rect -1195 19365 -1165 19395
rect -1035 19365 -1005 19395
rect -875 19365 -845 19395
rect -715 19365 -685 19395
rect -555 19365 -525 19395
rect -15515 19325 -15485 19355
rect -15355 19325 -15325 19355
rect -15195 19325 -15165 19355
rect -15035 19325 -15005 19355
rect -1675 19285 -1645 19315
rect -1515 19285 -1485 19315
rect -1355 19285 -1325 19315
rect -1195 19285 -1165 19315
rect -1035 19285 -1005 19315
rect -875 19285 -845 19315
rect -715 19285 -685 19315
rect -555 19285 -525 19315
rect -15515 19245 -15485 19275
rect -15355 19245 -15325 19275
rect -15195 19245 -15165 19275
rect -15035 19245 -15005 19275
rect -1675 19205 -1645 19235
rect -1515 19205 -1485 19235
rect -1355 19205 -1325 19235
rect -1195 19205 -1165 19235
rect -1035 19205 -1005 19235
rect -875 19205 -845 19235
rect -715 19205 -685 19235
rect -555 19205 -525 19235
rect -15515 19165 -15485 19195
rect -15355 19165 -15325 19195
rect -15195 19165 -15165 19195
rect -15035 19165 -15005 19195
rect -1675 19125 -1645 19155
rect -1515 19125 -1485 19155
rect -1355 19125 -1325 19155
rect -1195 19125 -1165 19155
rect -1035 19125 -1005 19155
rect -875 19125 -845 19155
rect -715 19125 -685 19155
rect -555 19125 -525 19155
rect -15515 19085 -15485 19115
rect -15355 19085 -15325 19115
rect -15195 19085 -15165 19115
rect -15035 19085 -15005 19115
rect -1675 19045 -1645 19075
rect -1515 19045 -1485 19075
rect -1355 19045 -1325 19075
rect -1195 19045 -1165 19075
rect -1035 19045 -1005 19075
rect -875 19045 -845 19075
rect -715 19045 -685 19075
rect -555 19045 -525 19075
rect -15515 19005 -15485 19035
rect -15355 19005 -15325 19035
rect -15195 19005 -15165 19035
rect -15035 19005 -15005 19035
rect -1675 18965 -1645 18995
rect -1515 18965 -1485 18995
rect -1355 18965 -1325 18995
rect -1195 18965 -1165 18995
rect -1035 18965 -1005 18995
rect -875 18965 -845 18995
rect -715 18965 -685 18995
rect -555 18965 -525 18995
rect -15515 18925 -15485 18955
rect -15355 18925 -15325 18955
rect -15195 18925 -15165 18955
rect -15035 18925 -15005 18955
rect -1675 18885 -1645 18915
rect -1515 18885 -1485 18915
rect -1355 18885 -1325 18915
rect -1195 18885 -1165 18915
rect -1035 18885 -1005 18915
rect -875 18885 -845 18915
rect -715 18885 -685 18915
rect -555 18885 -525 18915
rect -16555 18845 -16525 18875
rect -16475 18845 -16445 18875
rect -16395 18845 -16365 18875
rect -16315 18845 -16285 18875
rect -16235 18845 -16205 18875
rect -16155 18845 -16125 18875
rect -16075 18845 -16045 18875
rect -15995 18845 -15965 18875
rect -15915 18845 -15885 18875
rect -15835 18845 -15805 18875
rect -15755 18845 -15725 18875
rect -15675 18845 -15645 18875
rect -15595 18845 -15565 18875
rect -15515 18845 -15485 18875
rect -15355 18845 -15325 18875
rect -15195 18845 -15165 18875
rect -15035 18845 -15005 18875
rect -1675 18805 -1645 18835
rect -1515 18805 -1485 18835
rect -1355 18805 -1325 18835
rect -1195 18805 -1165 18835
rect -1035 18805 -1005 18835
rect -875 18805 -845 18835
rect -715 18805 -685 18835
rect -635 18805 -605 18835
rect -15435 18765 -15405 18795
rect -15275 18765 -15245 18795
rect -1675 18725 -1645 18755
rect -1515 18725 -1485 18755
rect -1355 18725 -1325 18755
rect -1195 18725 -1165 18755
rect -1035 18725 -1005 18755
rect -875 18725 -845 18755
rect -715 18725 -685 18755
rect -555 18725 -525 18755
rect -16555 18685 -16525 18715
rect -16475 18685 -16445 18715
rect -16395 18685 -16365 18715
rect -16315 18685 -16285 18715
rect -16235 18685 -16205 18715
rect -16155 18685 -16125 18715
rect -16075 18685 -16045 18715
rect -15995 18685 -15965 18715
rect -15915 18685 -15885 18715
rect -15835 18685 -15805 18715
rect -15755 18685 -15725 18715
rect -15675 18685 -15645 18715
rect -15595 18685 -15565 18715
rect -15515 18685 -15485 18715
rect -15355 18685 -15325 18715
rect -15195 18685 -15165 18715
rect -15035 18685 -15005 18715
rect -1675 18645 -1645 18675
rect -1515 18645 -1485 18675
rect -1355 18645 -1325 18675
rect -1195 18645 -1165 18675
rect -1035 18645 -1005 18675
rect -875 18645 -845 18675
rect -715 18645 -685 18675
rect -555 18645 -525 18675
rect -15435 18605 -15405 18635
rect -15115 18605 -15085 18635
rect -1675 18565 -1645 18595
rect -1515 18565 -1485 18595
rect -1355 18565 -1325 18595
rect -1195 18565 -1165 18595
rect -1035 18565 -1005 18595
rect -875 18565 -845 18595
rect -715 18565 -685 18595
rect -555 18565 -525 18595
rect -16555 18525 -16525 18555
rect -16475 18525 -16445 18555
rect -16395 18525 -16365 18555
rect -16315 18525 -16285 18555
rect -16235 18525 -16205 18555
rect -16155 18525 -16125 18555
rect -16075 18525 -16045 18555
rect -15995 18525 -15965 18555
rect -15915 18525 -15885 18555
rect -15835 18525 -15805 18555
rect -15755 18525 -15725 18555
rect -15675 18525 -15645 18555
rect -15595 18525 -15565 18555
rect -15515 18525 -15485 18555
rect -15355 18525 -15325 18555
rect -15195 18525 -15165 18555
rect -15035 18525 -15005 18555
rect -1675 18485 -1645 18515
rect -1515 18485 -1485 18515
rect -1355 18485 -1325 18515
rect -1195 18485 -1165 18515
rect -1035 18485 -1005 18515
rect -875 18485 -845 18515
rect -715 18485 -685 18515
rect -555 18485 -525 18515
rect -15515 18445 -15485 18475
rect -15355 18445 -15325 18475
rect -15195 18445 -15165 18475
rect -15035 18445 -15005 18475
rect -1675 18405 -1645 18435
rect -1515 18405 -1485 18435
rect -1355 18405 -1325 18435
rect -1195 18405 -1165 18435
rect -1035 18405 -1005 18435
rect -875 18405 -845 18435
rect -715 18405 -685 18435
rect -555 18405 -525 18435
rect -15515 18365 -15485 18395
rect -15355 18365 -15325 18395
rect -15195 18365 -15165 18395
rect -15035 18365 -15005 18395
rect -1675 18325 -1645 18355
rect -1515 18325 -1485 18355
rect -1355 18325 -1325 18355
rect -1195 18325 -1165 18355
rect -1035 18325 -1005 18355
rect -875 18325 -845 18355
rect -715 18325 -685 18355
rect -555 18325 -525 18355
rect -15515 18285 -15485 18315
rect -15355 18285 -15325 18315
rect -15195 18285 -15165 18315
rect -15035 18285 -15005 18315
rect -1675 18245 -1645 18275
rect -1515 18245 -1485 18275
rect -1355 18245 -1325 18275
rect -1195 18245 -1165 18275
rect -1035 18245 -1005 18275
rect -875 18245 -845 18275
rect -715 18245 -685 18275
rect -555 18245 -525 18275
rect -15515 18205 -15485 18235
rect -15355 18205 -15325 18235
rect -15195 18205 -15165 18235
rect -15035 18205 -15005 18235
rect -1675 18165 -1645 18195
rect -1515 18165 -1485 18195
rect -1355 18165 -1325 18195
rect -1195 18165 -1165 18195
rect -1035 18165 -1005 18195
rect -875 18165 -845 18195
rect -715 18165 -685 18195
rect -555 18165 -525 18195
rect -15515 18125 -15485 18155
rect -15355 18125 -15325 18155
rect -15195 18125 -15165 18155
rect -15035 18125 -15005 18155
rect -1675 18085 -1645 18115
rect -1515 18085 -1485 18115
rect -1435 18085 -1405 18115
rect -955 18085 -925 18115
rect -15515 18045 -15485 18075
rect -15355 18045 -15325 18075
rect -15195 18045 -15165 18075
rect -15035 18045 -15005 18075
rect -1675 18005 -1645 18035
rect -1515 18005 -1485 18035
rect -1355 18005 -1325 18035
rect -1195 18005 -1165 18035
rect -1035 18005 -1005 18035
rect -875 18005 -845 18035
rect -715 18005 -685 18035
rect -555 18005 -525 18035
rect 20525 18005 20555 18035
rect 20605 18005 20635 18035
rect 20685 18005 20715 18035
rect 20765 18005 20795 18035
rect 20845 18005 20875 18035
rect 20925 18005 20955 18035
rect 21005 18005 21035 18035
rect 21085 18005 21115 18035
rect 21165 18005 21195 18035
rect 21245 18005 21275 18035
rect 21325 18005 21355 18035
rect 21405 18005 21435 18035
rect 21485 18005 21515 18035
rect 21565 18005 21595 18035
rect -15515 17965 -15485 17995
rect -15355 17965 -15325 17995
rect -15195 17965 -15165 17995
rect -15035 17965 -15005 17995
rect -1595 17925 -1565 17955
rect -795 17925 -765 17955
rect -15515 17885 -15485 17915
rect -15355 17885 -15325 17915
rect -15195 17885 -15165 17915
rect -15035 17885 -15005 17915
rect -1675 17845 -1645 17875
rect -1515 17845 -1485 17875
rect -1355 17845 -1325 17875
rect -1195 17845 -1165 17875
rect -1035 17845 -1005 17875
rect -875 17845 -845 17875
rect -715 17845 -685 17875
rect -555 17845 -525 17875
rect 20525 17845 20555 17875
rect 20605 17845 20635 17875
rect 20685 17845 20715 17875
rect 20765 17845 20795 17875
rect 20845 17845 20875 17875
rect 20925 17845 20955 17875
rect 21005 17845 21035 17875
rect 21085 17845 21115 17875
rect 21165 17845 21195 17875
rect 21245 17845 21275 17875
rect 21325 17845 21355 17875
rect 21405 17845 21435 17875
rect 21485 17845 21515 17875
rect 21565 17845 21595 17875
rect -15515 17805 -15485 17835
rect -15355 17805 -15325 17835
rect -15195 17805 -15165 17835
rect -15035 17805 -15005 17835
rect -1675 17765 -1645 17795
rect -1515 17765 -1485 17795
rect -1355 17765 -1325 17795
rect -1195 17765 -1165 17795
rect -1035 17765 -1005 17795
rect -875 17765 -845 17795
rect -715 17765 -685 17795
rect -555 17765 -525 17795
rect -15515 17725 -15485 17755
rect -15355 17725 -15325 17755
rect -15195 17725 -15165 17755
rect -15035 17725 -15005 17755
rect -1675 17685 -1645 17715
rect -1515 17685 -1485 17715
rect -1355 17685 -1325 17715
rect -1195 17685 -1165 17715
rect -1035 17685 -1005 17715
rect -875 17685 -845 17715
rect -715 17685 -685 17715
rect -555 17685 -525 17715
rect -15515 17645 -15485 17675
rect -15355 17645 -15325 17675
rect -15195 17645 -15165 17675
rect -15035 17645 -15005 17675
rect -1675 17605 -1645 17635
rect -1515 17605 -1485 17635
rect -1355 17605 -1325 17635
rect -1195 17605 -1165 17635
rect -1035 17605 -1005 17635
rect -875 17605 -845 17635
rect -715 17605 -685 17635
rect -555 17605 -525 17635
rect -15515 17565 -15485 17595
rect -15355 17565 -15325 17595
rect -15195 17565 -15165 17595
rect -15035 17565 -15005 17595
rect -1675 17525 -1645 17555
rect -1515 17525 -1485 17555
rect -1355 17525 -1325 17555
rect -1195 17525 -1165 17555
rect -1035 17525 -1005 17555
rect -875 17525 -845 17555
rect -715 17525 -685 17555
rect -555 17525 -525 17555
rect -15515 17485 -15485 17515
rect -15355 17485 -15325 17515
rect -15195 17485 -15165 17515
rect -15035 17485 -15005 17515
rect -1675 17445 -1645 17475
rect -1515 17445 -1485 17475
rect -1355 17445 -1325 17475
rect -1195 17445 -1165 17475
rect -1035 17445 -1005 17475
rect -875 17445 -845 17475
rect -715 17445 -685 17475
rect -555 17445 -525 17475
rect -15515 17405 -15485 17435
rect -15355 17405 -15325 17435
rect -15195 17405 -15165 17435
rect -15035 17405 -15005 17435
rect -1675 17365 -1645 17395
rect -1515 17365 -1485 17395
rect -1355 17365 -1325 17395
rect -1195 17365 -1165 17395
rect -1035 17365 -1005 17395
rect -875 17365 -845 17395
rect -715 17365 -685 17395
rect -555 17365 -525 17395
rect -16555 17325 -16525 17355
rect -16475 17325 -16445 17355
rect -16395 17325 -16365 17355
rect -16315 17325 -16285 17355
rect -16235 17325 -16205 17355
rect -16155 17325 -16125 17355
rect -16075 17325 -16045 17355
rect -15995 17325 -15965 17355
rect -15915 17325 -15885 17355
rect -15835 17325 -15805 17355
rect -15755 17325 -15725 17355
rect -15675 17325 -15645 17355
rect -15595 17325 -15565 17355
rect -15515 17325 -15485 17355
rect -15355 17325 -15325 17355
rect -15195 17325 -15165 17355
rect -15035 17325 -15005 17355
rect -14955 17325 -14925 17355
rect -14875 17325 -14845 17355
rect -14795 17325 -14765 17355
rect -14715 17325 -14685 17355
rect -14635 17325 -14605 17355
rect -14555 17325 -14525 17355
rect -14475 17325 -14445 17355
rect -14395 17325 -14365 17355
rect -14315 17325 -14285 17355
rect -14235 17325 -14205 17355
rect -14155 17325 -14125 17355
rect -14075 17325 -14045 17355
rect -13995 17325 -13965 17355
rect -13915 17325 -13885 17355
rect -13835 17325 -13805 17355
rect -13755 17325 -13725 17355
rect -13675 17325 -13645 17355
rect -13595 17325 -13565 17355
rect -13515 17325 -13485 17355
rect -13435 17325 -13405 17355
rect -13355 17325 -13325 17355
rect -13275 17325 -13245 17355
rect -13195 17325 -13165 17355
rect -13115 17325 -13085 17355
rect -13035 17325 -13005 17355
rect -12955 17325 -12925 17355
rect -12875 17325 -12845 17355
rect -12795 17325 -12765 17355
rect -12715 17325 -12685 17355
rect -12635 17325 -12605 17355
rect -12555 17325 -12525 17355
rect -12475 17325 -12445 17355
rect -12395 17325 -12365 17355
rect -12315 17325 -12285 17355
rect -12235 17325 -12205 17355
rect -12155 17325 -12125 17355
rect -12075 17325 -12045 17355
rect -11995 17325 -11965 17355
rect -11915 17325 -11885 17355
rect -11835 17325 -11805 17355
rect -11755 17325 -11725 17355
rect -11675 17325 -11645 17355
rect -11595 17325 -11565 17355
rect -11515 17325 -11485 17355
rect -11435 17325 -11405 17355
rect -11355 17325 -11325 17355
rect -11275 17325 -11245 17355
rect -11195 17325 -11165 17355
rect -11115 17325 -11085 17355
rect -11035 17325 -11005 17355
rect -10955 17325 -10925 17355
rect -10875 17325 -10845 17355
rect -10795 17325 -10765 17355
rect -10715 17325 -10685 17355
rect -10635 17325 -10605 17355
rect -10555 17325 -10525 17355
rect -10475 17325 -10445 17355
rect -10395 17325 -10365 17355
rect -10315 17325 -10285 17355
rect -10235 17325 -10205 17355
rect -10155 17325 -10125 17355
rect -10075 17325 -10045 17355
rect -9995 17325 -9965 17355
rect -9915 17325 -9885 17355
rect -9835 17325 -9805 17355
rect -9755 17325 -9725 17355
rect -9675 17325 -9645 17355
rect -9595 17325 -9565 17355
rect -9515 17325 -9485 17355
rect -9435 17325 -9405 17355
rect -9355 17325 -9325 17355
rect -9275 17325 -9245 17355
rect -9195 17325 -9165 17355
rect -9115 17325 -9085 17355
rect -9035 17325 -9005 17355
rect -8955 17325 -8925 17355
rect -8875 17325 -8845 17355
rect -8795 17325 -8765 17355
rect -8715 17325 -8685 17355
rect -8635 17325 -8605 17355
rect -8555 17325 -8525 17355
rect -8475 17325 -8445 17355
rect -8395 17325 -8365 17355
rect -8315 17325 -8285 17355
rect -8235 17325 -8205 17355
rect -8155 17325 -8125 17355
rect -8075 17325 -8045 17355
rect -7995 17325 -7965 17355
rect -7915 17325 -7885 17355
rect -7835 17325 -7805 17355
rect -7755 17325 -7725 17355
rect -7675 17325 -7645 17355
rect -7595 17325 -7565 17355
rect -7515 17325 -7485 17355
rect -7435 17325 -7405 17355
rect -7355 17325 -7325 17355
rect -7275 17325 -7245 17355
rect -7195 17325 -7165 17355
rect -7115 17325 -7085 17355
rect -7035 17325 -7005 17355
rect -6955 17325 -6925 17355
rect -6875 17325 -6845 17355
rect -6795 17325 -6765 17355
rect -6715 17325 -6685 17355
rect -6635 17325 -6605 17355
rect -6555 17325 -6525 17355
rect -6475 17325 -6445 17355
rect -6395 17325 -6365 17355
rect -6315 17325 -6285 17355
rect -6235 17325 -6205 17355
rect -6155 17325 -6125 17355
rect -6075 17325 -6045 17355
rect -5995 17325 -5965 17355
rect -5915 17325 -5885 17355
rect -5835 17325 -5805 17355
rect -5755 17325 -5725 17355
rect -5595 17325 -5565 17355
rect -5435 17325 -5405 17355
rect -5275 17325 -5245 17355
rect -1675 17285 -1645 17315
rect -1515 17285 -1485 17315
rect -1355 17285 -1325 17315
rect -1195 17285 -1165 17315
rect -1035 17285 -1005 17315
rect -875 17285 -845 17315
rect -715 17285 -685 17315
rect -555 17285 -525 17315
rect -5355 17245 -5325 17275
rect -1675 17205 -1645 17235
rect -1515 17205 -1485 17235
rect -1355 17205 -1325 17235
rect -1195 17205 -1165 17235
rect -1035 17205 -1005 17235
rect -875 17205 -845 17235
rect -715 17205 -685 17235
rect -555 17205 -525 17235
rect -16555 17165 -16525 17195
rect -16475 17165 -16445 17195
rect -16395 17165 -16365 17195
rect -16315 17165 -16285 17195
rect -16235 17165 -16205 17195
rect -16155 17165 -16125 17195
rect -16075 17165 -16045 17195
rect -15995 17165 -15965 17195
rect -15915 17165 -15885 17195
rect -15835 17165 -15805 17195
rect -15755 17165 -15725 17195
rect -15675 17165 -15645 17195
rect -15595 17165 -15565 17195
rect -15515 17165 -15485 17195
rect -15355 17165 -15325 17195
rect -15195 17165 -15165 17195
rect -15035 17165 -15005 17195
rect -14955 17165 -14925 17195
rect -14875 17165 -14845 17195
rect -14795 17165 -14765 17195
rect -14715 17165 -14685 17195
rect -14635 17165 -14605 17195
rect -14555 17165 -14525 17195
rect -14475 17165 -14445 17195
rect -14395 17165 -14365 17195
rect -14315 17165 -14285 17195
rect -14235 17165 -14205 17195
rect -14155 17165 -14125 17195
rect -14075 17165 -14045 17195
rect -13995 17165 -13965 17195
rect -13915 17165 -13885 17195
rect -13835 17165 -13805 17195
rect -13755 17165 -13725 17195
rect -13675 17165 -13645 17195
rect -13595 17165 -13565 17195
rect -13515 17165 -13485 17195
rect -13435 17165 -13405 17195
rect -13355 17165 -13325 17195
rect -13275 17165 -13245 17195
rect -13195 17165 -13165 17195
rect -13115 17165 -13085 17195
rect -13035 17165 -13005 17195
rect -12955 17165 -12925 17195
rect -12875 17165 -12845 17195
rect -12795 17165 -12765 17195
rect -12715 17165 -12685 17195
rect -12635 17165 -12605 17195
rect -12555 17165 -12525 17195
rect -12475 17165 -12445 17195
rect -12395 17165 -12365 17195
rect -12315 17165 -12285 17195
rect -12235 17165 -12205 17195
rect -12155 17165 -12125 17195
rect -12075 17165 -12045 17195
rect -11995 17165 -11965 17195
rect -11915 17165 -11885 17195
rect -11835 17165 -11805 17195
rect -11755 17165 -11725 17195
rect -11675 17165 -11645 17195
rect -11595 17165 -11565 17195
rect -11515 17165 -11485 17195
rect -11435 17165 -11405 17195
rect -11355 17165 -11325 17195
rect -11275 17165 -11245 17195
rect -11195 17165 -11165 17195
rect -11115 17165 -11085 17195
rect -11035 17165 -11005 17195
rect -10955 17165 -10925 17195
rect -10875 17165 -10845 17195
rect -10795 17165 -10765 17195
rect -10715 17165 -10685 17195
rect -10635 17165 -10605 17195
rect -10555 17165 -10525 17195
rect -10475 17165 -10445 17195
rect -10395 17165 -10365 17195
rect -10315 17165 -10285 17195
rect -10235 17165 -10205 17195
rect -10155 17165 -10125 17195
rect -10075 17165 -10045 17195
rect -9995 17165 -9965 17195
rect -9915 17165 -9885 17195
rect -9835 17165 -9805 17195
rect -9755 17165 -9725 17195
rect -9675 17165 -9645 17195
rect -9595 17165 -9565 17195
rect -9515 17165 -9485 17195
rect -9435 17165 -9405 17195
rect -9355 17165 -9325 17195
rect -9275 17165 -9245 17195
rect -9195 17165 -9165 17195
rect -9115 17165 -9085 17195
rect -9035 17165 -9005 17195
rect -8955 17165 -8925 17195
rect -8875 17165 -8845 17195
rect -8795 17165 -8765 17195
rect -8715 17165 -8685 17195
rect -8635 17165 -8605 17195
rect -8555 17165 -8525 17195
rect -8475 17165 -8445 17195
rect -8395 17165 -8365 17195
rect -8315 17165 -8285 17195
rect -8235 17165 -8205 17195
rect -8155 17165 -8125 17195
rect -8075 17165 -8045 17195
rect -7995 17165 -7965 17195
rect -7915 17165 -7885 17195
rect -7835 17165 -7805 17195
rect -7755 17165 -7725 17195
rect -7675 17165 -7645 17195
rect -7595 17165 -7565 17195
rect -7515 17165 -7485 17195
rect -7435 17165 -7405 17195
rect -7355 17165 -7325 17195
rect -7275 17165 -7245 17195
rect -7195 17165 -7165 17195
rect -7115 17165 -7085 17195
rect -7035 17165 -7005 17195
rect -6955 17165 -6925 17195
rect -6875 17165 -6845 17195
rect -6795 17165 -6765 17195
rect -6715 17165 -6685 17195
rect -6635 17165 -6605 17195
rect -6555 17165 -6525 17195
rect -6475 17165 -6445 17195
rect -6395 17165 -6365 17195
rect -6315 17165 -6285 17195
rect -6235 17165 -6205 17195
rect -6155 17165 -6125 17195
rect -6075 17165 -6045 17195
rect -5995 17165 -5965 17195
rect -5915 17165 -5885 17195
rect -5835 17165 -5805 17195
rect -5755 17165 -5725 17195
rect -5595 17165 -5565 17195
rect -5435 17165 -5405 17195
rect -5275 17165 -5245 17195
rect -1675 17125 -1645 17155
rect -1515 17125 -1485 17155
rect -1355 17125 -1325 17155
rect -1195 17125 -1165 17155
rect -1035 17125 -1005 17155
rect -875 17125 -845 17155
rect -715 17125 -685 17155
rect -555 17125 -525 17155
rect -15515 17085 -15485 17115
rect -15355 17085 -15325 17115
rect -15195 17085 -15165 17115
rect -15035 17085 -15005 17115
rect -1675 17045 -1645 17075
rect -1515 17045 -1485 17075
rect -1355 17045 -1325 17075
rect -1195 17045 -1165 17075
rect -1035 17045 -1005 17075
rect -875 17045 -845 17075
rect -715 17045 -685 17075
rect -555 17045 -525 17075
rect -15515 17005 -15485 17035
rect -15355 17005 -15325 17035
rect -15195 17005 -15165 17035
rect -15035 17005 -15005 17035
rect -1675 16965 -1645 16995
rect -1515 16965 -1485 16995
rect -1355 16965 -1325 16995
rect -1195 16965 -1165 16995
rect -1035 16965 -1005 16995
rect -875 16965 -845 16995
rect -715 16965 -685 16995
rect -555 16965 -525 16995
rect -15515 16925 -15485 16955
rect -15355 16925 -15325 16955
rect -15195 16925 -15165 16955
rect -15035 16925 -15005 16955
rect -1675 16885 -1645 16915
rect -1515 16885 -1485 16915
rect -1355 16885 -1325 16915
rect -1195 16885 -1165 16915
rect -1035 16885 -1005 16915
rect -875 16885 -845 16915
rect -715 16885 -685 16915
rect -555 16885 -525 16915
rect -15515 16845 -15485 16875
rect -15355 16845 -15325 16875
rect -15195 16845 -15165 16875
rect -15035 16845 -15005 16875
rect -1675 16805 -1645 16835
rect -1515 16805 -1485 16835
rect -1355 16805 -1325 16835
rect -1195 16805 -1165 16835
rect -1035 16805 -1005 16835
rect -875 16805 -845 16835
rect -715 16805 -685 16835
rect -555 16805 -525 16835
rect -15515 16765 -15485 16795
rect -15355 16765 -15325 16795
rect -15195 16765 -15165 16795
rect -15035 16765 -15005 16795
rect -1675 16725 -1645 16755
rect -1515 16725 -1485 16755
rect -1355 16725 -1325 16755
rect -1195 16725 -1165 16755
rect -1035 16725 -1005 16755
rect -875 16725 -845 16755
rect -715 16725 -685 16755
rect -555 16725 -525 16755
rect -15515 16685 -15485 16715
rect -15355 16685 -15325 16715
rect -15195 16685 -15165 16715
rect -15035 16685 -15005 16715
rect -15515 16605 -15485 16635
rect -15355 16605 -15325 16635
rect -15195 16605 -15165 16635
rect -15035 16605 -15005 16635
rect -1675 16605 -1645 16635
rect -1515 16605 -1485 16635
rect -1355 16605 -1325 16635
rect -1195 16605 -1165 16635
rect -1035 16605 -1005 16635
rect -875 16605 -845 16635
rect -715 16605 -685 16635
rect -555 16605 -525 16635
rect -15515 16525 -15485 16555
rect -15355 16525 -15325 16555
rect -15195 16525 -15165 16555
rect -15035 16525 -15005 16555
rect -1675 16525 -1645 16555
rect -1515 16525 -1485 16555
rect -1355 16525 -1325 16555
rect -1195 16525 -1165 16555
rect -1035 16525 -1005 16555
rect -875 16525 -845 16555
rect -715 16525 -685 16555
rect -555 16525 -525 16555
rect -15515 16445 -15485 16475
rect -15355 16445 -15325 16475
rect -15195 16445 -15165 16475
rect -15035 16445 -15005 16475
rect -14955 16445 -14925 16475
rect -14875 16445 -14845 16475
rect -14795 16445 -14765 16475
rect -14715 16445 -14685 16475
rect -14635 16445 -14605 16475
rect -14555 16445 -14525 16475
rect -14475 16445 -14445 16475
rect -14395 16445 -14365 16475
rect -14315 16445 -14285 16475
rect -14235 16445 -14205 16475
rect -14155 16445 -14125 16475
rect -14075 16445 -14045 16475
rect -13995 16445 -13965 16475
rect -13915 16445 -13885 16475
rect -13835 16445 -13805 16475
rect -13755 16445 -13725 16475
rect -13675 16445 -13645 16475
rect -13595 16445 -13565 16475
rect -13515 16445 -13485 16475
rect -13435 16445 -13405 16475
rect -13355 16445 -13325 16475
rect -13275 16445 -13245 16475
rect -13195 16445 -13165 16475
rect -13115 16445 -13085 16475
rect -13035 16445 -13005 16475
rect -12955 16445 -12925 16475
rect -12875 16445 -12845 16475
rect -12795 16445 -12765 16475
rect -12715 16445 -12685 16475
rect -12635 16445 -12605 16475
rect -12555 16445 -12525 16475
rect -12475 16445 -12445 16475
rect -12395 16445 -12365 16475
rect -12315 16445 -12285 16475
rect -12235 16445 -12205 16475
rect -12155 16445 -12125 16475
rect -12075 16445 -12045 16475
rect -11995 16445 -11965 16475
rect -11915 16445 -11885 16475
rect -11835 16445 -11805 16475
rect -11755 16445 -11725 16475
rect -11675 16445 -11645 16475
rect -11595 16445 -11565 16475
rect -11515 16445 -11485 16475
rect -11435 16445 -11405 16475
rect -11355 16445 -11325 16475
rect -11275 16445 -11245 16475
rect -11195 16445 -11165 16475
rect -11115 16445 -11085 16475
rect -11035 16445 -11005 16475
rect -10955 16445 -10925 16475
rect -10875 16445 -10845 16475
rect -10795 16445 -10765 16475
rect -10715 16445 -10685 16475
rect -10635 16445 -10605 16475
rect -10555 16445 -10525 16475
rect -10475 16445 -10445 16475
rect -10395 16445 -10365 16475
rect -10315 16445 -10285 16475
rect -10235 16445 -10205 16475
rect -10155 16445 -10125 16475
rect -10075 16445 -10045 16475
rect -9995 16445 -9965 16475
rect -9915 16445 -9885 16475
rect -9835 16445 -9805 16475
rect -9755 16445 -9725 16475
rect -9675 16445 -9645 16475
rect -9595 16445 -9565 16475
rect -9515 16445 -9485 16475
rect -9435 16445 -9405 16475
rect -9355 16445 -9325 16475
rect -9275 16445 -9245 16475
rect -9195 16445 -9165 16475
rect -9115 16445 -9085 16475
rect -9035 16445 -9005 16475
rect -8955 16445 -8925 16475
rect -8875 16445 -8845 16475
rect -8795 16445 -8765 16475
rect -8715 16445 -8685 16475
rect -8635 16445 -8605 16475
rect -8555 16445 -8525 16475
rect -8475 16445 -8445 16475
rect -8395 16445 -8365 16475
rect -8315 16445 -8285 16475
rect -8235 16445 -8205 16475
rect -8155 16445 -8125 16475
rect -8075 16445 -8045 16475
rect -7995 16445 -7965 16475
rect -7915 16445 -7885 16475
rect -7835 16445 -7805 16475
rect -7755 16445 -7725 16475
rect -7675 16445 -7645 16475
rect -7595 16445 -7565 16475
rect -7515 16445 -7485 16475
rect -7435 16445 -7405 16475
rect -7355 16445 -7325 16475
rect -7275 16445 -7245 16475
rect -7195 16445 -7165 16475
rect -7115 16445 -7085 16475
rect -7035 16445 -7005 16475
rect -6955 16445 -6925 16475
rect -6875 16445 -6845 16475
rect -6795 16445 -6765 16475
rect -6715 16445 -6685 16475
rect -6635 16445 -6605 16475
rect -6555 16445 -6525 16475
rect -6475 16445 -6445 16475
rect -6395 16445 -6365 16475
rect -6315 16445 -6285 16475
rect -6235 16445 -6205 16475
rect -6155 16445 -6125 16475
rect -6075 16445 -6045 16475
rect -5995 16445 -5965 16475
rect -5915 16445 -5885 16475
rect -5835 16445 -5805 16475
rect -5755 16445 -5725 16475
rect -5595 16445 -5565 16475
rect -5435 16445 -5405 16475
rect -5355 16445 -5325 16475
rect -5275 16445 -5245 16475
rect -5195 16445 -5165 16475
rect -5115 16445 -5085 16475
rect -5035 16445 -5005 16475
rect -4955 16445 -4925 16475
rect -4875 16445 -4845 16475
rect -4795 16445 -4765 16475
rect -4715 16445 -4685 16475
rect -4635 16445 -4605 16475
rect -4555 16445 -4525 16475
rect -4475 16445 -4445 16475
rect -4395 16445 -4365 16475
rect -4315 16445 -4285 16475
rect -4235 16445 -4205 16475
rect -4155 16445 -4125 16475
rect -4075 16445 -4045 16475
rect -3995 16445 -3965 16475
rect -3915 16445 -3885 16475
rect -3835 16445 -3805 16475
rect -3755 16445 -3725 16475
rect -3675 16445 -3645 16475
rect -3595 16445 -3565 16475
rect -3515 16445 -3485 16475
rect -3435 16445 -3405 16475
rect -3355 16445 -3325 16475
rect -3275 16445 -3245 16475
rect -3195 16445 -3165 16475
rect -3115 16445 -3085 16475
rect -3035 16445 -3005 16475
rect -2955 16445 -2925 16475
rect -2875 16445 -2845 16475
rect -2795 16445 -2765 16475
rect -2715 16445 -2685 16475
rect -2635 16445 -2605 16475
rect -2555 16445 -2525 16475
rect -2475 16445 -2445 16475
rect -2395 16445 -2365 16475
rect -2315 16445 -2285 16475
rect -2235 16445 -2205 16475
rect -2155 16445 -2125 16475
rect -2075 16445 -2045 16475
rect -1995 16445 -1965 16475
rect -1835 16445 -1805 16475
rect -1755 16445 -1725 16475
rect -1675 16445 -1645 16475
rect -1595 16445 -1565 16475
rect -1515 16445 -1485 16475
rect -1435 16445 -1405 16475
rect -1355 16445 -1325 16475
rect -1195 16445 -1165 16475
rect -1035 16445 -1005 16475
rect -875 16445 -845 16475
rect -715 16445 -685 16475
rect -555 16445 -525 16475
rect -15515 16365 -15485 16395
rect -15355 16365 -15325 16395
rect -15275 16365 -15245 16395
rect -635 16365 -605 16395
rect -15515 16285 -15485 16315
rect -15355 16285 -15325 16315
rect -15195 16285 -15165 16315
rect -15035 16285 -15005 16315
rect -14955 16285 -14925 16315
rect -14875 16285 -14845 16315
rect -14795 16285 -14765 16315
rect -14715 16285 -14685 16315
rect -14635 16285 -14605 16315
rect -14555 16285 -14525 16315
rect -14475 16285 -14445 16315
rect -14395 16285 -14365 16315
rect -14315 16285 -14285 16315
rect -14235 16285 -14205 16315
rect -14155 16285 -14125 16315
rect -14075 16285 -14045 16315
rect -13995 16285 -13965 16315
rect -13915 16285 -13885 16315
rect -13835 16285 -13805 16315
rect -13755 16285 -13725 16315
rect -13675 16285 -13645 16315
rect -13595 16285 -13565 16315
rect -13515 16285 -13485 16315
rect -13435 16285 -13405 16315
rect -13355 16285 -13325 16315
rect -13275 16285 -13245 16315
rect -13195 16285 -13165 16315
rect -13115 16285 -13085 16315
rect -13035 16285 -13005 16315
rect -12955 16285 -12925 16315
rect -12875 16285 -12845 16315
rect -12795 16285 -12765 16315
rect -12715 16285 -12685 16315
rect -12635 16285 -12605 16315
rect -12555 16285 -12525 16315
rect -12475 16285 -12445 16315
rect -12395 16285 -12365 16315
rect -12315 16285 -12285 16315
rect -12235 16285 -12205 16315
rect -12155 16285 -12125 16315
rect -12075 16285 -12045 16315
rect -11995 16285 -11965 16315
rect -11915 16285 -11885 16315
rect -11835 16285 -11805 16315
rect -11755 16285 -11725 16315
rect -11675 16285 -11645 16315
rect -11595 16285 -11565 16315
rect -11515 16285 -11485 16315
rect -11435 16285 -11405 16315
rect -11355 16285 -11325 16315
rect -11275 16285 -11245 16315
rect -11195 16285 -11165 16315
rect -11115 16285 -11085 16315
rect -11035 16285 -11005 16315
rect -10955 16285 -10925 16315
rect -10875 16285 -10845 16315
rect -10795 16285 -10765 16315
rect -10715 16285 -10685 16315
rect -10635 16285 -10605 16315
rect -10555 16285 -10525 16315
rect -10475 16285 -10445 16315
rect -10395 16285 -10365 16315
rect -10315 16285 -10285 16315
rect -10235 16285 -10205 16315
rect -10155 16285 -10125 16315
rect -10075 16285 -10045 16315
rect -9995 16285 -9965 16315
rect -9915 16285 -9885 16315
rect -9835 16285 -9805 16315
rect -9755 16285 -9725 16315
rect -9675 16285 -9645 16315
rect -9595 16285 -9565 16315
rect -9515 16285 -9485 16315
rect -9435 16285 -9405 16315
rect -9355 16285 -9325 16315
rect -9275 16285 -9245 16315
rect -9195 16285 -9165 16315
rect -9115 16285 -9085 16315
rect -9035 16285 -9005 16315
rect -8955 16285 -8925 16315
rect -8875 16285 -8845 16315
rect -8795 16285 -8765 16315
rect -8715 16285 -8685 16315
rect -8635 16285 -8605 16315
rect -8555 16285 -8525 16315
rect -8475 16285 -8445 16315
rect -8395 16285 -8365 16315
rect -8315 16285 -8285 16315
rect -8235 16285 -8205 16315
rect -8155 16285 -8125 16315
rect -8075 16285 -8045 16315
rect -7995 16285 -7965 16315
rect -7915 16285 -7885 16315
rect -7835 16285 -7805 16315
rect -7755 16285 -7725 16315
rect -7675 16285 -7645 16315
rect -7595 16285 -7565 16315
rect -7515 16285 -7485 16315
rect -7435 16285 -7405 16315
rect -7355 16285 -7325 16315
rect -7275 16285 -7245 16315
rect -7195 16285 -7165 16315
rect -7115 16285 -7085 16315
rect -7035 16285 -7005 16315
rect -6955 16285 -6925 16315
rect -6875 16285 -6845 16315
rect -6795 16285 -6765 16315
rect -6715 16285 -6685 16315
rect -6635 16285 -6605 16315
rect -6555 16285 -6525 16315
rect -6475 16285 -6445 16315
rect -6395 16285 -6365 16315
rect -6315 16285 -6285 16315
rect -6235 16285 -6205 16315
rect -6155 16285 -6125 16315
rect -6075 16285 -6045 16315
rect -5995 16285 -5965 16315
rect -5915 16285 -5885 16315
rect -5835 16285 -5805 16315
rect -5755 16285 -5725 16315
rect -5595 16285 -5565 16315
rect -5435 16285 -5405 16315
rect -5355 16285 -5325 16315
rect -5275 16285 -5245 16315
rect -5195 16285 -5165 16315
rect -5115 16285 -5085 16315
rect -5035 16285 -5005 16315
rect -4955 16285 -4925 16315
rect -4875 16285 -4845 16315
rect -4795 16285 -4765 16315
rect -4715 16285 -4685 16315
rect -4635 16285 -4605 16315
rect -4555 16285 -4525 16315
rect -4475 16285 -4445 16315
rect -4395 16285 -4365 16315
rect -4315 16285 -4285 16315
rect -4235 16285 -4205 16315
rect -4155 16285 -4125 16315
rect -4075 16285 -4045 16315
rect -3995 16285 -3965 16315
rect -3915 16285 -3885 16315
rect -3835 16285 -3805 16315
rect -3755 16285 -3725 16315
rect -3675 16285 -3645 16315
rect -3595 16285 -3565 16315
rect -3515 16285 -3485 16315
rect -3435 16285 -3405 16315
rect -3355 16285 -3325 16315
rect -3275 16285 -3245 16315
rect -3195 16285 -3165 16315
rect -3115 16285 -3085 16315
rect -3035 16285 -3005 16315
rect -2955 16285 -2925 16315
rect -2875 16285 -2845 16315
rect -2795 16285 -2765 16315
rect -2715 16285 -2685 16315
rect -2635 16285 -2605 16315
rect -2555 16285 -2525 16315
rect -2475 16285 -2445 16315
rect -2395 16285 -2365 16315
rect -2315 16285 -2285 16315
rect -2235 16285 -2205 16315
rect -2155 16285 -2125 16315
rect -2075 16285 -2045 16315
rect -1995 16285 -1965 16315
rect -1835 16285 -1805 16315
rect -1755 16285 -1725 16315
rect -1675 16285 -1645 16315
rect -1595 16285 -1565 16315
rect -1515 16285 -1485 16315
rect -1435 16285 -1405 16315
rect -1355 16285 -1325 16315
rect -1195 16285 -1165 16315
rect -1035 16285 -1005 16315
rect -875 16285 -845 16315
rect -715 16285 -685 16315
rect -555 16285 -525 16315
rect -15515 16205 -15485 16235
rect -15355 16205 -15325 16235
rect -15115 16205 -15085 16235
rect -5675 16205 -5645 16235
rect -1275 16205 -1245 16235
rect -15515 16125 -15485 16155
rect -15355 16125 -15325 16155
rect -15195 16125 -15165 16155
rect -15035 16125 -15005 16155
rect -14955 16125 -14925 16155
rect -14875 16125 -14845 16155
rect -14795 16125 -14765 16155
rect -14715 16125 -14685 16155
rect -14635 16125 -14605 16155
rect -14555 16125 -14525 16155
rect -14475 16125 -14445 16155
rect -14395 16125 -14365 16155
rect -14315 16125 -14285 16155
rect -14235 16125 -14205 16155
rect -14155 16125 -14125 16155
rect -14075 16125 -14045 16155
rect -13995 16125 -13965 16155
rect -13915 16125 -13885 16155
rect -13835 16125 -13805 16155
rect -13755 16125 -13725 16155
rect -13675 16125 -13645 16155
rect -13595 16125 -13565 16155
rect -13515 16125 -13485 16155
rect -13435 16125 -13405 16155
rect -13355 16125 -13325 16155
rect -13275 16125 -13245 16155
rect -13195 16125 -13165 16155
rect -13115 16125 -13085 16155
rect -13035 16125 -13005 16155
rect -12955 16125 -12925 16155
rect -12875 16125 -12845 16155
rect -12795 16125 -12765 16155
rect -12715 16125 -12685 16155
rect -12635 16125 -12605 16155
rect -12555 16125 -12525 16155
rect -12475 16125 -12445 16155
rect -12395 16125 -12365 16155
rect -12315 16125 -12285 16155
rect -12235 16125 -12205 16155
rect -12155 16125 -12125 16155
rect -12075 16125 -12045 16155
rect -11995 16125 -11965 16155
rect -11915 16125 -11885 16155
rect -11835 16125 -11805 16155
rect -11755 16125 -11725 16155
rect -11675 16125 -11645 16155
rect -11595 16125 -11565 16155
rect -11515 16125 -11485 16155
rect -11435 16125 -11405 16155
rect -11355 16125 -11325 16155
rect -11275 16125 -11245 16155
rect -11195 16125 -11165 16155
rect -11115 16125 -11085 16155
rect -11035 16125 -11005 16155
rect -10955 16125 -10925 16155
rect -10875 16125 -10845 16155
rect -10795 16125 -10765 16155
rect -10715 16125 -10685 16155
rect -10635 16125 -10605 16155
rect -10555 16125 -10525 16155
rect -10475 16125 -10445 16155
rect -10395 16125 -10365 16155
rect -10315 16125 -10285 16155
rect -10235 16125 -10205 16155
rect -10155 16125 -10125 16155
rect -10075 16125 -10045 16155
rect -9995 16125 -9965 16155
rect -9915 16125 -9885 16155
rect -9835 16125 -9805 16155
rect -9755 16125 -9725 16155
rect -9675 16125 -9645 16155
rect -9595 16125 -9565 16155
rect -9515 16125 -9485 16155
rect -9435 16125 -9405 16155
rect -9355 16125 -9325 16155
rect -9275 16125 -9245 16155
rect -9195 16125 -9165 16155
rect -9115 16125 -9085 16155
rect -9035 16125 -9005 16155
rect -8955 16125 -8925 16155
rect -8875 16125 -8845 16155
rect -8795 16125 -8765 16155
rect -8715 16125 -8685 16155
rect -8635 16125 -8605 16155
rect -8555 16125 -8525 16155
rect -8475 16125 -8445 16155
rect -8395 16125 -8365 16155
rect -8315 16125 -8285 16155
rect -8235 16125 -8205 16155
rect -8155 16125 -8125 16155
rect -8075 16125 -8045 16155
rect -7995 16125 -7965 16155
rect -7915 16125 -7885 16155
rect -7835 16125 -7805 16155
rect -7755 16125 -7725 16155
rect -7675 16125 -7645 16155
rect -7595 16125 -7565 16155
rect -7515 16125 -7485 16155
rect -7435 16125 -7405 16155
rect -7355 16125 -7325 16155
rect -7275 16125 -7245 16155
rect -7195 16125 -7165 16155
rect -7115 16125 -7085 16155
rect -7035 16125 -7005 16155
rect -6955 16125 -6925 16155
rect -6875 16125 -6845 16155
rect -6795 16125 -6765 16155
rect -6715 16125 -6685 16155
rect -6635 16125 -6605 16155
rect -6555 16125 -6525 16155
rect -6475 16125 -6445 16155
rect -6395 16125 -6365 16155
rect -6315 16125 -6285 16155
rect -6235 16125 -6205 16155
rect -6155 16125 -6125 16155
rect -6075 16125 -6045 16155
rect -5995 16125 -5965 16155
rect -5915 16125 -5885 16155
rect -5835 16125 -5805 16155
rect -5755 16125 -5725 16155
rect -5675 16125 -5645 16155
rect -5595 16125 -5565 16155
rect -5435 16125 -5405 16155
rect -5355 16125 -5325 16155
rect -5275 16125 -5245 16155
rect -5195 16125 -5165 16155
rect -5115 16125 -5085 16155
rect -5035 16125 -5005 16155
rect -4955 16125 -4925 16155
rect -4875 16125 -4845 16155
rect -4795 16125 -4765 16155
rect -4715 16125 -4685 16155
rect -4635 16125 -4605 16155
rect -4555 16125 -4525 16155
rect -4475 16125 -4445 16155
rect -4395 16125 -4365 16155
rect -4315 16125 -4285 16155
rect -4235 16125 -4205 16155
rect -4155 16125 -4125 16155
rect -4075 16125 -4045 16155
rect -3995 16125 -3965 16155
rect -3915 16125 -3885 16155
rect -3835 16125 -3805 16155
rect -3755 16125 -3725 16155
rect -3675 16125 -3645 16155
rect -3595 16125 -3565 16155
rect -3515 16125 -3485 16155
rect -3435 16125 -3405 16155
rect -3355 16125 -3325 16155
rect -3275 16125 -3245 16155
rect -3195 16125 -3165 16155
rect -3115 16125 -3085 16155
rect -3035 16125 -3005 16155
rect -2955 16125 -2925 16155
rect -2875 16125 -2845 16155
rect -2795 16125 -2765 16155
rect -2715 16125 -2685 16155
rect -2635 16125 -2605 16155
rect -2555 16125 -2525 16155
rect -2475 16125 -2445 16155
rect -2395 16125 -2365 16155
rect -2315 16125 -2285 16155
rect -2235 16125 -2205 16155
rect -2155 16125 -2125 16155
rect -2075 16125 -2045 16155
rect -1995 16125 -1965 16155
rect -1835 16125 -1805 16155
rect -1755 16125 -1725 16155
rect -1675 16125 -1645 16155
rect -1595 16125 -1565 16155
rect -1515 16125 -1485 16155
rect -1435 16125 -1405 16155
rect -1355 16125 -1325 16155
rect -1195 16125 -1165 16155
rect -1035 16125 -1005 16155
rect -875 16125 -845 16155
rect -715 16125 -685 16155
rect -555 16125 -525 16155
rect -15515 16045 -15485 16075
rect -15355 16045 -15325 16075
rect -15275 16045 -15245 16075
rect -5515 16045 -5485 16075
rect -1115 16045 -1085 16075
rect -15515 15965 -15485 15995
rect -15355 15965 -15325 15995
rect -15195 15965 -15165 15995
rect -15035 15965 -15005 15995
rect -14955 15965 -14925 15995
rect -14875 15965 -14845 15995
rect -14795 15965 -14765 15995
rect -14715 15965 -14685 15995
rect -14635 15965 -14605 15995
rect -14555 15965 -14525 15995
rect -14475 15965 -14445 15995
rect -14395 15965 -14365 15995
rect -14315 15965 -14285 15995
rect -14235 15965 -14205 15995
rect -14155 15965 -14125 15995
rect -14075 15965 -14045 15995
rect -13995 15965 -13965 15995
rect -13915 15965 -13885 15995
rect -13835 15965 -13805 15995
rect -13755 15965 -13725 15995
rect -13675 15965 -13645 15995
rect -13595 15965 -13565 15995
rect -13515 15965 -13485 15995
rect -13435 15965 -13405 15995
rect -13355 15965 -13325 15995
rect -13275 15965 -13245 15995
rect -13195 15965 -13165 15995
rect -13115 15965 -13085 15995
rect -13035 15965 -13005 15995
rect -12955 15965 -12925 15995
rect -12875 15965 -12845 15995
rect -12795 15965 -12765 15995
rect -12715 15965 -12685 15995
rect -12635 15965 -12605 15995
rect -12555 15965 -12525 15995
rect -12475 15965 -12445 15995
rect -12395 15965 -12365 15995
rect -12315 15965 -12285 15995
rect -12235 15965 -12205 15995
rect -12155 15965 -12125 15995
rect -12075 15965 -12045 15995
rect -11995 15965 -11965 15995
rect -11915 15965 -11885 15995
rect -11835 15965 -11805 15995
rect -11755 15965 -11725 15995
rect -11675 15965 -11645 15995
rect -11595 15965 -11565 15995
rect -11515 15965 -11485 15995
rect -11435 15965 -11405 15995
rect -11355 15965 -11325 15995
rect -11275 15965 -11245 15995
rect -11195 15965 -11165 15995
rect -11115 15965 -11085 15995
rect -11035 15965 -11005 15995
rect -10955 15965 -10925 15995
rect -10875 15965 -10845 15995
rect -10795 15965 -10765 15995
rect -10715 15965 -10685 15995
rect -10635 15965 -10605 15995
rect -10555 15965 -10525 15995
rect -10475 15965 -10445 15995
rect -10395 15965 -10365 15995
rect -10315 15965 -10285 15995
rect -10235 15965 -10205 15995
rect -10155 15965 -10125 15995
rect -10075 15965 -10045 15995
rect -9995 15965 -9965 15995
rect -9915 15965 -9885 15995
rect -9835 15965 -9805 15995
rect -9755 15965 -9725 15995
rect -9675 15965 -9645 15995
rect -9595 15965 -9565 15995
rect -9515 15965 -9485 15995
rect -9435 15965 -9405 15995
rect -9355 15965 -9325 15995
rect -9275 15965 -9245 15995
rect -9195 15965 -9165 15995
rect -9115 15965 -9085 15995
rect -9035 15965 -9005 15995
rect -8955 15965 -8925 15995
rect -8875 15965 -8845 15995
rect -8795 15965 -8765 15995
rect -8715 15965 -8685 15995
rect -8635 15965 -8605 15995
rect -8555 15965 -8525 15995
rect -8475 15965 -8445 15995
rect -8395 15965 -8365 15995
rect -8315 15965 -8285 15995
rect -8235 15965 -8205 15995
rect -8155 15965 -8125 15995
rect -8075 15965 -8045 15995
rect -7995 15965 -7965 15995
rect -7915 15965 -7885 15995
rect -7835 15965 -7805 15995
rect -7755 15965 -7725 15995
rect -7675 15965 -7645 15995
rect -7595 15965 -7565 15995
rect -7515 15965 -7485 15995
rect -7435 15965 -7405 15995
rect -7355 15965 -7325 15995
rect -7275 15965 -7245 15995
rect -7195 15965 -7165 15995
rect -7115 15965 -7085 15995
rect -7035 15965 -7005 15995
rect -6955 15965 -6925 15995
rect -6875 15965 -6845 15995
rect -6795 15965 -6765 15995
rect -6715 15965 -6685 15995
rect -6635 15965 -6605 15995
rect -6555 15965 -6525 15995
rect -6475 15965 -6445 15995
rect -6395 15965 -6365 15995
rect -6315 15965 -6285 15995
rect -6235 15965 -6205 15995
rect -6155 15965 -6125 15995
rect -6075 15965 -6045 15995
rect -5995 15965 -5965 15995
rect -5915 15965 -5885 15995
rect -5835 15965 -5805 15995
rect -5755 15965 -5725 15995
rect -5675 15965 -5645 15995
rect -5595 15965 -5565 15995
rect -5435 15965 -5405 15995
rect -5355 15965 -5325 15995
rect -5275 15965 -5245 15995
rect -5195 15965 -5165 15995
rect -5115 15965 -5085 15995
rect -5035 15965 -5005 15995
rect -4955 15965 -4925 15995
rect -4875 15965 -4845 15995
rect -4795 15965 -4765 15995
rect -4715 15965 -4685 15995
rect -4635 15965 -4605 15995
rect -4555 15965 -4525 15995
rect -4475 15965 -4445 15995
rect -4395 15965 -4365 15995
rect -4315 15965 -4285 15995
rect -4235 15965 -4205 15995
rect -4155 15965 -4125 15995
rect -4075 15965 -4045 15995
rect -3995 15965 -3965 15995
rect -3915 15965 -3885 15995
rect -3835 15965 -3805 15995
rect -3755 15965 -3725 15995
rect -3675 15965 -3645 15995
rect -3595 15965 -3565 15995
rect -3515 15965 -3485 15995
rect -3435 15965 -3405 15995
rect -3355 15965 -3325 15995
rect -3275 15965 -3245 15995
rect -3195 15965 -3165 15995
rect -3115 15965 -3085 15995
rect -3035 15965 -3005 15995
rect -2955 15965 -2925 15995
rect -2875 15965 -2845 15995
rect -2795 15965 -2765 15995
rect -2715 15965 -2685 15995
rect -2635 15965 -2605 15995
rect -2555 15965 -2525 15995
rect -2475 15965 -2445 15995
rect -2395 15965 -2365 15995
rect -2315 15965 -2285 15995
rect -2235 15965 -2205 15995
rect -2155 15965 -2125 15995
rect -2075 15965 -2045 15995
rect -1995 15965 -1965 15995
rect -1835 15965 -1805 15995
rect -1755 15965 -1725 15995
rect -1675 15965 -1645 15995
rect -1595 15965 -1565 15995
rect -1515 15965 -1485 15995
rect -1435 15965 -1405 15995
rect -1355 15965 -1325 15995
rect -1195 15965 -1165 15995
rect -1035 15965 -1005 15995
rect -875 15965 -845 15995
rect -715 15965 -685 15995
rect -555 15965 -525 15995
<< metal3 >>
rect 15880 37560 16880 37640
rect -15520 21435 -15480 21480
rect -15520 21405 -15515 21435
rect -15485 21405 -15480 21435
rect -15520 21355 -15480 21405
rect -15520 21325 -15515 21355
rect -15485 21325 -15480 21355
rect -15520 21275 -15480 21325
rect -15520 21245 -15515 21275
rect -15485 21245 -15480 21275
rect -15520 21195 -15480 21245
rect -15520 21165 -15515 21195
rect -15485 21165 -15480 21195
rect -15520 21115 -15480 21165
rect -15520 21085 -15515 21115
rect -15485 21085 -15480 21115
rect -15520 21035 -15480 21085
rect -15520 21005 -15515 21035
rect -15485 21005 -15480 21035
rect -15520 20955 -15480 21005
rect -15520 20925 -15515 20955
rect -15485 20925 -15480 20955
rect -15520 20876 -15480 20925
rect -15520 20844 -15516 20876
rect -15484 20844 -15480 20876
rect -15520 20796 -15480 20844
rect -15520 20764 -15516 20796
rect -15484 20764 -15480 20796
rect -16560 20675 -16520 20680
rect -16560 20645 -16555 20675
rect -16525 20645 -16520 20675
rect -16560 20515 -16520 20645
rect -16560 20485 -16555 20515
rect -16525 20485 -16520 20515
rect -16560 20480 -16520 20485
rect -16480 20675 -16440 20680
rect -16480 20645 -16475 20675
rect -16445 20645 -16440 20675
rect -16480 20515 -16440 20645
rect -16480 20485 -16475 20515
rect -16445 20485 -16440 20515
rect -16480 20480 -16440 20485
rect -16400 20675 -16360 20680
rect -16400 20645 -16395 20675
rect -16365 20645 -16360 20675
rect -16400 20515 -16360 20645
rect -16400 20485 -16395 20515
rect -16365 20485 -16360 20515
rect -16400 20480 -16360 20485
rect -16320 20675 -16280 20680
rect -16320 20645 -16315 20675
rect -16285 20645 -16280 20675
rect -16320 20515 -16280 20645
rect -16320 20485 -16315 20515
rect -16285 20485 -16280 20515
rect -16320 20480 -16280 20485
rect -16240 20675 -16200 20680
rect -16240 20645 -16235 20675
rect -16205 20645 -16200 20675
rect -16240 20515 -16200 20645
rect -16240 20485 -16235 20515
rect -16205 20485 -16200 20515
rect -16240 20480 -16200 20485
rect -16160 20675 -16120 20680
rect -16160 20645 -16155 20675
rect -16125 20645 -16120 20675
rect -16160 20515 -16120 20645
rect -16160 20485 -16155 20515
rect -16125 20485 -16120 20515
rect -16160 20480 -16120 20485
rect -16080 20675 -16040 20680
rect -16080 20645 -16075 20675
rect -16045 20645 -16040 20675
rect -16080 20515 -16040 20645
rect -16080 20485 -16075 20515
rect -16045 20485 -16040 20515
rect -16080 20480 -16040 20485
rect -16000 20675 -15960 20680
rect -16000 20645 -15995 20675
rect -15965 20645 -15960 20675
rect -16000 20515 -15960 20645
rect -16000 20485 -15995 20515
rect -15965 20485 -15960 20515
rect -16000 20480 -15960 20485
rect -15920 20675 -15880 20680
rect -15920 20645 -15915 20675
rect -15885 20645 -15880 20675
rect -15920 20515 -15880 20645
rect -15920 20485 -15915 20515
rect -15885 20485 -15880 20515
rect -15920 20480 -15880 20485
rect -15840 20675 -15800 20680
rect -15840 20645 -15835 20675
rect -15805 20645 -15800 20675
rect -15840 20515 -15800 20645
rect -15840 20485 -15835 20515
rect -15805 20485 -15800 20515
rect -15840 20480 -15800 20485
rect -15760 20675 -15720 20680
rect -15760 20645 -15755 20675
rect -15725 20645 -15720 20675
rect -15760 20515 -15720 20645
rect -15760 20485 -15755 20515
rect -15725 20485 -15720 20515
rect -15760 20480 -15720 20485
rect -15680 20675 -15640 20680
rect -15680 20645 -15675 20675
rect -15645 20645 -15640 20675
rect -15680 20515 -15640 20645
rect -15680 20485 -15675 20515
rect -15645 20485 -15640 20515
rect -15680 20480 -15640 20485
rect -15600 20675 -15560 20680
rect -15600 20645 -15595 20675
rect -15565 20645 -15560 20675
rect -15600 20515 -15560 20645
rect -15600 20485 -15595 20515
rect -15565 20485 -15560 20515
rect -15600 20480 -15560 20485
rect -15520 20396 -15480 20764
rect -15520 20364 -15516 20396
rect -15484 20364 -15480 20396
rect -15520 20316 -15480 20364
rect -15520 20284 -15516 20316
rect -15484 20284 -15480 20316
rect -15520 20236 -15480 20284
rect -15520 20204 -15516 20236
rect -15484 20204 -15480 20236
rect -15520 20156 -15480 20204
rect -15520 20124 -15516 20156
rect -15484 20124 -15480 20156
rect -15520 20076 -15480 20124
rect -15520 20044 -15516 20076
rect -15484 20044 -15480 20076
rect -15520 19996 -15480 20044
rect -15520 19964 -15516 19996
rect -15484 19964 -15480 19996
rect -15520 19916 -15480 19964
rect -15520 19884 -15516 19916
rect -15484 19884 -15480 19916
rect -15520 19836 -15480 19884
rect -15520 19804 -15516 19836
rect -15484 19804 -15480 19836
rect -15520 19756 -15480 19804
rect -15520 19724 -15516 19756
rect -15484 19724 -15480 19756
rect -15520 19676 -15480 19724
rect -15520 19644 -15516 19676
rect -15484 19644 -15480 19676
rect -15520 19596 -15480 19644
rect -15520 19564 -15516 19596
rect -15484 19564 -15480 19596
rect -15520 19516 -15480 19564
rect -15520 19484 -15516 19516
rect -15484 19484 -15480 19516
rect -15520 19436 -15480 19484
rect -15520 19404 -15516 19436
rect -15484 19404 -15480 19436
rect -15520 19356 -15480 19404
rect -15520 19324 -15516 19356
rect -15484 19324 -15480 19356
rect -15520 19276 -15480 19324
rect -15520 19244 -15516 19276
rect -15484 19244 -15480 19276
rect -15520 19196 -15480 19244
rect -15520 19164 -15516 19196
rect -15484 19164 -15480 19196
rect -15520 19116 -15480 19164
rect -15520 19084 -15516 19116
rect -15484 19084 -15480 19116
rect -15520 19036 -15480 19084
rect -15520 19004 -15516 19036
rect -15484 19004 -15480 19036
rect -15520 18956 -15480 19004
rect -15520 18924 -15516 18956
rect -15484 18924 -15480 18956
rect -16560 18875 -16520 18880
rect -16560 18845 -16555 18875
rect -16525 18845 -16520 18875
rect -16560 18715 -16520 18845
rect -16560 18685 -16555 18715
rect -16525 18685 -16520 18715
rect -16560 18555 -16520 18685
rect -16560 18525 -16555 18555
rect -16525 18525 -16520 18555
rect -16560 18520 -16520 18525
rect -16480 18875 -16440 18880
rect -16480 18845 -16475 18875
rect -16445 18845 -16440 18875
rect -16480 18715 -16440 18845
rect -16480 18685 -16475 18715
rect -16445 18685 -16440 18715
rect -16480 18555 -16440 18685
rect -16480 18525 -16475 18555
rect -16445 18525 -16440 18555
rect -16480 18520 -16440 18525
rect -16400 18875 -16360 18880
rect -16400 18845 -16395 18875
rect -16365 18845 -16360 18875
rect -16400 18715 -16360 18845
rect -16400 18685 -16395 18715
rect -16365 18685 -16360 18715
rect -16400 18555 -16360 18685
rect -16400 18525 -16395 18555
rect -16365 18525 -16360 18555
rect -16400 18520 -16360 18525
rect -16320 18875 -16280 18880
rect -16320 18845 -16315 18875
rect -16285 18845 -16280 18875
rect -16320 18715 -16280 18845
rect -16320 18685 -16315 18715
rect -16285 18685 -16280 18715
rect -16320 18555 -16280 18685
rect -16320 18525 -16315 18555
rect -16285 18525 -16280 18555
rect -16320 18520 -16280 18525
rect -16240 18875 -16200 18880
rect -16240 18845 -16235 18875
rect -16205 18845 -16200 18875
rect -16240 18715 -16200 18845
rect -16240 18685 -16235 18715
rect -16205 18685 -16200 18715
rect -16240 18555 -16200 18685
rect -16240 18525 -16235 18555
rect -16205 18525 -16200 18555
rect -16240 18520 -16200 18525
rect -16160 18875 -16120 18880
rect -16160 18845 -16155 18875
rect -16125 18845 -16120 18875
rect -16160 18715 -16120 18845
rect -16160 18685 -16155 18715
rect -16125 18685 -16120 18715
rect -16160 18555 -16120 18685
rect -16160 18525 -16155 18555
rect -16125 18525 -16120 18555
rect -16160 18520 -16120 18525
rect -16080 18875 -16040 18880
rect -16080 18845 -16075 18875
rect -16045 18845 -16040 18875
rect -16080 18715 -16040 18845
rect -16080 18685 -16075 18715
rect -16045 18685 -16040 18715
rect -16080 18555 -16040 18685
rect -16080 18525 -16075 18555
rect -16045 18525 -16040 18555
rect -16080 18520 -16040 18525
rect -16000 18875 -15960 18880
rect -16000 18845 -15995 18875
rect -15965 18845 -15960 18875
rect -16000 18715 -15960 18845
rect -16000 18685 -15995 18715
rect -15965 18685 -15960 18715
rect -16000 18555 -15960 18685
rect -16000 18525 -15995 18555
rect -15965 18525 -15960 18555
rect -16000 18520 -15960 18525
rect -15920 18875 -15880 18880
rect -15920 18845 -15915 18875
rect -15885 18845 -15880 18875
rect -15920 18715 -15880 18845
rect -15920 18685 -15915 18715
rect -15885 18685 -15880 18715
rect -15920 18555 -15880 18685
rect -15920 18525 -15915 18555
rect -15885 18525 -15880 18555
rect -15920 18520 -15880 18525
rect -15840 18875 -15800 18880
rect -15840 18845 -15835 18875
rect -15805 18845 -15800 18875
rect -15840 18715 -15800 18845
rect -15840 18685 -15835 18715
rect -15805 18685 -15800 18715
rect -15840 18555 -15800 18685
rect -15840 18525 -15835 18555
rect -15805 18525 -15800 18555
rect -15840 18520 -15800 18525
rect -15760 18875 -15720 18880
rect -15760 18845 -15755 18875
rect -15725 18845 -15720 18875
rect -15760 18715 -15720 18845
rect -15760 18685 -15755 18715
rect -15725 18685 -15720 18715
rect -15760 18555 -15720 18685
rect -15760 18525 -15755 18555
rect -15725 18525 -15720 18555
rect -15760 18520 -15720 18525
rect -15680 18875 -15640 18880
rect -15680 18845 -15675 18875
rect -15645 18845 -15640 18875
rect -15680 18715 -15640 18845
rect -15680 18685 -15675 18715
rect -15645 18685 -15640 18715
rect -15680 18555 -15640 18685
rect -15680 18525 -15675 18555
rect -15645 18525 -15640 18555
rect -15680 18520 -15640 18525
rect -15600 18875 -15560 18880
rect -15600 18845 -15595 18875
rect -15565 18845 -15560 18875
rect -15600 18715 -15560 18845
rect -15600 18685 -15595 18715
rect -15565 18685 -15560 18715
rect -15600 18555 -15560 18685
rect -15600 18525 -15595 18555
rect -15565 18525 -15560 18555
rect -15600 18520 -15560 18525
rect -15520 18876 -15480 18924
rect -15520 18844 -15516 18876
rect -15484 18844 -15480 18876
rect -15520 18715 -15480 18844
rect -15440 18795 -15400 21480
rect -15440 18765 -15435 18795
rect -15405 18765 -15400 18795
rect -15440 18760 -15400 18765
rect -15360 21435 -15320 21480
rect -15360 21405 -15355 21435
rect -15325 21405 -15320 21435
rect -15360 21355 -15320 21405
rect -15360 21325 -15355 21355
rect -15325 21325 -15320 21355
rect -15360 21275 -15320 21325
rect -15360 21245 -15355 21275
rect -15325 21245 -15320 21275
rect -15360 21195 -15320 21245
rect -15360 21165 -15355 21195
rect -15325 21165 -15320 21195
rect -15360 21115 -15320 21165
rect -15280 21195 -15240 21480
rect -15280 21165 -15275 21195
rect -15245 21165 -15240 21195
rect -15280 21160 -15240 21165
rect -15200 21435 -15160 21480
rect -15200 21405 -15195 21435
rect -15165 21405 -15160 21435
rect -15200 21355 -15160 21405
rect -15200 21325 -15195 21355
rect -15165 21325 -15160 21355
rect -15200 21275 -15160 21325
rect -15120 21355 -15080 21480
rect -15120 21325 -15115 21355
rect -15085 21325 -15080 21355
rect -15120 21320 -15080 21325
rect -15040 21435 -15000 21480
rect -15040 21405 -15035 21435
rect -15005 21405 -15000 21435
rect -15200 21245 -15195 21275
rect -15165 21245 -15160 21275
rect -15360 21085 -15355 21115
rect -15325 21085 -15320 21115
rect -15360 21035 -15320 21085
rect -15360 21005 -15355 21035
rect -15325 21005 -15320 21035
rect -15360 20955 -15320 21005
rect -15360 20925 -15355 20955
rect -15325 20925 -15320 20955
rect -15360 20876 -15320 20925
rect -15360 20844 -15356 20876
rect -15324 20844 -15320 20876
rect -15360 20796 -15320 20844
rect -15360 20764 -15356 20796
rect -15324 20764 -15320 20796
rect -15360 20396 -15320 20764
rect -15360 20364 -15356 20396
rect -15324 20364 -15320 20396
rect -15360 20316 -15320 20364
rect -15360 20284 -15356 20316
rect -15324 20284 -15320 20316
rect -15360 20236 -15320 20284
rect -15360 20204 -15356 20236
rect -15324 20204 -15320 20236
rect -15360 20156 -15320 20204
rect -15360 20124 -15356 20156
rect -15324 20124 -15320 20156
rect -15360 20076 -15320 20124
rect -15360 20044 -15356 20076
rect -15324 20044 -15320 20076
rect -15360 19996 -15320 20044
rect -15360 19964 -15356 19996
rect -15324 19964 -15320 19996
rect -15360 19916 -15320 19964
rect -15360 19884 -15356 19916
rect -15324 19884 -15320 19916
rect -15360 19836 -15320 19884
rect -15360 19804 -15356 19836
rect -15324 19804 -15320 19836
rect -15360 19756 -15320 19804
rect -15360 19724 -15356 19756
rect -15324 19724 -15320 19756
rect -15360 19676 -15320 19724
rect -15360 19644 -15356 19676
rect -15324 19644 -15320 19676
rect -15360 19596 -15320 19644
rect -15360 19564 -15356 19596
rect -15324 19564 -15320 19596
rect -15360 19516 -15320 19564
rect -15360 19484 -15356 19516
rect -15324 19484 -15320 19516
rect -15360 19436 -15320 19484
rect -15360 19404 -15356 19436
rect -15324 19404 -15320 19436
rect -15360 19356 -15320 19404
rect -15360 19324 -15356 19356
rect -15324 19324 -15320 19356
rect -15360 19276 -15320 19324
rect -15360 19244 -15356 19276
rect -15324 19244 -15320 19276
rect -15360 19196 -15320 19244
rect -15360 19164 -15356 19196
rect -15324 19164 -15320 19196
rect -15360 19116 -15320 19164
rect -15360 19084 -15356 19116
rect -15324 19084 -15320 19116
rect -15360 19036 -15320 19084
rect -15360 19004 -15356 19036
rect -15324 19004 -15320 19036
rect -15360 18956 -15320 19004
rect -15360 18924 -15356 18956
rect -15324 18924 -15320 18956
rect -15360 18876 -15320 18924
rect -15360 18844 -15356 18876
rect -15324 18844 -15320 18876
rect -15520 18685 -15515 18715
rect -15485 18685 -15480 18715
rect -15520 18556 -15480 18685
rect -15360 18715 -15320 18844
rect -15200 21115 -15160 21245
rect -15200 21085 -15195 21115
rect -15165 21085 -15160 21115
rect -15200 21035 -15160 21085
rect -15040 21275 -15000 21405
rect -15040 21245 -15035 21275
rect -15005 21245 -15000 21275
rect -15040 21115 -15000 21245
rect -15040 21085 -15035 21115
rect -15005 21085 -15000 21115
rect -15200 21005 -15195 21035
rect -15165 21005 -15160 21035
rect -15200 20955 -15160 21005
rect -15200 20925 -15195 20955
rect -15165 20925 -15160 20955
rect -15200 20876 -15160 20925
rect -15200 20844 -15196 20876
rect -15164 20844 -15160 20876
rect -15200 20796 -15160 20844
rect -15200 20764 -15196 20796
rect -15164 20764 -15160 20796
rect -15200 20396 -15160 20764
rect -15200 20364 -15196 20396
rect -15164 20364 -15160 20396
rect -15200 20316 -15160 20364
rect -15200 20284 -15196 20316
rect -15164 20284 -15160 20316
rect -15200 20236 -15160 20284
rect -15200 20204 -15196 20236
rect -15164 20204 -15160 20236
rect -15200 20156 -15160 20204
rect -15200 20124 -15196 20156
rect -15164 20124 -15160 20156
rect -15200 20076 -15160 20124
rect -15200 20044 -15196 20076
rect -15164 20044 -15160 20076
rect -15200 19996 -15160 20044
rect -15200 19964 -15196 19996
rect -15164 19964 -15160 19996
rect -15200 19916 -15160 19964
rect -15200 19884 -15196 19916
rect -15164 19884 -15160 19916
rect -15200 19836 -15160 19884
rect -15200 19804 -15196 19836
rect -15164 19804 -15160 19836
rect -15200 19756 -15160 19804
rect -15200 19724 -15196 19756
rect -15164 19724 -15160 19756
rect -15200 19676 -15160 19724
rect -15200 19644 -15196 19676
rect -15164 19644 -15160 19676
rect -15200 19596 -15160 19644
rect -15200 19564 -15196 19596
rect -15164 19564 -15160 19596
rect -15200 19516 -15160 19564
rect -15200 19484 -15196 19516
rect -15164 19484 -15160 19516
rect -15200 19436 -15160 19484
rect -15200 19404 -15196 19436
rect -15164 19404 -15160 19436
rect -15200 19356 -15160 19404
rect -15200 19324 -15196 19356
rect -15164 19324 -15160 19356
rect -15200 19276 -15160 19324
rect -15200 19244 -15196 19276
rect -15164 19244 -15160 19276
rect -15200 19196 -15160 19244
rect -15200 19164 -15196 19196
rect -15164 19164 -15160 19196
rect -15200 19116 -15160 19164
rect -15200 19084 -15196 19116
rect -15164 19084 -15160 19116
rect -15200 19036 -15160 19084
rect -15200 19004 -15196 19036
rect -15164 19004 -15160 19036
rect -15200 18956 -15160 19004
rect -15200 18924 -15196 18956
rect -15164 18924 -15160 18956
rect -15200 18876 -15160 18924
rect -15200 18844 -15196 18876
rect -15164 18844 -15160 18876
rect -15360 18685 -15355 18715
rect -15325 18685 -15320 18715
rect -15520 18524 -15516 18556
rect -15484 18524 -15480 18556
rect -15520 18476 -15480 18524
rect -15520 18444 -15516 18476
rect -15484 18444 -15480 18476
rect -15520 18396 -15480 18444
rect -15520 18364 -15516 18396
rect -15484 18364 -15480 18396
rect -15520 18316 -15480 18364
rect -15520 18284 -15516 18316
rect -15484 18284 -15480 18316
rect -15520 18236 -15480 18284
rect -15520 18204 -15516 18236
rect -15484 18204 -15480 18236
rect -15520 18156 -15480 18204
rect -15520 18124 -15516 18156
rect -15484 18124 -15480 18156
rect -15520 18076 -15480 18124
rect -15520 18044 -15516 18076
rect -15484 18044 -15480 18076
rect -15520 17996 -15480 18044
rect -15520 17964 -15516 17996
rect -15484 17964 -15480 17996
rect -15520 17916 -15480 17964
rect -15520 17884 -15516 17916
rect -15484 17884 -15480 17916
rect -15520 17836 -15480 17884
rect -15520 17804 -15516 17836
rect -15484 17804 -15480 17836
rect -15520 17756 -15480 17804
rect -15520 17724 -15516 17756
rect -15484 17724 -15480 17756
rect -15520 17676 -15480 17724
rect -15520 17644 -15516 17676
rect -15484 17644 -15480 17676
rect -15520 17596 -15480 17644
rect -15520 17564 -15516 17596
rect -15484 17564 -15480 17596
rect -15520 17516 -15480 17564
rect -15520 17484 -15516 17516
rect -15484 17484 -15480 17516
rect -15520 17436 -15480 17484
rect -15520 17404 -15516 17436
rect -15484 17404 -15480 17436
rect -16560 17355 -16520 17360
rect -16560 17325 -16555 17355
rect -16525 17325 -16520 17355
rect -16560 17195 -16520 17325
rect -16560 17165 -16555 17195
rect -16525 17165 -16520 17195
rect -16560 17160 -16520 17165
rect -16480 17355 -16440 17360
rect -16480 17325 -16475 17355
rect -16445 17325 -16440 17355
rect -16480 17195 -16440 17325
rect -16480 17165 -16475 17195
rect -16445 17165 -16440 17195
rect -16480 17160 -16440 17165
rect -16400 17355 -16360 17360
rect -16400 17325 -16395 17355
rect -16365 17325 -16360 17355
rect -16400 17195 -16360 17325
rect -16400 17165 -16395 17195
rect -16365 17165 -16360 17195
rect -16400 17160 -16360 17165
rect -16320 17355 -16280 17360
rect -16320 17325 -16315 17355
rect -16285 17325 -16280 17355
rect -16320 17195 -16280 17325
rect -16320 17165 -16315 17195
rect -16285 17165 -16280 17195
rect -16320 17160 -16280 17165
rect -16240 17355 -16200 17360
rect -16240 17325 -16235 17355
rect -16205 17325 -16200 17355
rect -16240 17195 -16200 17325
rect -16240 17165 -16235 17195
rect -16205 17165 -16200 17195
rect -16240 17160 -16200 17165
rect -16160 17355 -16120 17360
rect -16160 17325 -16155 17355
rect -16125 17325 -16120 17355
rect -16160 17195 -16120 17325
rect -16160 17165 -16155 17195
rect -16125 17165 -16120 17195
rect -16160 17160 -16120 17165
rect -16080 17355 -16040 17360
rect -16080 17325 -16075 17355
rect -16045 17325 -16040 17355
rect -16080 17195 -16040 17325
rect -16080 17165 -16075 17195
rect -16045 17165 -16040 17195
rect -16080 17160 -16040 17165
rect -16000 17355 -15960 17360
rect -16000 17325 -15995 17355
rect -15965 17325 -15960 17355
rect -16000 17195 -15960 17325
rect -16000 17165 -15995 17195
rect -15965 17165 -15960 17195
rect -16000 17160 -15960 17165
rect -15920 17355 -15880 17360
rect -15920 17325 -15915 17355
rect -15885 17325 -15880 17355
rect -15920 17195 -15880 17325
rect -15920 17165 -15915 17195
rect -15885 17165 -15880 17195
rect -15920 17160 -15880 17165
rect -15840 17355 -15800 17360
rect -15840 17325 -15835 17355
rect -15805 17325 -15800 17355
rect -15840 17195 -15800 17325
rect -15840 17165 -15835 17195
rect -15805 17165 -15800 17195
rect -15840 17160 -15800 17165
rect -15760 17355 -15720 17360
rect -15760 17325 -15755 17355
rect -15725 17325 -15720 17355
rect -15760 17195 -15720 17325
rect -15760 17165 -15755 17195
rect -15725 17165 -15720 17195
rect -15760 17160 -15720 17165
rect -15680 17355 -15640 17360
rect -15680 17325 -15675 17355
rect -15645 17325 -15640 17355
rect -15680 17195 -15640 17325
rect -15680 17165 -15675 17195
rect -15645 17165 -15640 17195
rect -15680 17160 -15640 17165
rect -15600 17355 -15560 17360
rect -15600 17325 -15595 17355
rect -15565 17325 -15560 17355
rect -15600 17195 -15560 17325
rect -15600 17165 -15595 17195
rect -15565 17165 -15560 17195
rect -15600 17160 -15560 17165
rect -15520 17355 -15480 17404
rect -15520 17325 -15515 17355
rect -15485 17325 -15480 17355
rect -15520 17195 -15480 17325
rect -15520 17165 -15515 17195
rect -15485 17165 -15480 17195
rect -15520 17116 -15480 17165
rect -15520 17084 -15516 17116
rect -15484 17084 -15480 17116
rect -15520 17036 -15480 17084
rect -15520 17004 -15516 17036
rect -15484 17004 -15480 17036
rect -15520 16956 -15480 17004
rect -15520 16924 -15516 16956
rect -15484 16924 -15480 16956
rect -15520 16876 -15480 16924
rect -15520 16844 -15516 16876
rect -15484 16844 -15480 16876
rect -15520 16796 -15480 16844
rect -15520 16764 -15516 16796
rect -15484 16764 -15480 16796
rect -15520 16716 -15480 16764
rect -15520 16684 -15516 16716
rect -15484 16684 -15480 16716
rect -15520 16636 -15480 16684
rect -15520 16604 -15516 16636
rect -15484 16604 -15480 16636
rect -15520 16556 -15480 16604
rect -15520 16524 -15516 16556
rect -15484 16524 -15480 16556
rect -15520 16476 -15480 16524
rect -15520 16444 -15516 16476
rect -15484 16444 -15480 16476
rect -15520 16395 -15480 16444
rect -15520 16365 -15515 16395
rect -15485 16365 -15480 16395
rect -15520 16315 -15480 16365
rect -15520 16285 -15515 16315
rect -15485 16285 -15480 16315
rect -15520 16235 -15480 16285
rect -15520 16205 -15515 16235
rect -15485 16205 -15480 16235
rect -15520 16155 -15480 16205
rect -15520 16125 -15515 16155
rect -15485 16125 -15480 16155
rect -15520 16075 -15480 16125
rect -15520 16045 -15515 16075
rect -15485 16045 -15480 16075
rect -15520 15995 -15480 16045
rect -15520 15965 -15515 15995
rect -15485 15965 -15480 15995
rect -15520 15920 -15480 15965
rect -15440 18635 -15400 18640
rect -15440 18605 -15435 18635
rect -15405 18605 -15400 18635
rect -15440 15920 -15400 18605
rect -15360 18556 -15320 18685
rect -15360 18524 -15356 18556
rect -15324 18524 -15320 18556
rect -15360 18476 -15320 18524
rect -15360 18444 -15356 18476
rect -15324 18444 -15320 18476
rect -15360 18396 -15320 18444
rect -15360 18364 -15356 18396
rect -15324 18364 -15320 18396
rect -15360 18316 -15320 18364
rect -15360 18284 -15356 18316
rect -15324 18284 -15320 18316
rect -15360 18236 -15320 18284
rect -15360 18204 -15356 18236
rect -15324 18204 -15320 18236
rect -15360 18156 -15320 18204
rect -15360 18124 -15356 18156
rect -15324 18124 -15320 18156
rect -15360 18076 -15320 18124
rect -15360 18044 -15356 18076
rect -15324 18044 -15320 18076
rect -15360 17996 -15320 18044
rect -15360 17964 -15356 17996
rect -15324 17964 -15320 17996
rect -15360 17916 -15320 17964
rect -15360 17884 -15356 17916
rect -15324 17884 -15320 17916
rect -15360 17836 -15320 17884
rect -15360 17804 -15356 17836
rect -15324 17804 -15320 17836
rect -15360 17756 -15320 17804
rect -15360 17724 -15356 17756
rect -15324 17724 -15320 17756
rect -15360 17676 -15320 17724
rect -15360 17644 -15356 17676
rect -15324 17644 -15320 17676
rect -15360 17596 -15320 17644
rect -15360 17564 -15356 17596
rect -15324 17564 -15320 17596
rect -15360 17516 -15320 17564
rect -15360 17484 -15356 17516
rect -15324 17484 -15320 17516
rect -15360 17436 -15320 17484
rect -15360 17404 -15356 17436
rect -15324 17404 -15320 17436
rect -15360 17355 -15320 17404
rect -15360 17325 -15355 17355
rect -15325 17325 -15320 17355
rect -15360 17195 -15320 17325
rect -15360 17165 -15355 17195
rect -15325 17165 -15320 17195
rect -15360 17116 -15320 17165
rect -15360 17084 -15356 17116
rect -15324 17084 -15320 17116
rect -15360 17036 -15320 17084
rect -15360 17004 -15356 17036
rect -15324 17004 -15320 17036
rect -15360 16956 -15320 17004
rect -15360 16924 -15356 16956
rect -15324 16924 -15320 16956
rect -15360 16876 -15320 16924
rect -15360 16844 -15356 16876
rect -15324 16844 -15320 16876
rect -15360 16796 -15320 16844
rect -15360 16764 -15356 16796
rect -15324 16764 -15320 16796
rect -15360 16716 -15320 16764
rect -15360 16684 -15356 16716
rect -15324 16684 -15320 16716
rect -15360 16636 -15320 16684
rect -15360 16604 -15356 16636
rect -15324 16604 -15320 16636
rect -15360 16556 -15320 16604
rect -15360 16524 -15356 16556
rect -15324 16524 -15320 16556
rect -15360 16476 -15320 16524
rect -15360 16444 -15356 16476
rect -15324 16444 -15320 16476
rect -15360 16395 -15320 16444
rect -15360 16365 -15355 16395
rect -15325 16365 -15320 16395
rect -15360 16315 -15320 16365
rect -15280 18795 -15240 18800
rect -15280 18765 -15275 18795
rect -15245 18765 -15240 18795
rect -15280 16395 -15240 18765
rect -15280 16365 -15275 16395
rect -15245 16365 -15240 16395
rect -15280 16360 -15240 16365
rect -15200 18715 -15160 18844
rect -15200 18685 -15195 18715
rect -15165 18685 -15160 18715
rect -15200 18556 -15160 18685
rect -15120 21035 -15080 21040
rect -15120 21005 -15115 21035
rect -15085 21005 -15080 21035
rect -15120 18635 -15080 21005
rect -15120 18605 -15115 18635
rect -15085 18605 -15080 18635
rect -15120 18600 -15080 18605
rect -15040 20955 -15000 21085
rect -15040 20925 -15035 20955
rect -15005 20925 -15000 20955
rect -15040 20876 -15000 20925
rect -14960 21435 -14920 21440
rect -14960 21405 -14955 21435
rect -14925 21405 -14920 21435
rect -14960 21275 -14920 21405
rect -14960 21245 -14955 21275
rect -14925 21245 -14920 21275
rect -14960 21115 -14920 21245
rect -14960 21085 -14955 21115
rect -14925 21085 -14920 21115
rect -14960 20955 -14920 21085
rect -14960 20925 -14955 20955
rect -14925 20925 -14920 20955
rect -14960 20920 -14920 20925
rect -14880 21435 -14840 21440
rect -14880 21405 -14875 21435
rect -14845 21405 -14840 21435
rect -14880 21275 -14840 21405
rect -14880 21245 -14875 21275
rect -14845 21245 -14840 21275
rect -14880 21115 -14840 21245
rect -14880 21085 -14875 21115
rect -14845 21085 -14840 21115
rect -14880 20955 -14840 21085
rect -14880 20925 -14875 20955
rect -14845 20925 -14840 20955
rect -14880 20920 -14840 20925
rect -14800 21435 -14760 21440
rect -14800 21405 -14795 21435
rect -14765 21405 -14760 21435
rect -14800 21275 -14760 21405
rect -14800 21245 -14795 21275
rect -14765 21245 -14760 21275
rect -14800 21115 -14760 21245
rect -14800 21085 -14795 21115
rect -14765 21085 -14760 21115
rect -14800 20955 -14760 21085
rect -14800 20925 -14795 20955
rect -14765 20925 -14760 20955
rect -14800 20920 -14760 20925
rect -14720 21435 -14680 21440
rect -14720 21405 -14715 21435
rect -14685 21405 -14680 21435
rect -14720 21275 -14680 21405
rect -14720 21245 -14715 21275
rect -14685 21245 -14680 21275
rect -14720 21115 -14680 21245
rect -14720 21085 -14715 21115
rect -14685 21085 -14680 21115
rect -14720 20955 -14680 21085
rect -14720 20925 -14715 20955
rect -14685 20925 -14680 20955
rect -14720 20920 -14680 20925
rect -14640 21435 -14600 21440
rect -14640 21405 -14635 21435
rect -14605 21405 -14600 21435
rect -14640 21275 -14600 21405
rect -14640 21245 -14635 21275
rect -14605 21245 -14600 21275
rect -14640 21115 -14600 21245
rect -14640 21085 -14635 21115
rect -14605 21085 -14600 21115
rect -14640 20955 -14600 21085
rect -14640 20925 -14635 20955
rect -14605 20925 -14600 20955
rect -14640 20920 -14600 20925
rect -14560 21435 -14520 21440
rect -14560 21405 -14555 21435
rect -14525 21405 -14520 21435
rect -14560 21275 -14520 21405
rect -14560 21245 -14555 21275
rect -14525 21245 -14520 21275
rect -14560 21115 -14520 21245
rect -14560 21085 -14555 21115
rect -14525 21085 -14520 21115
rect -14560 20955 -14520 21085
rect -14560 20925 -14555 20955
rect -14525 20925 -14520 20955
rect -14560 20920 -14520 20925
rect -14480 21435 -14440 21440
rect -14480 21405 -14475 21435
rect -14445 21405 -14440 21435
rect -14480 21275 -14440 21405
rect -14480 21245 -14475 21275
rect -14445 21245 -14440 21275
rect -14480 21115 -14440 21245
rect -14480 21085 -14475 21115
rect -14445 21085 -14440 21115
rect -14480 20955 -14440 21085
rect -14480 20925 -14475 20955
rect -14445 20925 -14440 20955
rect -14480 20920 -14440 20925
rect -14400 21435 -14360 21440
rect -14400 21405 -14395 21435
rect -14365 21405 -14360 21435
rect -14400 21275 -14360 21405
rect -14400 21245 -14395 21275
rect -14365 21245 -14360 21275
rect -14400 21115 -14360 21245
rect -14400 21085 -14395 21115
rect -14365 21085 -14360 21115
rect -14400 20955 -14360 21085
rect -14400 20925 -14395 20955
rect -14365 20925 -14360 20955
rect -14400 20920 -14360 20925
rect -14320 21435 -14280 21440
rect -14320 21405 -14315 21435
rect -14285 21405 -14280 21435
rect -14320 21275 -14280 21405
rect -14320 21245 -14315 21275
rect -14285 21245 -14280 21275
rect -14320 21115 -14280 21245
rect -14320 21085 -14315 21115
rect -14285 21085 -14280 21115
rect -14320 20955 -14280 21085
rect -14320 20925 -14315 20955
rect -14285 20925 -14280 20955
rect -14320 20920 -14280 20925
rect -14240 21435 -14200 21440
rect -14240 21405 -14235 21435
rect -14205 21405 -14200 21435
rect -14240 21275 -14200 21405
rect -14240 21245 -14235 21275
rect -14205 21245 -14200 21275
rect -14240 21115 -14200 21245
rect -14240 21085 -14235 21115
rect -14205 21085 -14200 21115
rect -14240 20955 -14200 21085
rect -14240 20925 -14235 20955
rect -14205 20925 -14200 20955
rect -14240 20920 -14200 20925
rect -14160 21435 -14120 21440
rect -14160 21405 -14155 21435
rect -14125 21405 -14120 21435
rect -14160 21275 -14120 21405
rect -14160 21245 -14155 21275
rect -14125 21245 -14120 21275
rect -14160 21115 -14120 21245
rect -14160 21085 -14155 21115
rect -14125 21085 -14120 21115
rect -14160 20955 -14120 21085
rect -14160 20925 -14155 20955
rect -14125 20925 -14120 20955
rect -14160 20920 -14120 20925
rect -14080 21435 -14040 21440
rect -14080 21405 -14075 21435
rect -14045 21405 -14040 21435
rect -14080 21275 -14040 21405
rect -14080 21245 -14075 21275
rect -14045 21245 -14040 21275
rect -14080 21115 -14040 21245
rect -14080 21085 -14075 21115
rect -14045 21085 -14040 21115
rect -14080 20955 -14040 21085
rect -14080 20925 -14075 20955
rect -14045 20925 -14040 20955
rect -14080 20920 -14040 20925
rect -14000 21435 -13960 21440
rect -14000 21405 -13995 21435
rect -13965 21405 -13960 21435
rect -14000 21275 -13960 21405
rect -14000 21245 -13995 21275
rect -13965 21245 -13960 21275
rect -14000 21115 -13960 21245
rect -14000 21085 -13995 21115
rect -13965 21085 -13960 21115
rect -14000 20955 -13960 21085
rect -14000 20925 -13995 20955
rect -13965 20925 -13960 20955
rect -14000 20920 -13960 20925
rect -13920 21435 -13880 21440
rect -13920 21405 -13915 21435
rect -13885 21405 -13880 21435
rect -13920 21275 -13880 21405
rect -13920 21245 -13915 21275
rect -13885 21245 -13880 21275
rect -13920 21115 -13880 21245
rect -13920 21085 -13915 21115
rect -13885 21085 -13880 21115
rect -13920 20955 -13880 21085
rect -13920 20925 -13915 20955
rect -13885 20925 -13880 20955
rect -13920 20920 -13880 20925
rect -13840 21435 -13800 21440
rect -13840 21405 -13835 21435
rect -13805 21405 -13800 21435
rect -13840 21275 -13800 21405
rect -13840 21245 -13835 21275
rect -13805 21245 -13800 21275
rect -13840 21115 -13800 21245
rect -13840 21085 -13835 21115
rect -13805 21085 -13800 21115
rect -13840 20955 -13800 21085
rect -13840 20925 -13835 20955
rect -13805 20925 -13800 20955
rect -13840 20920 -13800 20925
rect -13760 21435 -13720 21440
rect -13760 21405 -13755 21435
rect -13725 21405 -13720 21435
rect -13760 21275 -13720 21405
rect -13760 21245 -13755 21275
rect -13725 21245 -13720 21275
rect -13760 21115 -13720 21245
rect -13760 21085 -13755 21115
rect -13725 21085 -13720 21115
rect -13760 20955 -13720 21085
rect -13760 20925 -13755 20955
rect -13725 20925 -13720 20955
rect -13760 20920 -13720 20925
rect -13680 21435 -13640 21440
rect -13680 21405 -13675 21435
rect -13645 21405 -13640 21435
rect -13680 21275 -13640 21405
rect -13680 21245 -13675 21275
rect -13645 21245 -13640 21275
rect -13680 21115 -13640 21245
rect -13680 21085 -13675 21115
rect -13645 21085 -13640 21115
rect -13680 20955 -13640 21085
rect -13680 20925 -13675 20955
rect -13645 20925 -13640 20955
rect -13680 20920 -13640 20925
rect -13600 21435 -13560 21440
rect -13600 21405 -13595 21435
rect -13565 21405 -13560 21435
rect -13600 21275 -13560 21405
rect -13600 21245 -13595 21275
rect -13565 21245 -13560 21275
rect -13600 21115 -13560 21245
rect -13600 21085 -13595 21115
rect -13565 21085 -13560 21115
rect -13600 20955 -13560 21085
rect -13600 20925 -13595 20955
rect -13565 20925 -13560 20955
rect -13600 20920 -13560 20925
rect -13520 21435 -13480 21440
rect -13520 21405 -13515 21435
rect -13485 21405 -13480 21435
rect -13520 21275 -13480 21405
rect -13520 21245 -13515 21275
rect -13485 21245 -13480 21275
rect -13520 21115 -13480 21245
rect -13520 21085 -13515 21115
rect -13485 21085 -13480 21115
rect -13520 20955 -13480 21085
rect -13520 20925 -13515 20955
rect -13485 20925 -13480 20955
rect -13520 20920 -13480 20925
rect -13440 21435 -13400 21440
rect -13440 21405 -13435 21435
rect -13405 21405 -13400 21435
rect -13440 21275 -13400 21405
rect -13440 21245 -13435 21275
rect -13405 21245 -13400 21275
rect -13440 21115 -13400 21245
rect -13440 21085 -13435 21115
rect -13405 21085 -13400 21115
rect -13440 20955 -13400 21085
rect -13440 20925 -13435 20955
rect -13405 20925 -13400 20955
rect -13440 20920 -13400 20925
rect -13360 21435 -13320 21440
rect -13360 21405 -13355 21435
rect -13325 21405 -13320 21435
rect -13360 21275 -13320 21405
rect -13360 21245 -13355 21275
rect -13325 21245 -13320 21275
rect -13360 21115 -13320 21245
rect -13360 21085 -13355 21115
rect -13325 21085 -13320 21115
rect -13360 20955 -13320 21085
rect -13360 20925 -13355 20955
rect -13325 20925 -13320 20955
rect -13360 20920 -13320 20925
rect -13280 21435 -13240 21440
rect -13280 21405 -13275 21435
rect -13245 21405 -13240 21435
rect -13280 21275 -13240 21405
rect -13280 21245 -13275 21275
rect -13245 21245 -13240 21275
rect -13280 21115 -13240 21245
rect -13280 21085 -13275 21115
rect -13245 21085 -13240 21115
rect -13280 20955 -13240 21085
rect -13280 20925 -13275 20955
rect -13245 20925 -13240 20955
rect -13280 20920 -13240 20925
rect -13200 21435 -13160 21440
rect -13200 21405 -13195 21435
rect -13165 21405 -13160 21435
rect -13200 21275 -13160 21405
rect -13200 21245 -13195 21275
rect -13165 21245 -13160 21275
rect -13200 21115 -13160 21245
rect -13200 21085 -13195 21115
rect -13165 21085 -13160 21115
rect -13200 20955 -13160 21085
rect -13200 20925 -13195 20955
rect -13165 20925 -13160 20955
rect -13200 20920 -13160 20925
rect -13120 21435 -13080 21440
rect -13120 21405 -13115 21435
rect -13085 21405 -13080 21435
rect -13120 21275 -13080 21405
rect -13120 21245 -13115 21275
rect -13085 21245 -13080 21275
rect -13120 21115 -13080 21245
rect -13120 21085 -13115 21115
rect -13085 21085 -13080 21115
rect -13120 20955 -13080 21085
rect -13120 20925 -13115 20955
rect -13085 20925 -13080 20955
rect -13120 20920 -13080 20925
rect -13040 21435 -13000 21440
rect -13040 21405 -13035 21435
rect -13005 21405 -13000 21435
rect -13040 21275 -13000 21405
rect -13040 21245 -13035 21275
rect -13005 21245 -13000 21275
rect -13040 21115 -13000 21245
rect -13040 21085 -13035 21115
rect -13005 21085 -13000 21115
rect -13040 20955 -13000 21085
rect -13040 20925 -13035 20955
rect -13005 20925 -13000 20955
rect -13040 20920 -13000 20925
rect -12960 21435 -12920 21440
rect -12960 21405 -12955 21435
rect -12925 21405 -12920 21435
rect -12960 21275 -12920 21405
rect -12960 21245 -12955 21275
rect -12925 21245 -12920 21275
rect -12960 21115 -12920 21245
rect -12960 21085 -12955 21115
rect -12925 21085 -12920 21115
rect -12960 20955 -12920 21085
rect -12960 20925 -12955 20955
rect -12925 20925 -12920 20955
rect -12960 20920 -12920 20925
rect -12880 21435 -12840 21440
rect -12880 21405 -12875 21435
rect -12845 21405 -12840 21435
rect -12880 21275 -12840 21405
rect -12880 21245 -12875 21275
rect -12845 21245 -12840 21275
rect -12880 21115 -12840 21245
rect -12880 21085 -12875 21115
rect -12845 21085 -12840 21115
rect -12880 20955 -12840 21085
rect -12880 20925 -12875 20955
rect -12845 20925 -12840 20955
rect -12880 20920 -12840 20925
rect -12800 21435 -12760 21440
rect -12800 21405 -12795 21435
rect -12765 21405 -12760 21435
rect -12800 21275 -12760 21405
rect -12800 21245 -12795 21275
rect -12765 21245 -12760 21275
rect -12800 21115 -12760 21245
rect -12800 21085 -12795 21115
rect -12765 21085 -12760 21115
rect -12800 20955 -12760 21085
rect -12800 20925 -12795 20955
rect -12765 20925 -12760 20955
rect -12800 20920 -12760 20925
rect -12720 21435 -12680 21440
rect -12720 21405 -12715 21435
rect -12685 21405 -12680 21435
rect -12720 21275 -12680 21405
rect -12720 21245 -12715 21275
rect -12685 21245 -12680 21275
rect -12720 21115 -12680 21245
rect -12720 21085 -12715 21115
rect -12685 21085 -12680 21115
rect -12720 20955 -12680 21085
rect -12720 20925 -12715 20955
rect -12685 20925 -12680 20955
rect -12720 20920 -12680 20925
rect -12640 21435 -12600 21440
rect -12640 21405 -12635 21435
rect -12605 21405 -12600 21435
rect -12640 21275 -12600 21405
rect -12640 21245 -12635 21275
rect -12605 21245 -12600 21275
rect -12640 21115 -12600 21245
rect -12640 21085 -12635 21115
rect -12605 21085 -12600 21115
rect -12640 20955 -12600 21085
rect -12640 20925 -12635 20955
rect -12605 20925 -12600 20955
rect -12640 20920 -12600 20925
rect -12560 21435 -12520 21440
rect -12560 21405 -12555 21435
rect -12525 21405 -12520 21435
rect -12560 21275 -12520 21405
rect -12560 21245 -12555 21275
rect -12525 21245 -12520 21275
rect -12560 21115 -12520 21245
rect -12560 21085 -12555 21115
rect -12525 21085 -12520 21115
rect -12560 20955 -12520 21085
rect -12560 20925 -12555 20955
rect -12525 20925 -12520 20955
rect -12560 20920 -12520 20925
rect -12480 21435 -12440 21440
rect -12480 21405 -12475 21435
rect -12445 21405 -12440 21435
rect -12480 21275 -12440 21405
rect -12480 21245 -12475 21275
rect -12445 21245 -12440 21275
rect -12480 21115 -12440 21245
rect -12480 21085 -12475 21115
rect -12445 21085 -12440 21115
rect -12480 20955 -12440 21085
rect -12480 20925 -12475 20955
rect -12445 20925 -12440 20955
rect -12480 20920 -12440 20925
rect -12400 21435 -12360 21440
rect -12400 21405 -12395 21435
rect -12365 21405 -12360 21435
rect -12400 21275 -12360 21405
rect -12400 21245 -12395 21275
rect -12365 21245 -12360 21275
rect -12400 21115 -12360 21245
rect -12400 21085 -12395 21115
rect -12365 21085 -12360 21115
rect -12400 20955 -12360 21085
rect -12400 20925 -12395 20955
rect -12365 20925 -12360 20955
rect -12400 20920 -12360 20925
rect -12320 21435 -12280 21440
rect -12320 21405 -12315 21435
rect -12285 21405 -12280 21435
rect -12320 21275 -12280 21405
rect -12320 21245 -12315 21275
rect -12285 21245 -12280 21275
rect -12320 21115 -12280 21245
rect -12320 21085 -12315 21115
rect -12285 21085 -12280 21115
rect -12320 20955 -12280 21085
rect -12320 20925 -12315 20955
rect -12285 20925 -12280 20955
rect -12320 20920 -12280 20925
rect -12240 21435 -12200 21440
rect -12240 21405 -12235 21435
rect -12205 21405 -12200 21435
rect -12240 21275 -12200 21405
rect -12240 21245 -12235 21275
rect -12205 21245 -12200 21275
rect -12240 21115 -12200 21245
rect -12240 21085 -12235 21115
rect -12205 21085 -12200 21115
rect -12240 20955 -12200 21085
rect -12240 20925 -12235 20955
rect -12205 20925 -12200 20955
rect -12240 20920 -12200 20925
rect -12160 21435 -12120 21440
rect -12160 21405 -12155 21435
rect -12125 21405 -12120 21435
rect -12160 21275 -12120 21405
rect -12160 21245 -12155 21275
rect -12125 21245 -12120 21275
rect -12160 21115 -12120 21245
rect -12160 21085 -12155 21115
rect -12125 21085 -12120 21115
rect -12160 20955 -12120 21085
rect -12160 20925 -12155 20955
rect -12125 20925 -12120 20955
rect -12160 20920 -12120 20925
rect -12080 21435 -12040 21440
rect -12080 21405 -12075 21435
rect -12045 21405 -12040 21435
rect -12080 21275 -12040 21405
rect -12080 21245 -12075 21275
rect -12045 21245 -12040 21275
rect -12080 21115 -12040 21245
rect -12080 21085 -12075 21115
rect -12045 21085 -12040 21115
rect -12080 20955 -12040 21085
rect -12080 20925 -12075 20955
rect -12045 20925 -12040 20955
rect -12080 20920 -12040 20925
rect -12000 21435 -11960 21440
rect -12000 21405 -11995 21435
rect -11965 21405 -11960 21435
rect -12000 21275 -11960 21405
rect -12000 21245 -11995 21275
rect -11965 21245 -11960 21275
rect -12000 21115 -11960 21245
rect -12000 21085 -11995 21115
rect -11965 21085 -11960 21115
rect -12000 20955 -11960 21085
rect -12000 20925 -11995 20955
rect -11965 20925 -11960 20955
rect -12000 20920 -11960 20925
rect -11920 21435 -11880 21440
rect -11920 21405 -11915 21435
rect -11885 21405 -11880 21435
rect -11920 21275 -11880 21405
rect -11920 21245 -11915 21275
rect -11885 21245 -11880 21275
rect -11920 21115 -11880 21245
rect -11920 21085 -11915 21115
rect -11885 21085 -11880 21115
rect -11920 20955 -11880 21085
rect -11920 20925 -11915 20955
rect -11885 20925 -11880 20955
rect -11920 20920 -11880 20925
rect -11840 21435 -11800 21440
rect -11840 21405 -11835 21435
rect -11805 21405 -11800 21435
rect -11840 21275 -11800 21405
rect -11840 21245 -11835 21275
rect -11805 21245 -11800 21275
rect -11840 21115 -11800 21245
rect -11840 21085 -11835 21115
rect -11805 21085 -11800 21115
rect -11840 20955 -11800 21085
rect -11840 20925 -11835 20955
rect -11805 20925 -11800 20955
rect -11840 20920 -11800 20925
rect -11760 21435 -11720 21440
rect -11760 21405 -11755 21435
rect -11725 21405 -11720 21435
rect -11760 21275 -11720 21405
rect -11760 21245 -11755 21275
rect -11725 21245 -11720 21275
rect -11760 21115 -11720 21245
rect -11760 21085 -11755 21115
rect -11725 21085 -11720 21115
rect -11760 20955 -11720 21085
rect -11760 20925 -11755 20955
rect -11725 20925 -11720 20955
rect -11760 20920 -11720 20925
rect -11680 21435 -11640 21440
rect -11680 21405 -11675 21435
rect -11645 21405 -11640 21435
rect -11680 21275 -11640 21405
rect -11680 21245 -11675 21275
rect -11645 21245 -11640 21275
rect -11680 21115 -11640 21245
rect -11680 21085 -11675 21115
rect -11645 21085 -11640 21115
rect -11680 20955 -11640 21085
rect -11680 20925 -11675 20955
rect -11645 20925 -11640 20955
rect -11680 20920 -11640 20925
rect -11600 21435 -11560 21440
rect -11600 21405 -11595 21435
rect -11565 21405 -11560 21435
rect -11600 21275 -11560 21405
rect -11600 21245 -11595 21275
rect -11565 21245 -11560 21275
rect -11600 21115 -11560 21245
rect -11600 21085 -11595 21115
rect -11565 21085 -11560 21115
rect -11600 20955 -11560 21085
rect -11600 20925 -11595 20955
rect -11565 20925 -11560 20955
rect -11600 20920 -11560 20925
rect -11520 21435 -11480 21440
rect -11520 21405 -11515 21435
rect -11485 21405 -11480 21435
rect -11520 21275 -11480 21405
rect -11520 21245 -11515 21275
rect -11485 21245 -11480 21275
rect -11520 21115 -11480 21245
rect -11520 21085 -11515 21115
rect -11485 21085 -11480 21115
rect -11520 20955 -11480 21085
rect -11520 20925 -11515 20955
rect -11485 20925 -11480 20955
rect -11520 20920 -11480 20925
rect -11440 21435 -11400 21440
rect -11440 21405 -11435 21435
rect -11405 21405 -11400 21435
rect -11440 21275 -11400 21405
rect -11440 21245 -11435 21275
rect -11405 21245 -11400 21275
rect -11440 21115 -11400 21245
rect -11440 21085 -11435 21115
rect -11405 21085 -11400 21115
rect -11440 20955 -11400 21085
rect -11440 20925 -11435 20955
rect -11405 20925 -11400 20955
rect -11440 20920 -11400 20925
rect -11360 21435 -11320 21440
rect -11360 21405 -11355 21435
rect -11325 21405 -11320 21435
rect -11360 21275 -11320 21405
rect -11360 21245 -11355 21275
rect -11325 21245 -11320 21275
rect -11360 21115 -11320 21245
rect -11360 21085 -11355 21115
rect -11325 21085 -11320 21115
rect -11360 20955 -11320 21085
rect -11360 20925 -11355 20955
rect -11325 20925 -11320 20955
rect -11360 20920 -11320 20925
rect -11280 21435 -11240 21440
rect -11280 21405 -11275 21435
rect -11245 21405 -11240 21435
rect -11280 21275 -11240 21405
rect -11280 21245 -11275 21275
rect -11245 21245 -11240 21275
rect -11280 21115 -11240 21245
rect -11280 21085 -11275 21115
rect -11245 21085 -11240 21115
rect -11280 20955 -11240 21085
rect -11280 20925 -11275 20955
rect -11245 20925 -11240 20955
rect -11280 20920 -11240 20925
rect -11200 21435 -11160 21440
rect -11200 21405 -11195 21435
rect -11165 21405 -11160 21435
rect -11200 21275 -11160 21405
rect -11200 21245 -11195 21275
rect -11165 21245 -11160 21275
rect -11200 21115 -11160 21245
rect -11200 21085 -11195 21115
rect -11165 21085 -11160 21115
rect -11200 20955 -11160 21085
rect -11200 20925 -11195 20955
rect -11165 20925 -11160 20955
rect -11200 20920 -11160 20925
rect -11120 21435 -11080 21440
rect -11120 21405 -11115 21435
rect -11085 21405 -11080 21435
rect -11120 21275 -11080 21405
rect -11120 21245 -11115 21275
rect -11085 21245 -11080 21275
rect -11120 21115 -11080 21245
rect -11120 21085 -11115 21115
rect -11085 21085 -11080 21115
rect -11120 20955 -11080 21085
rect -11120 20925 -11115 20955
rect -11085 20925 -11080 20955
rect -11120 20920 -11080 20925
rect -11040 21435 -11000 21440
rect -11040 21405 -11035 21435
rect -11005 21405 -11000 21435
rect -11040 21275 -11000 21405
rect -11040 21245 -11035 21275
rect -11005 21245 -11000 21275
rect -11040 21115 -11000 21245
rect -11040 21085 -11035 21115
rect -11005 21085 -11000 21115
rect -11040 20955 -11000 21085
rect -11040 20925 -11035 20955
rect -11005 20925 -11000 20955
rect -11040 20920 -11000 20925
rect -10960 21435 -10920 21440
rect -10960 21405 -10955 21435
rect -10925 21405 -10920 21435
rect -10960 21275 -10920 21405
rect -10960 21245 -10955 21275
rect -10925 21245 -10920 21275
rect -10960 21115 -10920 21245
rect -10960 21085 -10955 21115
rect -10925 21085 -10920 21115
rect -10960 20955 -10920 21085
rect -10960 20925 -10955 20955
rect -10925 20925 -10920 20955
rect -10960 20920 -10920 20925
rect -10880 21435 -10840 21440
rect -10880 21405 -10875 21435
rect -10845 21405 -10840 21435
rect -10880 21275 -10840 21405
rect -10880 21245 -10875 21275
rect -10845 21245 -10840 21275
rect -10880 21115 -10840 21245
rect -10880 21085 -10875 21115
rect -10845 21085 -10840 21115
rect -10880 20955 -10840 21085
rect -10880 20925 -10875 20955
rect -10845 20925 -10840 20955
rect -10880 20920 -10840 20925
rect -10800 21435 -10760 21440
rect -10800 21405 -10795 21435
rect -10765 21405 -10760 21435
rect -10800 21275 -10760 21405
rect -10800 21245 -10795 21275
rect -10765 21245 -10760 21275
rect -10800 21115 -10760 21245
rect -10800 21085 -10795 21115
rect -10765 21085 -10760 21115
rect -10800 20955 -10760 21085
rect -10800 20925 -10795 20955
rect -10765 20925 -10760 20955
rect -10800 20920 -10760 20925
rect -10720 21435 -10680 21440
rect -10720 21405 -10715 21435
rect -10685 21405 -10680 21435
rect -10720 21275 -10680 21405
rect -10720 21245 -10715 21275
rect -10685 21245 -10680 21275
rect -10720 21115 -10680 21245
rect -10720 21085 -10715 21115
rect -10685 21085 -10680 21115
rect -10720 20955 -10680 21085
rect -10720 20925 -10715 20955
rect -10685 20925 -10680 20955
rect -10720 20920 -10680 20925
rect -10640 21435 -10600 21440
rect -10640 21405 -10635 21435
rect -10605 21405 -10600 21435
rect -10640 21275 -10600 21405
rect -10640 21245 -10635 21275
rect -10605 21245 -10600 21275
rect -10640 21115 -10600 21245
rect -10640 21085 -10635 21115
rect -10605 21085 -10600 21115
rect -10640 20955 -10600 21085
rect -10640 20925 -10635 20955
rect -10605 20925 -10600 20955
rect -10640 20920 -10600 20925
rect -10560 21435 -10520 21440
rect -10560 21405 -10555 21435
rect -10525 21405 -10520 21435
rect -10560 21275 -10520 21405
rect -10560 21245 -10555 21275
rect -10525 21245 -10520 21275
rect -10560 21115 -10520 21245
rect -10560 21085 -10555 21115
rect -10525 21085 -10520 21115
rect -10560 20955 -10520 21085
rect -10560 20925 -10555 20955
rect -10525 20925 -10520 20955
rect -10560 20920 -10520 20925
rect -10480 21435 -10440 21440
rect -10480 21405 -10475 21435
rect -10445 21405 -10440 21435
rect -10480 21275 -10440 21405
rect -10480 21245 -10475 21275
rect -10445 21245 -10440 21275
rect -10480 21115 -10440 21245
rect -10480 21085 -10475 21115
rect -10445 21085 -10440 21115
rect -10480 20955 -10440 21085
rect -10480 20925 -10475 20955
rect -10445 20925 -10440 20955
rect -10480 20920 -10440 20925
rect -10400 21435 -10360 21440
rect -10400 21405 -10395 21435
rect -10365 21405 -10360 21435
rect -10400 21275 -10360 21405
rect -10400 21245 -10395 21275
rect -10365 21245 -10360 21275
rect -10400 21115 -10360 21245
rect -10400 21085 -10395 21115
rect -10365 21085 -10360 21115
rect -10400 20955 -10360 21085
rect -10400 20925 -10395 20955
rect -10365 20925 -10360 20955
rect -10400 20920 -10360 20925
rect -10320 21435 -10280 21440
rect -10320 21405 -10315 21435
rect -10285 21405 -10280 21435
rect -10320 21275 -10280 21405
rect -10320 21245 -10315 21275
rect -10285 21245 -10280 21275
rect -10320 21115 -10280 21245
rect -10320 21085 -10315 21115
rect -10285 21085 -10280 21115
rect -10320 20955 -10280 21085
rect -10320 20925 -10315 20955
rect -10285 20925 -10280 20955
rect -10320 20920 -10280 20925
rect -10240 21435 -10200 21440
rect -10240 21405 -10235 21435
rect -10205 21405 -10200 21435
rect -10240 21275 -10200 21405
rect -10240 21245 -10235 21275
rect -10205 21245 -10200 21275
rect -10240 21115 -10200 21245
rect -10240 21085 -10235 21115
rect -10205 21085 -10200 21115
rect -10240 20955 -10200 21085
rect -10240 20925 -10235 20955
rect -10205 20925 -10200 20955
rect -10240 20920 -10200 20925
rect -10160 21435 -10120 21440
rect -10160 21405 -10155 21435
rect -10125 21405 -10120 21435
rect -10160 21275 -10120 21405
rect -10160 21245 -10155 21275
rect -10125 21245 -10120 21275
rect -10160 21115 -10120 21245
rect -10160 21085 -10155 21115
rect -10125 21085 -10120 21115
rect -10160 20955 -10120 21085
rect -10160 20925 -10155 20955
rect -10125 20925 -10120 20955
rect -10160 20920 -10120 20925
rect -10080 21435 -10040 21440
rect -10080 21405 -10075 21435
rect -10045 21405 -10040 21435
rect -10080 21275 -10040 21405
rect -10080 21245 -10075 21275
rect -10045 21245 -10040 21275
rect -10080 21115 -10040 21245
rect -10080 21085 -10075 21115
rect -10045 21085 -10040 21115
rect -10080 20955 -10040 21085
rect -10080 20925 -10075 20955
rect -10045 20925 -10040 20955
rect -10080 20920 -10040 20925
rect -10000 21435 -9960 21440
rect -10000 21405 -9995 21435
rect -9965 21405 -9960 21435
rect -10000 21275 -9960 21405
rect -10000 21245 -9995 21275
rect -9965 21245 -9960 21275
rect -10000 21115 -9960 21245
rect -10000 21085 -9995 21115
rect -9965 21085 -9960 21115
rect -10000 20955 -9960 21085
rect -10000 20925 -9995 20955
rect -9965 20925 -9960 20955
rect -10000 20920 -9960 20925
rect -9920 21435 -9880 21440
rect -9920 21405 -9915 21435
rect -9885 21405 -9880 21435
rect -9920 21275 -9880 21405
rect -9920 21245 -9915 21275
rect -9885 21245 -9880 21275
rect -9920 21115 -9880 21245
rect -9920 21085 -9915 21115
rect -9885 21085 -9880 21115
rect -9920 20955 -9880 21085
rect -9920 20925 -9915 20955
rect -9885 20925 -9880 20955
rect -9920 20920 -9880 20925
rect -9840 21435 -9800 21440
rect -9840 21405 -9835 21435
rect -9805 21405 -9800 21435
rect -9840 21275 -9800 21405
rect -9840 21245 -9835 21275
rect -9805 21245 -9800 21275
rect -9840 21115 -9800 21245
rect -9840 21085 -9835 21115
rect -9805 21085 -9800 21115
rect -9840 20955 -9800 21085
rect -9840 20925 -9835 20955
rect -9805 20925 -9800 20955
rect -9840 20920 -9800 20925
rect -9760 21435 -9720 21440
rect -9760 21405 -9755 21435
rect -9725 21405 -9720 21435
rect -9760 21275 -9720 21405
rect -9760 21245 -9755 21275
rect -9725 21245 -9720 21275
rect -9760 21115 -9720 21245
rect -9760 21085 -9755 21115
rect -9725 21085 -9720 21115
rect -9760 20955 -9720 21085
rect -9760 20925 -9755 20955
rect -9725 20925 -9720 20955
rect -9760 20920 -9720 20925
rect -9680 21435 -9640 21440
rect -9680 21405 -9675 21435
rect -9645 21405 -9640 21435
rect -9680 21275 -9640 21405
rect -9680 21245 -9675 21275
rect -9645 21245 -9640 21275
rect -9680 21115 -9640 21245
rect -9680 21085 -9675 21115
rect -9645 21085 -9640 21115
rect -9680 20955 -9640 21085
rect -9680 20925 -9675 20955
rect -9645 20925 -9640 20955
rect -9680 20920 -9640 20925
rect -9600 21435 -9560 21440
rect -9600 21405 -9595 21435
rect -9565 21405 -9560 21435
rect -9600 21275 -9560 21405
rect -9600 21245 -9595 21275
rect -9565 21245 -9560 21275
rect -9600 21115 -9560 21245
rect -9600 21085 -9595 21115
rect -9565 21085 -9560 21115
rect -9600 20955 -9560 21085
rect -9600 20925 -9595 20955
rect -9565 20925 -9560 20955
rect -9600 20920 -9560 20925
rect -9520 21435 -9480 21440
rect -9520 21405 -9515 21435
rect -9485 21405 -9480 21435
rect -9520 21275 -9480 21405
rect -9520 21245 -9515 21275
rect -9485 21245 -9480 21275
rect -9520 21115 -9480 21245
rect -9520 21085 -9515 21115
rect -9485 21085 -9480 21115
rect -9520 20955 -9480 21085
rect -9520 20925 -9515 20955
rect -9485 20925 -9480 20955
rect -9520 20920 -9480 20925
rect -9440 21435 -9400 21440
rect -9440 21405 -9435 21435
rect -9405 21405 -9400 21435
rect -9440 21275 -9400 21405
rect -9440 21245 -9435 21275
rect -9405 21245 -9400 21275
rect -9440 21115 -9400 21245
rect -9440 21085 -9435 21115
rect -9405 21085 -9400 21115
rect -9440 20955 -9400 21085
rect -9440 20925 -9435 20955
rect -9405 20925 -9400 20955
rect -9440 20920 -9400 20925
rect -9360 21435 -9320 21440
rect -9360 21405 -9355 21435
rect -9325 21405 -9320 21435
rect -9360 21275 -9320 21405
rect -9360 21245 -9355 21275
rect -9325 21245 -9320 21275
rect -9360 21115 -9320 21245
rect -9360 21085 -9355 21115
rect -9325 21085 -9320 21115
rect -9360 20955 -9320 21085
rect -9360 20925 -9355 20955
rect -9325 20925 -9320 20955
rect -9360 20920 -9320 20925
rect -9280 21435 -9240 21440
rect -9280 21405 -9275 21435
rect -9245 21405 -9240 21435
rect -9280 21275 -9240 21405
rect -9280 21245 -9275 21275
rect -9245 21245 -9240 21275
rect -9280 21115 -9240 21245
rect -9280 21085 -9275 21115
rect -9245 21085 -9240 21115
rect -9280 20955 -9240 21085
rect -9280 20925 -9275 20955
rect -9245 20925 -9240 20955
rect -9280 20920 -9240 20925
rect -9200 21435 -9160 21440
rect -9200 21405 -9195 21435
rect -9165 21405 -9160 21435
rect -9200 21275 -9160 21405
rect -9200 21245 -9195 21275
rect -9165 21245 -9160 21275
rect -9200 21115 -9160 21245
rect -9200 21085 -9195 21115
rect -9165 21085 -9160 21115
rect -9200 20955 -9160 21085
rect -9200 20925 -9195 20955
rect -9165 20925 -9160 20955
rect -9200 20920 -9160 20925
rect -9120 21435 -9080 21440
rect -9120 21405 -9115 21435
rect -9085 21405 -9080 21435
rect -9120 21275 -9080 21405
rect -9120 21245 -9115 21275
rect -9085 21245 -9080 21275
rect -9120 21115 -9080 21245
rect -9120 21085 -9115 21115
rect -9085 21085 -9080 21115
rect -9120 20955 -9080 21085
rect -9120 20925 -9115 20955
rect -9085 20925 -9080 20955
rect -9120 20920 -9080 20925
rect -9040 21435 -9000 21440
rect -9040 21405 -9035 21435
rect -9005 21405 -9000 21435
rect -9040 21275 -9000 21405
rect -9040 21245 -9035 21275
rect -9005 21245 -9000 21275
rect -9040 21115 -9000 21245
rect -9040 21085 -9035 21115
rect -9005 21085 -9000 21115
rect -9040 20955 -9000 21085
rect -9040 20925 -9035 20955
rect -9005 20925 -9000 20955
rect -9040 20920 -9000 20925
rect -8960 21435 -8920 21440
rect -8960 21405 -8955 21435
rect -8925 21405 -8920 21435
rect -8960 21275 -8920 21405
rect -8960 21245 -8955 21275
rect -8925 21245 -8920 21275
rect -8960 21115 -8920 21245
rect -8960 21085 -8955 21115
rect -8925 21085 -8920 21115
rect -8960 20955 -8920 21085
rect -8960 20925 -8955 20955
rect -8925 20925 -8920 20955
rect -8960 20920 -8920 20925
rect -8880 21435 -8840 21440
rect -8880 21405 -8875 21435
rect -8845 21405 -8840 21435
rect -8880 21275 -8840 21405
rect -8880 21245 -8875 21275
rect -8845 21245 -8840 21275
rect -8880 21115 -8840 21245
rect -8880 21085 -8875 21115
rect -8845 21085 -8840 21115
rect -8880 20955 -8840 21085
rect -8880 20925 -8875 20955
rect -8845 20925 -8840 20955
rect -8880 20920 -8840 20925
rect -8800 21435 -8760 21440
rect -8800 21405 -8795 21435
rect -8765 21405 -8760 21435
rect -8800 21275 -8760 21405
rect -8800 21245 -8795 21275
rect -8765 21245 -8760 21275
rect -8800 21115 -8760 21245
rect -8800 21085 -8795 21115
rect -8765 21085 -8760 21115
rect -8800 20955 -8760 21085
rect -8800 20925 -8795 20955
rect -8765 20925 -8760 20955
rect -8800 20920 -8760 20925
rect -8720 21435 -8680 21440
rect -8720 21405 -8715 21435
rect -8685 21405 -8680 21435
rect -8720 21275 -8680 21405
rect -8720 21245 -8715 21275
rect -8685 21245 -8680 21275
rect -8720 21115 -8680 21245
rect -8720 21085 -8715 21115
rect -8685 21085 -8680 21115
rect -8720 20955 -8680 21085
rect -8720 20925 -8715 20955
rect -8685 20925 -8680 20955
rect -8720 20920 -8680 20925
rect -8640 21435 -8600 21440
rect -8640 21405 -8635 21435
rect -8605 21405 -8600 21435
rect -8640 21275 -8600 21405
rect -8640 21245 -8635 21275
rect -8605 21245 -8600 21275
rect -8640 21115 -8600 21245
rect -8640 21085 -8635 21115
rect -8605 21085 -8600 21115
rect -8640 20955 -8600 21085
rect -8640 20925 -8635 20955
rect -8605 20925 -8600 20955
rect -8640 20920 -8600 20925
rect -8560 21435 -8520 21440
rect -8560 21405 -8555 21435
rect -8525 21405 -8520 21435
rect -8560 21275 -8520 21405
rect -8560 21245 -8555 21275
rect -8525 21245 -8520 21275
rect -8560 21115 -8520 21245
rect -8560 21085 -8555 21115
rect -8525 21085 -8520 21115
rect -8560 20955 -8520 21085
rect -8560 20925 -8555 20955
rect -8525 20925 -8520 20955
rect -8560 20920 -8520 20925
rect -8480 21435 -8440 21440
rect -8480 21405 -8475 21435
rect -8445 21405 -8440 21435
rect -8480 21275 -8440 21405
rect -8480 21245 -8475 21275
rect -8445 21245 -8440 21275
rect -8480 21115 -8440 21245
rect -8480 21085 -8475 21115
rect -8445 21085 -8440 21115
rect -8480 20955 -8440 21085
rect -8480 20925 -8475 20955
rect -8445 20925 -8440 20955
rect -8480 20920 -8440 20925
rect -8400 21435 -8360 21440
rect -8400 21405 -8395 21435
rect -8365 21405 -8360 21435
rect -8400 21275 -8360 21405
rect -8400 21245 -8395 21275
rect -8365 21245 -8360 21275
rect -8400 21115 -8360 21245
rect -8400 21085 -8395 21115
rect -8365 21085 -8360 21115
rect -8400 20955 -8360 21085
rect -8400 20925 -8395 20955
rect -8365 20925 -8360 20955
rect -8400 20920 -8360 20925
rect -8320 21435 -8280 21440
rect -8320 21405 -8315 21435
rect -8285 21405 -8280 21435
rect -8320 21275 -8280 21405
rect -8320 21245 -8315 21275
rect -8285 21245 -8280 21275
rect -8320 21115 -8280 21245
rect -8320 21085 -8315 21115
rect -8285 21085 -8280 21115
rect -8320 20955 -8280 21085
rect -8320 20925 -8315 20955
rect -8285 20925 -8280 20955
rect -8320 20920 -8280 20925
rect -8240 21435 -8200 21440
rect -8240 21405 -8235 21435
rect -8205 21405 -8200 21435
rect -8240 21275 -8200 21405
rect -8240 21245 -8235 21275
rect -8205 21245 -8200 21275
rect -8240 21115 -8200 21245
rect -8240 21085 -8235 21115
rect -8205 21085 -8200 21115
rect -8240 20955 -8200 21085
rect -8240 20925 -8235 20955
rect -8205 20925 -8200 20955
rect -8240 20920 -8200 20925
rect -8160 21435 -8120 21440
rect -8160 21405 -8155 21435
rect -8125 21405 -8120 21435
rect -8160 21275 -8120 21405
rect -8160 21245 -8155 21275
rect -8125 21245 -8120 21275
rect -8160 21115 -8120 21245
rect -8160 21085 -8155 21115
rect -8125 21085 -8120 21115
rect -8160 20955 -8120 21085
rect -8160 20925 -8155 20955
rect -8125 20925 -8120 20955
rect -8160 20920 -8120 20925
rect -8080 21435 -8040 21440
rect -8080 21405 -8075 21435
rect -8045 21405 -8040 21435
rect -8080 21275 -8040 21405
rect -8080 21245 -8075 21275
rect -8045 21245 -8040 21275
rect -8080 21115 -8040 21245
rect -8080 21085 -8075 21115
rect -8045 21085 -8040 21115
rect -8080 20955 -8040 21085
rect -8080 20925 -8075 20955
rect -8045 20925 -8040 20955
rect -8080 20920 -8040 20925
rect -8000 21435 -7960 21440
rect -8000 21405 -7995 21435
rect -7965 21405 -7960 21435
rect -8000 21275 -7960 21405
rect -8000 21245 -7995 21275
rect -7965 21245 -7960 21275
rect -8000 21115 -7960 21245
rect -8000 21085 -7995 21115
rect -7965 21085 -7960 21115
rect -8000 20955 -7960 21085
rect -8000 20925 -7995 20955
rect -7965 20925 -7960 20955
rect -8000 20920 -7960 20925
rect -7920 21435 -7880 21440
rect -7920 21405 -7915 21435
rect -7885 21405 -7880 21435
rect -7920 21275 -7880 21405
rect -7920 21245 -7915 21275
rect -7885 21245 -7880 21275
rect -7920 21115 -7880 21245
rect -7920 21085 -7915 21115
rect -7885 21085 -7880 21115
rect -7920 20955 -7880 21085
rect -7920 20925 -7915 20955
rect -7885 20925 -7880 20955
rect -7920 20920 -7880 20925
rect -7840 21435 -7800 21440
rect -7840 21405 -7835 21435
rect -7805 21405 -7800 21435
rect -7840 21275 -7800 21405
rect -7840 21245 -7835 21275
rect -7805 21245 -7800 21275
rect -7840 21115 -7800 21245
rect -7840 21085 -7835 21115
rect -7805 21085 -7800 21115
rect -7840 20955 -7800 21085
rect -7840 20925 -7835 20955
rect -7805 20925 -7800 20955
rect -7840 20920 -7800 20925
rect -7760 21435 -7720 21440
rect -7760 21405 -7755 21435
rect -7725 21405 -7720 21435
rect -7760 21275 -7720 21405
rect -7760 21245 -7755 21275
rect -7725 21245 -7720 21275
rect -7760 21115 -7720 21245
rect -7760 21085 -7755 21115
rect -7725 21085 -7720 21115
rect -7760 20955 -7720 21085
rect -7760 20925 -7755 20955
rect -7725 20925 -7720 20955
rect -7760 20920 -7720 20925
rect -7680 21435 -7640 21440
rect -7680 21405 -7675 21435
rect -7645 21405 -7640 21435
rect -7680 21275 -7640 21405
rect -7680 21245 -7675 21275
rect -7645 21245 -7640 21275
rect -7680 21115 -7640 21245
rect -7680 21085 -7675 21115
rect -7645 21085 -7640 21115
rect -7680 20955 -7640 21085
rect -7680 20925 -7675 20955
rect -7645 20925 -7640 20955
rect -7680 20920 -7640 20925
rect -7600 21435 -7560 21440
rect -7600 21405 -7595 21435
rect -7565 21405 -7560 21435
rect -7600 21275 -7560 21405
rect -7600 21245 -7595 21275
rect -7565 21245 -7560 21275
rect -7600 21115 -7560 21245
rect -7600 21085 -7595 21115
rect -7565 21085 -7560 21115
rect -7600 20955 -7560 21085
rect -7600 20925 -7595 20955
rect -7565 20925 -7560 20955
rect -7600 20920 -7560 20925
rect -7520 21435 -7480 21440
rect -7520 21405 -7515 21435
rect -7485 21405 -7480 21435
rect -7520 21275 -7480 21405
rect -7520 21245 -7515 21275
rect -7485 21245 -7480 21275
rect -7520 21115 -7480 21245
rect -7520 21085 -7515 21115
rect -7485 21085 -7480 21115
rect -7520 20955 -7480 21085
rect -7520 20925 -7515 20955
rect -7485 20925 -7480 20955
rect -7520 20920 -7480 20925
rect -7440 21435 -7400 21440
rect -7440 21405 -7435 21435
rect -7405 21405 -7400 21435
rect -7440 21275 -7400 21405
rect -7440 21245 -7435 21275
rect -7405 21245 -7400 21275
rect -7440 21115 -7400 21245
rect -7440 21085 -7435 21115
rect -7405 21085 -7400 21115
rect -7440 20955 -7400 21085
rect -7440 20925 -7435 20955
rect -7405 20925 -7400 20955
rect -7440 20920 -7400 20925
rect -7360 21435 -7320 21440
rect -7360 21405 -7355 21435
rect -7325 21405 -7320 21435
rect -7360 21275 -7320 21405
rect -7360 21245 -7355 21275
rect -7325 21245 -7320 21275
rect -7360 21115 -7320 21245
rect -7360 21085 -7355 21115
rect -7325 21085 -7320 21115
rect -7360 20955 -7320 21085
rect -7360 20925 -7355 20955
rect -7325 20925 -7320 20955
rect -7360 20920 -7320 20925
rect -7280 21435 -7240 21440
rect -7280 21405 -7275 21435
rect -7245 21405 -7240 21435
rect -7280 21275 -7240 21405
rect -7280 21245 -7275 21275
rect -7245 21245 -7240 21275
rect -7280 21115 -7240 21245
rect -7280 21085 -7275 21115
rect -7245 21085 -7240 21115
rect -7280 20955 -7240 21085
rect -7280 20925 -7275 20955
rect -7245 20925 -7240 20955
rect -7280 20920 -7240 20925
rect -7200 21435 -7160 21440
rect -7200 21405 -7195 21435
rect -7165 21405 -7160 21435
rect -7200 21275 -7160 21405
rect -7200 21245 -7195 21275
rect -7165 21245 -7160 21275
rect -7200 21115 -7160 21245
rect -7200 21085 -7195 21115
rect -7165 21085 -7160 21115
rect -7200 20955 -7160 21085
rect -7200 20925 -7195 20955
rect -7165 20925 -7160 20955
rect -7200 20920 -7160 20925
rect -7120 21435 -7080 21440
rect -7120 21405 -7115 21435
rect -7085 21405 -7080 21435
rect -7120 21275 -7080 21405
rect -7120 21245 -7115 21275
rect -7085 21245 -7080 21275
rect -7120 21115 -7080 21245
rect -7120 21085 -7115 21115
rect -7085 21085 -7080 21115
rect -7120 20955 -7080 21085
rect -7120 20925 -7115 20955
rect -7085 20925 -7080 20955
rect -7120 20920 -7080 20925
rect -7040 21435 -7000 21440
rect -7040 21405 -7035 21435
rect -7005 21405 -7000 21435
rect -7040 21275 -7000 21405
rect -7040 21245 -7035 21275
rect -7005 21245 -7000 21275
rect -7040 21115 -7000 21245
rect -7040 21085 -7035 21115
rect -7005 21085 -7000 21115
rect -7040 20955 -7000 21085
rect -7040 20925 -7035 20955
rect -7005 20925 -7000 20955
rect -7040 20920 -7000 20925
rect -6960 21435 -6920 21440
rect -6960 21405 -6955 21435
rect -6925 21405 -6920 21435
rect -6960 21275 -6920 21405
rect -6960 21245 -6955 21275
rect -6925 21245 -6920 21275
rect -6960 21115 -6920 21245
rect -6960 21085 -6955 21115
rect -6925 21085 -6920 21115
rect -6960 20955 -6920 21085
rect -6960 20925 -6955 20955
rect -6925 20925 -6920 20955
rect -6960 20920 -6920 20925
rect -6880 21435 -6840 21440
rect -6880 21405 -6875 21435
rect -6845 21405 -6840 21435
rect -6880 21275 -6840 21405
rect -6880 21245 -6875 21275
rect -6845 21245 -6840 21275
rect -6880 21115 -6840 21245
rect -6880 21085 -6875 21115
rect -6845 21085 -6840 21115
rect -6880 20955 -6840 21085
rect -6880 20925 -6875 20955
rect -6845 20925 -6840 20955
rect -6880 20920 -6840 20925
rect -6800 21435 -6760 21440
rect -6800 21405 -6795 21435
rect -6765 21405 -6760 21435
rect -6800 21275 -6760 21405
rect -6800 21245 -6795 21275
rect -6765 21245 -6760 21275
rect -6800 21115 -6760 21245
rect -6800 21085 -6795 21115
rect -6765 21085 -6760 21115
rect -6800 20955 -6760 21085
rect -6800 20925 -6795 20955
rect -6765 20925 -6760 20955
rect -6800 20920 -6760 20925
rect -6720 21435 -6680 21440
rect -6720 21405 -6715 21435
rect -6685 21405 -6680 21435
rect -6720 21275 -6680 21405
rect -6720 21245 -6715 21275
rect -6685 21245 -6680 21275
rect -6720 21115 -6680 21245
rect -6720 21085 -6715 21115
rect -6685 21085 -6680 21115
rect -6720 20955 -6680 21085
rect -6720 20925 -6715 20955
rect -6685 20925 -6680 20955
rect -6720 20920 -6680 20925
rect -6640 21435 -6600 21440
rect -6640 21405 -6635 21435
rect -6605 21405 -6600 21435
rect -6640 21275 -6600 21405
rect -6640 21245 -6635 21275
rect -6605 21245 -6600 21275
rect -6640 21115 -6600 21245
rect -6640 21085 -6635 21115
rect -6605 21085 -6600 21115
rect -6640 20955 -6600 21085
rect -6640 20925 -6635 20955
rect -6605 20925 -6600 20955
rect -6640 20920 -6600 20925
rect -6560 21435 -6520 21440
rect -6560 21405 -6555 21435
rect -6525 21405 -6520 21435
rect -6560 21275 -6520 21405
rect -6560 21245 -6555 21275
rect -6525 21245 -6520 21275
rect -6560 21115 -6520 21245
rect -6560 21085 -6555 21115
rect -6525 21085 -6520 21115
rect -6560 20955 -6520 21085
rect -6560 20925 -6555 20955
rect -6525 20925 -6520 20955
rect -6560 20920 -6520 20925
rect -6480 21435 -6440 21440
rect -6480 21405 -6475 21435
rect -6445 21405 -6440 21435
rect -6480 21275 -6440 21405
rect -6480 21245 -6475 21275
rect -6445 21245 -6440 21275
rect -6480 21115 -6440 21245
rect -6480 21085 -6475 21115
rect -6445 21085 -6440 21115
rect -6480 20955 -6440 21085
rect -6480 20925 -6475 20955
rect -6445 20925 -6440 20955
rect -6480 20920 -6440 20925
rect -6400 21435 -6360 21440
rect -6400 21405 -6395 21435
rect -6365 21405 -6360 21435
rect -6400 21275 -6360 21405
rect -6400 21245 -6395 21275
rect -6365 21245 -6360 21275
rect -6400 21115 -6360 21245
rect -6400 21085 -6395 21115
rect -6365 21085 -6360 21115
rect -6400 20955 -6360 21085
rect -6400 20925 -6395 20955
rect -6365 20925 -6360 20955
rect -6400 20920 -6360 20925
rect -6320 21435 -6280 21440
rect -6320 21405 -6315 21435
rect -6285 21405 -6280 21435
rect -6320 21275 -6280 21405
rect -6320 21245 -6315 21275
rect -6285 21245 -6280 21275
rect -6320 21115 -6280 21245
rect -6320 21085 -6315 21115
rect -6285 21085 -6280 21115
rect -6320 20955 -6280 21085
rect -6320 20925 -6315 20955
rect -6285 20925 -6280 20955
rect -6320 20920 -6280 20925
rect -6240 21435 -6200 21440
rect -6240 21405 -6235 21435
rect -6205 21405 -6200 21435
rect -6240 21275 -6200 21405
rect -6240 21245 -6235 21275
rect -6205 21245 -6200 21275
rect -6240 21115 -6200 21245
rect -6240 21085 -6235 21115
rect -6205 21085 -6200 21115
rect -6240 20955 -6200 21085
rect -6240 20925 -6235 20955
rect -6205 20925 -6200 20955
rect -6240 20920 -6200 20925
rect -6160 21435 -6120 21440
rect -6160 21405 -6155 21435
rect -6125 21405 -6120 21435
rect -6160 21275 -6120 21405
rect -6160 21245 -6155 21275
rect -6125 21245 -6120 21275
rect -6160 21115 -6120 21245
rect -6160 21085 -6155 21115
rect -6125 21085 -6120 21115
rect -6160 20955 -6120 21085
rect -6160 20925 -6155 20955
rect -6125 20925 -6120 20955
rect -6160 20920 -6120 20925
rect -6080 21435 -6040 21440
rect -6080 21405 -6075 21435
rect -6045 21405 -6040 21435
rect -6080 21275 -6040 21405
rect -5920 21435 -5880 21440
rect -5920 21405 -5915 21435
rect -5885 21405 -5880 21435
rect -6080 21245 -6075 21275
rect -6045 21245 -6040 21275
rect -6080 21115 -6040 21245
rect -6080 21085 -6075 21115
rect -6045 21085 -6040 21115
rect -6080 20955 -6040 21085
rect -6080 20925 -6075 20955
rect -6045 20925 -6040 20955
rect -15040 20844 -15036 20876
rect -15004 20844 -15000 20876
rect -15040 20796 -15000 20844
rect -15040 20764 -15036 20796
rect -15004 20764 -15000 20796
rect -15040 20396 -15000 20764
rect -6080 20875 -6040 20925
rect -6080 20845 -6075 20875
rect -6045 20845 -6040 20875
rect -6080 20795 -6040 20845
rect -6080 20765 -6075 20795
rect -6045 20765 -6040 20795
rect -14960 20675 -14920 20680
rect -14960 20645 -14955 20675
rect -14925 20645 -14920 20675
rect -14960 20515 -14920 20645
rect -14960 20485 -14955 20515
rect -14925 20485 -14920 20515
rect -14960 20480 -14920 20485
rect -14880 20675 -14840 20680
rect -14880 20645 -14875 20675
rect -14845 20645 -14840 20675
rect -14880 20515 -14840 20645
rect -14880 20485 -14875 20515
rect -14845 20485 -14840 20515
rect -14880 20480 -14840 20485
rect -14800 20675 -14760 20680
rect -14800 20645 -14795 20675
rect -14765 20645 -14760 20675
rect -14800 20515 -14760 20645
rect -14800 20485 -14795 20515
rect -14765 20485 -14760 20515
rect -14800 20480 -14760 20485
rect -14720 20675 -14680 20680
rect -14720 20645 -14715 20675
rect -14685 20645 -14680 20675
rect -14720 20515 -14680 20645
rect -14720 20485 -14715 20515
rect -14685 20485 -14680 20515
rect -14720 20480 -14680 20485
rect -14640 20675 -14600 20680
rect -14640 20645 -14635 20675
rect -14605 20645 -14600 20675
rect -14640 20515 -14600 20645
rect -14640 20485 -14635 20515
rect -14605 20485 -14600 20515
rect -14640 20480 -14600 20485
rect -14560 20675 -14520 20680
rect -14560 20645 -14555 20675
rect -14525 20645 -14520 20675
rect -14560 20515 -14520 20645
rect -14560 20485 -14555 20515
rect -14525 20485 -14520 20515
rect -14560 20480 -14520 20485
rect -14480 20675 -14440 20680
rect -14480 20645 -14475 20675
rect -14445 20645 -14440 20675
rect -14480 20515 -14440 20645
rect -14480 20485 -14475 20515
rect -14445 20485 -14440 20515
rect -14480 20480 -14440 20485
rect -14400 20675 -14360 20680
rect -14400 20645 -14395 20675
rect -14365 20645 -14360 20675
rect -14400 20515 -14360 20645
rect -14400 20485 -14395 20515
rect -14365 20485 -14360 20515
rect -14400 20480 -14360 20485
rect -14320 20675 -14280 20680
rect -14320 20645 -14315 20675
rect -14285 20645 -14280 20675
rect -14320 20515 -14280 20645
rect -14320 20485 -14315 20515
rect -14285 20485 -14280 20515
rect -14320 20480 -14280 20485
rect -14240 20675 -14200 20680
rect -14240 20645 -14235 20675
rect -14205 20645 -14200 20675
rect -14240 20515 -14200 20645
rect -14240 20485 -14235 20515
rect -14205 20485 -14200 20515
rect -14240 20480 -14200 20485
rect -14160 20675 -14120 20680
rect -14160 20645 -14155 20675
rect -14125 20645 -14120 20675
rect -14160 20515 -14120 20645
rect -14160 20485 -14155 20515
rect -14125 20485 -14120 20515
rect -14160 20480 -14120 20485
rect -14080 20675 -14040 20680
rect -14080 20645 -14075 20675
rect -14045 20645 -14040 20675
rect -14080 20515 -14040 20645
rect -14080 20485 -14075 20515
rect -14045 20485 -14040 20515
rect -14080 20480 -14040 20485
rect -14000 20675 -13960 20680
rect -14000 20645 -13995 20675
rect -13965 20645 -13960 20675
rect -14000 20515 -13960 20645
rect -14000 20485 -13995 20515
rect -13965 20485 -13960 20515
rect -14000 20480 -13960 20485
rect -13920 20675 -13880 20680
rect -13920 20645 -13915 20675
rect -13885 20645 -13880 20675
rect -13920 20515 -13880 20645
rect -13920 20485 -13915 20515
rect -13885 20485 -13880 20515
rect -13920 20480 -13880 20485
rect -13840 20675 -13800 20680
rect -13840 20645 -13835 20675
rect -13805 20645 -13800 20675
rect -13840 20515 -13800 20645
rect -13840 20485 -13835 20515
rect -13805 20485 -13800 20515
rect -13840 20480 -13800 20485
rect -13760 20675 -13720 20680
rect -13760 20645 -13755 20675
rect -13725 20645 -13720 20675
rect -13760 20515 -13720 20645
rect -13760 20485 -13755 20515
rect -13725 20485 -13720 20515
rect -13760 20480 -13720 20485
rect -13680 20675 -13640 20680
rect -13680 20645 -13675 20675
rect -13645 20645 -13640 20675
rect -13680 20515 -13640 20645
rect -13680 20485 -13675 20515
rect -13645 20485 -13640 20515
rect -13680 20480 -13640 20485
rect -13600 20675 -13560 20680
rect -13600 20645 -13595 20675
rect -13565 20645 -13560 20675
rect -13600 20515 -13560 20645
rect -13600 20485 -13595 20515
rect -13565 20485 -13560 20515
rect -13600 20480 -13560 20485
rect -13520 20675 -13480 20680
rect -13520 20645 -13515 20675
rect -13485 20645 -13480 20675
rect -13520 20515 -13480 20645
rect -13520 20485 -13515 20515
rect -13485 20485 -13480 20515
rect -13520 20480 -13480 20485
rect -13440 20675 -13400 20680
rect -13440 20645 -13435 20675
rect -13405 20645 -13400 20675
rect -13440 20515 -13400 20645
rect -13440 20485 -13435 20515
rect -13405 20485 -13400 20515
rect -13440 20480 -13400 20485
rect -13360 20675 -13320 20680
rect -13360 20645 -13355 20675
rect -13325 20645 -13320 20675
rect -13360 20515 -13320 20645
rect -13360 20485 -13355 20515
rect -13325 20485 -13320 20515
rect -13360 20480 -13320 20485
rect -13280 20675 -13240 20680
rect -13280 20645 -13275 20675
rect -13245 20645 -13240 20675
rect -13280 20515 -13240 20645
rect -13280 20485 -13275 20515
rect -13245 20485 -13240 20515
rect -13280 20480 -13240 20485
rect -13200 20675 -13160 20680
rect -13200 20645 -13195 20675
rect -13165 20645 -13160 20675
rect -13200 20515 -13160 20645
rect -13200 20485 -13195 20515
rect -13165 20485 -13160 20515
rect -13200 20480 -13160 20485
rect -13120 20675 -13080 20680
rect -13120 20645 -13115 20675
rect -13085 20645 -13080 20675
rect -13120 20515 -13080 20645
rect -13120 20485 -13115 20515
rect -13085 20485 -13080 20515
rect -13120 20480 -13080 20485
rect -13040 20675 -13000 20680
rect -13040 20645 -13035 20675
rect -13005 20645 -13000 20675
rect -13040 20515 -13000 20645
rect -13040 20485 -13035 20515
rect -13005 20485 -13000 20515
rect -13040 20480 -13000 20485
rect -12960 20675 -12920 20680
rect -12960 20645 -12955 20675
rect -12925 20645 -12920 20675
rect -12960 20515 -12920 20645
rect -12960 20485 -12955 20515
rect -12925 20485 -12920 20515
rect -12960 20480 -12920 20485
rect -12880 20675 -12840 20680
rect -12880 20645 -12875 20675
rect -12845 20645 -12840 20675
rect -12880 20515 -12840 20645
rect -12880 20485 -12875 20515
rect -12845 20485 -12840 20515
rect -12880 20480 -12840 20485
rect -12800 20675 -12760 20680
rect -12800 20645 -12795 20675
rect -12765 20645 -12760 20675
rect -12800 20515 -12760 20645
rect -12800 20485 -12795 20515
rect -12765 20485 -12760 20515
rect -12800 20480 -12760 20485
rect -12720 20675 -12680 20680
rect -12720 20645 -12715 20675
rect -12685 20645 -12680 20675
rect -12720 20515 -12680 20645
rect -12720 20485 -12715 20515
rect -12685 20485 -12680 20515
rect -12720 20480 -12680 20485
rect -12640 20675 -12600 20680
rect -12640 20645 -12635 20675
rect -12605 20645 -12600 20675
rect -12640 20515 -12600 20645
rect -12640 20485 -12635 20515
rect -12605 20485 -12600 20515
rect -12640 20480 -12600 20485
rect -12560 20675 -12520 20680
rect -12560 20645 -12555 20675
rect -12525 20645 -12520 20675
rect -12560 20515 -12520 20645
rect -12560 20485 -12555 20515
rect -12525 20485 -12520 20515
rect -12560 20480 -12520 20485
rect -12480 20675 -12440 20680
rect -12480 20645 -12475 20675
rect -12445 20645 -12440 20675
rect -12480 20515 -12440 20645
rect -12480 20485 -12475 20515
rect -12445 20485 -12440 20515
rect -12480 20480 -12440 20485
rect -12400 20675 -12360 20680
rect -12400 20645 -12395 20675
rect -12365 20645 -12360 20675
rect -12400 20515 -12360 20645
rect -12400 20485 -12395 20515
rect -12365 20485 -12360 20515
rect -12400 20480 -12360 20485
rect -12320 20675 -12280 20680
rect -12320 20645 -12315 20675
rect -12285 20645 -12280 20675
rect -12320 20515 -12280 20645
rect -12320 20485 -12315 20515
rect -12285 20485 -12280 20515
rect -12320 20480 -12280 20485
rect -12240 20675 -12200 20680
rect -12240 20645 -12235 20675
rect -12205 20645 -12200 20675
rect -12240 20515 -12200 20645
rect -12240 20485 -12235 20515
rect -12205 20485 -12200 20515
rect -12240 20480 -12200 20485
rect -12160 20675 -12120 20680
rect -12160 20645 -12155 20675
rect -12125 20645 -12120 20675
rect -12160 20515 -12120 20645
rect -12160 20485 -12155 20515
rect -12125 20485 -12120 20515
rect -12160 20480 -12120 20485
rect -12080 20675 -12040 20680
rect -12080 20645 -12075 20675
rect -12045 20645 -12040 20675
rect -12080 20515 -12040 20645
rect -12080 20485 -12075 20515
rect -12045 20485 -12040 20515
rect -12080 20480 -12040 20485
rect -12000 20675 -11960 20680
rect -12000 20645 -11995 20675
rect -11965 20645 -11960 20675
rect -12000 20515 -11960 20645
rect -12000 20485 -11995 20515
rect -11965 20485 -11960 20515
rect -12000 20480 -11960 20485
rect -11920 20675 -11880 20680
rect -11920 20645 -11915 20675
rect -11885 20645 -11880 20675
rect -11920 20515 -11880 20645
rect -11920 20485 -11915 20515
rect -11885 20485 -11880 20515
rect -11920 20480 -11880 20485
rect -11840 20675 -11800 20680
rect -11840 20645 -11835 20675
rect -11805 20645 -11800 20675
rect -11840 20515 -11800 20645
rect -11840 20485 -11835 20515
rect -11805 20485 -11800 20515
rect -11840 20480 -11800 20485
rect -11760 20675 -11720 20680
rect -11760 20645 -11755 20675
rect -11725 20645 -11720 20675
rect -11760 20515 -11720 20645
rect -11760 20485 -11755 20515
rect -11725 20485 -11720 20515
rect -11760 20480 -11720 20485
rect -11680 20675 -11640 20680
rect -11680 20645 -11675 20675
rect -11645 20645 -11640 20675
rect -11680 20515 -11640 20645
rect -11680 20485 -11675 20515
rect -11645 20485 -11640 20515
rect -11680 20480 -11640 20485
rect -11600 20675 -11560 20680
rect -11600 20645 -11595 20675
rect -11565 20645 -11560 20675
rect -11600 20515 -11560 20645
rect -11600 20485 -11595 20515
rect -11565 20485 -11560 20515
rect -11600 20480 -11560 20485
rect -11520 20675 -11480 20680
rect -11520 20645 -11515 20675
rect -11485 20645 -11480 20675
rect -11520 20515 -11480 20645
rect -11520 20485 -11515 20515
rect -11485 20485 -11480 20515
rect -11520 20480 -11480 20485
rect -11440 20675 -11400 20680
rect -11440 20645 -11435 20675
rect -11405 20645 -11400 20675
rect -11440 20515 -11400 20645
rect -11440 20485 -11435 20515
rect -11405 20485 -11400 20515
rect -11440 20480 -11400 20485
rect -11360 20675 -11320 20680
rect -11360 20645 -11355 20675
rect -11325 20645 -11320 20675
rect -11360 20515 -11320 20645
rect -11360 20485 -11355 20515
rect -11325 20485 -11320 20515
rect -11360 20480 -11320 20485
rect -11280 20675 -11240 20680
rect -11280 20645 -11275 20675
rect -11245 20645 -11240 20675
rect -11280 20515 -11240 20645
rect -11280 20485 -11275 20515
rect -11245 20485 -11240 20515
rect -11280 20480 -11240 20485
rect -11200 20675 -11160 20680
rect -11200 20645 -11195 20675
rect -11165 20645 -11160 20675
rect -11200 20515 -11160 20645
rect -11200 20485 -11195 20515
rect -11165 20485 -11160 20515
rect -11200 20480 -11160 20485
rect -11120 20675 -11080 20680
rect -11120 20645 -11115 20675
rect -11085 20645 -11080 20675
rect -11120 20515 -11080 20645
rect -11120 20485 -11115 20515
rect -11085 20485 -11080 20515
rect -11120 20480 -11080 20485
rect -11040 20675 -11000 20680
rect -11040 20645 -11035 20675
rect -11005 20645 -11000 20675
rect -11040 20515 -11000 20645
rect -11040 20485 -11035 20515
rect -11005 20485 -11000 20515
rect -11040 20480 -11000 20485
rect -10960 20675 -10920 20680
rect -10960 20645 -10955 20675
rect -10925 20645 -10920 20675
rect -10960 20515 -10920 20645
rect -10960 20485 -10955 20515
rect -10925 20485 -10920 20515
rect -10960 20480 -10920 20485
rect -10880 20675 -10840 20680
rect -10880 20645 -10875 20675
rect -10845 20645 -10840 20675
rect -10880 20515 -10840 20645
rect -10880 20485 -10875 20515
rect -10845 20485 -10840 20515
rect -10880 20480 -10840 20485
rect -10800 20675 -10760 20680
rect -10800 20645 -10795 20675
rect -10765 20645 -10760 20675
rect -10800 20515 -10760 20645
rect -10800 20485 -10795 20515
rect -10765 20485 -10760 20515
rect -10800 20480 -10760 20485
rect -10720 20675 -10680 20680
rect -10720 20645 -10715 20675
rect -10685 20645 -10680 20675
rect -10720 20515 -10680 20645
rect -10720 20485 -10715 20515
rect -10685 20485 -10680 20515
rect -10720 20480 -10680 20485
rect -10640 20675 -10600 20680
rect -10640 20645 -10635 20675
rect -10605 20645 -10600 20675
rect -10640 20515 -10600 20645
rect -10640 20485 -10635 20515
rect -10605 20485 -10600 20515
rect -10640 20480 -10600 20485
rect -10560 20675 -10520 20680
rect -10560 20645 -10555 20675
rect -10525 20645 -10520 20675
rect -10560 20515 -10520 20645
rect -10560 20485 -10555 20515
rect -10525 20485 -10520 20515
rect -10560 20480 -10520 20485
rect -10480 20675 -10440 20680
rect -10480 20645 -10475 20675
rect -10445 20645 -10440 20675
rect -10480 20515 -10440 20645
rect -10480 20485 -10475 20515
rect -10445 20485 -10440 20515
rect -10480 20480 -10440 20485
rect -10400 20675 -10360 20680
rect -10400 20645 -10395 20675
rect -10365 20645 -10360 20675
rect -10400 20515 -10360 20645
rect -10400 20485 -10395 20515
rect -10365 20485 -10360 20515
rect -10400 20480 -10360 20485
rect -10320 20675 -10280 20680
rect -10320 20645 -10315 20675
rect -10285 20645 -10280 20675
rect -10320 20515 -10280 20645
rect -10320 20485 -10315 20515
rect -10285 20485 -10280 20515
rect -10320 20480 -10280 20485
rect -10240 20675 -10200 20680
rect -10240 20645 -10235 20675
rect -10205 20645 -10200 20675
rect -10240 20515 -10200 20645
rect -10240 20485 -10235 20515
rect -10205 20485 -10200 20515
rect -10240 20480 -10200 20485
rect -10160 20675 -10120 20680
rect -10160 20645 -10155 20675
rect -10125 20645 -10120 20675
rect -10160 20515 -10120 20645
rect -10160 20485 -10155 20515
rect -10125 20485 -10120 20515
rect -10160 20480 -10120 20485
rect -10080 20675 -10040 20680
rect -10080 20645 -10075 20675
rect -10045 20645 -10040 20675
rect -10080 20515 -10040 20645
rect -10080 20485 -10075 20515
rect -10045 20485 -10040 20515
rect -10080 20480 -10040 20485
rect -10000 20675 -9960 20680
rect -10000 20645 -9995 20675
rect -9965 20645 -9960 20675
rect -10000 20515 -9960 20645
rect -10000 20485 -9995 20515
rect -9965 20485 -9960 20515
rect -10000 20480 -9960 20485
rect -9920 20675 -9880 20680
rect -9920 20645 -9915 20675
rect -9885 20645 -9880 20675
rect -9920 20515 -9880 20645
rect -9920 20485 -9915 20515
rect -9885 20485 -9880 20515
rect -9920 20480 -9880 20485
rect -9840 20675 -9800 20680
rect -9840 20645 -9835 20675
rect -9805 20645 -9800 20675
rect -9840 20515 -9800 20645
rect -9840 20485 -9835 20515
rect -9805 20485 -9800 20515
rect -9840 20480 -9800 20485
rect -9760 20675 -9720 20680
rect -9760 20645 -9755 20675
rect -9725 20645 -9720 20675
rect -9760 20515 -9720 20645
rect -9760 20485 -9755 20515
rect -9725 20485 -9720 20515
rect -9760 20480 -9720 20485
rect -9680 20675 -9640 20680
rect -9680 20645 -9675 20675
rect -9645 20645 -9640 20675
rect -9680 20515 -9640 20645
rect -9680 20485 -9675 20515
rect -9645 20485 -9640 20515
rect -9680 20480 -9640 20485
rect -9600 20675 -9560 20680
rect -9600 20645 -9595 20675
rect -9565 20645 -9560 20675
rect -9600 20515 -9560 20645
rect -9600 20485 -9595 20515
rect -9565 20485 -9560 20515
rect -9600 20480 -9560 20485
rect -9520 20675 -9480 20680
rect -9520 20645 -9515 20675
rect -9485 20645 -9480 20675
rect -9520 20515 -9480 20645
rect -9520 20485 -9515 20515
rect -9485 20485 -9480 20515
rect -9520 20480 -9480 20485
rect -9440 20675 -9400 20680
rect -9440 20645 -9435 20675
rect -9405 20645 -9400 20675
rect -9440 20515 -9400 20645
rect -9440 20485 -9435 20515
rect -9405 20485 -9400 20515
rect -9440 20480 -9400 20485
rect -9360 20675 -9320 20680
rect -9360 20645 -9355 20675
rect -9325 20645 -9320 20675
rect -9360 20515 -9320 20645
rect -9360 20485 -9355 20515
rect -9325 20485 -9320 20515
rect -9360 20480 -9320 20485
rect -9280 20675 -9240 20680
rect -9280 20645 -9275 20675
rect -9245 20645 -9240 20675
rect -9280 20515 -9240 20645
rect -9280 20485 -9275 20515
rect -9245 20485 -9240 20515
rect -9280 20480 -9240 20485
rect -9200 20675 -9160 20680
rect -9200 20645 -9195 20675
rect -9165 20645 -9160 20675
rect -9200 20515 -9160 20645
rect -9200 20485 -9195 20515
rect -9165 20485 -9160 20515
rect -9200 20480 -9160 20485
rect -9120 20675 -9080 20680
rect -9120 20645 -9115 20675
rect -9085 20645 -9080 20675
rect -9120 20515 -9080 20645
rect -9120 20485 -9115 20515
rect -9085 20485 -9080 20515
rect -9120 20480 -9080 20485
rect -9040 20675 -9000 20680
rect -9040 20645 -9035 20675
rect -9005 20645 -9000 20675
rect -9040 20515 -9000 20645
rect -9040 20485 -9035 20515
rect -9005 20485 -9000 20515
rect -9040 20480 -9000 20485
rect -8960 20675 -8920 20680
rect -8960 20645 -8955 20675
rect -8925 20645 -8920 20675
rect -8960 20515 -8920 20645
rect -8960 20485 -8955 20515
rect -8925 20485 -8920 20515
rect -8960 20480 -8920 20485
rect -8880 20675 -8840 20680
rect -8880 20645 -8875 20675
rect -8845 20645 -8840 20675
rect -8880 20515 -8840 20645
rect -8880 20485 -8875 20515
rect -8845 20485 -8840 20515
rect -8880 20480 -8840 20485
rect -8800 20675 -8760 20680
rect -8800 20645 -8795 20675
rect -8765 20645 -8760 20675
rect -8800 20515 -8760 20645
rect -8800 20485 -8795 20515
rect -8765 20485 -8760 20515
rect -8800 20480 -8760 20485
rect -8720 20675 -8680 20680
rect -8720 20645 -8715 20675
rect -8685 20645 -8680 20675
rect -8720 20515 -8680 20645
rect -8720 20485 -8715 20515
rect -8685 20485 -8680 20515
rect -8720 20480 -8680 20485
rect -8640 20675 -8600 20680
rect -8640 20645 -8635 20675
rect -8605 20645 -8600 20675
rect -8640 20515 -8600 20645
rect -8640 20485 -8635 20515
rect -8605 20485 -8600 20515
rect -8640 20480 -8600 20485
rect -8560 20675 -8520 20680
rect -8560 20645 -8555 20675
rect -8525 20645 -8520 20675
rect -8560 20515 -8520 20645
rect -8560 20485 -8555 20515
rect -8525 20485 -8520 20515
rect -8560 20480 -8520 20485
rect -8480 20675 -8440 20680
rect -8480 20645 -8475 20675
rect -8445 20645 -8440 20675
rect -8480 20515 -8440 20645
rect -8480 20485 -8475 20515
rect -8445 20485 -8440 20515
rect -8480 20480 -8440 20485
rect -8400 20675 -8360 20680
rect -8400 20645 -8395 20675
rect -8365 20645 -8360 20675
rect -8400 20515 -8360 20645
rect -8400 20485 -8395 20515
rect -8365 20485 -8360 20515
rect -8400 20480 -8360 20485
rect -8320 20675 -8280 20680
rect -8320 20645 -8315 20675
rect -8285 20645 -8280 20675
rect -8320 20515 -8280 20645
rect -8320 20485 -8315 20515
rect -8285 20485 -8280 20515
rect -8320 20480 -8280 20485
rect -8240 20675 -8200 20680
rect -8240 20645 -8235 20675
rect -8205 20645 -8200 20675
rect -8240 20515 -8200 20645
rect -8240 20485 -8235 20515
rect -8205 20485 -8200 20515
rect -8240 20480 -8200 20485
rect -8160 20675 -8120 20680
rect -8160 20645 -8155 20675
rect -8125 20645 -8120 20675
rect -8160 20515 -8120 20645
rect -8160 20485 -8155 20515
rect -8125 20485 -8120 20515
rect -8160 20480 -8120 20485
rect -8080 20675 -8040 20680
rect -8080 20645 -8075 20675
rect -8045 20645 -8040 20675
rect -8080 20515 -8040 20645
rect -8080 20485 -8075 20515
rect -8045 20485 -8040 20515
rect -8080 20480 -8040 20485
rect -8000 20675 -7960 20680
rect -8000 20645 -7995 20675
rect -7965 20645 -7960 20675
rect -8000 20515 -7960 20645
rect -8000 20485 -7995 20515
rect -7965 20485 -7960 20515
rect -8000 20480 -7960 20485
rect -7920 20675 -7880 20680
rect -7920 20645 -7915 20675
rect -7885 20645 -7880 20675
rect -7920 20515 -7880 20645
rect -7920 20485 -7915 20515
rect -7885 20485 -7880 20515
rect -7920 20480 -7880 20485
rect -7840 20675 -7800 20680
rect -7840 20645 -7835 20675
rect -7805 20645 -7800 20675
rect -7840 20515 -7800 20645
rect -7840 20485 -7835 20515
rect -7805 20485 -7800 20515
rect -7840 20480 -7800 20485
rect -7760 20675 -7720 20680
rect -7760 20645 -7755 20675
rect -7725 20645 -7720 20675
rect -7760 20515 -7720 20645
rect -7760 20485 -7755 20515
rect -7725 20485 -7720 20515
rect -7760 20480 -7720 20485
rect -7680 20675 -7640 20680
rect -7680 20645 -7675 20675
rect -7645 20645 -7640 20675
rect -7680 20515 -7640 20645
rect -7680 20485 -7675 20515
rect -7645 20485 -7640 20515
rect -7680 20480 -7640 20485
rect -7600 20675 -7560 20680
rect -7600 20645 -7595 20675
rect -7565 20645 -7560 20675
rect -7600 20515 -7560 20645
rect -7600 20485 -7595 20515
rect -7565 20485 -7560 20515
rect -7600 20480 -7560 20485
rect -7520 20675 -7480 20680
rect -7520 20645 -7515 20675
rect -7485 20645 -7480 20675
rect -7520 20515 -7480 20645
rect -7520 20485 -7515 20515
rect -7485 20485 -7480 20515
rect -7520 20480 -7480 20485
rect -7440 20675 -7400 20680
rect -7440 20645 -7435 20675
rect -7405 20645 -7400 20675
rect -7440 20515 -7400 20645
rect -7440 20485 -7435 20515
rect -7405 20485 -7400 20515
rect -7440 20480 -7400 20485
rect -7360 20675 -7320 20680
rect -7360 20645 -7355 20675
rect -7325 20645 -7320 20675
rect -7360 20515 -7320 20645
rect -7360 20485 -7355 20515
rect -7325 20485 -7320 20515
rect -7360 20480 -7320 20485
rect -7280 20675 -7240 20680
rect -7280 20645 -7275 20675
rect -7245 20645 -7240 20675
rect -7280 20515 -7240 20645
rect -7280 20485 -7275 20515
rect -7245 20485 -7240 20515
rect -7280 20480 -7240 20485
rect -7200 20675 -7160 20680
rect -7200 20645 -7195 20675
rect -7165 20645 -7160 20675
rect -7200 20515 -7160 20645
rect -7200 20485 -7195 20515
rect -7165 20485 -7160 20515
rect -7200 20480 -7160 20485
rect -7120 20675 -7080 20680
rect -7120 20645 -7115 20675
rect -7085 20645 -7080 20675
rect -7120 20515 -7080 20645
rect -7120 20485 -7115 20515
rect -7085 20485 -7080 20515
rect -7120 20480 -7080 20485
rect -7040 20675 -7000 20680
rect -7040 20645 -7035 20675
rect -7005 20645 -7000 20675
rect -7040 20515 -7000 20645
rect -7040 20485 -7035 20515
rect -7005 20485 -7000 20515
rect -7040 20480 -7000 20485
rect -6960 20675 -6920 20680
rect -6960 20645 -6955 20675
rect -6925 20645 -6920 20675
rect -6960 20515 -6920 20645
rect -6960 20485 -6955 20515
rect -6925 20485 -6920 20515
rect -6960 20480 -6920 20485
rect -6880 20675 -6840 20680
rect -6880 20645 -6875 20675
rect -6845 20645 -6840 20675
rect -6880 20515 -6840 20645
rect -6880 20485 -6875 20515
rect -6845 20485 -6840 20515
rect -6880 20480 -6840 20485
rect -6800 20675 -6760 20680
rect -6800 20645 -6795 20675
rect -6765 20645 -6760 20675
rect -6800 20515 -6760 20645
rect -6800 20485 -6795 20515
rect -6765 20485 -6760 20515
rect -6800 20480 -6760 20485
rect -6720 20675 -6680 20680
rect -6720 20645 -6715 20675
rect -6685 20645 -6680 20675
rect -6720 20515 -6680 20645
rect -6720 20485 -6715 20515
rect -6685 20485 -6680 20515
rect -6720 20480 -6680 20485
rect -6640 20675 -6600 20680
rect -6640 20645 -6635 20675
rect -6605 20645 -6600 20675
rect -6640 20515 -6600 20645
rect -6640 20485 -6635 20515
rect -6605 20485 -6600 20515
rect -6640 20480 -6600 20485
rect -6560 20675 -6520 20680
rect -6560 20645 -6555 20675
rect -6525 20645 -6520 20675
rect -6560 20515 -6520 20645
rect -6560 20485 -6555 20515
rect -6525 20485 -6520 20515
rect -6560 20480 -6520 20485
rect -6480 20675 -6440 20680
rect -6480 20645 -6475 20675
rect -6445 20645 -6440 20675
rect -6480 20515 -6440 20645
rect -6480 20485 -6475 20515
rect -6445 20485 -6440 20515
rect -6480 20480 -6440 20485
rect -6400 20675 -6360 20680
rect -6400 20645 -6395 20675
rect -6365 20645 -6360 20675
rect -6400 20515 -6360 20645
rect -6400 20485 -6395 20515
rect -6365 20485 -6360 20515
rect -6400 20480 -6360 20485
rect -6320 20675 -6280 20680
rect -6320 20645 -6315 20675
rect -6285 20645 -6280 20675
rect -6320 20515 -6280 20645
rect -6320 20485 -6315 20515
rect -6285 20485 -6280 20515
rect -6320 20480 -6280 20485
rect -6240 20675 -6200 20680
rect -6240 20645 -6235 20675
rect -6205 20645 -6200 20675
rect -6240 20515 -6200 20645
rect -6240 20485 -6235 20515
rect -6205 20485 -6200 20515
rect -6240 20480 -6200 20485
rect -6160 20675 -6120 20680
rect -6160 20645 -6155 20675
rect -6125 20645 -6120 20675
rect -6160 20515 -6120 20645
rect -6160 20485 -6155 20515
rect -6125 20485 -6120 20515
rect -6160 20480 -6120 20485
rect -15040 20364 -15036 20396
rect -15004 20364 -15000 20396
rect -15040 20316 -15000 20364
rect -15040 20284 -15036 20316
rect -15004 20284 -15000 20316
rect -15040 20236 -15000 20284
rect -15040 20204 -15036 20236
rect -15004 20204 -15000 20236
rect -15040 20156 -15000 20204
rect -6080 20435 -6040 20765
rect -6080 20405 -6075 20435
rect -6045 20405 -6040 20435
rect -6080 20355 -6040 20405
rect -6080 20325 -6075 20355
rect -6045 20325 -6040 20355
rect -6080 20195 -6040 20325
rect -6080 20165 -6075 20195
rect -6045 20165 -6040 20195
rect -6080 20160 -6040 20165
rect -6000 21355 -5960 21360
rect -6000 21325 -5995 21355
rect -5965 21325 -5960 21355
rect -15040 20124 -15036 20156
rect -15004 20124 -15000 20156
rect -15040 20076 -15000 20124
rect -15040 20044 -15036 20076
rect -15004 20044 -15000 20076
rect -15040 19996 -15000 20044
rect -15040 19964 -15036 19996
rect -15004 19964 -15000 19996
rect -15040 19916 -15000 19964
rect -6000 19960 -5960 21325
rect -5920 21275 -5880 21405
rect -5920 21245 -5915 21275
rect -5885 21245 -5880 21275
rect -5920 21115 -5880 21245
rect -5760 21435 -5720 21440
rect -5760 21405 -5755 21435
rect -5725 21405 -5720 21435
rect -5760 21275 -5720 21405
rect -5760 21245 -5755 21275
rect -5725 21245 -5720 21275
rect -5920 21085 -5915 21115
rect -5885 21085 -5880 21115
rect -5920 20955 -5880 21085
rect -5920 20925 -5915 20955
rect -5885 20925 -5880 20955
rect -5920 20875 -5880 20925
rect -5920 20845 -5915 20875
rect -5885 20845 -5880 20875
rect -5920 20795 -5880 20845
rect -5920 20765 -5915 20795
rect -5885 20765 -5880 20795
rect -5920 20435 -5880 20765
rect -5920 20405 -5915 20435
rect -5885 20405 -5880 20435
rect -5920 20355 -5880 20405
rect -5920 20325 -5915 20355
rect -5885 20325 -5880 20355
rect -5920 20195 -5880 20325
rect -5920 20165 -5915 20195
rect -5885 20165 -5880 20195
rect -5920 20160 -5880 20165
rect -5840 21195 -5800 21200
rect -5840 21165 -5835 21195
rect -5805 21165 -5800 21195
rect -5840 19960 -5800 21165
rect -5760 21115 -5720 21245
rect -5760 21085 -5755 21115
rect -5725 21085 -5720 21115
rect -5760 20955 -5720 21085
rect -5760 20925 -5755 20955
rect -5725 20925 -5720 20955
rect -5760 20875 -5720 20925
rect -5680 21435 -5640 21440
rect -5680 21405 -5675 21435
rect -5645 21405 -5640 21435
rect -5680 21275 -5640 21405
rect -5680 21245 -5675 21275
rect -5645 21245 -5640 21275
rect -5680 21115 -5640 21245
rect -5680 21085 -5675 21115
rect -5645 21085 -5640 21115
rect -5680 20955 -5640 21085
rect -5680 20925 -5675 20955
rect -5645 20925 -5640 20955
rect -5680 20920 -5640 20925
rect -5600 21435 -5560 21440
rect -5600 21405 -5595 21435
rect -5565 21405 -5560 21435
rect -5600 21275 -5560 21405
rect -5600 21245 -5595 21275
rect -5565 21245 -5560 21275
rect -5600 21115 -5560 21245
rect -5600 21085 -5595 21115
rect -5565 21085 -5560 21115
rect -5600 20955 -5560 21085
rect -5600 20925 -5595 20955
rect -5565 20925 -5560 20955
rect -5600 20920 -5560 20925
rect -5520 21435 -5480 21440
rect -5520 21405 -5515 21435
rect -5485 21405 -5480 21435
rect -5520 21275 -5480 21405
rect -5520 21245 -5515 21275
rect -5485 21245 -5480 21275
rect -5520 21115 -5480 21245
rect -5520 21085 -5515 21115
rect -5485 21085 -5480 21115
rect -5520 20955 -5480 21085
rect -5520 20925 -5515 20955
rect -5485 20925 -5480 20955
rect -5520 20920 -5480 20925
rect -5440 21435 -5400 21440
rect -5440 21405 -5435 21435
rect -5405 21405 -5400 21435
rect -5440 21275 -5400 21405
rect -5440 21245 -5435 21275
rect -5405 21245 -5400 21275
rect -5440 21115 -5400 21245
rect -5440 21085 -5435 21115
rect -5405 21085 -5400 21115
rect -5440 20955 -5400 21085
rect -5440 20925 -5435 20955
rect -5405 20925 -5400 20955
rect -5440 20920 -5400 20925
rect -5360 21435 -5320 21440
rect -5360 21405 -5355 21435
rect -5325 21405 -5320 21435
rect -5360 21275 -5320 21405
rect -5360 21245 -5355 21275
rect -5325 21245 -5320 21275
rect -5360 21115 -5320 21245
rect -5360 21085 -5355 21115
rect -5325 21085 -5320 21115
rect -5360 20955 -5320 21085
rect -5360 20925 -5355 20955
rect -5325 20925 -5320 20955
rect -5360 20920 -5320 20925
rect -5280 21435 -5240 21440
rect -5280 21405 -5275 21435
rect -5245 21405 -5240 21435
rect -5280 21275 -5240 21405
rect -5280 21245 -5275 21275
rect -5245 21245 -5240 21275
rect -5280 21115 -5240 21245
rect -5280 21085 -5275 21115
rect -5245 21085 -5240 21115
rect -5280 20955 -5240 21085
rect -5280 20925 -5275 20955
rect -5245 20925 -5240 20955
rect -5280 20920 -5240 20925
rect -5200 21435 -5160 21440
rect -5200 21405 -5195 21435
rect -5165 21405 -5160 21435
rect -5200 21275 -5160 21405
rect -5200 21245 -5195 21275
rect -5165 21245 -5160 21275
rect -5200 21115 -5160 21245
rect -5200 21085 -5195 21115
rect -5165 21085 -5160 21115
rect -5200 20955 -5160 21085
rect -5200 20925 -5195 20955
rect -5165 20925 -5160 20955
rect -5200 20920 -5160 20925
rect -5120 21435 -5080 21440
rect -5120 21405 -5115 21435
rect -5085 21405 -5080 21435
rect -5120 21275 -5080 21405
rect -5120 21245 -5115 21275
rect -5085 21245 -5080 21275
rect -5120 21115 -5080 21245
rect -5120 21085 -5115 21115
rect -5085 21085 -5080 21115
rect -5120 20955 -5080 21085
rect -5120 20925 -5115 20955
rect -5085 20925 -5080 20955
rect -5120 20920 -5080 20925
rect -5040 21435 -5000 21440
rect -5040 21405 -5035 21435
rect -5005 21405 -5000 21435
rect -5040 21275 -5000 21405
rect -5040 21245 -5035 21275
rect -5005 21245 -5000 21275
rect -5040 21115 -5000 21245
rect -5040 21085 -5035 21115
rect -5005 21085 -5000 21115
rect -5040 20955 -5000 21085
rect -5040 20925 -5035 20955
rect -5005 20925 -5000 20955
rect -5040 20920 -5000 20925
rect -4960 21435 -4920 21440
rect -4960 21405 -4955 21435
rect -4925 21405 -4920 21435
rect -4960 21275 -4920 21405
rect -4960 21245 -4955 21275
rect -4925 21245 -4920 21275
rect -4960 21115 -4920 21245
rect -4960 21085 -4955 21115
rect -4925 21085 -4920 21115
rect -4960 20955 -4920 21085
rect -4960 20925 -4955 20955
rect -4925 20925 -4920 20955
rect -4960 20920 -4920 20925
rect -4880 21435 -4840 21440
rect -4880 21405 -4875 21435
rect -4845 21405 -4840 21435
rect -4880 21275 -4840 21405
rect -4880 21245 -4875 21275
rect -4845 21245 -4840 21275
rect -4880 21115 -4840 21245
rect -4880 21085 -4875 21115
rect -4845 21085 -4840 21115
rect -4880 20955 -4840 21085
rect -4880 20925 -4875 20955
rect -4845 20925 -4840 20955
rect -4880 20920 -4840 20925
rect -4800 21435 -4760 21440
rect -4800 21405 -4795 21435
rect -4765 21405 -4760 21435
rect -4800 21275 -4760 21405
rect -4800 21245 -4795 21275
rect -4765 21245 -4760 21275
rect -4800 21115 -4760 21245
rect -4800 21085 -4795 21115
rect -4765 21085 -4760 21115
rect -4800 20955 -4760 21085
rect -4800 20925 -4795 20955
rect -4765 20925 -4760 20955
rect -4800 20920 -4760 20925
rect -4720 21435 -4680 21440
rect -4720 21405 -4715 21435
rect -4685 21405 -4680 21435
rect -4720 21275 -4680 21405
rect -4720 21245 -4715 21275
rect -4685 21245 -4680 21275
rect -4720 21115 -4680 21245
rect -4720 21085 -4715 21115
rect -4685 21085 -4680 21115
rect -4720 20955 -4680 21085
rect -4720 20925 -4715 20955
rect -4685 20925 -4680 20955
rect -4720 20920 -4680 20925
rect -4640 21435 -4600 21440
rect -4640 21405 -4635 21435
rect -4605 21405 -4600 21435
rect -4640 21275 -4600 21405
rect -4640 21245 -4635 21275
rect -4605 21245 -4600 21275
rect -4640 21115 -4600 21245
rect -4640 21085 -4635 21115
rect -4605 21085 -4600 21115
rect -4640 20955 -4600 21085
rect -4640 20925 -4635 20955
rect -4605 20925 -4600 20955
rect -4640 20920 -4600 20925
rect -4560 21435 -4520 21440
rect -4560 21405 -4555 21435
rect -4525 21405 -4520 21435
rect -4560 21275 -4520 21405
rect -4560 21245 -4555 21275
rect -4525 21245 -4520 21275
rect -4560 21115 -4520 21245
rect -4560 21085 -4555 21115
rect -4525 21085 -4520 21115
rect -4560 20955 -4520 21085
rect -4560 20925 -4555 20955
rect -4525 20925 -4520 20955
rect -4560 20920 -4520 20925
rect -4480 21435 -4440 21440
rect -4480 21405 -4475 21435
rect -4445 21405 -4440 21435
rect -4480 21275 -4440 21405
rect -4480 21245 -4475 21275
rect -4445 21245 -4440 21275
rect -4480 21115 -4440 21245
rect -4480 21085 -4475 21115
rect -4445 21085 -4440 21115
rect -4480 20955 -4440 21085
rect -4480 20925 -4475 20955
rect -4445 20925 -4440 20955
rect -4480 20920 -4440 20925
rect -4400 21435 -4360 21440
rect -4400 21405 -4395 21435
rect -4365 21405 -4360 21435
rect -4400 21275 -4360 21405
rect -4400 21245 -4395 21275
rect -4365 21245 -4360 21275
rect -4400 21115 -4360 21245
rect -4400 21085 -4395 21115
rect -4365 21085 -4360 21115
rect -4400 20955 -4360 21085
rect -4400 20925 -4395 20955
rect -4365 20925 -4360 20955
rect -4400 20920 -4360 20925
rect -4320 21435 -4280 21440
rect -4320 21405 -4315 21435
rect -4285 21405 -4280 21435
rect -4320 21275 -4280 21405
rect -4320 21245 -4315 21275
rect -4285 21245 -4280 21275
rect -4320 21115 -4280 21245
rect -4320 21085 -4315 21115
rect -4285 21085 -4280 21115
rect -4320 20955 -4280 21085
rect -4320 20925 -4315 20955
rect -4285 20925 -4280 20955
rect -4320 20920 -4280 20925
rect -4240 21435 -4200 21440
rect -4240 21405 -4235 21435
rect -4205 21405 -4200 21435
rect -4240 21275 -4200 21405
rect -4240 21245 -4235 21275
rect -4205 21245 -4200 21275
rect -4240 21115 -4200 21245
rect -4240 21085 -4235 21115
rect -4205 21085 -4200 21115
rect -4240 20955 -4200 21085
rect -4240 20925 -4235 20955
rect -4205 20925 -4200 20955
rect -4240 20920 -4200 20925
rect -4160 21435 -4120 21440
rect -4160 21405 -4155 21435
rect -4125 21405 -4120 21435
rect -4160 21275 -4120 21405
rect -4160 21245 -4155 21275
rect -4125 21245 -4120 21275
rect -4160 21115 -4120 21245
rect -4160 21085 -4155 21115
rect -4125 21085 -4120 21115
rect -4160 20955 -4120 21085
rect -4160 20925 -4155 20955
rect -4125 20925 -4120 20955
rect -4160 20920 -4120 20925
rect -4080 21435 -4040 21440
rect -4080 21405 -4075 21435
rect -4045 21405 -4040 21435
rect -4080 21275 -4040 21405
rect -4080 21245 -4075 21275
rect -4045 21245 -4040 21275
rect -4080 21115 -4040 21245
rect -4080 21085 -4075 21115
rect -4045 21085 -4040 21115
rect -4080 20955 -4040 21085
rect -4080 20925 -4075 20955
rect -4045 20925 -4040 20955
rect -4080 20920 -4040 20925
rect -4000 21435 -3960 21440
rect -4000 21405 -3995 21435
rect -3965 21405 -3960 21435
rect -4000 21275 -3960 21405
rect -4000 21245 -3995 21275
rect -3965 21245 -3960 21275
rect -4000 21115 -3960 21245
rect -4000 21085 -3995 21115
rect -3965 21085 -3960 21115
rect -4000 20955 -3960 21085
rect -4000 20925 -3995 20955
rect -3965 20925 -3960 20955
rect -4000 20920 -3960 20925
rect -3920 21435 -3880 21440
rect -3920 21405 -3915 21435
rect -3885 21405 -3880 21435
rect -3920 21275 -3880 21405
rect -3920 21245 -3915 21275
rect -3885 21245 -3880 21275
rect -3920 21115 -3880 21245
rect -3920 21085 -3915 21115
rect -3885 21085 -3880 21115
rect -3920 20955 -3880 21085
rect -3920 20925 -3915 20955
rect -3885 20925 -3880 20955
rect -3920 20920 -3880 20925
rect -3840 21435 -3800 21440
rect -3840 21405 -3835 21435
rect -3805 21405 -3800 21435
rect -3840 21275 -3800 21405
rect -3840 21245 -3835 21275
rect -3805 21245 -3800 21275
rect -3840 21115 -3800 21245
rect -3840 21085 -3835 21115
rect -3805 21085 -3800 21115
rect -3840 20955 -3800 21085
rect -3840 20925 -3835 20955
rect -3805 20925 -3800 20955
rect -3840 20920 -3800 20925
rect -3760 21435 -3720 21440
rect -3760 21405 -3755 21435
rect -3725 21405 -3720 21435
rect -3760 21275 -3720 21405
rect -3760 21245 -3755 21275
rect -3725 21245 -3720 21275
rect -3760 21115 -3720 21245
rect -3760 21085 -3755 21115
rect -3725 21085 -3720 21115
rect -3760 20955 -3720 21085
rect -3760 20925 -3755 20955
rect -3725 20925 -3720 20955
rect -3760 20920 -3720 20925
rect -3680 21435 -3640 21440
rect -3680 21405 -3675 21435
rect -3645 21405 -3640 21435
rect -3680 21275 -3640 21405
rect -3680 21245 -3675 21275
rect -3645 21245 -3640 21275
rect -3680 21115 -3640 21245
rect -3680 21085 -3675 21115
rect -3645 21085 -3640 21115
rect -3680 20955 -3640 21085
rect -3680 20925 -3675 20955
rect -3645 20925 -3640 20955
rect -3680 20920 -3640 20925
rect -3600 21435 -3560 21440
rect -3600 21405 -3595 21435
rect -3565 21405 -3560 21435
rect -3600 21275 -3560 21405
rect -3600 21245 -3595 21275
rect -3565 21245 -3560 21275
rect -3600 21115 -3560 21245
rect -3600 21085 -3595 21115
rect -3565 21085 -3560 21115
rect -3600 20955 -3560 21085
rect -3600 20925 -3595 20955
rect -3565 20925 -3560 20955
rect -3600 20920 -3560 20925
rect -3520 21435 -3480 21440
rect -3520 21405 -3515 21435
rect -3485 21405 -3480 21435
rect -3520 21275 -3480 21405
rect -3520 21245 -3515 21275
rect -3485 21245 -3480 21275
rect -3520 21115 -3480 21245
rect -3520 21085 -3515 21115
rect -3485 21085 -3480 21115
rect -3520 20955 -3480 21085
rect -3520 20925 -3515 20955
rect -3485 20925 -3480 20955
rect -3520 20920 -3480 20925
rect -3440 21435 -3400 21440
rect -3440 21405 -3435 21435
rect -3405 21405 -3400 21435
rect -3440 21275 -3400 21405
rect -3440 21245 -3435 21275
rect -3405 21245 -3400 21275
rect -3440 21115 -3400 21245
rect -3440 21085 -3435 21115
rect -3405 21085 -3400 21115
rect -3440 20955 -3400 21085
rect -3440 20925 -3435 20955
rect -3405 20925 -3400 20955
rect -3440 20920 -3400 20925
rect -3360 21435 -3320 21440
rect -3360 21405 -3355 21435
rect -3325 21405 -3320 21435
rect -3360 21275 -3320 21405
rect -3360 21245 -3355 21275
rect -3325 21245 -3320 21275
rect -3360 21115 -3320 21245
rect -3360 21085 -3355 21115
rect -3325 21085 -3320 21115
rect -3360 20955 -3320 21085
rect -3360 20925 -3355 20955
rect -3325 20925 -3320 20955
rect -3360 20920 -3320 20925
rect -3280 21435 -3240 21440
rect -3280 21405 -3275 21435
rect -3245 21405 -3240 21435
rect -3280 21275 -3240 21405
rect -3280 21245 -3275 21275
rect -3245 21245 -3240 21275
rect -3280 21115 -3240 21245
rect -3280 21085 -3275 21115
rect -3245 21085 -3240 21115
rect -3280 20955 -3240 21085
rect -3280 20925 -3275 20955
rect -3245 20925 -3240 20955
rect -3280 20920 -3240 20925
rect -3200 21435 -3160 21440
rect -3200 21405 -3195 21435
rect -3165 21405 -3160 21435
rect -3200 21275 -3160 21405
rect -3200 21245 -3195 21275
rect -3165 21245 -3160 21275
rect -3200 21115 -3160 21245
rect -3200 21085 -3195 21115
rect -3165 21085 -3160 21115
rect -3200 20955 -3160 21085
rect -3200 20925 -3195 20955
rect -3165 20925 -3160 20955
rect -3200 20920 -3160 20925
rect -3120 21435 -3080 21440
rect -3120 21405 -3115 21435
rect -3085 21405 -3080 21435
rect -3120 21275 -3080 21405
rect -3120 21245 -3115 21275
rect -3085 21245 -3080 21275
rect -3120 21115 -3080 21245
rect -3120 21085 -3115 21115
rect -3085 21085 -3080 21115
rect -3120 20955 -3080 21085
rect -3120 20925 -3115 20955
rect -3085 20925 -3080 20955
rect -3120 20920 -3080 20925
rect -3040 21435 -3000 21440
rect -3040 21405 -3035 21435
rect -3005 21405 -3000 21435
rect -3040 21275 -3000 21405
rect -3040 21245 -3035 21275
rect -3005 21245 -3000 21275
rect -3040 21115 -3000 21245
rect -3040 21085 -3035 21115
rect -3005 21085 -3000 21115
rect -3040 20955 -3000 21085
rect -3040 20925 -3035 20955
rect -3005 20925 -3000 20955
rect -3040 20920 -3000 20925
rect -2960 21435 -2920 21440
rect -2960 21405 -2955 21435
rect -2925 21405 -2920 21435
rect -2960 21275 -2920 21405
rect -2960 21245 -2955 21275
rect -2925 21245 -2920 21275
rect -2960 21115 -2920 21245
rect -2960 21085 -2955 21115
rect -2925 21085 -2920 21115
rect -2960 20955 -2920 21085
rect -2960 20925 -2955 20955
rect -2925 20925 -2920 20955
rect -2960 20920 -2920 20925
rect -2880 21435 -2840 21440
rect -2880 21405 -2875 21435
rect -2845 21405 -2840 21435
rect -2880 21275 -2840 21405
rect -2880 21245 -2875 21275
rect -2845 21245 -2840 21275
rect -2880 21115 -2840 21245
rect -2880 21085 -2875 21115
rect -2845 21085 -2840 21115
rect -2880 20955 -2840 21085
rect -2880 20925 -2875 20955
rect -2845 20925 -2840 20955
rect -2880 20920 -2840 20925
rect -2800 21435 -2760 21440
rect -2800 21405 -2795 21435
rect -2765 21405 -2760 21435
rect -2800 21275 -2760 21405
rect -2800 21245 -2795 21275
rect -2765 21245 -2760 21275
rect -2800 21115 -2760 21245
rect -2800 21085 -2795 21115
rect -2765 21085 -2760 21115
rect -2800 20955 -2760 21085
rect -2800 20925 -2795 20955
rect -2765 20925 -2760 20955
rect -2800 20920 -2760 20925
rect -2720 21435 -2680 21440
rect -2720 21405 -2715 21435
rect -2685 21405 -2680 21435
rect -2720 21275 -2680 21405
rect -2720 21245 -2715 21275
rect -2685 21245 -2680 21275
rect -2720 21115 -2680 21245
rect -2720 21085 -2715 21115
rect -2685 21085 -2680 21115
rect -2720 20955 -2680 21085
rect -2720 20925 -2715 20955
rect -2685 20925 -2680 20955
rect -2720 20920 -2680 20925
rect -2640 21435 -2600 21440
rect -2640 21405 -2635 21435
rect -2605 21405 -2600 21435
rect -2640 21275 -2600 21405
rect -2640 21245 -2635 21275
rect -2605 21245 -2600 21275
rect -2640 21115 -2600 21245
rect -2640 21085 -2635 21115
rect -2605 21085 -2600 21115
rect -2640 20955 -2600 21085
rect -2640 20925 -2635 20955
rect -2605 20925 -2600 20955
rect -2640 20920 -2600 20925
rect -2560 21435 -2520 21440
rect -2560 21405 -2555 21435
rect -2525 21405 -2520 21435
rect -2560 21275 -2520 21405
rect -2560 21245 -2555 21275
rect -2525 21245 -2520 21275
rect -2560 21115 -2520 21245
rect -2560 21085 -2555 21115
rect -2525 21085 -2520 21115
rect -2560 20955 -2520 21085
rect -2560 20925 -2555 20955
rect -2525 20925 -2520 20955
rect -2560 20920 -2520 20925
rect -2480 21435 -2440 21440
rect -2480 21405 -2475 21435
rect -2445 21405 -2440 21435
rect -2480 21275 -2440 21405
rect -2480 21245 -2475 21275
rect -2445 21245 -2440 21275
rect -2480 21115 -2440 21245
rect -2480 21085 -2475 21115
rect -2445 21085 -2440 21115
rect -2480 20955 -2440 21085
rect -2480 20925 -2475 20955
rect -2445 20925 -2440 20955
rect -2480 20920 -2440 20925
rect -2400 21435 -2360 21440
rect -2400 21405 -2395 21435
rect -2365 21405 -2360 21435
rect -2400 21275 -2360 21405
rect -2400 21245 -2395 21275
rect -2365 21245 -2360 21275
rect -2400 21115 -2360 21245
rect -2400 21085 -2395 21115
rect -2365 21085 -2360 21115
rect -2400 20955 -2360 21085
rect -2400 20925 -2395 20955
rect -2365 20925 -2360 20955
rect -2400 20920 -2360 20925
rect -2320 21435 -2280 21440
rect -2320 21405 -2315 21435
rect -2285 21405 -2280 21435
rect -2320 21275 -2280 21405
rect -2320 21245 -2315 21275
rect -2285 21245 -2280 21275
rect -2320 21115 -2280 21245
rect -2320 21085 -2315 21115
rect -2285 21085 -2280 21115
rect -2320 20955 -2280 21085
rect -2320 20925 -2315 20955
rect -2285 20925 -2280 20955
rect -2320 20920 -2280 20925
rect -2240 21435 -2200 21440
rect -2240 21405 -2235 21435
rect -2205 21405 -2200 21435
rect -2240 21275 -2200 21405
rect -2240 21245 -2235 21275
rect -2205 21245 -2200 21275
rect -2240 21115 -2200 21245
rect -2240 21085 -2235 21115
rect -2205 21085 -2200 21115
rect -2240 20955 -2200 21085
rect -2240 20925 -2235 20955
rect -2205 20925 -2200 20955
rect -2240 20920 -2200 20925
rect -2160 21435 -2120 21440
rect -2160 21405 -2155 21435
rect -2125 21405 -2120 21435
rect -2160 21275 -2120 21405
rect -2160 21245 -2155 21275
rect -2125 21245 -2120 21275
rect -2160 21115 -2120 21245
rect -2160 21085 -2155 21115
rect -2125 21085 -2120 21115
rect -2160 20955 -2120 21085
rect -2160 20925 -2155 20955
rect -2125 20925 -2120 20955
rect -2160 20920 -2120 20925
rect -2080 21435 -2040 21440
rect -2080 21405 -2075 21435
rect -2045 21405 -2040 21435
rect -2080 21275 -2040 21405
rect -2080 21245 -2075 21275
rect -2045 21245 -2040 21275
rect -2080 21115 -2040 21245
rect -2080 21085 -2075 21115
rect -2045 21085 -2040 21115
rect -2080 20955 -2040 21085
rect -2080 20925 -2075 20955
rect -2045 20925 -2040 20955
rect -2080 20920 -2040 20925
rect -2000 21435 -1960 21440
rect -2000 21405 -1995 21435
rect -1965 21405 -1960 21435
rect -2000 21275 -1960 21405
rect -2000 21245 -1995 21275
rect -1965 21245 -1960 21275
rect -2000 21115 -1960 21245
rect -2000 21085 -1995 21115
rect -1965 21085 -1960 21115
rect -2000 20955 -1960 21085
rect -2000 20925 -1995 20955
rect -1965 20925 -1960 20955
rect -2000 20920 -1960 20925
rect -1840 21435 -1800 21440
rect -1840 21405 -1835 21435
rect -1805 21405 -1800 21435
rect -1840 21275 -1800 21405
rect -1840 21245 -1835 21275
rect -1805 21245 -1800 21275
rect -1840 21115 -1800 21245
rect -1840 21085 -1835 21115
rect -1805 21085 -1800 21115
rect -1840 20955 -1800 21085
rect -1840 20925 -1835 20955
rect -1805 20925 -1800 20955
rect -1840 20920 -1800 20925
rect -1760 21435 -1720 21440
rect -1760 21405 -1755 21435
rect -1725 21405 -1720 21435
rect -1760 21275 -1720 21405
rect -1760 21245 -1755 21275
rect -1725 21245 -1720 21275
rect -1760 21115 -1720 21245
rect -1760 21085 -1755 21115
rect -1725 21085 -1720 21115
rect -1760 20955 -1720 21085
rect -1760 20925 -1755 20955
rect -1725 20925 -1720 20955
rect -1760 20920 -1720 20925
rect -1680 21435 -1640 21440
rect -1680 21405 -1675 21435
rect -1645 21405 -1640 21435
rect -1680 21275 -1640 21405
rect -1680 21245 -1675 21275
rect -1645 21245 -1640 21275
rect -1680 21115 -1640 21245
rect -1600 21435 -1560 21440
rect -1600 21405 -1595 21435
rect -1565 21405 -1560 21435
rect -1600 21275 -1560 21405
rect -1600 21245 -1595 21275
rect -1565 21245 -1560 21275
rect -1600 21240 -1560 21245
rect -1520 21435 -1480 21440
rect -1520 21405 -1515 21435
rect -1485 21405 -1480 21435
rect -1520 21275 -1480 21405
rect -1360 21435 -1320 21440
rect -1360 21405 -1355 21435
rect -1325 21405 -1320 21435
rect -1520 21245 -1515 21275
rect -1485 21245 -1480 21275
rect -1680 21085 -1675 21115
rect -1645 21085 -1640 21115
rect -1680 20955 -1640 21085
rect -1680 20925 -1675 20955
rect -1645 20925 -1640 20955
rect -5760 20845 -5755 20875
rect -5725 20845 -5720 20875
rect -5760 20795 -5720 20845
rect -5760 20765 -5755 20795
rect -5725 20765 -5720 20795
rect -5760 20435 -5720 20765
rect -1680 20875 -1640 20925
rect -1680 20845 -1675 20875
rect -1645 20845 -1640 20875
rect -1680 20795 -1640 20845
rect -1680 20765 -1675 20795
rect -1645 20765 -1640 20795
rect -5680 20675 -5640 20680
rect -5680 20645 -5675 20675
rect -5645 20645 -5640 20675
rect -5680 20515 -5640 20645
rect -5680 20485 -5675 20515
rect -5645 20485 -5640 20515
rect -5680 20480 -5640 20485
rect -5600 20675 -5560 20680
rect -5600 20645 -5595 20675
rect -5565 20645 -5560 20675
rect -5600 20515 -5560 20645
rect -5600 20485 -5595 20515
rect -5565 20485 -5560 20515
rect -5600 20480 -5560 20485
rect -5520 20675 -5480 20680
rect -5520 20645 -5515 20675
rect -5485 20645 -5480 20675
rect -5520 20515 -5480 20645
rect -5520 20485 -5515 20515
rect -5485 20485 -5480 20515
rect -5520 20480 -5480 20485
rect -5440 20675 -5400 20680
rect -5440 20645 -5435 20675
rect -5405 20645 -5400 20675
rect -5440 20515 -5400 20645
rect -5440 20485 -5435 20515
rect -5405 20485 -5400 20515
rect -5440 20480 -5400 20485
rect -5360 20675 -5320 20680
rect -5360 20645 -5355 20675
rect -5325 20645 -5320 20675
rect -5360 20515 -5320 20645
rect -5360 20485 -5355 20515
rect -5325 20485 -5320 20515
rect -5360 20480 -5320 20485
rect -5280 20675 -5240 20680
rect -5280 20645 -5275 20675
rect -5245 20645 -5240 20675
rect -5280 20515 -5240 20645
rect -5280 20485 -5275 20515
rect -5245 20485 -5240 20515
rect -5280 20480 -5240 20485
rect -5200 20675 -5160 20680
rect -5200 20645 -5195 20675
rect -5165 20645 -5160 20675
rect -5200 20515 -5160 20645
rect -5200 20485 -5195 20515
rect -5165 20485 -5160 20515
rect -5200 20480 -5160 20485
rect -5120 20675 -5080 20680
rect -5120 20645 -5115 20675
rect -5085 20645 -5080 20675
rect -5120 20515 -5080 20645
rect -5120 20485 -5115 20515
rect -5085 20485 -5080 20515
rect -5120 20480 -5080 20485
rect -5040 20675 -5000 20680
rect -5040 20645 -5035 20675
rect -5005 20645 -5000 20675
rect -5040 20515 -5000 20645
rect -5040 20485 -5035 20515
rect -5005 20485 -5000 20515
rect -5040 20480 -5000 20485
rect -4960 20675 -4920 20680
rect -4960 20645 -4955 20675
rect -4925 20645 -4920 20675
rect -4960 20515 -4920 20645
rect -4960 20485 -4955 20515
rect -4925 20485 -4920 20515
rect -4960 20480 -4920 20485
rect -4880 20675 -4840 20680
rect -4880 20645 -4875 20675
rect -4845 20645 -4840 20675
rect -4880 20515 -4840 20645
rect -4880 20485 -4875 20515
rect -4845 20485 -4840 20515
rect -4880 20480 -4840 20485
rect -4800 20675 -4760 20680
rect -4800 20645 -4795 20675
rect -4765 20645 -4760 20675
rect -4800 20515 -4760 20645
rect -4800 20485 -4795 20515
rect -4765 20485 -4760 20515
rect -4800 20480 -4760 20485
rect -4720 20675 -4680 20680
rect -4720 20645 -4715 20675
rect -4685 20645 -4680 20675
rect -4720 20515 -4680 20645
rect -4720 20485 -4715 20515
rect -4685 20485 -4680 20515
rect -4720 20480 -4680 20485
rect -4640 20675 -4600 20680
rect -4640 20645 -4635 20675
rect -4605 20645 -4600 20675
rect -4640 20515 -4600 20645
rect -4640 20485 -4635 20515
rect -4605 20485 -4600 20515
rect -4640 20480 -4600 20485
rect -4560 20675 -4520 20680
rect -4560 20645 -4555 20675
rect -4525 20645 -4520 20675
rect -4560 20515 -4520 20645
rect -4560 20485 -4555 20515
rect -4525 20485 -4520 20515
rect -4560 20480 -4520 20485
rect -4480 20675 -4440 20680
rect -4480 20645 -4475 20675
rect -4445 20645 -4440 20675
rect -4480 20515 -4440 20645
rect -4480 20485 -4475 20515
rect -4445 20485 -4440 20515
rect -4480 20480 -4440 20485
rect -4400 20675 -4360 20680
rect -4400 20645 -4395 20675
rect -4365 20645 -4360 20675
rect -4400 20515 -4360 20645
rect -4400 20485 -4395 20515
rect -4365 20485 -4360 20515
rect -4400 20480 -4360 20485
rect -4320 20675 -4280 20680
rect -4320 20645 -4315 20675
rect -4285 20645 -4280 20675
rect -4320 20515 -4280 20645
rect -4320 20485 -4315 20515
rect -4285 20485 -4280 20515
rect -4320 20480 -4280 20485
rect -4240 20675 -4200 20680
rect -4240 20645 -4235 20675
rect -4205 20645 -4200 20675
rect -4240 20515 -4200 20645
rect -4240 20485 -4235 20515
rect -4205 20485 -4200 20515
rect -4240 20480 -4200 20485
rect -4160 20675 -4120 20680
rect -4160 20645 -4155 20675
rect -4125 20645 -4120 20675
rect -4160 20515 -4120 20645
rect -4160 20485 -4155 20515
rect -4125 20485 -4120 20515
rect -4160 20480 -4120 20485
rect -4080 20675 -4040 20680
rect -4080 20645 -4075 20675
rect -4045 20645 -4040 20675
rect -4080 20515 -4040 20645
rect -4080 20485 -4075 20515
rect -4045 20485 -4040 20515
rect -4080 20480 -4040 20485
rect -4000 20675 -3960 20680
rect -4000 20645 -3995 20675
rect -3965 20645 -3960 20675
rect -4000 20515 -3960 20645
rect -4000 20485 -3995 20515
rect -3965 20485 -3960 20515
rect -4000 20480 -3960 20485
rect -3920 20675 -3880 20680
rect -3920 20645 -3915 20675
rect -3885 20645 -3880 20675
rect -3920 20515 -3880 20645
rect -3920 20485 -3915 20515
rect -3885 20485 -3880 20515
rect -3920 20480 -3880 20485
rect -3840 20675 -3800 20680
rect -3840 20645 -3835 20675
rect -3805 20645 -3800 20675
rect -3840 20515 -3800 20645
rect -3840 20485 -3835 20515
rect -3805 20485 -3800 20515
rect -3840 20480 -3800 20485
rect -3760 20675 -3720 20680
rect -3760 20645 -3755 20675
rect -3725 20645 -3720 20675
rect -3760 20515 -3720 20645
rect -3760 20485 -3755 20515
rect -3725 20485 -3720 20515
rect -3760 20480 -3720 20485
rect -3680 20675 -3640 20680
rect -3680 20645 -3675 20675
rect -3645 20645 -3640 20675
rect -3680 20515 -3640 20645
rect -3680 20485 -3675 20515
rect -3645 20485 -3640 20515
rect -3680 20480 -3640 20485
rect -3600 20675 -3560 20680
rect -3600 20645 -3595 20675
rect -3565 20645 -3560 20675
rect -3600 20515 -3560 20645
rect -3600 20485 -3595 20515
rect -3565 20485 -3560 20515
rect -3600 20480 -3560 20485
rect -3520 20675 -3480 20680
rect -3520 20645 -3515 20675
rect -3485 20645 -3480 20675
rect -3520 20515 -3480 20645
rect -3520 20485 -3515 20515
rect -3485 20485 -3480 20515
rect -3520 20480 -3480 20485
rect -3440 20675 -3400 20680
rect -3440 20645 -3435 20675
rect -3405 20645 -3400 20675
rect -3440 20515 -3400 20645
rect -3440 20485 -3435 20515
rect -3405 20485 -3400 20515
rect -3440 20480 -3400 20485
rect -3360 20675 -3320 20680
rect -3360 20645 -3355 20675
rect -3325 20645 -3320 20675
rect -3360 20515 -3320 20645
rect -3360 20485 -3355 20515
rect -3325 20485 -3320 20515
rect -3360 20480 -3320 20485
rect -3280 20675 -3240 20680
rect -3280 20645 -3275 20675
rect -3245 20645 -3240 20675
rect -3280 20515 -3240 20645
rect -3280 20485 -3275 20515
rect -3245 20485 -3240 20515
rect -3280 20480 -3240 20485
rect -3200 20675 -3160 20680
rect -3200 20645 -3195 20675
rect -3165 20645 -3160 20675
rect -3200 20515 -3160 20645
rect -3200 20485 -3195 20515
rect -3165 20485 -3160 20515
rect -3200 20480 -3160 20485
rect -3120 20675 -3080 20680
rect -3120 20645 -3115 20675
rect -3085 20645 -3080 20675
rect -3120 20515 -3080 20645
rect -3120 20485 -3115 20515
rect -3085 20485 -3080 20515
rect -3120 20480 -3080 20485
rect -3040 20675 -3000 20680
rect -3040 20645 -3035 20675
rect -3005 20645 -3000 20675
rect -3040 20515 -3000 20645
rect -3040 20485 -3035 20515
rect -3005 20485 -3000 20515
rect -3040 20480 -3000 20485
rect -2960 20675 -2920 20680
rect -2960 20645 -2955 20675
rect -2925 20645 -2920 20675
rect -2960 20515 -2920 20645
rect -2960 20485 -2955 20515
rect -2925 20485 -2920 20515
rect -2960 20480 -2920 20485
rect -2880 20675 -2840 20680
rect -2880 20645 -2875 20675
rect -2845 20645 -2840 20675
rect -2880 20515 -2840 20645
rect -2880 20485 -2875 20515
rect -2845 20485 -2840 20515
rect -2880 20480 -2840 20485
rect -2800 20675 -2760 20680
rect -2800 20645 -2795 20675
rect -2765 20645 -2760 20675
rect -2800 20515 -2760 20645
rect -2800 20485 -2795 20515
rect -2765 20485 -2760 20515
rect -2800 20480 -2760 20485
rect -2720 20675 -2680 20680
rect -2720 20645 -2715 20675
rect -2685 20645 -2680 20675
rect -2720 20515 -2680 20645
rect -2720 20485 -2715 20515
rect -2685 20485 -2680 20515
rect -2720 20480 -2680 20485
rect -2640 20675 -2600 20680
rect -2640 20645 -2635 20675
rect -2605 20645 -2600 20675
rect -2640 20515 -2600 20645
rect -2640 20485 -2635 20515
rect -2605 20485 -2600 20515
rect -2640 20480 -2600 20485
rect -2560 20675 -2520 20680
rect -2560 20645 -2555 20675
rect -2525 20645 -2520 20675
rect -2560 20515 -2520 20645
rect -2560 20485 -2555 20515
rect -2525 20485 -2520 20515
rect -2560 20480 -2520 20485
rect -2480 20675 -2440 20680
rect -2480 20645 -2475 20675
rect -2445 20645 -2440 20675
rect -2480 20515 -2440 20645
rect -2480 20485 -2475 20515
rect -2445 20485 -2440 20515
rect -2480 20480 -2440 20485
rect -2400 20675 -2360 20680
rect -2400 20645 -2395 20675
rect -2365 20645 -2360 20675
rect -2400 20515 -2360 20645
rect -2400 20485 -2395 20515
rect -2365 20485 -2360 20515
rect -2400 20480 -2360 20485
rect -2320 20675 -2280 20680
rect -2320 20645 -2315 20675
rect -2285 20645 -2280 20675
rect -2320 20515 -2280 20645
rect -2320 20485 -2315 20515
rect -2285 20485 -2280 20515
rect -2320 20480 -2280 20485
rect -2240 20675 -2200 20680
rect -2240 20645 -2235 20675
rect -2205 20645 -2200 20675
rect -2240 20515 -2200 20645
rect -2240 20485 -2235 20515
rect -2205 20485 -2200 20515
rect -2240 20480 -2200 20485
rect -2160 20675 -2120 20680
rect -2160 20645 -2155 20675
rect -2125 20645 -2120 20675
rect -2160 20515 -2120 20645
rect -2160 20485 -2155 20515
rect -2125 20485 -2120 20515
rect -2160 20480 -2120 20485
rect -2080 20675 -2040 20680
rect -2080 20645 -2075 20675
rect -2045 20645 -2040 20675
rect -2080 20515 -2040 20645
rect -2080 20485 -2075 20515
rect -2045 20485 -2040 20515
rect -2080 20480 -2040 20485
rect -2000 20675 -1960 20680
rect -2000 20645 -1995 20675
rect -1965 20645 -1960 20675
rect -2000 20515 -1960 20645
rect -2000 20485 -1995 20515
rect -1965 20485 -1960 20515
rect -2000 20480 -1960 20485
rect -1920 20675 -1880 20680
rect -1920 20645 -1915 20675
rect -1885 20645 -1880 20675
rect -1920 20515 -1880 20645
rect -1920 20485 -1915 20515
rect -1885 20485 -1880 20515
rect -1920 20480 -1880 20485
rect -1840 20675 -1800 20680
rect -1840 20645 -1835 20675
rect -1805 20645 -1800 20675
rect -1840 20515 -1800 20645
rect -1840 20485 -1835 20515
rect -1805 20485 -1800 20515
rect -1840 20480 -1800 20485
rect -1760 20675 -1720 20680
rect -1760 20645 -1755 20675
rect -1725 20645 -1720 20675
rect -1760 20515 -1720 20645
rect -1760 20485 -1755 20515
rect -1725 20485 -1720 20515
rect -1760 20480 -1720 20485
rect -5760 20405 -5755 20435
rect -5725 20405 -5720 20435
rect -5760 20355 -5720 20405
rect -1680 20435 -1640 20765
rect -1680 20405 -1675 20435
rect -1645 20405 -1640 20435
rect -5760 20325 -5755 20355
rect -5725 20325 -5720 20355
rect -5760 20195 -5720 20325
rect -5760 20165 -5755 20195
rect -5725 20165 -5720 20195
rect -5760 20160 -5720 20165
rect -5280 20355 -5240 20360
rect -5280 20325 -5275 20355
rect -5245 20325 -5240 20355
rect -5280 20195 -5240 20325
rect -5120 20355 -5080 20360
rect -5120 20325 -5115 20355
rect -5085 20325 -5080 20355
rect -5280 20165 -5275 20195
rect -5245 20165 -5240 20195
rect -5280 20160 -5240 20165
rect -5200 20275 -5160 20280
rect -5200 20245 -5195 20275
rect -5165 20245 -5160 20275
rect -5200 19960 -5160 20245
rect -5120 20195 -5080 20325
rect -5120 20165 -5115 20195
rect -5085 20165 -5080 20195
rect -5120 20160 -5080 20165
rect -5040 20355 -5000 20360
rect -5040 20325 -5035 20355
rect -5005 20325 -5000 20355
rect -5040 20195 -5000 20325
rect -5040 20165 -5035 20195
rect -5005 20165 -5000 20195
rect -5040 20160 -5000 20165
rect -4960 20355 -4920 20360
rect -4960 20325 -4955 20355
rect -4925 20325 -4920 20355
rect -4960 20195 -4920 20325
rect -4960 20165 -4955 20195
rect -4925 20165 -4920 20195
rect -4960 20160 -4920 20165
rect -4880 20355 -4840 20360
rect -4880 20325 -4875 20355
rect -4845 20325 -4840 20355
rect -4880 20195 -4840 20325
rect -4880 20165 -4875 20195
rect -4845 20165 -4840 20195
rect -4880 20160 -4840 20165
rect -4800 20355 -4760 20360
rect -4800 20325 -4795 20355
rect -4765 20325 -4760 20355
rect -4800 20195 -4760 20325
rect -4800 20165 -4795 20195
rect -4765 20165 -4760 20195
rect -4800 20160 -4760 20165
rect -4720 20355 -4680 20360
rect -4720 20325 -4715 20355
rect -4685 20325 -4680 20355
rect -4720 20195 -4680 20325
rect -4720 20165 -4715 20195
rect -4685 20165 -4680 20195
rect -4720 20160 -4680 20165
rect -4640 20355 -4600 20360
rect -4640 20325 -4635 20355
rect -4605 20325 -4600 20355
rect -4640 20195 -4600 20325
rect -4640 20165 -4635 20195
rect -4605 20165 -4600 20195
rect -4640 20160 -4600 20165
rect -4560 20355 -4520 20360
rect -4560 20325 -4555 20355
rect -4525 20325 -4520 20355
rect -4560 20195 -4520 20325
rect -4560 20165 -4555 20195
rect -4525 20165 -4520 20195
rect -4560 20160 -4520 20165
rect -4480 20355 -4440 20360
rect -4480 20325 -4475 20355
rect -4445 20325 -4440 20355
rect -4480 20195 -4440 20325
rect -4480 20165 -4475 20195
rect -4445 20165 -4440 20195
rect -4480 20160 -4440 20165
rect -4400 20355 -4360 20360
rect -4400 20325 -4395 20355
rect -4365 20325 -4360 20355
rect -4400 20195 -4360 20325
rect -4400 20165 -4395 20195
rect -4365 20165 -4360 20195
rect -4400 20160 -4360 20165
rect -4320 20355 -4280 20360
rect -4320 20325 -4315 20355
rect -4285 20325 -4280 20355
rect -4320 20195 -4280 20325
rect -4320 20165 -4315 20195
rect -4285 20165 -4280 20195
rect -4320 20160 -4280 20165
rect -4240 20355 -4200 20360
rect -4240 20325 -4235 20355
rect -4205 20325 -4200 20355
rect -4240 20195 -4200 20325
rect -4240 20165 -4235 20195
rect -4205 20165 -4200 20195
rect -4240 20160 -4200 20165
rect -4160 20355 -4120 20360
rect -4160 20325 -4155 20355
rect -4125 20325 -4120 20355
rect -4160 20195 -4120 20325
rect -4160 20165 -4155 20195
rect -4125 20165 -4120 20195
rect -4160 20160 -4120 20165
rect -4080 20355 -4040 20360
rect -4080 20325 -4075 20355
rect -4045 20325 -4040 20355
rect -4080 20195 -4040 20325
rect -4080 20165 -4075 20195
rect -4045 20165 -4040 20195
rect -4080 20160 -4040 20165
rect -4000 20355 -3960 20360
rect -4000 20325 -3995 20355
rect -3965 20325 -3960 20355
rect -4000 20195 -3960 20325
rect -4000 20165 -3995 20195
rect -3965 20165 -3960 20195
rect -4000 20160 -3960 20165
rect -3920 20355 -3880 20360
rect -3920 20325 -3915 20355
rect -3885 20325 -3880 20355
rect -3920 20195 -3880 20325
rect -3920 20165 -3915 20195
rect -3885 20165 -3880 20195
rect -3920 20160 -3880 20165
rect -3840 20355 -3800 20360
rect -3840 20325 -3835 20355
rect -3805 20325 -3800 20355
rect -3840 20195 -3800 20325
rect -3840 20165 -3835 20195
rect -3805 20165 -3800 20195
rect -3840 20160 -3800 20165
rect -3760 20355 -3720 20360
rect -3760 20325 -3755 20355
rect -3725 20325 -3720 20355
rect -3760 20195 -3720 20325
rect -3760 20165 -3755 20195
rect -3725 20165 -3720 20195
rect -3760 20160 -3720 20165
rect -3680 20355 -3640 20360
rect -3680 20325 -3675 20355
rect -3645 20325 -3640 20355
rect -3680 20195 -3640 20325
rect -3680 20165 -3675 20195
rect -3645 20165 -3640 20195
rect -3680 20160 -3640 20165
rect -3600 20355 -3560 20360
rect -3600 20325 -3595 20355
rect -3565 20325 -3560 20355
rect -3600 20195 -3560 20325
rect -3600 20165 -3595 20195
rect -3565 20165 -3560 20195
rect -3600 20160 -3560 20165
rect -3520 20355 -3480 20360
rect -3520 20325 -3515 20355
rect -3485 20325 -3480 20355
rect -3520 20195 -3480 20325
rect -3520 20165 -3515 20195
rect -3485 20165 -3480 20195
rect -3520 20160 -3480 20165
rect -3440 20355 -3400 20360
rect -3440 20325 -3435 20355
rect -3405 20325 -3400 20355
rect -3440 20195 -3400 20325
rect -3440 20165 -3435 20195
rect -3405 20165 -3400 20195
rect -3440 20160 -3400 20165
rect -3360 20355 -3320 20360
rect -3360 20325 -3355 20355
rect -3325 20325 -3320 20355
rect -3360 20195 -3320 20325
rect -3360 20165 -3355 20195
rect -3325 20165 -3320 20195
rect -3360 20160 -3320 20165
rect -3280 20355 -3240 20360
rect -3280 20325 -3275 20355
rect -3245 20325 -3240 20355
rect -3280 20195 -3240 20325
rect -3280 20165 -3275 20195
rect -3245 20165 -3240 20195
rect -3280 20160 -3240 20165
rect -3200 20355 -3160 20360
rect -3200 20325 -3195 20355
rect -3165 20325 -3160 20355
rect -3200 20195 -3160 20325
rect -3200 20165 -3195 20195
rect -3165 20165 -3160 20195
rect -3200 20160 -3160 20165
rect -3120 20355 -3080 20360
rect -3120 20325 -3115 20355
rect -3085 20325 -3080 20355
rect -3120 20195 -3080 20325
rect -3120 20165 -3115 20195
rect -3085 20165 -3080 20195
rect -3120 20160 -3080 20165
rect -3040 20355 -3000 20360
rect -3040 20325 -3035 20355
rect -3005 20325 -3000 20355
rect -3040 20195 -3000 20325
rect -3040 20165 -3035 20195
rect -3005 20165 -3000 20195
rect -3040 20160 -3000 20165
rect -2960 20355 -2920 20360
rect -2960 20325 -2955 20355
rect -2925 20325 -2920 20355
rect -2960 20195 -2920 20325
rect -2960 20165 -2955 20195
rect -2925 20165 -2920 20195
rect -2960 20160 -2920 20165
rect -2880 20355 -2840 20360
rect -2880 20325 -2875 20355
rect -2845 20325 -2840 20355
rect -2880 20195 -2840 20325
rect -2880 20165 -2875 20195
rect -2845 20165 -2840 20195
rect -2880 20160 -2840 20165
rect -2800 20355 -2760 20360
rect -2800 20325 -2795 20355
rect -2765 20325 -2760 20355
rect -2800 20195 -2760 20325
rect -2800 20165 -2795 20195
rect -2765 20165 -2760 20195
rect -2800 20160 -2760 20165
rect -2720 20355 -2680 20360
rect -2720 20325 -2715 20355
rect -2685 20325 -2680 20355
rect -2720 20195 -2680 20325
rect -2720 20165 -2715 20195
rect -2685 20165 -2680 20195
rect -2720 20160 -2680 20165
rect -2640 20355 -2600 20360
rect -2640 20325 -2635 20355
rect -2605 20325 -2600 20355
rect -2640 20195 -2600 20325
rect -2640 20165 -2635 20195
rect -2605 20165 -2600 20195
rect -2640 20160 -2600 20165
rect -2560 20355 -2520 20360
rect -2560 20325 -2555 20355
rect -2525 20325 -2520 20355
rect -2560 20195 -2520 20325
rect -2560 20165 -2555 20195
rect -2525 20165 -2520 20195
rect -2560 20160 -2520 20165
rect -2480 20355 -2440 20360
rect -2480 20325 -2475 20355
rect -2445 20325 -2440 20355
rect -2480 20195 -2440 20325
rect -2480 20165 -2475 20195
rect -2445 20165 -2440 20195
rect -2480 20160 -2440 20165
rect -2400 20355 -2360 20360
rect -2400 20325 -2395 20355
rect -2365 20325 -2360 20355
rect -2400 20195 -2360 20325
rect -2400 20165 -2395 20195
rect -2365 20165 -2360 20195
rect -2400 20160 -2360 20165
rect -2320 20355 -2280 20360
rect -2320 20325 -2315 20355
rect -2285 20325 -2280 20355
rect -2320 20195 -2280 20325
rect -2320 20165 -2315 20195
rect -2285 20165 -2280 20195
rect -2320 20160 -2280 20165
rect -2240 20355 -2200 20360
rect -2240 20325 -2235 20355
rect -2205 20325 -2200 20355
rect -2240 20195 -2200 20325
rect -2240 20165 -2235 20195
rect -2205 20165 -2200 20195
rect -2240 20160 -2200 20165
rect -2160 20355 -2120 20360
rect -2160 20325 -2155 20355
rect -2125 20325 -2120 20355
rect -2160 20195 -2120 20325
rect -2160 20165 -2155 20195
rect -2125 20165 -2120 20195
rect -2160 20160 -2120 20165
rect -2080 20355 -2040 20360
rect -2080 20325 -2075 20355
rect -2045 20325 -2040 20355
rect -2080 20195 -2040 20325
rect -2080 20165 -2075 20195
rect -2045 20165 -2040 20195
rect -2080 20160 -2040 20165
rect -2000 20355 -1960 20360
rect -2000 20325 -1995 20355
rect -1965 20325 -1960 20355
rect -2000 20195 -1960 20325
rect -2000 20165 -1995 20195
rect -1965 20165 -1960 20195
rect -2000 20160 -1960 20165
rect -1840 20355 -1800 20360
rect -1840 20325 -1835 20355
rect -1805 20325 -1800 20355
rect -1840 20195 -1800 20325
rect -1840 20165 -1835 20195
rect -1805 20165 -1800 20195
rect -1840 20160 -1800 20165
rect -1760 20355 -1720 20360
rect -1760 20325 -1755 20355
rect -1725 20325 -1720 20355
rect -1760 20195 -1720 20325
rect -1760 20165 -1755 20195
rect -1725 20165 -1720 20195
rect -1760 20160 -1720 20165
rect -1680 20355 -1640 20405
rect -1680 20325 -1675 20355
rect -1645 20325 -1640 20355
rect -1680 20195 -1640 20325
rect -1680 20165 -1675 20195
rect -1645 20165 -1640 20195
rect -1680 20115 -1640 20165
rect -1680 20085 -1675 20115
rect -1645 20085 -1640 20115
rect -1680 20035 -1640 20085
rect -1680 20005 -1675 20035
rect -1645 20005 -1640 20035
rect -15040 19884 -15036 19916
rect -15004 19884 -15000 19916
rect -15040 19836 -15000 19884
rect -15040 19804 -15036 19836
rect -15004 19804 -15000 19836
rect -15040 19756 -15000 19804
rect -15040 19724 -15036 19756
rect -15004 19724 -15000 19756
rect -15040 19676 -15000 19724
rect -15040 19644 -15036 19676
rect -15004 19644 -15000 19676
rect -15040 19596 -15000 19644
rect -15040 19564 -15036 19596
rect -15004 19564 -15000 19596
rect -15040 19516 -15000 19564
rect -15040 19484 -15036 19516
rect -15004 19484 -15000 19516
rect -15040 19436 -15000 19484
rect -15040 19404 -15036 19436
rect -15004 19404 -15000 19436
rect -15040 19356 -15000 19404
rect -15040 19324 -15036 19356
rect -15004 19324 -15000 19356
rect -15040 19276 -15000 19324
rect -15040 19244 -15036 19276
rect -15004 19244 -15000 19276
rect -15040 19196 -15000 19244
rect -15040 19164 -15036 19196
rect -15004 19164 -15000 19196
rect -15040 19116 -15000 19164
rect -15040 19084 -15036 19116
rect -15004 19084 -15000 19116
rect -15040 19036 -15000 19084
rect -15040 19004 -15036 19036
rect -15004 19004 -15000 19036
rect -15040 18956 -15000 19004
rect -15040 18924 -15036 18956
rect -15004 18924 -15000 18956
rect -15040 18876 -15000 18924
rect -15040 18844 -15036 18876
rect -15004 18844 -15000 18876
rect -15040 18715 -15000 18844
rect -15040 18685 -15035 18715
rect -15005 18685 -15000 18715
rect -15200 18524 -15196 18556
rect -15164 18524 -15160 18556
rect -15200 18476 -15160 18524
rect -15200 18444 -15196 18476
rect -15164 18444 -15160 18476
rect -15200 18396 -15160 18444
rect -15200 18364 -15196 18396
rect -15164 18364 -15160 18396
rect -15200 18316 -15160 18364
rect -15200 18284 -15196 18316
rect -15164 18284 -15160 18316
rect -15200 18236 -15160 18284
rect -15200 18204 -15196 18236
rect -15164 18204 -15160 18236
rect -15200 18156 -15160 18204
rect -15200 18124 -15196 18156
rect -15164 18124 -15160 18156
rect -15200 18076 -15160 18124
rect -15200 18044 -15196 18076
rect -15164 18044 -15160 18076
rect -15200 17996 -15160 18044
rect -15200 17964 -15196 17996
rect -15164 17964 -15160 17996
rect -15200 17916 -15160 17964
rect -15200 17884 -15196 17916
rect -15164 17884 -15160 17916
rect -15200 17836 -15160 17884
rect -15120 17880 -15080 18560
rect -15040 18556 -15000 18685
rect -15040 18524 -15036 18556
rect -15004 18524 -15000 18556
rect -15040 18476 -15000 18524
rect -15040 18444 -15036 18476
rect -15004 18444 -15000 18476
rect -15040 18396 -15000 18444
rect -15040 18364 -15036 18396
rect -15004 18364 -15000 18396
rect -15040 18316 -15000 18364
rect -15040 18284 -15036 18316
rect -15004 18284 -15000 18316
rect -15040 18236 -15000 18284
rect -15040 18204 -15036 18236
rect -15004 18204 -15000 18236
rect -15040 18156 -15000 18204
rect -15040 18124 -15036 18156
rect -15004 18124 -15000 18156
rect -15040 18076 -15000 18124
rect -15040 18044 -15036 18076
rect -15004 18044 -15000 18076
rect -15040 17996 -15000 18044
rect -15040 17964 -15036 17996
rect -15004 17964 -15000 17996
rect -15040 17916 -15000 17964
rect -15040 17884 -15036 17916
rect -15004 17884 -15000 17916
rect -15200 17804 -15196 17836
rect -15164 17804 -15160 17836
rect -15200 17756 -15160 17804
rect -15200 17724 -15196 17756
rect -15164 17724 -15160 17756
rect -15200 17676 -15160 17724
rect -15200 17644 -15196 17676
rect -15164 17644 -15160 17676
rect -15200 17596 -15160 17644
rect -15200 17564 -15196 17596
rect -15164 17564 -15160 17596
rect -15200 17516 -15160 17564
rect -15200 17484 -15196 17516
rect -15164 17484 -15160 17516
rect -15200 17436 -15160 17484
rect -15200 17404 -15196 17436
rect -15164 17404 -15160 17436
rect -15200 17355 -15160 17404
rect -15120 17400 -15080 17840
rect -15040 17836 -15000 17884
rect -15040 17804 -15036 17836
rect -15004 17804 -15000 17836
rect -15040 17756 -15000 17804
rect -15040 17724 -15036 17756
rect -15004 17724 -15000 17756
rect -15040 17676 -15000 17724
rect -15040 17644 -15036 17676
rect -15004 17644 -15000 17676
rect -15040 17596 -15000 17644
rect -15040 17564 -15036 17596
rect -15004 17564 -15000 17596
rect -15040 17516 -15000 17564
rect -15040 17484 -15036 17516
rect -15004 17484 -15000 17516
rect -15040 17436 -15000 17484
rect -1680 19955 -1640 20005
rect -1680 19925 -1675 19955
rect -1645 19925 -1640 19955
rect -1680 19876 -1640 19925
rect -1680 19844 -1676 19876
rect -1644 19844 -1640 19876
rect -1680 19796 -1640 19844
rect -1680 19764 -1676 19796
rect -1644 19764 -1640 19796
rect -1680 19716 -1640 19764
rect -1680 19684 -1676 19716
rect -1644 19684 -1640 19716
rect -1680 19636 -1640 19684
rect -1680 19604 -1676 19636
rect -1644 19604 -1640 19636
rect -1680 19556 -1640 19604
rect -1680 19524 -1676 19556
rect -1644 19524 -1640 19556
rect -1680 19476 -1640 19524
rect -1680 19444 -1676 19476
rect -1644 19444 -1640 19476
rect -1680 19396 -1640 19444
rect -1680 19364 -1676 19396
rect -1644 19364 -1640 19396
rect -1680 19316 -1640 19364
rect -1680 19284 -1676 19316
rect -1644 19284 -1640 19316
rect -1680 19236 -1640 19284
rect -1680 19204 -1676 19236
rect -1644 19204 -1640 19236
rect -1680 19156 -1640 19204
rect -1680 19124 -1676 19156
rect -1644 19124 -1640 19156
rect -1680 19076 -1640 19124
rect -1680 19044 -1676 19076
rect -1644 19044 -1640 19076
rect -1680 18996 -1640 19044
rect -1680 18964 -1676 18996
rect -1644 18964 -1640 18996
rect -1680 18916 -1640 18964
rect -1680 18884 -1676 18916
rect -1644 18884 -1640 18916
rect -1680 18835 -1640 18884
rect -1680 18805 -1675 18835
rect -1645 18805 -1640 18835
rect -1680 18756 -1640 18805
rect -1680 18724 -1676 18756
rect -1644 18724 -1640 18756
rect -1680 18676 -1640 18724
rect -1680 18644 -1676 18676
rect -1644 18644 -1640 18676
rect -1680 18596 -1640 18644
rect -1680 18564 -1676 18596
rect -1644 18564 -1640 18596
rect -1680 18516 -1640 18564
rect -1680 18484 -1676 18516
rect -1644 18484 -1640 18516
rect -1680 18436 -1640 18484
rect -1680 18404 -1676 18436
rect -1644 18404 -1640 18436
rect -1680 18356 -1640 18404
rect -1680 18324 -1676 18356
rect -1644 18324 -1640 18356
rect -1680 18276 -1640 18324
rect -1680 18244 -1676 18276
rect -1644 18244 -1640 18276
rect -1680 18196 -1640 18244
rect -1680 18164 -1676 18196
rect -1644 18164 -1640 18196
rect -1680 18115 -1640 18164
rect -1680 18085 -1675 18115
rect -1645 18085 -1640 18115
rect -1680 18035 -1640 18085
rect -1680 18005 -1675 18035
rect -1645 18005 -1640 18035
rect -1680 17876 -1640 18005
rect -1600 21195 -1560 21200
rect -1600 21165 -1595 21195
rect -1565 21165 -1560 21195
rect -1600 17955 -1560 21165
rect -1600 17925 -1595 17955
rect -1565 17925 -1560 17955
rect -1600 17920 -1560 17925
rect -1520 21115 -1480 21245
rect -1520 21085 -1515 21115
rect -1485 21085 -1480 21115
rect -1520 20955 -1480 21085
rect -1520 20925 -1515 20955
rect -1485 20925 -1480 20955
rect -1520 20875 -1480 20925
rect -1520 20845 -1515 20875
rect -1485 20845 -1480 20875
rect -1520 20795 -1480 20845
rect -1520 20765 -1515 20795
rect -1485 20765 -1480 20795
rect -1520 20435 -1480 20765
rect -1520 20405 -1515 20435
rect -1485 20405 -1480 20435
rect -1520 20355 -1480 20405
rect -1520 20325 -1515 20355
rect -1485 20325 -1480 20355
rect -1520 20195 -1480 20325
rect -1520 20165 -1515 20195
rect -1485 20165 -1480 20195
rect -1520 20115 -1480 20165
rect -1520 20085 -1515 20115
rect -1485 20085 -1480 20115
rect -1520 20035 -1480 20085
rect -1520 20005 -1515 20035
rect -1485 20005 -1480 20035
rect -1520 19955 -1480 20005
rect -1520 19925 -1515 19955
rect -1485 19925 -1480 19955
rect -1520 19876 -1480 19925
rect -1520 19844 -1516 19876
rect -1484 19844 -1480 19876
rect -1520 19796 -1480 19844
rect -1520 19764 -1516 19796
rect -1484 19764 -1480 19796
rect -1520 19716 -1480 19764
rect -1520 19684 -1516 19716
rect -1484 19684 -1480 19716
rect -1520 19636 -1480 19684
rect -1520 19604 -1516 19636
rect -1484 19604 -1480 19636
rect -1520 19556 -1480 19604
rect -1520 19524 -1516 19556
rect -1484 19524 -1480 19556
rect -1520 19476 -1480 19524
rect -1520 19444 -1516 19476
rect -1484 19444 -1480 19476
rect -1520 19396 -1480 19444
rect -1520 19364 -1516 19396
rect -1484 19364 -1480 19396
rect -1520 19316 -1480 19364
rect -1520 19284 -1516 19316
rect -1484 19284 -1480 19316
rect -1520 19236 -1480 19284
rect -1520 19204 -1516 19236
rect -1484 19204 -1480 19236
rect -1520 19156 -1480 19204
rect -1520 19124 -1516 19156
rect -1484 19124 -1480 19156
rect -1520 19076 -1480 19124
rect -1520 19044 -1516 19076
rect -1484 19044 -1480 19076
rect -1520 18996 -1480 19044
rect -1520 18964 -1516 18996
rect -1484 18964 -1480 18996
rect -1520 18916 -1480 18964
rect -1520 18884 -1516 18916
rect -1484 18884 -1480 18916
rect -1520 18835 -1480 18884
rect -1520 18805 -1515 18835
rect -1485 18805 -1480 18835
rect -1520 18756 -1480 18805
rect -1520 18724 -1516 18756
rect -1484 18724 -1480 18756
rect -1520 18676 -1480 18724
rect -1520 18644 -1516 18676
rect -1484 18644 -1480 18676
rect -1520 18596 -1480 18644
rect -1520 18564 -1516 18596
rect -1484 18564 -1480 18596
rect -1520 18516 -1480 18564
rect -1520 18484 -1516 18516
rect -1484 18484 -1480 18516
rect -1520 18436 -1480 18484
rect -1520 18404 -1516 18436
rect -1484 18404 -1480 18436
rect -1520 18356 -1480 18404
rect -1520 18324 -1516 18356
rect -1484 18324 -1480 18356
rect -1520 18276 -1480 18324
rect -1520 18244 -1516 18276
rect -1484 18244 -1480 18276
rect -1520 18196 -1480 18244
rect -1520 18164 -1516 18196
rect -1484 18164 -1480 18196
rect -1520 18115 -1480 18164
rect -1520 18085 -1515 18115
rect -1485 18085 -1480 18115
rect -1520 18035 -1480 18085
rect -1440 21355 -1400 21360
rect -1440 21325 -1435 21355
rect -1405 21325 -1400 21355
rect -1440 18115 -1400 21325
rect -1440 18085 -1435 18115
rect -1405 18085 -1400 18115
rect -1440 18080 -1400 18085
rect -1360 21275 -1320 21405
rect -1360 21245 -1355 21275
rect -1325 21245 -1320 21275
rect -1360 21115 -1320 21245
rect -1360 21085 -1355 21115
rect -1325 21085 -1320 21115
rect -1360 20955 -1320 21085
rect -1360 20925 -1355 20955
rect -1325 20925 -1320 20955
rect -1360 20875 -1320 20925
rect -1280 21435 -1240 21440
rect -1280 21405 -1275 21435
rect -1245 21405 -1240 21435
rect -1280 21275 -1240 21405
rect -1280 21245 -1275 21275
rect -1245 21245 -1240 21275
rect -1280 21115 -1240 21245
rect -1280 21085 -1275 21115
rect -1245 21085 -1240 21115
rect -1280 20955 -1240 21085
rect -1280 20925 -1275 20955
rect -1245 20925 -1240 20955
rect -1280 20920 -1240 20925
rect -1200 21435 -1160 21440
rect -1200 21405 -1195 21435
rect -1165 21405 -1160 21435
rect -1200 21275 -1160 21405
rect -1200 21245 -1195 21275
rect -1165 21245 -1160 21275
rect -1200 21115 -1160 21245
rect -1200 21085 -1195 21115
rect -1165 21085 -1160 21115
rect -1200 20955 -1160 21085
rect -1200 20925 -1195 20955
rect -1165 20925 -1160 20955
rect -1360 20845 -1355 20875
rect -1325 20845 -1320 20875
rect -1360 20795 -1320 20845
rect -1360 20765 -1355 20795
rect -1325 20765 -1320 20795
rect -1360 20435 -1320 20765
rect -1360 20405 -1355 20435
rect -1325 20405 -1320 20435
rect -1360 20355 -1320 20405
rect -1360 20325 -1355 20355
rect -1325 20325 -1320 20355
rect -1360 20195 -1320 20325
rect -1360 20165 -1355 20195
rect -1325 20165 -1320 20195
rect -1360 20115 -1320 20165
rect -1200 20875 -1160 20925
rect -1120 21435 -1080 21440
rect -1120 21405 -1115 21435
rect -1085 21405 -1080 21435
rect -1120 21275 -1080 21405
rect -1120 21245 -1115 21275
rect -1085 21245 -1080 21275
rect -1120 21115 -1080 21245
rect -1120 21085 -1115 21115
rect -1085 21085 -1080 21115
rect -1120 20955 -1080 21085
rect -1120 20925 -1115 20955
rect -1085 20925 -1080 20955
rect -1120 20920 -1080 20925
rect -1040 21435 -1000 21480
rect -1040 21405 -1035 21435
rect -1005 21405 -1000 21435
rect -1040 21275 -1000 21405
rect -1040 21245 -1035 21275
rect -1005 21245 -1000 21275
rect -1040 21115 -1000 21245
rect -1040 21085 -1035 21115
rect -1005 21085 -1000 21115
rect -1040 20955 -1000 21085
rect -1040 20925 -1035 20955
rect -1005 20925 -1000 20955
rect -1200 20845 -1195 20875
rect -1165 20845 -1160 20875
rect -1200 20795 -1160 20845
rect -1200 20765 -1195 20795
rect -1165 20765 -1160 20795
rect -1200 20435 -1160 20765
rect -1200 20405 -1195 20435
rect -1165 20405 -1160 20435
rect -1200 20355 -1160 20405
rect -1200 20325 -1195 20355
rect -1165 20325 -1160 20355
rect -1200 20195 -1160 20325
rect -1200 20165 -1195 20195
rect -1165 20165 -1160 20195
rect -1360 20085 -1355 20115
rect -1325 20085 -1320 20115
rect -1360 20035 -1320 20085
rect -1360 20005 -1355 20035
rect -1325 20005 -1320 20035
rect -1360 19955 -1320 20005
rect -1360 19925 -1355 19955
rect -1325 19925 -1320 19955
rect -1360 19876 -1320 19925
rect -1360 19844 -1356 19876
rect -1324 19844 -1320 19876
rect -1360 19796 -1320 19844
rect -1360 19764 -1356 19796
rect -1324 19764 -1320 19796
rect -1360 19716 -1320 19764
rect -1360 19684 -1356 19716
rect -1324 19684 -1320 19716
rect -1360 19636 -1320 19684
rect -1360 19604 -1356 19636
rect -1324 19604 -1320 19636
rect -1360 19556 -1320 19604
rect -1360 19524 -1356 19556
rect -1324 19524 -1320 19556
rect -1360 19476 -1320 19524
rect -1360 19444 -1356 19476
rect -1324 19444 -1320 19476
rect -1360 19396 -1320 19444
rect -1360 19364 -1356 19396
rect -1324 19364 -1320 19396
rect -1360 19316 -1320 19364
rect -1360 19284 -1356 19316
rect -1324 19284 -1320 19316
rect -1360 19236 -1320 19284
rect -1360 19204 -1356 19236
rect -1324 19204 -1320 19236
rect -1360 19156 -1320 19204
rect -1360 19124 -1356 19156
rect -1324 19124 -1320 19156
rect -1360 19076 -1320 19124
rect -1360 19044 -1356 19076
rect -1324 19044 -1320 19076
rect -1360 18996 -1320 19044
rect -1360 18964 -1356 18996
rect -1324 18964 -1320 18996
rect -1360 18916 -1320 18964
rect -1360 18884 -1356 18916
rect -1324 18884 -1320 18916
rect -1360 18835 -1320 18884
rect -1360 18805 -1355 18835
rect -1325 18805 -1320 18835
rect -1360 18756 -1320 18805
rect -1360 18724 -1356 18756
rect -1324 18724 -1320 18756
rect -1360 18676 -1320 18724
rect -1360 18644 -1356 18676
rect -1324 18644 -1320 18676
rect -1360 18596 -1320 18644
rect -1360 18564 -1356 18596
rect -1324 18564 -1320 18596
rect -1360 18516 -1320 18564
rect -1360 18484 -1356 18516
rect -1324 18484 -1320 18516
rect -1360 18436 -1320 18484
rect -1360 18404 -1356 18436
rect -1324 18404 -1320 18436
rect -1360 18356 -1320 18404
rect -1360 18324 -1356 18356
rect -1324 18324 -1320 18356
rect -1360 18276 -1320 18324
rect -1360 18244 -1356 18276
rect -1324 18244 -1320 18276
rect -1360 18196 -1320 18244
rect -1360 18164 -1356 18196
rect -1324 18164 -1320 18196
rect -1520 18005 -1515 18035
rect -1485 18005 -1480 18035
rect -1680 17844 -1676 17876
rect -1644 17844 -1640 17876
rect -1680 17796 -1640 17844
rect -1680 17764 -1676 17796
rect -1644 17764 -1640 17796
rect -1680 17716 -1640 17764
rect -1680 17684 -1676 17716
rect -1644 17684 -1640 17716
rect -1680 17636 -1640 17684
rect -1680 17604 -1676 17636
rect -1644 17604 -1640 17636
rect -1680 17556 -1640 17604
rect -1680 17524 -1676 17556
rect -1644 17524 -1640 17556
rect -1680 17476 -1640 17524
rect -1680 17444 -1676 17476
rect -1644 17444 -1640 17476
rect -15040 17404 -15036 17436
rect -15004 17404 -15000 17436
rect -15200 17325 -15195 17355
rect -15165 17325 -15160 17355
rect -15200 17195 -15160 17325
rect -15200 17165 -15195 17195
rect -15165 17165 -15160 17195
rect -15200 17116 -15160 17165
rect -15040 17355 -15000 17404
rect -15040 17325 -15035 17355
rect -15005 17325 -15000 17355
rect -15040 17195 -15000 17325
rect -15040 17165 -15035 17195
rect -15005 17165 -15000 17195
rect -15200 17084 -15196 17116
rect -15164 17084 -15160 17116
rect -15200 17036 -15160 17084
rect -15200 17004 -15196 17036
rect -15164 17004 -15160 17036
rect -15200 16956 -15160 17004
rect -15200 16924 -15196 16956
rect -15164 16924 -15160 16956
rect -15200 16876 -15160 16924
rect -15200 16844 -15196 16876
rect -15164 16844 -15160 16876
rect -15200 16796 -15160 16844
rect -15200 16764 -15196 16796
rect -15164 16764 -15160 16796
rect -15200 16716 -15160 16764
rect -15200 16684 -15196 16716
rect -15164 16684 -15160 16716
rect -15200 16636 -15160 16684
rect -15200 16604 -15196 16636
rect -15164 16604 -15160 16636
rect -15200 16556 -15160 16604
rect -15200 16524 -15196 16556
rect -15164 16524 -15160 16556
rect -15200 16476 -15160 16524
rect -15200 16444 -15196 16476
rect -15164 16444 -15160 16476
rect -15360 16285 -15355 16315
rect -15325 16285 -15320 16315
rect -15360 16235 -15320 16285
rect -15360 16205 -15355 16235
rect -15325 16205 -15320 16235
rect -15360 16155 -15320 16205
rect -15360 16125 -15355 16155
rect -15325 16125 -15320 16155
rect -15360 16075 -15320 16125
rect -15200 16315 -15160 16444
rect -15120 16440 -15080 17120
rect -15040 17116 -15000 17165
rect -14960 17355 -14920 17360
rect -14960 17325 -14955 17355
rect -14925 17325 -14920 17355
rect -14960 17195 -14920 17325
rect -14960 17165 -14955 17195
rect -14925 17165 -14920 17195
rect -14960 17160 -14920 17165
rect -14880 17355 -14840 17360
rect -14880 17325 -14875 17355
rect -14845 17325 -14840 17355
rect -14880 17195 -14840 17325
rect -14880 17165 -14875 17195
rect -14845 17165 -14840 17195
rect -14880 17160 -14840 17165
rect -14800 17355 -14760 17360
rect -14800 17325 -14795 17355
rect -14765 17325 -14760 17355
rect -14800 17195 -14760 17325
rect -14800 17165 -14795 17195
rect -14765 17165 -14760 17195
rect -14800 17160 -14760 17165
rect -14720 17355 -14680 17360
rect -14720 17325 -14715 17355
rect -14685 17325 -14680 17355
rect -14720 17195 -14680 17325
rect -14720 17165 -14715 17195
rect -14685 17165 -14680 17195
rect -14720 17160 -14680 17165
rect -14640 17355 -14600 17360
rect -14640 17325 -14635 17355
rect -14605 17325 -14600 17355
rect -14640 17195 -14600 17325
rect -14640 17165 -14635 17195
rect -14605 17165 -14600 17195
rect -14640 17160 -14600 17165
rect -14560 17355 -14520 17360
rect -14560 17325 -14555 17355
rect -14525 17325 -14520 17355
rect -14560 17195 -14520 17325
rect -14560 17165 -14555 17195
rect -14525 17165 -14520 17195
rect -14560 17160 -14520 17165
rect -14480 17355 -14440 17360
rect -14480 17325 -14475 17355
rect -14445 17325 -14440 17355
rect -14480 17195 -14440 17325
rect -14480 17165 -14475 17195
rect -14445 17165 -14440 17195
rect -14480 17160 -14440 17165
rect -14400 17355 -14360 17360
rect -14400 17325 -14395 17355
rect -14365 17325 -14360 17355
rect -14400 17195 -14360 17325
rect -14400 17165 -14395 17195
rect -14365 17165 -14360 17195
rect -14400 17160 -14360 17165
rect -14320 17355 -14280 17360
rect -14320 17325 -14315 17355
rect -14285 17325 -14280 17355
rect -14320 17195 -14280 17325
rect -14320 17165 -14315 17195
rect -14285 17165 -14280 17195
rect -14320 17160 -14280 17165
rect -14240 17355 -14200 17360
rect -14240 17325 -14235 17355
rect -14205 17325 -14200 17355
rect -14240 17195 -14200 17325
rect -14240 17165 -14235 17195
rect -14205 17165 -14200 17195
rect -14240 17160 -14200 17165
rect -14160 17355 -14120 17360
rect -14160 17325 -14155 17355
rect -14125 17325 -14120 17355
rect -14160 17195 -14120 17325
rect -14160 17165 -14155 17195
rect -14125 17165 -14120 17195
rect -14160 17160 -14120 17165
rect -14080 17355 -14040 17360
rect -14080 17325 -14075 17355
rect -14045 17325 -14040 17355
rect -14080 17195 -14040 17325
rect -14080 17165 -14075 17195
rect -14045 17165 -14040 17195
rect -14080 17160 -14040 17165
rect -14000 17355 -13960 17360
rect -14000 17325 -13995 17355
rect -13965 17325 -13960 17355
rect -14000 17195 -13960 17325
rect -14000 17165 -13995 17195
rect -13965 17165 -13960 17195
rect -14000 17160 -13960 17165
rect -13920 17355 -13880 17360
rect -13920 17325 -13915 17355
rect -13885 17325 -13880 17355
rect -13920 17195 -13880 17325
rect -13920 17165 -13915 17195
rect -13885 17165 -13880 17195
rect -13920 17160 -13880 17165
rect -13840 17355 -13800 17360
rect -13840 17325 -13835 17355
rect -13805 17325 -13800 17355
rect -13840 17195 -13800 17325
rect -13840 17165 -13835 17195
rect -13805 17165 -13800 17195
rect -13840 17160 -13800 17165
rect -13760 17355 -13720 17360
rect -13760 17325 -13755 17355
rect -13725 17325 -13720 17355
rect -13760 17195 -13720 17325
rect -13760 17165 -13755 17195
rect -13725 17165 -13720 17195
rect -13760 17160 -13720 17165
rect -13680 17355 -13640 17360
rect -13680 17325 -13675 17355
rect -13645 17325 -13640 17355
rect -13680 17195 -13640 17325
rect -13680 17165 -13675 17195
rect -13645 17165 -13640 17195
rect -13680 17160 -13640 17165
rect -13600 17355 -13560 17360
rect -13600 17325 -13595 17355
rect -13565 17325 -13560 17355
rect -13600 17195 -13560 17325
rect -13600 17165 -13595 17195
rect -13565 17165 -13560 17195
rect -13600 17160 -13560 17165
rect -13520 17355 -13480 17360
rect -13520 17325 -13515 17355
rect -13485 17325 -13480 17355
rect -13520 17195 -13480 17325
rect -13520 17165 -13515 17195
rect -13485 17165 -13480 17195
rect -13520 17160 -13480 17165
rect -13440 17355 -13400 17360
rect -13440 17325 -13435 17355
rect -13405 17325 -13400 17355
rect -13440 17195 -13400 17325
rect -13440 17165 -13435 17195
rect -13405 17165 -13400 17195
rect -13440 17160 -13400 17165
rect -13360 17355 -13320 17360
rect -13360 17325 -13355 17355
rect -13325 17325 -13320 17355
rect -13360 17195 -13320 17325
rect -13360 17165 -13355 17195
rect -13325 17165 -13320 17195
rect -13360 17160 -13320 17165
rect -13280 17355 -13240 17360
rect -13280 17325 -13275 17355
rect -13245 17325 -13240 17355
rect -13280 17195 -13240 17325
rect -13280 17165 -13275 17195
rect -13245 17165 -13240 17195
rect -13280 17160 -13240 17165
rect -13200 17355 -13160 17360
rect -13200 17325 -13195 17355
rect -13165 17325 -13160 17355
rect -13200 17195 -13160 17325
rect -13200 17165 -13195 17195
rect -13165 17165 -13160 17195
rect -13200 17160 -13160 17165
rect -13120 17355 -13080 17360
rect -13120 17325 -13115 17355
rect -13085 17325 -13080 17355
rect -13120 17195 -13080 17325
rect -13120 17165 -13115 17195
rect -13085 17165 -13080 17195
rect -13120 17160 -13080 17165
rect -13040 17355 -13000 17360
rect -13040 17325 -13035 17355
rect -13005 17325 -13000 17355
rect -13040 17195 -13000 17325
rect -13040 17165 -13035 17195
rect -13005 17165 -13000 17195
rect -13040 17160 -13000 17165
rect -12960 17355 -12920 17360
rect -12960 17325 -12955 17355
rect -12925 17325 -12920 17355
rect -12960 17195 -12920 17325
rect -12960 17165 -12955 17195
rect -12925 17165 -12920 17195
rect -12960 17160 -12920 17165
rect -12880 17355 -12840 17360
rect -12880 17325 -12875 17355
rect -12845 17325 -12840 17355
rect -12880 17195 -12840 17325
rect -12880 17165 -12875 17195
rect -12845 17165 -12840 17195
rect -12880 17160 -12840 17165
rect -12800 17355 -12760 17360
rect -12800 17325 -12795 17355
rect -12765 17325 -12760 17355
rect -12800 17195 -12760 17325
rect -12800 17165 -12795 17195
rect -12765 17165 -12760 17195
rect -12800 17160 -12760 17165
rect -12720 17355 -12680 17360
rect -12720 17325 -12715 17355
rect -12685 17325 -12680 17355
rect -12720 17195 -12680 17325
rect -12720 17165 -12715 17195
rect -12685 17165 -12680 17195
rect -12720 17160 -12680 17165
rect -12640 17355 -12600 17360
rect -12640 17325 -12635 17355
rect -12605 17325 -12600 17355
rect -12640 17195 -12600 17325
rect -12640 17165 -12635 17195
rect -12605 17165 -12600 17195
rect -12640 17160 -12600 17165
rect -12560 17355 -12520 17360
rect -12560 17325 -12555 17355
rect -12525 17325 -12520 17355
rect -12560 17195 -12520 17325
rect -12560 17165 -12555 17195
rect -12525 17165 -12520 17195
rect -12560 17160 -12520 17165
rect -12480 17355 -12440 17360
rect -12480 17325 -12475 17355
rect -12445 17325 -12440 17355
rect -12480 17195 -12440 17325
rect -12480 17165 -12475 17195
rect -12445 17165 -12440 17195
rect -12480 17160 -12440 17165
rect -12400 17355 -12360 17360
rect -12400 17325 -12395 17355
rect -12365 17325 -12360 17355
rect -12400 17195 -12360 17325
rect -12400 17165 -12395 17195
rect -12365 17165 -12360 17195
rect -12400 17160 -12360 17165
rect -12320 17355 -12280 17360
rect -12320 17325 -12315 17355
rect -12285 17325 -12280 17355
rect -12320 17195 -12280 17325
rect -12320 17165 -12315 17195
rect -12285 17165 -12280 17195
rect -12320 17160 -12280 17165
rect -12240 17355 -12200 17360
rect -12240 17325 -12235 17355
rect -12205 17325 -12200 17355
rect -12240 17195 -12200 17325
rect -12240 17165 -12235 17195
rect -12205 17165 -12200 17195
rect -12240 17160 -12200 17165
rect -12160 17355 -12120 17360
rect -12160 17325 -12155 17355
rect -12125 17325 -12120 17355
rect -12160 17195 -12120 17325
rect -12160 17165 -12155 17195
rect -12125 17165 -12120 17195
rect -12160 17160 -12120 17165
rect -12080 17355 -12040 17360
rect -12080 17325 -12075 17355
rect -12045 17325 -12040 17355
rect -12080 17195 -12040 17325
rect -12080 17165 -12075 17195
rect -12045 17165 -12040 17195
rect -12080 17160 -12040 17165
rect -12000 17355 -11960 17360
rect -12000 17325 -11995 17355
rect -11965 17325 -11960 17355
rect -12000 17195 -11960 17325
rect -12000 17165 -11995 17195
rect -11965 17165 -11960 17195
rect -12000 17160 -11960 17165
rect -11920 17355 -11880 17360
rect -11920 17325 -11915 17355
rect -11885 17325 -11880 17355
rect -11920 17195 -11880 17325
rect -11920 17165 -11915 17195
rect -11885 17165 -11880 17195
rect -11920 17160 -11880 17165
rect -11840 17355 -11800 17360
rect -11840 17325 -11835 17355
rect -11805 17325 -11800 17355
rect -11840 17195 -11800 17325
rect -11840 17165 -11835 17195
rect -11805 17165 -11800 17195
rect -11840 17160 -11800 17165
rect -11760 17355 -11720 17360
rect -11760 17325 -11755 17355
rect -11725 17325 -11720 17355
rect -11760 17195 -11720 17325
rect -11760 17165 -11755 17195
rect -11725 17165 -11720 17195
rect -11760 17160 -11720 17165
rect -11680 17355 -11640 17360
rect -11680 17325 -11675 17355
rect -11645 17325 -11640 17355
rect -11680 17195 -11640 17325
rect -11680 17165 -11675 17195
rect -11645 17165 -11640 17195
rect -11680 17160 -11640 17165
rect -11600 17355 -11560 17360
rect -11600 17325 -11595 17355
rect -11565 17325 -11560 17355
rect -11600 17195 -11560 17325
rect -11600 17165 -11595 17195
rect -11565 17165 -11560 17195
rect -11600 17160 -11560 17165
rect -11520 17355 -11480 17360
rect -11520 17325 -11515 17355
rect -11485 17325 -11480 17355
rect -11520 17195 -11480 17325
rect -11520 17165 -11515 17195
rect -11485 17165 -11480 17195
rect -11520 17160 -11480 17165
rect -11440 17355 -11400 17360
rect -11440 17325 -11435 17355
rect -11405 17325 -11400 17355
rect -11440 17195 -11400 17325
rect -11440 17165 -11435 17195
rect -11405 17165 -11400 17195
rect -11440 17160 -11400 17165
rect -11360 17355 -11320 17360
rect -11360 17325 -11355 17355
rect -11325 17325 -11320 17355
rect -11360 17195 -11320 17325
rect -11360 17165 -11355 17195
rect -11325 17165 -11320 17195
rect -11360 17160 -11320 17165
rect -11280 17355 -11240 17360
rect -11280 17325 -11275 17355
rect -11245 17325 -11240 17355
rect -11280 17195 -11240 17325
rect -11280 17165 -11275 17195
rect -11245 17165 -11240 17195
rect -11280 17160 -11240 17165
rect -11200 17355 -11160 17360
rect -11200 17325 -11195 17355
rect -11165 17325 -11160 17355
rect -11200 17195 -11160 17325
rect -11200 17165 -11195 17195
rect -11165 17165 -11160 17195
rect -11200 17160 -11160 17165
rect -11120 17355 -11080 17360
rect -11120 17325 -11115 17355
rect -11085 17325 -11080 17355
rect -11120 17195 -11080 17325
rect -11120 17165 -11115 17195
rect -11085 17165 -11080 17195
rect -11120 17160 -11080 17165
rect -11040 17355 -11000 17360
rect -11040 17325 -11035 17355
rect -11005 17325 -11000 17355
rect -11040 17195 -11000 17325
rect -11040 17165 -11035 17195
rect -11005 17165 -11000 17195
rect -11040 17160 -11000 17165
rect -10960 17355 -10920 17360
rect -10960 17325 -10955 17355
rect -10925 17325 -10920 17355
rect -10960 17195 -10920 17325
rect -10960 17165 -10955 17195
rect -10925 17165 -10920 17195
rect -10960 17160 -10920 17165
rect -10880 17355 -10840 17360
rect -10880 17325 -10875 17355
rect -10845 17325 -10840 17355
rect -10880 17195 -10840 17325
rect -10880 17165 -10875 17195
rect -10845 17165 -10840 17195
rect -10880 17160 -10840 17165
rect -10800 17355 -10760 17360
rect -10800 17325 -10795 17355
rect -10765 17325 -10760 17355
rect -10800 17195 -10760 17325
rect -10800 17165 -10795 17195
rect -10765 17165 -10760 17195
rect -10800 17160 -10760 17165
rect -10720 17355 -10680 17360
rect -10720 17325 -10715 17355
rect -10685 17325 -10680 17355
rect -10720 17195 -10680 17325
rect -10720 17165 -10715 17195
rect -10685 17165 -10680 17195
rect -10720 17160 -10680 17165
rect -10640 17355 -10600 17360
rect -10640 17325 -10635 17355
rect -10605 17325 -10600 17355
rect -10640 17195 -10600 17325
rect -10640 17165 -10635 17195
rect -10605 17165 -10600 17195
rect -10640 17160 -10600 17165
rect -10560 17355 -10520 17360
rect -10560 17325 -10555 17355
rect -10525 17325 -10520 17355
rect -10560 17195 -10520 17325
rect -10560 17165 -10555 17195
rect -10525 17165 -10520 17195
rect -10560 17160 -10520 17165
rect -10480 17355 -10440 17360
rect -10480 17325 -10475 17355
rect -10445 17325 -10440 17355
rect -10480 17195 -10440 17325
rect -10480 17165 -10475 17195
rect -10445 17165 -10440 17195
rect -10480 17160 -10440 17165
rect -10400 17355 -10360 17360
rect -10400 17325 -10395 17355
rect -10365 17325 -10360 17355
rect -10400 17195 -10360 17325
rect -10400 17165 -10395 17195
rect -10365 17165 -10360 17195
rect -10400 17160 -10360 17165
rect -10320 17355 -10280 17360
rect -10320 17325 -10315 17355
rect -10285 17325 -10280 17355
rect -10320 17195 -10280 17325
rect -10320 17165 -10315 17195
rect -10285 17165 -10280 17195
rect -10320 17160 -10280 17165
rect -10240 17355 -10200 17360
rect -10240 17325 -10235 17355
rect -10205 17325 -10200 17355
rect -10240 17195 -10200 17325
rect -10240 17165 -10235 17195
rect -10205 17165 -10200 17195
rect -10240 17160 -10200 17165
rect -10160 17355 -10120 17360
rect -10160 17325 -10155 17355
rect -10125 17325 -10120 17355
rect -10160 17195 -10120 17325
rect -10160 17165 -10155 17195
rect -10125 17165 -10120 17195
rect -10160 17160 -10120 17165
rect -10080 17355 -10040 17360
rect -10080 17325 -10075 17355
rect -10045 17325 -10040 17355
rect -10080 17195 -10040 17325
rect -10080 17165 -10075 17195
rect -10045 17165 -10040 17195
rect -10080 17160 -10040 17165
rect -10000 17355 -9960 17360
rect -10000 17325 -9995 17355
rect -9965 17325 -9960 17355
rect -10000 17195 -9960 17325
rect -10000 17165 -9995 17195
rect -9965 17165 -9960 17195
rect -10000 17160 -9960 17165
rect -9920 17355 -9880 17360
rect -9920 17325 -9915 17355
rect -9885 17325 -9880 17355
rect -9920 17195 -9880 17325
rect -9920 17165 -9915 17195
rect -9885 17165 -9880 17195
rect -9920 17160 -9880 17165
rect -9840 17355 -9800 17360
rect -9840 17325 -9835 17355
rect -9805 17325 -9800 17355
rect -9840 17195 -9800 17325
rect -9840 17165 -9835 17195
rect -9805 17165 -9800 17195
rect -9840 17160 -9800 17165
rect -9760 17355 -9720 17360
rect -9760 17325 -9755 17355
rect -9725 17325 -9720 17355
rect -9760 17195 -9720 17325
rect -9760 17165 -9755 17195
rect -9725 17165 -9720 17195
rect -9760 17160 -9720 17165
rect -9680 17355 -9640 17360
rect -9680 17325 -9675 17355
rect -9645 17325 -9640 17355
rect -9680 17195 -9640 17325
rect -9680 17165 -9675 17195
rect -9645 17165 -9640 17195
rect -9680 17160 -9640 17165
rect -9600 17355 -9560 17360
rect -9600 17325 -9595 17355
rect -9565 17325 -9560 17355
rect -9600 17195 -9560 17325
rect -9600 17165 -9595 17195
rect -9565 17165 -9560 17195
rect -9600 17160 -9560 17165
rect -9520 17355 -9480 17360
rect -9520 17325 -9515 17355
rect -9485 17325 -9480 17355
rect -9520 17195 -9480 17325
rect -9520 17165 -9515 17195
rect -9485 17165 -9480 17195
rect -9520 17160 -9480 17165
rect -9440 17355 -9400 17360
rect -9440 17325 -9435 17355
rect -9405 17325 -9400 17355
rect -9440 17195 -9400 17325
rect -9440 17165 -9435 17195
rect -9405 17165 -9400 17195
rect -9440 17160 -9400 17165
rect -9360 17355 -9320 17360
rect -9360 17325 -9355 17355
rect -9325 17325 -9320 17355
rect -9360 17195 -9320 17325
rect -9360 17165 -9355 17195
rect -9325 17165 -9320 17195
rect -9360 17160 -9320 17165
rect -9280 17355 -9240 17360
rect -9280 17325 -9275 17355
rect -9245 17325 -9240 17355
rect -9280 17195 -9240 17325
rect -9280 17165 -9275 17195
rect -9245 17165 -9240 17195
rect -9280 17160 -9240 17165
rect -9200 17355 -9160 17360
rect -9200 17325 -9195 17355
rect -9165 17325 -9160 17355
rect -9200 17195 -9160 17325
rect -9200 17165 -9195 17195
rect -9165 17165 -9160 17195
rect -9200 17160 -9160 17165
rect -9120 17355 -9080 17360
rect -9120 17325 -9115 17355
rect -9085 17325 -9080 17355
rect -9120 17195 -9080 17325
rect -9120 17165 -9115 17195
rect -9085 17165 -9080 17195
rect -9120 17160 -9080 17165
rect -9040 17355 -9000 17360
rect -9040 17325 -9035 17355
rect -9005 17325 -9000 17355
rect -9040 17195 -9000 17325
rect -9040 17165 -9035 17195
rect -9005 17165 -9000 17195
rect -9040 17160 -9000 17165
rect -8960 17355 -8920 17360
rect -8960 17325 -8955 17355
rect -8925 17325 -8920 17355
rect -8960 17195 -8920 17325
rect -8960 17165 -8955 17195
rect -8925 17165 -8920 17195
rect -8960 17160 -8920 17165
rect -8880 17355 -8840 17360
rect -8880 17325 -8875 17355
rect -8845 17325 -8840 17355
rect -8880 17195 -8840 17325
rect -8880 17165 -8875 17195
rect -8845 17165 -8840 17195
rect -8880 17160 -8840 17165
rect -8800 17355 -8760 17360
rect -8800 17325 -8795 17355
rect -8765 17325 -8760 17355
rect -8800 17195 -8760 17325
rect -8800 17165 -8795 17195
rect -8765 17165 -8760 17195
rect -8800 17160 -8760 17165
rect -8720 17355 -8680 17360
rect -8720 17325 -8715 17355
rect -8685 17325 -8680 17355
rect -8720 17195 -8680 17325
rect -8720 17165 -8715 17195
rect -8685 17165 -8680 17195
rect -8720 17160 -8680 17165
rect -8640 17355 -8600 17360
rect -8640 17325 -8635 17355
rect -8605 17325 -8600 17355
rect -8640 17195 -8600 17325
rect -8640 17165 -8635 17195
rect -8605 17165 -8600 17195
rect -8640 17160 -8600 17165
rect -8560 17355 -8520 17360
rect -8560 17325 -8555 17355
rect -8525 17325 -8520 17355
rect -8560 17195 -8520 17325
rect -8560 17165 -8555 17195
rect -8525 17165 -8520 17195
rect -8560 17160 -8520 17165
rect -8480 17355 -8440 17360
rect -8480 17325 -8475 17355
rect -8445 17325 -8440 17355
rect -8480 17195 -8440 17325
rect -8480 17165 -8475 17195
rect -8445 17165 -8440 17195
rect -8480 17160 -8440 17165
rect -8400 17355 -8360 17360
rect -8400 17325 -8395 17355
rect -8365 17325 -8360 17355
rect -8400 17195 -8360 17325
rect -8400 17165 -8395 17195
rect -8365 17165 -8360 17195
rect -8400 17160 -8360 17165
rect -8320 17355 -8280 17360
rect -8320 17325 -8315 17355
rect -8285 17325 -8280 17355
rect -8320 17195 -8280 17325
rect -8320 17165 -8315 17195
rect -8285 17165 -8280 17195
rect -8320 17160 -8280 17165
rect -8240 17355 -8200 17360
rect -8240 17325 -8235 17355
rect -8205 17325 -8200 17355
rect -8240 17195 -8200 17325
rect -8240 17165 -8235 17195
rect -8205 17165 -8200 17195
rect -8240 17160 -8200 17165
rect -8160 17355 -8120 17360
rect -8160 17325 -8155 17355
rect -8125 17325 -8120 17355
rect -8160 17195 -8120 17325
rect -8160 17165 -8155 17195
rect -8125 17165 -8120 17195
rect -8160 17160 -8120 17165
rect -8080 17355 -8040 17360
rect -8080 17325 -8075 17355
rect -8045 17325 -8040 17355
rect -8080 17195 -8040 17325
rect -8080 17165 -8075 17195
rect -8045 17165 -8040 17195
rect -8080 17160 -8040 17165
rect -8000 17355 -7960 17360
rect -8000 17325 -7995 17355
rect -7965 17325 -7960 17355
rect -8000 17195 -7960 17325
rect -8000 17165 -7995 17195
rect -7965 17165 -7960 17195
rect -8000 17160 -7960 17165
rect -7920 17355 -7880 17360
rect -7920 17325 -7915 17355
rect -7885 17325 -7880 17355
rect -7920 17195 -7880 17325
rect -7920 17165 -7915 17195
rect -7885 17165 -7880 17195
rect -7920 17160 -7880 17165
rect -7840 17355 -7800 17360
rect -7840 17325 -7835 17355
rect -7805 17325 -7800 17355
rect -7840 17195 -7800 17325
rect -7840 17165 -7835 17195
rect -7805 17165 -7800 17195
rect -7840 17160 -7800 17165
rect -7760 17355 -7720 17360
rect -7760 17325 -7755 17355
rect -7725 17325 -7720 17355
rect -7760 17195 -7720 17325
rect -7760 17165 -7755 17195
rect -7725 17165 -7720 17195
rect -7760 17160 -7720 17165
rect -7680 17355 -7640 17360
rect -7680 17325 -7675 17355
rect -7645 17325 -7640 17355
rect -7680 17195 -7640 17325
rect -7680 17165 -7675 17195
rect -7645 17165 -7640 17195
rect -7680 17160 -7640 17165
rect -7600 17355 -7560 17360
rect -7600 17325 -7595 17355
rect -7565 17325 -7560 17355
rect -7600 17195 -7560 17325
rect -7600 17165 -7595 17195
rect -7565 17165 -7560 17195
rect -7600 17160 -7560 17165
rect -7520 17355 -7480 17360
rect -7520 17325 -7515 17355
rect -7485 17325 -7480 17355
rect -7520 17195 -7480 17325
rect -7520 17165 -7515 17195
rect -7485 17165 -7480 17195
rect -7520 17160 -7480 17165
rect -7440 17355 -7400 17360
rect -7440 17325 -7435 17355
rect -7405 17325 -7400 17355
rect -7440 17195 -7400 17325
rect -7440 17165 -7435 17195
rect -7405 17165 -7400 17195
rect -7440 17160 -7400 17165
rect -7360 17355 -7320 17360
rect -7360 17325 -7355 17355
rect -7325 17325 -7320 17355
rect -7360 17195 -7320 17325
rect -7360 17165 -7355 17195
rect -7325 17165 -7320 17195
rect -7360 17160 -7320 17165
rect -7280 17355 -7240 17360
rect -7280 17325 -7275 17355
rect -7245 17325 -7240 17355
rect -7280 17195 -7240 17325
rect -7280 17165 -7275 17195
rect -7245 17165 -7240 17195
rect -7280 17160 -7240 17165
rect -7200 17355 -7160 17360
rect -7200 17325 -7195 17355
rect -7165 17325 -7160 17355
rect -7200 17195 -7160 17325
rect -7200 17165 -7195 17195
rect -7165 17165 -7160 17195
rect -7200 17160 -7160 17165
rect -7120 17355 -7080 17360
rect -7120 17325 -7115 17355
rect -7085 17325 -7080 17355
rect -7120 17195 -7080 17325
rect -7120 17165 -7115 17195
rect -7085 17165 -7080 17195
rect -7120 17160 -7080 17165
rect -7040 17355 -7000 17360
rect -7040 17325 -7035 17355
rect -7005 17325 -7000 17355
rect -7040 17195 -7000 17325
rect -7040 17165 -7035 17195
rect -7005 17165 -7000 17195
rect -7040 17160 -7000 17165
rect -6960 17355 -6920 17360
rect -6960 17325 -6955 17355
rect -6925 17325 -6920 17355
rect -6960 17195 -6920 17325
rect -6960 17165 -6955 17195
rect -6925 17165 -6920 17195
rect -6960 17160 -6920 17165
rect -6880 17355 -6840 17360
rect -6880 17325 -6875 17355
rect -6845 17325 -6840 17355
rect -6880 17195 -6840 17325
rect -6880 17165 -6875 17195
rect -6845 17165 -6840 17195
rect -6880 17160 -6840 17165
rect -6800 17355 -6760 17360
rect -6800 17325 -6795 17355
rect -6765 17325 -6760 17355
rect -6800 17195 -6760 17325
rect -6800 17165 -6795 17195
rect -6765 17165 -6760 17195
rect -6800 17160 -6760 17165
rect -6720 17355 -6680 17360
rect -6720 17325 -6715 17355
rect -6685 17325 -6680 17355
rect -6720 17195 -6680 17325
rect -6720 17165 -6715 17195
rect -6685 17165 -6680 17195
rect -6720 17160 -6680 17165
rect -6640 17355 -6600 17360
rect -6640 17325 -6635 17355
rect -6605 17325 -6600 17355
rect -6640 17195 -6600 17325
rect -6640 17165 -6635 17195
rect -6605 17165 -6600 17195
rect -6640 17160 -6600 17165
rect -6560 17355 -6520 17360
rect -6560 17325 -6555 17355
rect -6525 17325 -6520 17355
rect -6560 17195 -6520 17325
rect -6560 17165 -6555 17195
rect -6525 17165 -6520 17195
rect -6560 17160 -6520 17165
rect -6480 17355 -6440 17360
rect -6480 17325 -6475 17355
rect -6445 17325 -6440 17355
rect -6480 17195 -6440 17325
rect -6480 17165 -6475 17195
rect -6445 17165 -6440 17195
rect -6480 17160 -6440 17165
rect -6400 17355 -6360 17360
rect -6400 17325 -6395 17355
rect -6365 17325 -6360 17355
rect -6400 17195 -6360 17325
rect -6400 17165 -6395 17195
rect -6365 17165 -6360 17195
rect -6400 17160 -6360 17165
rect -6320 17355 -6280 17360
rect -6320 17325 -6315 17355
rect -6285 17325 -6280 17355
rect -6320 17195 -6280 17325
rect -6320 17165 -6315 17195
rect -6285 17165 -6280 17195
rect -6320 17160 -6280 17165
rect -6240 17355 -6200 17360
rect -6240 17325 -6235 17355
rect -6205 17325 -6200 17355
rect -6240 17195 -6200 17325
rect -6240 17165 -6235 17195
rect -6205 17165 -6200 17195
rect -6240 17160 -6200 17165
rect -6160 17355 -6120 17360
rect -6160 17325 -6155 17355
rect -6125 17325 -6120 17355
rect -6160 17195 -6120 17325
rect -6160 17165 -6155 17195
rect -6125 17165 -6120 17195
rect -6160 17160 -6120 17165
rect -6080 17355 -6040 17440
rect -6080 17325 -6075 17355
rect -6045 17325 -6040 17355
rect -6080 17195 -6040 17325
rect -6080 17165 -6075 17195
rect -6045 17165 -6040 17195
rect -6080 17160 -6040 17165
rect -6000 17355 -5960 17360
rect -6000 17325 -5995 17355
rect -5965 17325 -5960 17355
rect -6000 17195 -5960 17325
rect -6000 17165 -5995 17195
rect -5965 17165 -5960 17195
rect -6000 17160 -5960 17165
rect -5920 17355 -5880 17440
rect -5920 17325 -5915 17355
rect -5885 17325 -5880 17355
rect -5920 17195 -5880 17325
rect -5920 17165 -5915 17195
rect -5885 17165 -5880 17195
rect -5920 17160 -5880 17165
rect -5840 17355 -5800 17360
rect -5840 17325 -5835 17355
rect -5805 17325 -5800 17355
rect -5840 17195 -5800 17325
rect -5840 17165 -5835 17195
rect -5805 17165 -5800 17195
rect -5840 17160 -5800 17165
rect -5760 17355 -5720 17440
rect -5760 17325 -5755 17355
rect -5725 17325 -5720 17355
rect -5760 17195 -5720 17325
rect -5760 17165 -5755 17195
rect -5725 17165 -5720 17195
rect -5760 17160 -5720 17165
rect -15040 17084 -15036 17116
rect -15004 17084 -15000 17116
rect -15040 17036 -15000 17084
rect -15040 17004 -15036 17036
rect -15004 17004 -15000 17036
rect -15040 16956 -15000 17004
rect -15040 16924 -15036 16956
rect -15004 16924 -15000 16956
rect -15040 16876 -15000 16924
rect -15040 16844 -15036 16876
rect -15004 16844 -15000 16876
rect -15040 16796 -15000 16844
rect -15040 16764 -15036 16796
rect -15004 16764 -15000 16796
rect -15040 16716 -15000 16764
rect -15040 16684 -15036 16716
rect -15004 16684 -15000 16716
rect -15040 16636 -15000 16684
rect -15040 16604 -15036 16636
rect -15004 16604 -15000 16636
rect -15040 16556 -15000 16604
rect -15040 16524 -15036 16556
rect -15004 16524 -15000 16556
rect -15040 16476 -15000 16524
rect -15040 16444 -15036 16476
rect -15004 16444 -15000 16476
rect -15200 16285 -15195 16315
rect -15165 16285 -15160 16315
rect -15200 16155 -15160 16285
rect -15040 16315 -15000 16444
rect -15040 16285 -15035 16315
rect -15005 16285 -15000 16315
rect -15200 16125 -15195 16155
rect -15165 16125 -15160 16155
rect -15360 16045 -15355 16075
rect -15325 16045 -15320 16075
rect -15360 15995 -15320 16045
rect -15360 15965 -15355 15995
rect -15325 15965 -15320 15995
rect -15360 15920 -15320 15965
rect -15280 16075 -15240 16080
rect -15280 16045 -15275 16075
rect -15245 16045 -15240 16075
rect -15280 15920 -15240 16045
rect -15200 15995 -15160 16125
rect -15200 15965 -15195 15995
rect -15165 15965 -15160 15995
rect -15200 15920 -15160 15965
rect -15120 16235 -15080 16240
rect -15120 16205 -15115 16235
rect -15085 16205 -15080 16235
rect -15120 15920 -15080 16205
rect -15040 16155 -15000 16285
rect -15040 16125 -15035 16155
rect -15005 16125 -15000 16155
rect -15040 15995 -15000 16125
rect -15040 15965 -15035 15995
rect -15005 15965 -15000 15995
rect -15040 15920 -15000 15965
rect -14960 16475 -14920 16480
rect -14960 16445 -14955 16475
rect -14925 16445 -14920 16475
rect -14960 16315 -14920 16445
rect -14960 16285 -14955 16315
rect -14925 16285 -14920 16315
rect -14960 16155 -14920 16285
rect -14960 16125 -14955 16155
rect -14925 16125 -14920 16155
rect -14960 15995 -14920 16125
rect -14960 15965 -14955 15995
rect -14925 15965 -14920 15995
rect -14960 15960 -14920 15965
rect -14880 16475 -14840 16480
rect -14880 16445 -14875 16475
rect -14845 16445 -14840 16475
rect -14880 16315 -14840 16445
rect -14880 16285 -14875 16315
rect -14845 16285 -14840 16315
rect -14880 16155 -14840 16285
rect -14880 16125 -14875 16155
rect -14845 16125 -14840 16155
rect -14880 15995 -14840 16125
rect -14880 15965 -14875 15995
rect -14845 15965 -14840 15995
rect -14880 15960 -14840 15965
rect -14800 16475 -14760 16480
rect -14800 16445 -14795 16475
rect -14765 16445 -14760 16475
rect -14800 16315 -14760 16445
rect -14800 16285 -14795 16315
rect -14765 16285 -14760 16315
rect -14800 16155 -14760 16285
rect -14800 16125 -14795 16155
rect -14765 16125 -14760 16155
rect -14800 15995 -14760 16125
rect -14800 15965 -14795 15995
rect -14765 15965 -14760 15995
rect -14800 15960 -14760 15965
rect -14720 16475 -14680 16480
rect -14720 16445 -14715 16475
rect -14685 16445 -14680 16475
rect -14720 16315 -14680 16445
rect -14720 16285 -14715 16315
rect -14685 16285 -14680 16315
rect -14720 16155 -14680 16285
rect -14720 16125 -14715 16155
rect -14685 16125 -14680 16155
rect -14720 15995 -14680 16125
rect -14720 15965 -14715 15995
rect -14685 15965 -14680 15995
rect -14720 15960 -14680 15965
rect -14640 16475 -14600 16480
rect -14640 16445 -14635 16475
rect -14605 16445 -14600 16475
rect -14640 16315 -14600 16445
rect -14640 16285 -14635 16315
rect -14605 16285 -14600 16315
rect -14640 16155 -14600 16285
rect -14640 16125 -14635 16155
rect -14605 16125 -14600 16155
rect -14640 15995 -14600 16125
rect -14640 15965 -14635 15995
rect -14605 15965 -14600 15995
rect -14640 15960 -14600 15965
rect -14560 16475 -14520 16480
rect -14560 16445 -14555 16475
rect -14525 16445 -14520 16475
rect -14560 16315 -14520 16445
rect -14560 16285 -14555 16315
rect -14525 16285 -14520 16315
rect -14560 16155 -14520 16285
rect -14560 16125 -14555 16155
rect -14525 16125 -14520 16155
rect -14560 15995 -14520 16125
rect -14560 15965 -14555 15995
rect -14525 15965 -14520 15995
rect -14560 15960 -14520 15965
rect -14480 16475 -14440 16480
rect -14480 16445 -14475 16475
rect -14445 16445 -14440 16475
rect -14480 16315 -14440 16445
rect -14480 16285 -14475 16315
rect -14445 16285 -14440 16315
rect -14480 16155 -14440 16285
rect -14480 16125 -14475 16155
rect -14445 16125 -14440 16155
rect -14480 15995 -14440 16125
rect -14480 15965 -14475 15995
rect -14445 15965 -14440 15995
rect -14480 15960 -14440 15965
rect -14400 16475 -14360 16480
rect -14400 16445 -14395 16475
rect -14365 16445 -14360 16475
rect -14400 16315 -14360 16445
rect -14400 16285 -14395 16315
rect -14365 16285 -14360 16315
rect -14400 16155 -14360 16285
rect -14400 16125 -14395 16155
rect -14365 16125 -14360 16155
rect -14400 15995 -14360 16125
rect -14400 15965 -14395 15995
rect -14365 15965 -14360 15995
rect -14400 15960 -14360 15965
rect -14320 16475 -14280 16480
rect -14320 16445 -14315 16475
rect -14285 16445 -14280 16475
rect -14320 16315 -14280 16445
rect -14320 16285 -14315 16315
rect -14285 16285 -14280 16315
rect -14320 16155 -14280 16285
rect -14320 16125 -14315 16155
rect -14285 16125 -14280 16155
rect -14320 15995 -14280 16125
rect -14320 15965 -14315 15995
rect -14285 15965 -14280 15995
rect -14320 15960 -14280 15965
rect -14240 16475 -14200 16480
rect -14240 16445 -14235 16475
rect -14205 16445 -14200 16475
rect -14240 16315 -14200 16445
rect -14240 16285 -14235 16315
rect -14205 16285 -14200 16315
rect -14240 16155 -14200 16285
rect -14240 16125 -14235 16155
rect -14205 16125 -14200 16155
rect -14240 15995 -14200 16125
rect -14240 15965 -14235 15995
rect -14205 15965 -14200 15995
rect -14240 15960 -14200 15965
rect -14160 16475 -14120 16480
rect -14160 16445 -14155 16475
rect -14125 16445 -14120 16475
rect -14160 16315 -14120 16445
rect -14160 16285 -14155 16315
rect -14125 16285 -14120 16315
rect -14160 16155 -14120 16285
rect -14160 16125 -14155 16155
rect -14125 16125 -14120 16155
rect -14160 15995 -14120 16125
rect -14160 15965 -14155 15995
rect -14125 15965 -14120 15995
rect -14160 15960 -14120 15965
rect -14080 16475 -14040 16480
rect -14080 16445 -14075 16475
rect -14045 16445 -14040 16475
rect -14080 16315 -14040 16445
rect -14080 16285 -14075 16315
rect -14045 16285 -14040 16315
rect -14080 16155 -14040 16285
rect -14080 16125 -14075 16155
rect -14045 16125 -14040 16155
rect -14080 15995 -14040 16125
rect -14080 15965 -14075 15995
rect -14045 15965 -14040 15995
rect -14080 15960 -14040 15965
rect -14000 16475 -13960 16480
rect -14000 16445 -13995 16475
rect -13965 16445 -13960 16475
rect -14000 16315 -13960 16445
rect -14000 16285 -13995 16315
rect -13965 16285 -13960 16315
rect -14000 16155 -13960 16285
rect -14000 16125 -13995 16155
rect -13965 16125 -13960 16155
rect -14000 15995 -13960 16125
rect -14000 15965 -13995 15995
rect -13965 15965 -13960 15995
rect -14000 15960 -13960 15965
rect -13920 16475 -13880 16480
rect -13920 16445 -13915 16475
rect -13885 16445 -13880 16475
rect -13920 16315 -13880 16445
rect -13920 16285 -13915 16315
rect -13885 16285 -13880 16315
rect -13920 16155 -13880 16285
rect -13920 16125 -13915 16155
rect -13885 16125 -13880 16155
rect -13920 15995 -13880 16125
rect -13920 15965 -13915 15995
rect -13885 15965 -13880 15995
rect -13920 15960 -13880 15965
rect -13840 16475 -13800 16480
rect -13840 16445 -13835 16475
rect -13805 16445 -13800 16475
rect -13840 16315 -13800 16445
rect -13840 16285 -13835 16315
rect -13805 16285 -13800 16315
rect -13840 16155 -13800 16285
rect -13840 16125 -13835 16155
rect -13805 16125 -13800 16155
rect -13840 15995 -13800 16125
rect -13840 15965 -13835 15995
rect -13805 15965 -13800 15995
rect -13840 15960 -13800 15965
rect -13760 16475 -13720 16480
rect -13760 16445 -13755 16475
rect -13725 16445 -13720 16475
rect -13760 16315 -13720 16445
rect -13760 16285 -13755 16315
rect -13725 16285 -13720 16315
rect -13760 16155 -13720 16285
rect -13760 16125 -13755 16155
rect -13725 16125 -13720 16155
rect -13760 15995 -13720 16125
rect -13760 15965 -13755 15995
rect -13725 15965 -13720 15995
rect -13760 15960 -13720 15965
rect -13680 16475 -13640 16480
rect -13680 16445 -13675 16475
rect -13645 16445 -13640 16475
rect -13680 16315 -13640 16445
rect -13680 16285 -13675 16315
rect -13645 16285 -13640 16315
rect -13680 16155 -13640 16285
rect -13680 16125 -13675 16155
rect -13645 16125 -13640 16155
rect -13680 15995 -13640 16125
rect -13680 15965 -13675 15995
rect -13645 15965 -13640 15995
rect -13680 15960 -13640 15965
rect -13600 16475 -13560 16480
rect -13600 16445 -13595 16475
rect -13565 16445 -13560 16475
rect -13600 16315 -13560 16445
rect -13600 16285 -13595 16315
rect -13565 16285 -13560 16315
rect -13600 16155 -13560 16285
rect -13600 16125 -13595 16155
rect -13565 16125 -13560 16155
rect -13600 15995 -13560 16125
rect -13600 15965 -13595 15995
rect -13565 15965 -13560 15995
rect -13600 15960 -13560 15965
rect -13520 16475 -13480 16480
rect -13520 16445 -13515 16475
rect -13485 16445 -13480 16475
rect -13520 16315 -13480 16445
rect -13520 16285 -13515 16315
rect -13485 16285 -13480 16315
rect -13520 16155 -13480 16285
rect -13520 16125 -13515 16155
rect -13485 16125 -13480 16155
rect -13520 15995 -13480 16125
rect -13520 15965 -13515 15995
rect -13485 15965 -13480 15995
rect -13520 15960 -13480 15965
rect -13440 16475 -13400 16480
rect -13440 16445 -13435 16475
rect -13405 16445 -13400 16475
rect -13440 16315 -13400 16445
rect -13440 16285 -13435 16315
rect -13405 16285 -13400 16315
rect -13440 16155 -13400 16285
rect -13440 16125 -13435 16155
rect -13405 16125 -13400 16155
rect -13440 15995 -13400 16125
rect -13440 15965 -13435 15995
rect -13405 15965 -13400 15995
rect -13440 15960 -13400 15965
rect -13360 16475 -13320 16480
rect -13360 16445 -13355 16475
rect -13325 16445 -13320 16475
rect -13360 16315 -13320 16445
rect -13360 16285 -13355 16315
rect -13325 16285 -13320 16315
rect -13360 16155 -13320 16285
rect -13360 16125 -13355 16155
rect -13325 16125 -13320 16155
rect -13360 15995 -13320 16125
rect -13360 15965 -13355 15995
rect -13325 15965 -13320 15995
rect -13360 15960 -13320 15965
rect -13280 16475 -13240 16480
rect -13280 16445 -13275 16475
rect -13245 16445 -13240 16475
rect -13280 16315 -13240 16445
rect -13280 16285 -13275 16315
rect -13245 16285 -13240 16315
rect -13280 16155 -13240 16285
rect -13280 16125 -13275 16155
rect -13245 16125 -13240 16155
rect -13280 15995 -13240 16125
rect -13280 15965 -13275 15995
rect -13245 15965 -13240 15995
rect -13280 15960 -13240 15965
rect -13200 16475 -13160 16480
rect -13200 16445 -13195 16475
rect -13165 16445 -13160 16475
rect -13200 16315 -13160 16445
rect -13200 16285 -13195 16315
rect -13165 16285 -13160 16315
rect -13200 16155 -13160 16285
rect -13200 16125 -13195 16155
rect -13165 16125 -13160 16155
rect -13200 15995 -13160 16125
rect -13200 15965 -13195 15995
rect -13165 15965 -13160 15995
rect -13200 15960 -13160 15965
rect -13120 16475 -13080 16480
rect -13120 16445 -13115 16475
rect -13085 16445 -13080 16475
rect -13120 16315 -13080 16445
rect -13120 16285 -13115 16315
rect -13085 16285 -13080 16315
rect -13120 16155 -13080 16285
rect -13120 16125 -13115 16155
rect -13085 16125 -13080 16155
rect -13120 15995 -13080 16125
rect -13120 15965 -13115 15995
rect -13085 15965 -13080 15995
rect -13120 15960 -13080 15965
rect -13040 16475 -13000 16480
rect -13040 16445 -13035 16475
rect -13005 16445 -13000 16475
rect -13040 16315 -13000 16445
rect -13040 16285 -13035 16315
rect -13005 16285 -13000 16315
rect -13040 16155 -13000 16285
rect -13040 16125 -13035 16155
rect -13005 16125 -13000 16155
rect -13040 15995 -13000 16125
rect -13040 15965 -13035 15995
rect -13005 15965 -13000 15995
rect -13040 15960 -13000 15965
rect -12960 16475 -12920 16480
rect -12960 16445 -12955 16475
rect -12925 16445 -12920 16475
rect -12960 16315 -12920 16445
rect -12960 16285 -12955 16315
rect -12925 16285 -12920 16315
rect -12960 16155 -12920 16285
rect -12960 16125 -12955 16155
rect -12925 16125 -12920 16155
rect -12960 15995 -12920 16125
rect -12960 15965 -12955 15995
rect -12925 15965 -12920 15995
rect -12960 15960 -12920 15965
rect -12880 16475 -12840 16480
rect -12880 16445 -12875 16475
rect -12845 16445 -12840 16475
rect -12880 16315 -12840 16445
rect -12880 16285 -12875 16315
rect -12845 16285 -12840 16315
rect -12880 16155 -12840 16285
rect -12880 16125 -12875 16155
rect -12845 16125 -12840 16155
rect -12880 15995 -12840 16125
rect -12880 15965 -12875 15995
rect -12845 15965 -12840 15995
rect -12880 15960 -12840 15965
rect -12800 16475 -12760 16480
rect -12800 16445 -12795 16475
rect -12765 16445 -12760 16475
rect -12800 16315 -12760 16445
rect -12800 16285 -12795 16315
rect -12765 16285 -12760 16315
rect -12800 16155 -12760 16285
rect -12800 16125 -12795 16155
rect -12765 16125 -12760 16155
rect -12800 15995 -12760 16125
rect -12800 15965 -12795 15995
rect -12765 15965 -12760 15995
rect -12800 15960 -12760 15965
rect -12720 16475 -12680 16480
rect -12720 16445 -12715 16475
rect -12685 16445 -12680 16475
rect -12720 16315 -12680 16445
rect -12720 16285 -12715 16315
rect -12685 16285 -12680 16315
rect -12720 16155 -12680 16285
rect -12720 16125 -12715 16155
rect -12685 16125 -12680 16155
rect -12720 15995 -12680 16125
rect -12720 15965 -12715 15995
rect -12685 15965 -12680 15995
rect -12720 15960 -12680 15965
rect -12640 16475 -12600 16480
rect -12640 16445 -12635 16475
rect -12605 16445 -12600 16475
rect -12640 16315 -12600 16445
rect -12640 16285 -12635 16315
rect -12605 16285 -12600 16315
rect -12640 16155 -12600 16285
rect -12640 16125 -12635 16155
rect -12605 16125 -12600 16155
rect -12640 15995 -12600 16125
rect -12640 15965 -12635 15995
rect -12605 15965 -12600 15995
rect -12640 15960 -12600 15965
rect -12560 16475 -12520 16480
rect -12560 16445 -12555 16475
rect -12525 16445 -12520 16475
rect -12560 16315 -12520 16445
rect -12560 16285 -12555 16315
rect -12525 16285 -12520 16315
rect -12560 16155 -12520 16285
rect -12560 16125 -12555 16155
rect -12525 16125 -12520 16155
rect -12560 15995 -12520 16125
rect -12560 15965 -12555 15995
rect -12525 15965 -12520 15995
rect -12560 15960 -12520 15965
rect -12480 16475 -12440 16480
rect -12480 16445 -12475 16475
rect -12445 16445 -12440 16475
rect -12480 16315 -12440 16445
rect -12480 16285 -12475 16315
rect -12445 16285 -12440 16315
rect -12480 16155 -12440 16285
rect -12480 16125 -12475 16155
rect -12445 16125 -12440 16155
rect -12480 15995 -12440 16125
rect -12480 15965 -12475 15995
rect -12445 15965 -12440 15995
rect -12480 15960 -12440 15965
rect -12400 16475 -12360 16480
rect -12400 16445 -12395 16475
rect -12365 16445 -12360 16475
rect -12400 16315 -12360 16445
rect -12400 16285 -12395 16315
rect -12365 16285 -12360 16315
rect -12400 16155 -12360 16285
rect -12400 16125 -12395 16155
rect -12365 16125 -12360 16155
rect -12400 15995 -12360 16125
rect -12400 15965 -12395 15995
rect -12365 15965 -12360 15995
rect -12400 15960 -12360 15965
rect -12320 16475 -12280 16480
rect -12320 16445 -12315 16475
rect -12285 16445 -12280 16475
rect -12320 16315 -12280 16445
rect -12320 16285 -12315 16315
rect -12285 16285 -12280 16315
rect -12320 16155 -12280 16285
rect -12320 16125 -12315 16155
rect -12285 16125 -12280 16155
rect -12320 15995 -12280 16125
rect -12320 15965 -12315 15995
rect -12285 15965 -12280 15995
rect -12320 15960 -12280 15965
rect -12240 16475 -12200 16480
rect -12240 16445 -12235 16475
rect -12205 16445 -12200 16475
rect -12240 16315 -12200 16445
rect -12240 16285 -12235 16315
rect -12205 16285 -12200 16315
rect -12240 16155 -12200 16285
rect -12240 16125 -12235 16155
rect -12205 16125 -12200 16155
rect -12240 15995 -12200 16125
rect -12240 15965 -12235 15995
rect -12205 15965 -12200 15995
rect -12240 15960 -12200 15965
rect -12160 16475 -12120 16480
rect -12160 16445 -12155 16475
rect -12125 16445 -12120 16475
rect -12160 16315 -12120 16445
rect -12160 16285 -12155 16315
rect -12125 16285 -12120 16315
rect -12160 16155 -12120 16285
rect -12160 16125 -12155 16155
rect -12125 16125 -12120 16155
rect -12160 15995 -12120 16125
rect -12160 15965 -12155 15995
rect -12125 15965 -12120 15995
rect -12160 15960 -12120 15965
rect -12080 16475 -12040 16480
rect -12080 16445 -12075 16475
rect -12045 16445 -12040 16475
rect -12080 16315 -12040 16445
rect -12080 16285 -12075 16315
rect -12045 16285 -12040 16315
rect -12080 16155 -12040 16285
rect -12080 16125 -12075 16155
rect -12045 16125 -12040 16155
rect -12080 15995 -12040 16125
rect -12080 15965 -12075 15995
rect -12045 15965 -12040 15995
rect -12080 15960 -12040 15965
rect -12000 16475 -11960 16480
rect -12000 16445 -11995 16475
rect -11965 16445 -11960 16475
rect -12000 16315 -11960 16445
rect -12000 16285 -11995 16315
rect -11965 16285 -11960 16315
rect -12000 16155 -11960 16285
rect -12000 16125 -11995 16155
rect -11965 16125 -11960 16155
rect -12000 15995 -11960 16125
rect -12000 15965 -11995 15995
rect -11965 15965 -11960 15995
rect -12000 15960 -11960 15965
rect -11920 16475 -11880 16480
rect -11920 16445 -11915 16475
rect -11885 16445 -11880 16475
rect -11920 16315 -11880 16445
rect -11920 16285 -11915 16315
rect -11885 16285 -11880 16315
rect -11920 16155 -11880 16285
rect -11920 16125 -11915 16155
rect -11885 16125 -11880 16155
rect -11920 15995 -11880 16125
rect -11920 15965 -11915 15995
rect -11885 15965 -11880 15995
rect -11920 15960 -11880 15965
rect -11840 16475 -11800 16480
rect -11840 16445 -11835 16475
rect -11805 16445 -11800 16475
rect -11840 16315 -11800 16445
rect -11840 16285 -11835 16315
rect -11805 16285 -11800 16315
rect -11840 16155 -11800 16285
rect -11840 16125 -11835 16155
rect -11805 16125 -11800 16155
rect -11840 15995 -11800 16125
rect -11840 15965 -11835 15995
rect -11805 15965 -11800 15995
rect -11840 15960 -11800 15965
rect -11760 16475 -11720 16480
rect -11760 16445 -11755 16475
rect -11725 16445 -11720 16475
rect -11760 16315 -11720 16445
rect -11760 16285 -11755 16315
rect -11725 16285 -11720 16315
rect -11760 16155 -11720 16285
rect -11760 16125 -11755 16155
rect -11725 16125 -11720 16155
rect -11760 15995 -11720 16125
rect -11760 15965 -11755 15995
rect -11725 15965 -11720 15995
rect -11760 15960 -11720 15965
rect -11680 16475 -11640 16480
rect -11680 16445 -11675 16475
rect -11645 16445 -11640 16475
rect -11680 16315 -11640 16445
rect -11680 16285 -11675 16315
rect -11645 16285 -11640 16315
rect -11680 16155 -11640 16285
rect -11680 16125 -11675 16155
rect -11645 16125 -11640 16155
rect -11680 15995 -11640 16125
rect -11680 15965 -11675 15995
rect -11645 15965 -11640 15995
rect -11680 15960 -11640 15965
rect -11600 16475 -11560 16480
rect -11600 16445 -11595 16475
rect -11565 16445 -11560 16475
rect -11600 16315 -11560 16445
rect -11600 16285 -11595 16315
rect -11565 16285 -11560 16315
rect -11600 16155 -11560 16285
rect -11600 16125 -11595 16155
rect -11565 16125 -11560 16155
rect -11600 15995 -11560 16125
rect -11600 15965 -11595 15995
rect -11565 15965 -11560 15995
rect -11600 15960 -11560 15965
rect -11520 16475 -11480 16480
rect -11520 16445 -11515 16475
rect -11485 16445 -11480 16475
rect -11520 16315 -11480 16445
rect -11520 16285 -11515 16315
rect -11485 16285 -11480 16315
rect -11520 16155 -11480 16285
rect -11520 16125 -11515 16155
rect -11485 16125 -11480 16155
rect -11520 15995 -11480 16125
rect -11520 15965 -11515 15995
rect -11485 15965 -11480 15995
rect -11520 15960 -11480 15965
rect -11440 16475 -11400 16480
rect -11440 16445 -11435 16475
rect -11405 16445 -11400 16475
rect -11440 16315 -11400 16445
rect -11440 16285 -11435 16315
rect -11405 16285 -11400 16315
rect -11440 16155 -11400 16285
rect -11440 16125 -11435 16155
rect -11405 16125 -11400 16155
rect -11440 15995 -11400 16125
rect -11440 15965 -11435 15995
rect -11405 15965 -11400 15995
rect -11440 15960 -11400 15965
rect -11360 16475 -11320 16480
rect -11360 16445 -11355 16475
rect -11325 16445 -11320 16475
rect -11360 16315 -11320 16445
rect -11360 16285 -11355 16315
rect -11325 16285 -11320 16315
rect -11360 16155 -11320 16285
rect -11360 16125 -11355 16155
rect -11325 16125 -11320 16155
rect -11360 15995 -11320 16125
rect -11360 15965 -11355 15995
rect -11325 15965 -11320 15995
rect -11360 15960 -11320 15965
rect -11280 16475 -11240 16480
rect -11280 16445 -11275 16475
rect -11245 16445 -11240 16475
rect -11280 16315 -11240 16445
rect -11280 16285 -11275 16315
rect -11245 16285 -11240 16315
rect -11280 16155 -11240 16285
rect -11280 16125 -11275 16155
rect -11245 16125 -11240 16155
rect -11280 15995 -11240 16125
rect -11280 15965 -11275 15995
rect -11245 15965 -11240 15995
rect -11280 15960 -11240 15965
rect -11200 16475 -11160 16480
rect -11200 16445 -11195 16475
rect -11165 16445 -11160 16475
rect -11200 16315 -11160 16445
rect -11200 16285 -11195 16315
rect -11165 16285 -11160 16315
rect -11200 16155 -11160 16285
rect -11200 16125 -11195 16155
rect -11165 16125 -11160 16155
rect -11200 15995 -11160 16125
rect -11200 15965 -11195 15995
rect -11165 15965 -11160 15995
rect -11200 15960 -11160 15965
rect -11120 16475 -11080 16480
rect -11120 16445 -11115 16475
rect -11085 16445 -11080 16475
rect -11120 16315 -11080 16445
rect -11120 16285 -11115 16315
rect -11085 16285 -11080 16315
rect -11120 16155 -11080 16285
rect -11120 16125 -11115 16155
rect -11085 16125 -11080 16155
rect -11120 15995 -11080 16125
rect -11120 15965 -11115 15995
rect -11085 15965 -11080 15995
rect -11120 15960 -11080 15965
rect -11040 16475 -11000 16480
rect -11040 16445 -11035 16475
rect -11005 16445 -11000 16475
rect -11040 16315 -11000 16445
rect -11040 16285 -11035 16315
rect -11005 16285 -11000 16315
rect -11040 16155 -11000 16285
rect -11040 16125 -11035 16155
rect -11005 16125 -11000 16155
rect -11040 15995 -11000 16125
rect -11040 15965 -11035 15995
rect -11005 15965 -11000 15995
rect -11040 15960 -11000 15965
rect -10960 16475 -10920 16480
rect -10960 16445 -10955 16475
rect -10925 16445 -10920 16475
rect -10960 16315 -10920 16445
rect -10960 16285 -10955 16315
rect -10925 16285 -10920 16315
rect -10960 16155 -10920 16285
rect -10960 16125 -10955 16155
rect -10925 16125 -10920 16155
rect -10960 15995 -10920 16125
rect -10960 15965 -10955 15995
rect -10925 15965 -10920 15995
rect -10960 15960 -10920 15965
rect -10880 16475 -10840 16480
rect -10880 16445 -10875 16475
rect -10845 16445 -10840 16475
rect -10880 16315 -10840 16445
rect -10880 16285 -10875 16315
rect -10845 16285 -10840 16315
rect -10880 16155 -10840 16285
rect -10880 16125 -10875 16155
rect -10845 16125 -10840 16155
rect -10880 15995 -10840 16125
rect -10880 15965 -10875 15995
rect -10845 15965 -10840 15995
rect -10880 15960 -10840 15965
rect -10800 16475 -10760 16480
rect -10800 16445 -10795 16475
rect -10765 16445 -10760 16475
rect -10800 16315 -10760 16445
rect -10800 16285 -10795 16315
rect -10765 16285 -10760 16315
rect -10800 16155 -10760 16285
rect -10800 16125 -10795 16155
rect -10765 16125 -10760 16155
rect -10800 15995 -10760 16125
rect -10800 15965 -10795 15995
rect -10765 15965 -10760 15995
rect -10800 15960 -10760 15965
rect -10720 16475 -10680 16480
rect -10720 16445 -10715 16475
rect -10685 16445 -10680 16475
rect -10720 16315 -10680 16445
rect -10720 16285 -10715 16315
rect -10685 16285 -10680 16315
rect -10720 16155 -10680 16285
rect -10720 16125 -10715 16155
rect -10685 16125 -10680 16155
rect -10720 15995 -10680 16125
rect -10720 15965 -10715 15995
rect -10685 15965 -10680 15995
rect -10720 15960 -10680 15965
rect -10640 16475 -10600 16480
rect -10640 16445 -10635 16475
rect -10605 16445 -10600 16475
rect -10640 16315 -10600 16445
rect -10640 16285 -10635 16315
rect -10605 16285 -10600 16315
rect -10640 16155 -10600 16285
rect -10640 16125 -10635 16155
rect -10605 16125 -10600 16155
rect -10640 15995 -10600 16125
rect -10640 15965 -10635 15995
rect -10605 15965 -10600 15995
rect -10640 15960 -10600 15965
rect -10560 16475 -10520 16480
rect -10560 16445 -10555 16475
rect -10525 16445 -10520 16475
rect -10560 16315 -10520 16445
rect -10560 16285 -10555 16315
rect -10525 16285 -10520 16315
rect -10560 16155 -10520 16285
rect -10560 16125 -10555 16155
rect -10525 16125 -10520 16155
rect -10560 15995 -10520 16125
rect -10560 15965 -10555 15995
rect -10525 15965 -10520 15995
rect -10560 15960 -10520 15965
rect -10480 16475 -10440 16480
rect -10480 16445 -10475 16475
rect -10445 16445 -10440 16475
rect -10480 16315 -10440 16445
rect -10480 16285 -10475 16315
rect -10445 16285 -10440 16315
rect -10480 16155 -10440 16285
rect -10480 16125 -10475 16155
rect -10445 16125 -10440 16155
rect -10480 15995 -10440 16125
rect -10480 15965 -10475 15995
rect -10445 15965 -10440 15995
rect -10480 15960 -10440 15965
rect -10400 16475 -10360 16480
rect -10400 16445 -10395 16475
rect -10365 16445 -10360 16475
rect -10400 16315 -10360 16445
rect -10400 16285 -10395 16315
rect -10365 16285 -10360 16315
rect -10400 16155 -10360 16285
rect -10400 16125 -10395 16155
rect -10365 16125 -10360 16155
rect -10400 15995 -10360 16125
rect -10400 15965 -10395 15995
rect -10365 15965 -10360 15995
rect -10400 15960 -10360 15965
rect -10320 16475 -10280 16480
rect -10320 16445 -10315 16475
rect -10285 16445 -10280 16475
rect -10320 16315 -10280 16445
rect -10320 16285 -10315 16315
rect -10285 16285 -10280 16315
rect -10320 16155 -10280 16285
rect -10320 16125 -10315 16155
rect -10285 16125 -10280 16155
rect -10320 15995 -10280 16125
rect -10320 15965 -10315 15995
rect -10285 15965 -10280 15995
rect -10320 15960 -10280 15965
rect -10240 16475 -10200 16480
rect -10240 16445 -10235 16475
rect -10205 16445 -10200 16475
rect -10240 16315 -10200 16445
rect -10240 16285 -10235 16315
rect -10205 16285 -10200 16315
rect -10240 16155 -10200 16285
rect -10240 16125 -10235 16155
rect -10205 16125 -10200 16155
rect -10240 15995 -10200 16125
rect -10240 15965 -10235 15995
rect -10205 15965 -10200 15995
rect -10240 15960 -10200 15965
rect -10160 16475 -10120 16480
rect -10160 16445 -10155 16475
rect -10125 16445 -10120 16475
rect -10160 16315 -10120 16445
rect -10160 16285 -10155 16315
rect -10125 16285 -10120 16315
rect -10160 16155 -10120 16285
rect -10160 16125 -10155 16155
rect -10125 16125 -10120 16155
rect -10160 15995 -10120 16125
rect -10160 15965 -10155 15995
rect -10125 15965 -10120 15995
rect -10160 15960 -10120 15965
rect -10080 16475 -10040 16480
rect -10080 16445 -10075 16475
rect -10045 16445 -10040 16475
rect -10080 16315 -10040 16445
rect -10080 16285 -10075 16315
rect -10045 16285 -10040 16315
rect -10080 16155 -10040 16285
rect -10080 16125 -10075 16155
rect -10045 16125 -10040 16155
rect -10080 15995 -10040 16125
rect -10080 15965 -10075 15995
rect -10045 15965 -10040 15995
rect -10080 15960 -10040 15965
rect -10000 16475 -9960 16480
rect -10000 16445 -9995 16475
rect -9965 16445 -9960 16475
rect -10000 16315 -9960 16445
rect -10000 16285 -9995 16315
rect -9965 16285 -9960 16315
rect -10000 16155 -9960 16285
rect -10000 16125 -9995 16155
rect -9965 16125 -9960 16155
rect -10000 15995 -9960 16125
rect -10000 15965 -9995 15995
rect -9965 15965 -9960 15995
rect -10000 15960 -9960 15965
rect -9920 16475 -9880 16480
rect -9920 16445 -9915 16475
rect -9885 16445 -9880 16475
rect -9920 16315 -9880 16445
rect -9920 16285 -9915 16315
rect -9885 16285 -9880 16315
rect -9920 16155 -9880 16285
rect -9920 16125 -9915 16155
rect -9885 16125 -9880 16155
rect -9920 15995 -9880 16125
rect -9920 15965 -9915 15995
rect -9885 15965 -9880 15995
rect -9920 15960 -9880 15965
rect -9840 16475 -9800 16480
rect -9840 16445 -9835 16475
rect -9805 16445 -9800 16475
rect -9840 16315 -9800 16445
rect -9840 16285 -9835 16315
rect -9805 16285 -9800 16315
rect -9840 16155 -9800 16285
rect -9840 16125 -9835 16155
rect -9805 16125 -9800 16155
rect -9840 15995 -9800 16125
rect -9840 15965 -9835 15995
rect -9805 15965 -9800 15995
rect -9840 15960 -9800 15965
rect -9760 16475 -9720 16480
rect -9760 16445 -9755 16475
rect -9725 16445 -9720 16475
rect -9760 16315 -9720 16445
rect -9760 16285 -9755 16315
rect -9725 16285 -9720 16315
rect -9760 16155 -9720 16285
rect -9760 16125 -9755 16155
rect -9725 16125 -9720 16155
rect -9760 15995 -9720 16125
rect -9760 15965 -9755 15995
rect -9725 15965 -9720 15995
rect -9760 15960 -9720 15965
rect -9680 16475 -9640 16480
rect -9680 16445 -9675 16475
rect -9645 16445 -9640 16475
rect -9680 16315 -9640 16445
rect -9680 16285 -9675 16315
rect -9645 16285 -9640 16315
rect -9680 16155 -9640 16285
rect -9680 16125 -9675 16155
rect -9645 16125 -9640 16155
rect -9680 15995 -9640 16125
rect -9680 15965 -9675 15995
rect -9645 15965 -9640 15995
rect -9680 15960 -9640 15965
rect -9600 16475 -9560 16480
rect -9600 16445 -9595 16475
rect -9565 16445 -9560 16475
rect -9600 16315 -9560 16445
rect -9600 16285 -9595 16315
rect -9565 16285 -9560 16315
rect -9600 16155 -9560 16285
rect -9600 16125 -9595 16155
rect -9565 16125 -9560 16155
rect -9600 15995 -9560 16125
rect -9600 15965 -9595 15995
rect -9565 15965 -9560 15995
rect -9600 15960 -9560 15965
rect -9520 16475 -9480 16480
rect -9520 16445 -9515 16475
rect -9485 16445 -9480 16475
rect -9520 16315 -9480 16445
rect -9520 16285 -9515 16315
rect -9485 16285 -9480 16315
rect -9520 16155 -9480 16285
rect -9520 16125 -9515 16155
rect -9485 16125 -9480 16155
rect -9520 15995 -9480 16125
rect -9520 15965 -9515 15995
rect -9485 15965 -9480 15995
rect -9520 15960 -9480 15965
rect -9440 16475 -9400 16480
rect -9440 16445 -9435 16475
rect -9405 16445 -9400 16475
rect -9440 16315 -9400 16445
rect -9440 16285 -9435 16315
rect -9405 16285 -9400 16315
rect -9440 16155 -9400 16285
rect -9440 16125 -9435 16155
rect -9405 16125 -9400 16155
rect -9440 15995 -9400 16125
rect -9440 15965 -9435 15995
rect -9405 15965 -9400 15995
rect -9440 15960 -9400 15965
rect -9360 16475 -9320 16480
rect -9360 16445 -9355 16475
rect -9325 16445 -9320 16475
rect -9360 16315 -9320 16445
rect -9360 16285 -9355 16315
rect -9325 16285 -9320 16315
rect -9360 16155 -9320 16285
rect -9360 16125 -9355 16155
rect -9325 16125 -9320 16155
rect -9360 15995 -9320 16125
rect -9360 15965 -9355 15995
rect -9325 15965 -9320 15995
rect -9360 15960 -9320 15965
rect -9280 16475 -9240 16480
rect -9280 16445 -9275 16475
rect -9245 16445 -9240 16475
rect -9280 16315 -9240 16445
rect -9280 16285 -9275 16315
rect -9245 16285 -9240 16315
rect -9280 16155 -9240 16285
rect -9280 16125 -9275 16155
rect -9245 16125 -9240 16155
rect -9280 15995 -9240 16125
rect -9280 15965 -9275 15995
rect -9245 15965 -9240 15995
rect -9280 15960 -9240 15965
rect -9200 16475 -9160 16480
rect -9200 16445 -9195 16475
rect -9165 16445 -9160 16475
rect -9200 16315 -9160 16445
rect -9200 16285 -9195 16315
rect -9165 16285 -9160 16315
rect -9200 16155 -9160 16285
rect -9200 16125 -9195 16155
rect -9165 16125 -9160 16155
rect -9200 15995 -9160 16125
rect -9200 15965 -9195 15995
rect -9165 15965 -9160 15995
rect -9200 15960 -9160 15965
rect -9120 16475 -9080 16480
rect -9120 16445 -9115 16475
rect -9085 16445 -9080 16475
rect -9120 16315 -9080 16445
rect -9120 16285 -9115 16315
rect -9085 16285 -9080 16315
rect -9120 16155 -9080 16285
rect -9120 16125 -9115 16155
rect -9085 16125 -9080 16155
rect -9120 15995 -9080 16125
rect -9120 15965 -9115 15995
rect -9085 15965 -9080 15995
rect -9120 15960 -9080 15965
rect -9040 16475 -9000 16480
rect -9040 16445 -9035 16475
rect -9005 16445 -9000 16475
rect -9040 16315 -9000 16445
rect -9040 16285 -9035 16315
rect -9005 16285 -9000 16315
rect -9040 16155 -9000 16285
rect -9040 16125 -9035 16155
rect -9005 16125 -9000 16155
rect -9040 15995 -9000 16125
rect -9040 15965 -9035 15995
rect -9005 15965 -9000 15995
rect -9040 15960 -9000 15965
rect -8960 16475 -8920 16480
rect -8960 16445 -8955 16475
rect -8925 16445 -8920 16475
rect -8960 16315 -8920 16445
rect -8960 16285 -8955 16315
rect -8925 16285 -8920 16315
rect -8960 16155 -8920 16285
rect -8960 16125 -8955 16155
rect -8925 16125 -8920 16155
rect -8960 15995 -8920 16125
rect -8960 15965 -8955 15995
rect -8925 15965 -8920 15995
rect -8960 15960 -8920 15965
rect -8880 16475 -8840 16480
rect -8880 16445 -8875 16475
rect -8845 16445 -8840 16475
rect -8880 16315 -8840 16445
rect -8880 16285 -8875 16315
rect -8845 16285 -8840 16315
rect -8880 16155 -8840 16285
rect -8880 16125 -8875 16155
rect -8845 16125 -8840 16155
rect -8880 15995 -8840 16125
rect -8880 15965 -8875 15995
rect -8845 15965 -8840 15995
rect -8880 15960 -8840 15965
rect -8800 16475 -8760 16480
rect -8800 16445 -8795 16475
rect -8765 16445 -8760 16475
rect -8800 16315 -8760 16445
rect -8800 16285 -8795 16315
rect -8765 16285 -8760 16315
rect -8800 16155 -8760 16285
rect -8800 16125 -8795 16155
rect -8765 16125 -8760 16155
rect -8800 15995 -8760 16125
rect -8800 15965 -8795 15995
rect -8765 15965 -8760 15995
rect -8800 15960 -8760 15965
rect -8720 16475 -8680 16480
rect -8720 16445 -8715 16475
rect -8685 16445 -8680 16475
rect -8720 16315 -8680 16445
rect -8720 16285 -8715 16315
rect -8685 16285 -8680 16315
rect -8720 16155 -8680 16285
rect -8720 16125 -8715 16155
rect -8685 16125 -8680 16155
rect -8720 15995 -8680 16125
rect -8720 15965 -8715 15995
rect -8685 15965 -8680 15995
rect -8720 15960 -8680 15965
rect -8640 16475 -8600 16480
rect -8640 16445 -8635 16475
rect -8605 16445 -8600 16475
rect -8640 16315 -8600 16445
rect -8640 16285 -8635 16315
rect -8605 16285 -8600 16315
rect -8640 16155 -8600 16285
rect -8640 16125 -8635 16155
rect -8605 16125 -8600 16155
rect -8640 15995 -8600 16125
rect -8640 15965 -8635 15995
rect -8605 15965 -8600 15995
rect -8640 15960 -8600 15965
rect -8560 16475 -8520 16480
rect -8560 16445 -8555 16475
rect -8525 16445 -8520 16475
rect -8560 16315 -8520 16445
rect -8560 16285 -8555 16315
rect -8525 16285 -8520 16315
rect -8560 16155 -8520 16285
rect -8560 16125 -8555 16155
rect -8525 16125 -8520 16155
rect -8560 15995 -8520 16125
rect -8560 15965 -8555 15995
rect -8525 15965 -8520 15995
rect -8560 15960 -8520 15965
rect -8480 16475 -8440 16480
rect -8480 16445 -8475 16475
rect -8445 16445 -8440 16475
rect -8480 16315 -8440 16445
rect -8480 16285 -8475 16315
rect -8445 16285 -8440 16315
rect -8480 16155 -8440 16285
rect -8480 16125 -8475 16155
rect -8445 16125 -8440 16155
rect -8480 15995 -8440 16125
rect -8480 15965 -8475 15995
rect -8445 15965 -8440 15995
rect -8480 15960 -8440 15965
rect -8400 16475 -8360 16480
rect -8400 16445 -8395 16475
rect -8365 16445 -8360 16475
rect -8400 16315 -8360 16445
rect -8400 16285 -8395 16315
rect -8365 16285 -8360 16315
rect -8400 16155 -8360 16285
rect -8400 16125 -8395 16155
rect -8365 16125 -8360 16155
rect -8400 15995 -8360 16125
rect -8400 15965 -8395 15995
rect -8365 15965 -8360 15995
rect -8400 15960 -8360 15965
rect -8320 16475 -8280 16480
rect -8320 16445 -8315 16475
rect -8285 16445 -8280 16475
rect -8320 16315 -8280 16445
rect -8320 16285 -8315 16315
rect -8285 16285 -8280 16315
rect -8320 16155 -8280 16285
rect -8320 16125 -8315 16155
rect -8285 16125 -8280 16155
rect -8320 15995 -8280 16125
rect -8320 15965 -8315 15995
rect -8285 15965 -8280 15995
rect -8320 15960 -8280 15965
rect -8240 16475 -8200 16480
rect -8240 16445 -8235 16475
rect -8205 16445 -8200 16475
rect -8240 16315 -8200 16445
rect -8240 16285 -8235 16315
rect -8205 16285 -8200 16315
rect -8240 16155 -8200 16285
rect -8240 16125 -8235 16155
rect -8205 16125 -8200 16155
rect -8240 15995 -8200 16125
rect -8240 15965 -8235 15995
rect -8205 15965 -8200 15995
rect -8240 15960 -8200 15965
rect -8160 16475 -8120 16480
rect -8160 16445 -8155 16475
rect -8125 16445 -8120 16475
rect -8160 16315 -8120 16445
rect -8160 16285 -8155 16315
rect -8125 16285 -8120 16315
rect -8160 16155 -8120 16285
rect -8160 16125 -8155 16155
rect -8125 16125 -8120 16155
rect -8160 15995 -8120 16125
rect -8160 15965 -8155 15995
rect -8125 15965 -8120 15995
rect -8160 15960 -8120 15965
rect -8080 16475 -8040 16480
rect -8080 16445 -8075 16475
rect -8045 16445 -8040 16475
rect -8080 16315 -8040 16445
rect -8080 16285 -8075 16315
rect -8045 16285 -8040 16315
rect -8080 16155 -8040 16285
rect -8080 16125 -8075 16155
rect -8045 16125 -8040 16155
rect -8080 15995 -8040 16125
rect -8080 15965 -8075 15995
rect -8045 15965 -8040 15995
rect -8080 15960 -8040 15965
rect -8000 16475 -7960 16480
rect -8000 16445 -7995 16475
rect -7965 16445 -7960 16475
rect -8000 16315 -7960 16445
rect -8000 16285 -7995 16315
rect -7965 16285 -7960 16315
rect -8000 16155 -7960 16285
rect -8000 16125 -7995 16155
rect -7965 16125 -7960 16155
rect -8000 15995 -7960 16125
rect -8000 15965 -7995 15995
rect -7965 15965 -7960 15995
rect -8000 15960 -7960 15965
rect -7920 16475 -7880 16480
rect -7920 16445 -7915 16475
rect -7885 16445 -7880 16475
rect -7920 16315 -7880 16445
rect -7920 16285 -7915 16315
rect -7885 16285 -7880 16315
rect -7920 16155 -7880 16285
rect -7920 16125 -7915 16155
rect -7885 16125 -7880 16155
rect -7920 15995 -7880 16125
rect -7920 15965 -7915 15995
rect -7885 15965 -7880 15995
rect -7920 15960 -7880 15965
rect -7840 16475 -7800 16480
rect -7840 16445 -7835 16475
rect -7805 16445 -7800 16475
rect -7840 16315 -7800 16445
rect -7840 16285 -7835 16315
rect -7805 16285 -7800 16315
rect -7840 16155 -7800 16285
rect -7840 16125 -7835 16155
rect -7805 16125 -7800 16155
rect -7840 15995 -7800 16125
rect -7840 15965 -7835 15995
rect -7805 15965 -7800 15995
rect -7840 15960 -7800 15965
rect -7760 16475 -7720 16480
rect -7760 16445 -7755 16475
rect -7725 16445 -7720 16475
rect -7760 16315 -7720 16445
rect -7760 16285 -7755 16315
rect -7725 16285 -7720 16315
rect -7760 16155 -7720 16285
rect -7760 16125 -7755 16155
rect -7725 16125 -7720 16155
rect -7760 15995 -7720 16125
rect -7760 15965 -7755 15995
rect -7725 15965 -7720 15995
rect -7760 15960 -7720 15965
rect -7680 16475 -7640 16480
rect -7680 16445 -7675 16475
rect -7645 16445 -7640 16475
rect -7680 16315 -7640 16445
rect -7680 16285 -7675 16315
rect -7645 16285 -7640 16315
rect -7680 16155 -7640 16285
rect -7680 16125 -7675 16155
rect -7645 16125 -7640 16155
rect -7680 15995 -7640 16125
rect -7680 15965 -7675 15995
rect -7645 15965 -7640 15995
rect -7680 15960 -7640 15965
rect -7600 16475 -7560 16480
rect -7600 16445 -7595 16475
rect -7565 16445 -7560 16475
rect -7600 16315 -7560 16445
rect -7600 16285 -7595 16315
rect -7565 16285 -7560 16315
rect -7600 16155 -7560 16285
rect -7600 16125 -7595 16155
rect -7565 16125 -7560 16155
rect -7600 15995 -7560 16125
rect -7600 15965 -7595 15995
rect -7565 15965 -7560 15995
rect -7600 15960 -7560 15965
rect -7520 16475 -7480 16480
rect -7520 16445 -7515 16475
rect -7485 16445 -7480 16475
rect -7520 16315 -7480 16445
rect -7520 16285 -7515 16315
rect -7485 16285 -7480 16315
rect -7520 16155 -7480 16285
rect -7520 16125 -7515 16155
rect -7485 16125 -7480 16155
rect -7520 15995 -7480 16125
rect -7520 15965 -7515 15995
rect -7485 15965 -7480 15995
rect -7520 15960 -7480 15965
rect -7440 16475 -7400 16480
rect -7440 16445 -7435 16475
rect -7405 16445 -7400 16475
rect -7440 16315 -7400 16445
rect -7440 16285 -7435 16315
rect -7405 16285 -7400 16315
rect -7440 16155 -7400 16285
rect -7440 16125 -7435 16155
rect -7405 16125 -7400 16155
rect -7440 15995 -7400 16125
rect -7440 15965 -7435 15995
rect -7405 15965 -7400 15995
rect -7440 15960 -7400 15965
rect -7360 16475 -7320 16480
rect -7360 16445 -7355 16475
rect -7325 16445 -7320 16475
rect -7360 16315 -7320 16445
rect -7360 16285 -7355 16315
rect -7325 16285 -7320 16315
rect -7360 16155 -7320 16285
rect -7360 16125 -7355 16155
rect -7325 16125 -7320 16155
rect -7360 15995 -7320 16125
rect -7360 15965 -7355 15995
rect -7325 15965 -7320 15995
rect -7360 15960 -7320 15965
rect -7280 16475 -7240 16480
rect -7280 16445 -7275 16475
rect -7245 16445 -7240 16475
rect -7280 16315 -7240 16445
rect -7280 16285 -7275 16315
rect -7245 16285 -7240 16315
rect -7280 16155 -7240 16285
rect -7280 16125 -7275 16155
rect -7245 16125 -7240 16155
rect -7280 15995 -7240 16125
rect -7280 15965 -7275 15995
rect -7245 15965 -7240 15995
rect -7280 15960 -7240 15965
rect -7200 16475 -7160 16480
rect -7200 16445 -7195 16475
rect -7165 16445 -7160 16475
rect -7200 16315 -7160 16445
rect -7200 16285 -7195 16315
rect -7165 16285 -7160 16315
rect -7200 16155 -7160 16285
rect -7200 16125 -7195 16155
rect -7165 16125 -7160 16155
rect -7200 15995 -7160 16125
rect -7200 15965 -7195 15995
rect -7165 15965 -7160 15995
rect -7200 15960 -7160 15965
rect -7120 16475 -7080 16480
rect -7120 16445 -7115 16475
rect -7085 16445 -7080 16475
rect -7120 16315 -7080 16445
rect -7120 16285 -7115 16315
rect -7085 16285 -7080 16315
rect -7120 16155 -7080 16285
rect -7120 16125 -7115 16155
rect -7085 16125 -7080 16155
rect -7120 15995 -7080 16125
rect -7120 15965 -7115 15995
rect -7085 15965 -7080 15995
rect -7120 15960 -7080 15965
rect -7040 16475 -7000 16480
rect -7040 16445 -7035 16475
rect -7005 16445 -7000 16475
rect -7040 16315 -7000 16445
rect -7040 16285 -7035 16315
rect -7005 16285 -7000 16315
rect -7040 16155 -7000 16285
rect -7040 16125 -7035 16155
rect -7005 16125 -7000 16155
rect -7040 15995 -7000 16125
rect -7040 15965 -7035 15995
rect -7005 15965 -7000 15995
rect -7040 15960 -7000 15965
rect -6960 16475 -6920 16480
rect -6960 16445 -6955 16475
rect -6925 16445 -6920 16475
rect -6960 16315 -6920 16445
rect -6960 16285 -6955 16315
rect -6925 16285 -6920 16315
rect -6960 16155 -6920 16285
rect -6960 16125 -6955 16155
rect -6925 16125 -6920 16155
rect -6960 15995 -6920 16125
rect -6960 15965 -6955 15995
rect -6925 15965 -6920 15995
rect -6960 15960 -6920 15965
rect -6880 16475 -6840 16480
rect -6880 16445 -6875 16475
rect -6845 16445 -6840 16475
rect -6880 16315 -6840 16445
rect -6880 16285 -6875 16315
rect -6845 16285 -6840 16315
rect -6880 16155 -6840 16285
rect -6880 16125 -6875 16155
rect -6845 16125 -6840 16155
rect -6880 15995 -6840 16125
rect -6880 15965 -6875 15995
rect -6845 15965 -6840 15995
rect -6880 15960 -6840 15965
rect -6800 16475 -6760 16480
rect -6800 16445 -6795 16475
rect -6765 16445 -6760 16475
rect -6800 16315 -6760 16445
rect -6800 16285 -6795 16315
rect -6765 16285 -6760 16315
rect -6800 16155 -6760 16285
rect -6800 16125 -6795 16155
rect -6765 16125 -6760 16155
rect -6800 15995 -6760 16125
rect -6800 15965 -6795 15995
rect -6765 15965 -6760 15995
rect -6800 15960 -6760 15965
rect -6720 16475 -6680 16480
rect -6720 16445 -6715 16475
rect -6685 16445 -6680 16475
rect -6720 16315 -6680 16445
rect -6720 16285 -6715 16315
rect -6685 16285 -6680 16315
rect -6720 16155 -6680 16285
rect -6720 16125 -6715 16155
rect -6685 16125 -6680 16155
rect -6720 15995 -6680 16125
rect -6720 15965 -6715 15995
rect -6685 15965 -6680 15995
rect -6720 15960 -6680 15965
rect -6640 16475 -6600 16480
rect -6640 16445 -6635 16475
rect -6605 16445 -6600 16475
rect -6640 16315 -6600 16445
rect -6640 16285 -6635 16315
rect -6605 16285 -6600 16315
rect -6640 16155 -6600 16285
rect -6640 16125 -6635 16155
rect -6605 16125 -6600 16155
rect -6640 15995 -6600 16125
rect -6640 15965 -6635 15995
rect -6605 15965 -6600 15995
rect -6640 15960 -6600 15965
rect -6560 16475 -6520 16480
rect -6560 16445 -6555 16475
rect -6525 16445 -6520 16475
rect -6560 16315 -6520 16445
rect -6560 16285 -6555 16315
rect -6525 16285 -6520 16315
rect -6560 16155 -6520 16285
rect -6560 16125 -6555 16155
rect -6525 16125 -6520 16155
rect -6560 15995 -6520 16125
rect -6560 15965 -6555 15995
rect -6525 15965 -6520 15995
rect -6560 15960 -6520 15965
rect -6480 16475 -6440 16480
rect -6480 16445 -6475 16475
rect -6445 16445 -6440 16475
rect -6480 16315 -6440 16445
rect -6480 16285 -6475 16315
rect -6445 16285 -6440 16315
rect -6480 16155 -6440 16285
rect -6480 16125 -6475 16155
rect -6445 16125 -6440 16155
rect -6480 15995 -6440 16125
rect -6480 15965 -6475 15995
rect -6445 15965 -6440 15995
rect -6480 15960 -6440 15965
rect -6400 16475 -6360 16480
rect -6400 16445 -6395 16475
rect -6365 16445 -6360 16475
rect -6400 16315 -6360 16445
rect -6400 16285 -6395 16315
rect -6365 16285 -6360 16315
rect -6400 16155 -6360 16285
rect -6400 16125 -6395 16155
rect -6365 16125 -6360 16155
rect -6400 15995 -6360 16125
rect -6400 15965 -6395 15995
rect -6365 15965 -6360 15995
rect -6400 15960 -6360 15965
rect -6320 16475 -6280 16480
rect -6320 16445 -6315 16475
rect -6285 16445 -6280 16475
rect -6320 16315 -6280 16445
rect -6320 16285 -6315 16315
rect -6285 16285 -6280 16315
rect -6320 16155 -6280 16285
rect -6320 16125 -6315 16155
rect -6285 16125 -6280 16155
rect -6320 15995 -6280 16125
rect -6320 15965 -6315 15995
rect -6285 15965 -6280 15995
rect -6320 15960 -6280 15965
rect -6240 16475 -6200 16480
rect -6240 16445 -6235 16475
rect -6205 16445 -6200 16475
rect -6240 16315 -6200 16445
rect -6240 16285 -6235 16315
rect -6205 16285 -6200 16315
rect -6240 16155 -6200 16285
rect -6240 16125 -6235 16155
rect -6205 16125 -6200 16155
rect -6240 15995 -6200 16125
rect -6240 15965 -6235 15995
rect -6205 15965 -6200 15995
rect -6240 15960 -6200 15965
rect -6160 16475 -6120 16480
rect -6160 16445 -6155 16475
rect -6125 16445 -6120 16475
rect -6160 16315 -6120 16445
rect -6160 16285 -6155 16315
rect -6125 16285 -6120 16315
rect -6160 16155 -6120 16285
rect -6160 16125 -6155 16155
rect -6125 16125 -6120 16155
rect -6160 15995 -6120 16125
rect -6160 15965 -6155 15995
rect -6125 15965 -6120 15995
rect -6160 15960 -6120 15965
rect -6080 16475 -6040 16480
rect -6080 16445 -6075 16475
rect -6045 16445 -6040 16475
rect -6080 16315 -6040 16445
rect -6080 16285 -6075 16315
rect -6045 16285 -6040 16315
rect -6080 16155 -6040 16285
rect -6080 16125 -6075 16155
rect -6045 16125 -6040 16155
rect -6080 15995 -6040 16125
rect -6080 15965 -6075 15995
rect -6045 15965 -6040 15995
rect -6080 15960 -6040 15965
rect -6000 16475 -5960 16480
rect -6000 16445 -5995 16475
rect -5965 16445 -5960 16475
rect -6000 16315 -5960 16445
rect -6000 16285 -5995 16315
rect -5965 16285 -5960 16315
rect -6000 16155 -5960 16285
rect -6000 16125 -5995 16155
rect -5965 16125 -5960 16155
rect -6000 15995 -5960 16125
rect -6000 15965 -5995 15995
rect -5965 15965 -5960 15995
rect -6000 15960 -5960 15965
rect -5920 16475 -5880 16480
rect -5920 16445 -5915 16475
rect -5885 16445 -5880 16475
rect -5920 16315 -5880 16445
rect -5920 16285 -5915 16315
rect -5885 16285 -5880 16315
rect -5920 16155 -5880 16285
rect -5920 16125 -5915 16155
rect -5885 16125 -5880 16155
rect -5920 15995 -5880 16125
rect -5920 15965 -5915 15995
rect -5885 15965 -5880 15995
rect -5920 15960 -5880 15965
rect -5840 16475 -5800 16480
rect -5840 16445 -5835 16475
rect -5805 16445 -5800 16475
rect -5840 16315 -5800 16445
rect -5840 16285 -5835 16315
rect -5805 16285 -5800 16315
rect -5840 16155 -5800 16285
rect -5840 16125 -5835 16155
rect -5805 16125 -5800 16155
rect -5840 15995 -5800 16125
rect -5840 15965 -5835 15995
rect -5805 15965 -5800 15995
rect -5840 15960 -5800 15965
rect -5760 16475 -5720 16480
rect -5760 16445 -5755 16475
rect -5725 16445 -5720 16475
rect -5760 16315 -5720 16445
rect -5760 16285 -5755 16315
rect -5725 16285 -5720 16315
rect -5760 16155 -5720 16285
rect -5680 16235 -5640 17440
rect -5680 16205 -5675 16235
rect -5645 16205 -5640 16235
rect -5680 16200 -5640 16205
rect -5600 17355 -5560 17440
rect -5600 17325 -5595 17355
rect -5565 17325 -5560 17355
rect -5600 17195 -5560 17325
rect -5600 17165 -5595 17195
rect -5565 17165 -5560 17195
rect -5600 16475 -5560 17165
rect -5600 16445 -5595 16475
rect -5565 16445 -5560 16475
rect -5600 16315 -5560 16445
rect -5600 16285 -5595 16315
rect -5565 16285 -5560 16315
rect -5760 16125 -5755 16155
rect -5725 16125 -5720 16155
rect -5760 15995 -5720 16125
rect -5760 15965 -5755 15995
rect -5725 15965 -5720 15995
rect -5760 15960 -5720 15965
rect -5680 16155 -5640 16160
rect -5680 16125 -5675 16155
rect -5645 16125 -5640 16155
rect -5680 15995 -5640 16125
rect -5680 15965 -5675 15995
rect -5645 15965 -5640 15995
rect -5680 15960 -5640 15965
rect -5600 16155 -5560 16285
rect -5600 16125 -5595 16155
rect -5565 16125 -5560 16155
rect -5600 15995 -5560 16125
rect -5520 16075 -5480 17440
rect -5440 17355 -5400 17440
rect -5440 17325 -5435 17355
rect -5405 17325 -5400 17355
rect -5440 17195 -5400 17325
rect -5360 17275 -5320 17440
rect -5360 17245 -5355 17275
rect -5325 17245 -5320 17275
rect -5360 17240 -5320 17245
rect -5280 17355 -5240 17440
rect -5280 17325 -5275 17355
rect -5245 17325 -5240 17355
rect -5440 17165 -5435 17195
rect -5405 17165 -5400 17195
rect -5440 17160 -5400 17165
rect -5280 17195 -5240 17325
rect -5280 17165 -5275 17195
rect -5245 17165 -5240 17195
rect -5280 17160 -5240 17165
rect -1680 17396 -1640 17444
rect -1680 17364 -1676 17396
rect -1644 17364 -1640 17396
rect -1680 17316 -1640 17364
rect -1680 17284 -1676 17316
rect -1644 17284 -1640 17316
rect -1680 17236 -1640 17284
rect -1680 17204 -1676 17236
rect -1644 17204 -1640 17236
rect -1680 17156 -1640 17204
rect -1680 17124 -1676 17156
rect -1644 17124 -1640 17156
rect -1680 17076 -1640 17124
rect -1680 17044 -1676 17076
rect -1644 17044 -1640 17076
rect -1680 16996 -1640 17044
rect -1680 16964 -1676 16996
rect -1644 16964 -1640 16996
rect -1680 16916 -1640 16964
rect -1680 16884 -1676 16916
rect -1644 16884 -1640 16916
rect -1680 16836 -1640 16884
rect -1680 16804 -1676 16836
rect -1644 16804 -1640 16836
rect -1680 16756 -1640 16804
rect -1680 16724 -1676 16756
rect -1644 16724 -1640 16756
rect -1680 16636 -1640 16724
rect -1680 16604 -1676 16636
rect -1644 16604 -1640 16636
rect -1680 16556 -1640 16604
rect -1680 16524 -1676 16556
rect -1644 16524 -1640 16556
rect -5520 16045 -5515 16075
rect -5485 16045 -5480 16075
rect -5520 16040 -5480 16045
rect -5440 16475 -5400 16480
rect -5440 16445 -5435 16475
rect -5405 16445 -5400 16475
rect -5440 16315 -5400 16445
rect -5440 16285 -5435 16315
rect -5405 16285 -5400 16315
rect -5440 16155 -5400 16285
rect -5440 16125 -5435 16155
rect -5405 16125 -5400 16155
rect -5600 15965 -5595 15995
rect -5565 15965 -5560 15995
rect -5600 15960 -5560 15965
rect -5440 15995 -5400 16125
rect -5440 15965 -5435 15995
rect -5405 15965 -5400 15995
rect -5440 15960 -5400 15965
rect -5360 16475 -5320 16480
rect -5360 16445 -5355 16475
rect -5325 16445 -5320 16475
rect -5360 16315 -5320 16445
rect -5360 16285 -5355 16315
rect -5325 16285 -5320 16315
rect -5360 16155 -5320 16285
rect -5360 16125 -5355 16155
rect -5325 16125 -5320 16155
rect -5360 15995 -5320 16125
rect -5360 15965 -5355 15995
rect -5325 15965 -5320 15995
rect -5360 15960 -5320 15965
rect -5280 16475 -5240 16480
rect -5280 16445 -5275 16475
rect -5245 16445 -5240 16475
rect -5280 16315 -5240 16445
rect -5280 16285 -5275 16315
rect -5245 16285 -5240 16315
rect -5280 16155 -5240 16285
rect -5280 16125 -5275 16155
rect -5245 16125 -5240 16155
rect -5280 15995 -5240 16125
rect -5280 15965 -5275 15995
rect -5245 15965 -5240 15995
rect -5280 15960 -5240 15965
rect -5200 16475 -5160 16480
rect -5200 16445 -5195 16475
rect -5165 16445 -5160 16475
rect -5200 16315 -5160 16445
rect -5200 16285 -5195 16315
rect -5165 16285 -5160 16315
rect -5200 16155 -5160 16285
rect -5200 16125 -5195 16155
rect -5165 16125 -5160 16155
rect -5200 15995 -5160 16125
rect -5200 15965 -5195 15995
rect -5165 15965 -5160 15995
rect -5200 15960 -5160 15965
rect -5120 16475 -5080 16480
rect -5120 16445 -5115 16475
rect -5085 16445 -5080 16475
rect -5120 16315 -5080 16445
rect -5120 16285 -5115 16315
rect -5085 16285 -5080 16315
rect -5120 16155 -5080 16285
rect -5120 16125 -5115 16155
rect -5085 16125 -5080 16155
rect -5120 15995 -5080 16125
rect -5120 15965 -5115 15995
rect -5085 15965 -5080 15995
rect -5120 15960 -5080 15965
rect -5040 16475 -5000 16480
rect -5040 16445 -5035 16475
rect -5005 16445 -5000 16475
rect -5040 16315 -5000 16445
rect -5040 16285 -5035 16315
rect -5005 16285 -5000 16315
rect -5040 16155 -5000 16285
rect -5040 16125 -5035 16155
rect -5005 16125 -5000 16155
rect -5040 15995 -5000 16125
rect -5040 15965 -5035 15995
rect -5005 15965 -5000 15995
rect -5040 15960 -5000 15965
rect -4960 16475 -4920 16480
rect -4960 16445 -4955 16475
rect -4925 16445 -4920 16475
rect -4960 16315 -4920 16445
rect -4960 16285 -4955 16315
rect -4925 16285 -4920 16315
rect -4960 16155 -4920 16285
rect -4960 16125 -4955 16155
rect -4925 16125 -4920 16155
rect -4960 15995 -4920 16125
rect -4960 15965 -4955 15995
rect -4925 15965 -4920 15995
rect -4960 15960 -4920 15965
rect -4880 16475 -4840 16480
rect -4880 16445 -4875 16475
rect -4845 16445 -4840 16475
rect -4880 16315 -4840 16445
rect -4880 16285 -4875 16315
rect -4845 16285 -4840 16315
rect -4880 16155 -4840 16285
rect -4880 16125 -4875 16155
rect -4845 16125 -4840 16155
rect -4880 15995 -4840 16125
rect -4880 15965 -4875 15995
rect -4845 15965 -4840 15995
rect -4880 15960 -4840 15965
rect -4800 16475 -4760 16480
rect -4800 16445 -4795 16475
rect -4765 16445 -4760 16475
rect -4800 16315 -4760 16445
rect -4800 16285 -4795 16315
rect -4765 16285 -4760 16315
rect -4800 16155 -4760 16285
rect -4800 16125 -4795 16155
rect -4765 16125 -4760 16155
rect -4800 15995 -4760 16125
rect -4800 15965 -4795 15995
rect -4765 15965 -4760 15995
rect -4800 15960 -4760 15965
rect -4720 16475 -4680 16480
rect -4720 16445 -4715 16475
rect -4685 16445 -4680 16475
rect -4720 16315 -4680 16445
rect -4720 16285 -4715 16315
rect -4685 16285 -4680 16315
rect -4720 16155 -4680 16285
rect -4720 16125 -4715 16155
rect -4685 16125 -4680 16155
rect -4720 15995 -4680 16125
rect -4720 15965 -4715 15995
rect -4685 15965 -4680 15995
rect -4720 15960 -4680 15965
rect -4640 16475 -4600 16480
rect -4640 16445 -4635 16475
rect -4605 16445 -4600 16475
rect -4640 16315 -4600 16445
rect -4640 16285 -4635 16315
rect -4605 16285 -4600 16315
rect -4640 16155 -4600 16285
rect -4640 16125 -4635 16155
rect -4605 16125 -4600 16155
rect -4640 15995 -4600 16125
rect -4640 15965 -4635 15995
rect -4605 15965 -4600 15995
rect -4640 15960 -4600 15965
rect -4560 16475 -4520 16480
rect -4560 16445 -4555 16475
rect -4525 16445 -4520 16475
rect -4560 16315 -4520 16445
rect -4560 16285 -4555 16315
rect -4525 16285 -4520 16315
rect -4560 16155 -4520 16285
rect -4560 16125 -4555 16155
rect -4525 16125 -4520 16155
rect -4560 15995 -4520 16125
rect -4560 15965 -4555 15995
rect -4525 15965 -4520 15995
rect -4560 15960 -4520 15965
rect -4480 16475 -4440 16480
rect -4480 16445 -4475 16475
rect -4445 16445 -4440 16475
rect -4480 16315 -4440 16445
rect -4480 16285 -4475 16315
rect -4445 16285 -4440 16315
rect -4480 16155 -4440 16285
rect -4480 16125 -4475 16155
rect -4445 16125 -4440 16155
rect -4480 15995 -4440 16125
rect -4480 15965 -4475 15995
rect -4445 15965 -4440 15995
rect -4480 15960 -4440 15965
rect -4400 16475 -4360 16480
rect -4400 16445 -4395 16475
rect -4365 16445 -4360 16475
rect -4400 16315 -4360 16445
rect -4400 16285 -4395 16315
rect -4365 16285 -4360 16315
rect -4400 16155 -4360 16285
rect -4400 16125 -4395 16155
rect -4365 16125 -4360 16155
rect -4400 15995 -4360 16125
rect -4400 15965 -4395 15995
rect -4365 15965 -4360 15995
rect -4400 15960 -4360 15965
rect -4320 16475 -4280 16480
rect -4320 16445 -4315 16475
rect -4285 16445 -4280 16475
rect -4320 16315 -4280 16445
rect -4320 16285 -4315 16315
rect -4285 16285 -4280 16315
rect -4320 16155 -4280 16285
rect -4320 16125 -4315 16155
rect -4285 16125 -4280 16155
rect -4320 15995 -4280 16125
rect -4320 15965 -4315 15995
rect -4285 15965 -4280 15995
rect -4320 15960 -4280 15965
rect -4240 16475 -4200 16480
rect -4240 16445 -4235 16475
rect -4205 16445 -4200 16475
rect -4240 16315 -4200 16445
rect -4240 16285 -4235 16315
rect -4205 16285 -4200 16315
rect -4240 16155 -4200 16285
rect -4240 16125 -4235 16155
rect -4205 16125 -4200 16155
rect -4240 15995 -4200 16125
rect -4240 15965 -4235 15995
rect -4205 15965 -4200 15995
rect -4240 15960 -4200 15965
rect -4160 16475 -4120 16480
rect -4160 16445 -4155 16475
rect -4125 16445 -4120 16475
rect -4160 16315 -4120 16445
rect -4160 16285 -4155 16315
rect -4125 16285 -4120 16315
rect -4160 16155 -4120 16285
rect -4160 16125 -4155 16155
rect -4125 16125 -4120 16155
rect -4160 15995 -4120 16125
rect -4160 15965 -4155 15995
rect -4125 15965 -4120 15995
rect -4160 15960 -4120 15965
rect -4080 16475 -4040 16480
rect -4080 16445 -4075 16475
rect -4045 16445 -4040 16475
rect -4080 16315 -4040 16445
rect -4080 16285 -4075 16315
rect -4045 16285 -4040 16315
rect -4080 16155 -4040 16285
rect -4080 16125 -4075 16155
rect -4045 16125 -4040 16155
rect -4080 15995 -4040 16125
rect -4080 15965 -4075 15995
rect -4045 15965 -4040 15995
rect -4080 15960 -4040 15965
rect -4000 16475 -3960 16480
rect -4000 16445 -3995 16475
rect -3965 16445 -3960 16475
rect -4000 16315 -3960 16445
rect -4000 16285 -3995 16315
rect -3965 16285 -3960 16315
rect -4000 16155 -3960 16285
rect -4000 16125 -3995 16155
rect -3965 16125 -3960 16155
rect -4000 15995 -3960 16125
rect -4000 15965 -3995 15995
rect -3965 15965 -3960 15995
rect -4000 15960 -3960 15965
rect -3920 16475 -3880 16480
rect -3920 16445 -3915 16475
rect -3885 16445 -3880 16475
rect -3920 16315 -3880 16445
rect -3920 16285 -3915 16315
rect -3885 16285 -3880 16315
rect -3920 16155 -3880 16285
rect -3920 16125 -3915 16155
rect -3885 16125 -3880 16155
rect -3920 15995 -3880 16125
rect -3920 15965 -3915 15995
rect -3885 15965 -3880 15995
rect -3920 15960 -3880 15965
rect -3840 16475 -3800 16480
rect -3840 16445 -3835 16475
rect -3805 16445 -3800 16475
rect -3840 16315 -3800 16445
rect -3840 16285 -3835 16315
rect -3805 16285 -3800 16315
rect -3840 16155 -3800 16285
rect -3840 16125 -3835 16155
rect -3805 16125 -3800 16155
rect -3840 15995 -3800 16125
rect -3840 15965 -3835 15995
rect -3805 15965 -3800 15995
rect -3840 15960 -3800 15965
rect -3760 16475 -3720 16480
rect -3760 16445 -3755 16475
rect -3725 16445 -3720 16475
rect -3760 16315 -3720 16445
rect -3760 16285 -3755 16315
rect -3725 16285 -3720 16315
rect -3760 16155 -3720 16285
rect -3760 16125 -3755 16155
rect -3725 16125 -3720 16155
rect -3760 15995 -3720 16125
rect -3760 15965 -3755 15995
rect -3725 15965 -3720 15995
rect -3760 15960 -3720 15965
rect -3680 16475 -3640 16480
rect -3680 16445 -3675 16475
rect -3645 16445 -3640 16475
rect -3680 16315 -3640 16445
rect -3680 16285 -3675 16315
rect -3645 16285 -3640 16315
rect -3680 16155 -3640 16285
rect -3680 16125 -3675 16155
rect -3645 16125 -3640 16155
rect -3680 15995 -3640 16125
rect -3680 15965 -3675 15995
rect -3645 15965 -3640 15995
rect -3680 15960 -3640 15965
rect -3600 16475 -3560 16480
rect -3600 16445 -3595 16475
rect -3565 16445 -3560 16475
rect -3600 16315 -3560 16445
rect -3600 16285 -3595 16315
rect -3565 16285 -3560 16315
rect -3600 16155 -3560 16285
rect -3600 16125 -3595 16155
rect -3565 16125 -3560 16155
rect -3600 15995 -3560 16125
rect -3600 15965 -3595 15995
rect -3565 15965 -3560 15995
rect -3600 15960 -3560 15965
rect -3520 16475 -3480 16480
rect -3520 16445 -3515 16475
rect -3485 16445 -3480 16475
rect -3520 16315 -3480 16445
rect -3520 16285 -3515 16315
rect -3485 16285 -3480 16315
rect -3520 16155 -3480 16285
rect -3520 16125 -3515 16155
rect -3485 16125 -3480 16155
rect -3520 15995 -3480 16125
rect -3520 15965 -3515 15995
rect -3485 15965 -3480 15995
rect -3520 15960 -3480 15965
rect -3440 16475 -3400 16480
rect -3440 16445 -3435 16475
rect -3405 16445 -3400 16475
rect -3440 16315 -3400 16445
rect -3440 16285 -3435 16315
rect -3405 16285 -3400 16315
rect -3440 16155 -3400 16285
rect -3440 16125 -3435 16155
rect -3405 16125 -3400 16155
rect -3440 15995 -3400 16125
rect -3440 15965 -3435 15995
rect -3405 15965 -3400 15995
rect -3440 15960 -3400 15965
rect -3360 16475 -3320 16480
rect -3360 16445 -3355 16475
rect -3325 16445 -3320 16475
rect -3360 16315 -3320 16445
rect -3360 16285 -3355 16315
rect -3325 16285 -3320 16315
rect -3360 16155 -3320 16285
rect -3360 16125 -3355 16155
rect -3325 16125 -3320 16155
rect -3360 15995 -3320 16125
rect -3360 15965 -3355 15995
rect -3325 15965 -3320 15995
rect -3360 15960 -3320 15965
rect -3280 16475 -3240 16480
rect -3280 16445 -3275 16475
rect -3245 16445 -3240 16475
rect -3280 16315 -3240 16445
rect -3280 16285 -3275 16315
rect -3245 16285 -3240 16315
rect -3280 16155 -3240 16285
rect -3280 16125 -3275 16155
rect -3245 16125 -3240 16155
rect -3280 15995 -3240 16125
rect -3280 15965 -3275 15995
rect -3245 15965 -3240 15995
rect -3280 15960 -3240 15965
rect -3200 16475 -3160 16480
rect -3200 16445 -3195 16475
rect -3165 16445 -3160 16475
rect -3200 16315 -3160 16445
rect -3200 16285 -3195 16315
rect -3165 16285 -3160 16315
rect -3200 16155 -3160 16285
rect -3200 16125 -3195 16155
rect -3165 16125 -3160 16155
rect -3200 15995 -3160 16125
rect -3200 15965 -3195 15995
rect -3165 15965 -3160 15995
rect -3200 15960 -3160 15965
rect -3120 16475 -3080 16480
rect -3120 16445 -3115 16475
rect -3085 16445 -3080 16475
rect -3120 16315 -3080 16445
rect -3120 16285 -3115 16315
rect -3085 16285 -3080 16315
rect -3120 16155 -3080 16285
rect -3120 16125 -3115 16155
rect -3085 16125 -3080 16155
rect -3120 15995 -3080 16125
rect -3120 15965 -3115 15995
rect -3085 15965 -3080 15995
rect -3120 15960 -3080 15965
rect -3040 16475 -3000 16480
rect -3040 16445 -3035 16475
rect -3005 16445 -3000 16475
rect -3040 16315 -3000 16445
rect -3040 16285 -3035 16315
rect -3005 16285 -3000 16315
rect -3040 16155 -3000 16285
rect -3040 16125 -3035 16155
rect -3005 16125 -3000 16155
rect -3040 15995 -3000 16125
rect -3040 15965 -3035 15995
rect -3005 15965 -3000 15995
rect -3040 15960 -3000 15965
rect -2960 16475 -2920 16480
rect -2960 16445 -2955 16475
rect -2925 16445 -2920 16475
rect -2960 16315 -2920 16445
rect -2960 16285 -2955 16315
rect -2925 16285 -2920 16315
rect -2960 16155 -2920 16285
rect -2960 16125 -2955 16155
rect -2925 16125 -2920 16155
rect -2960 15995 -2920 16125
rect -2960 15965 -2955 15995
rect -2925 15965 -2920 15995
rect -2960 15960 -2920 15965
rect -2880 16475 -2840 16480
rect -2880 16445 -2875 16475
rect -2845 16445 -2840 16475
rect -2880 16315 -2840 16445
rect -2880 16285 -2875 16315
rect -2845 16285 -2840 16315
rect -2880 16155 -2840 16285
rect -2880 16125 -2875 16155
rect -2845 16125 -2840 16155
rect -2880 15995 -2840 16125
rect -2880 15965 -2875 15995
rect -2845 15965 -2840 15995
rect -2880 15960 -2840 15965
rect -2800 16475 -2760 16480
rect -2800 16445 -2795 16475
rect -2765 16445 -2760 16475
rect -2800 16315 -2760 16445
rect -2800 16285 -2795 16315
rect -2765 16285 -2760 16315
rect -2800 16155 -2760 16285
rect -2800 16125 -2795 16155
rect -2765 16125 -2760 16155
rect -2800 15995 -2760 16125
rect -2800 15965 -2795 15995
rect -2765 15965 -2760 15995
rect -2800 15960 -2760 15965
rect -2720 16475 -2680 16480
rect -2720 16445 -2715 16475
rect -2685 16445 -2680 16475
rect -2720 16315 -2680 16445
rect -2720 16285 -2715 16315
rect -2685 16285 -2680 16315
rect -2720 16155 -2680 16285
rect -2720 16125 -2715 16155
rect -2685 16125 -2680 16155
rect -2720 15995 -2680 16125
rect -2720 15965 -2715 15995
rect -2685 15965 -2680 15995
rect -2720 15960 -2680 15965
rect -2640 16475 -2600 16480
rect -2640 16445 -2635 16475
rect -2605 16445 -2600 16475
rect -2640 16315 -2600 16445
rect -2640 16285 -2635 16315
rect -2605 16285 -2600 16315
rect -2640 16155 -2600 16285
rect -2640 16125 -2635 16155
rect -2605 16125 -2600 16155
rect -2640 15995 -2600 16125
rect -2640 15965 -2635 15995
rect -2605 15965 -2600 15995
rect -2640 15960 -2600 15965
rect -2560 16475 -2520 16480
rect -2560 16445 -2555 16475
rect -2525 16445 -2520 16475
rect -2560 16315 -2520 16445
rect -2560 16285 -2555 16315
rect -2525 16285 -2520 16315
rect -2560 16155 -2520 16285
rect -2560 16125 -2555 16155
rect -2525 16125 -2520 16155
rect -2560 15995 -2520 16125
rect -2560 15965 -2555 15995
rect -2525 15965 -2520 15995
rect -2560 15960 -2520 15965
rect -2480 16475 -2440 16480
rect -2480 16445 -2475 16475
rect -2445 16445 -2440 16475
rect -2480 16315 -2440 16445
rect -2480 16285 -2475 16315
rect -2445 16285 -2440 16315
rect -2480 16155 -2440 16285
rect -2480 16125 -2475 16155
rect -2445 16125 -2440 16155
rect -2480 15995 -2440 16125
rect -2480 15965 -2475 15995
rect -2445 15965 -2440 15995
rect -2480 15960 -2440 15965
rect -2400 16475 -2360 16480
rect -2400 16445 -2395 16475
rect -2365 16445 -2360 16475
rect -2400 16315 -2360 16445
rect -2400 16285 -2395 16315
rect -2365 16285 -2360 16315
rect -2400 16155 -2360 16285
rect -2400 16125 -2395 16155
rect -2365 16125 -2360 16155
rect -2400 15995 -2360 16125
rect -2400 15965 -2395 15995
rect -2365 15965 -2360 15995
rect -2400 15960 -2360 15965
rect -2320 16475 -2280 16480
rect -2320 16445 -2315 16475
rect -2285 16445 -2280 16475
rect -2320 16315 -2280 16445
rect -2320 16285 -2315 16315
rect -2285 16285 -2280 16315
rect -2320 16155 -2280 16285
rect -2320 16125 -2315 16155
rect -2285 16125 -2280 16155
rect -2320 15995 -2280 16125
rect -2320 15965 -2315 15995
rect -2285 15965 -2280 15995
rect -2320 15960 -2280 15965
rect -2240 16475 -2200 16480
rect -2240 16445 -2235 16475
rect -2205 16445 -2200 16475
rect -2240 16315 -2200 16445
rect -2240 16285 -2235 16315
rect -2205 16285 -2200 16315
rect -2240 16155 -2200 16285
rect -2240 16125 -2235 16155
rect -2205 16125 -2200 16155
rect -2240 15995 -2200 16125
rect -2240 15965 -2235 15995
rect -2205 15965 -2200 15995
rect -2240 15960 -2200 15965
rect -2160 16475 -2120 16480
rect -2160 16445 -2155 16475
rect -2125 16445 -2120 16475
rect -2160 16315 -2120 16445
rect -2160 16285 -2155 16315
rect -2125 16285 -2120 16315
rect -2160 16155 -2120 16285
rect -2160 16125 -2155 16155
rect -2125 16125 -2120 16155
rect -2160 15995 -2120 16125
rect -2160 15965 -2155 15995
rect -2125 15965 -2120 15995
rect -2160 15960 -2120 15965
rect -2080 16475 -2040 16480
rect -2080 16445 -2075 16475
rect -2045 16445 -2040 16475
rect -2080 16315 -2040 16445
rect -2080 16285 -2075 16315
rect -2045 16285 -2040 16315
rect -2080 16155 -2040 16285
rect -2080 16125 -2075 16155
rect -2045 16125 -2040 16155
rect -2080 15995 -2040 16125
rect -2080 15965 -2075 15995
rect -2045 15965 -2040 15995
rect -2080 15960 -2040 15965
rect -2000 16475 -1960 16480
rect -2000 16445 -1995 16475
rect -1965 16445 -1960 16475
rect -2000 16315 -1960 16445
rect -2000 16285 -1995 16315
rect -1965 16285 -1960 16315
rect -2000 16155 -1960 16285
rect -2000 16125 -1995 16155
rect -1965 16125 -1960 16155
rect -2000 15995 -1960 16125
rect -2000 15965 -1995 15995
rect -1965 15965 -1960 15995
rect -2000 15960 -1960 15965
rect -1840 16475 -1800 16480
rect -1840 16445 -1835 16475
rect -1805 16445 -1800 16475
rect -1840 16315 -1800 16445
rect -1840 16285 -1835 16315
rect -1805 16285 -1800 16315
rect -1840 16155 -1800 16285
rect -1840 16125 -1835 16155
rect -1805 16125 -1800 16155
rect -1840 15995 -1800 16125
rect -1840 15965 -1835 15995
rect -1805 15965 -1800 15995
rect -1840 15960 -1800 15965
rect -1760 16475 -1720 16480
rect -1760 16445 -1755 16475
rect -1725 16445 -1720 16475
rect -1760 16315 -1720 16445
rect -1760 16285 -1755 16315
rect -1725 16285 -1720 16315
rect -1760 16155 -1720 16285
rect -1760 16125 -1755 16155
rect -1725 16125 -1720 16155
rect -1760 15995 -1720 16125
rect -1760 15965 -1755 15995
rect -1725 15965 -1720 15995
rect -1760 15960 -1720 15965
rect -1680 16475 -1640 16524
rect -1520 17876 -1480 18005
rect -1520 17844 -1516 17876
rect -1484 17844 -1480 17876
rect -1520 17796 -1480 17844
rect -1520 17764 -1516 17796
rect -1484 17764 -1480 17796
rect -1520 17716 -1480 17764
rect -1520 17684 -1516 17716
rect -1484 17684 -1480 17716
rect -1520 17636 -1480 17684
rect -1520 17604 -1516 17636
rect -1484 17604 -1480 17636
rect -1520 17556 -1480 17604
rect -1520 17524 -1516 17556
rect -1484 17524 -1480 17556
rect -1520 17476 -1480 17524
rect -1520 17444 -1516 17476
rect -1484 17444 -1480 17476
rect -1520 17396 -1480 17444
rect -1520 17364 -1516 17396
rect -1484 17364 -1480 17396
rect -1520 17316 -1480 17364
rect -1520 17284 -1516 17316
rect -1484 17284 -1480 17316
rect -1520 17236 -1480 17284
rect -1520 17204 -1516 17236
rect -1484 17204 -1480 17236
rect -1520 17156 -1480 17204
rect -1520 17124 -1516 17156
rect -1484 17124 -1480 17156
rect -1520 17076 -1480 17124
rect -1520 17044 -1516 17076
rect -1484 17044 -1480 17076
rect -1520 16996 -1480 17044
rect -1520 16964 -1516 16996
rect -1484 16964 -1480 16996
rect -1520 16916 -1480 16964
rect -1520 16884 -1516 16916
rect -1484 16884 -1480 16916
rect -1520 16836 -1480 16884
rect -1520 16804 -1516 16836
rect -1484 16804 -1480 16836
rect -1520 16756 -1480 16804
rect -1520 16724 -1516 16756
rect -1484 16724 -1480 16756
rect -1520 16636 -1480 16724
rect -1520 16604 -1516 16636
rect -1484 16604 -1480 16636
rect -1520 16556 -1480 16604
rect -1520 16524 -1516 16556
rect -1484 16524 -1480 16556
rect -1680 16445 -1675 16475
rect -1645 16445 -1640 16475
rect -1680 16315 -1640 16445
rect -1680 16285 -1675 16315
rect -1645 16285 -1640 16315
rect -1680 16155 -1640 16285
rect -1680 16125 -1675 16155
rect -1645 16125 -1640 16155
rect -1680 15995 -1640 16125
rect -1680 15965 -1675 15995
rect -1645 15965 -1640 15995
rect -1680 15960 -1640 15965
rect -1600 16475 -1560 16480
rect -1600 16445 -1595 16475
rect -1565 16445 -1560 16475
rect -1600 16315 -1560 16445
rect -1600 16285 -1595 16315
rect -1565 16285 -1560 16315
rect -1600 16155 -1560 16285
rect -1600 16125 -1595 16155
rect -1565 16125 -1560 16155
rect -1600 15995 -1560 16125
rect -1600 15965 -1595 15995
rect -1565 15965 -1560 15995
rect -1600 15960 -1560 15965
rect -1520 16475 -1480 16524
rect -1360 18035 -1320 18164
rect -1360 18005 -1355 18035
rect -1325 18005 -1320 18035
rect -1360 17876 -1320 18005
rect -1360 17844 -1356 17876
rect -1324 17844 -1320 17876
rect -1360 17796 -1320 17844
rect -1360 17764 -1356 17796
rect -1324 17764 -1320 17796
rect -1360 17716 -1320 17764
rect -1360 17684 -1356 17716
rect -1324 17684 -1320 17716
rect -1360 17636 -1320 17684
rect -1360 17604 -1356 17636
rect -1324 17604 -1320 17636
rect -1360 17556 -1320 17604
rect -1360 17524 -1356 17556
rect -1324 17524 -1320 17556
rect -1360 17476 -1320 17524
rect -1360 17444 -1356 17476
rect -1324 17444 -1320 17476
rect -1360 17396 -1320 17444
rect -1360 17364 -1356 17396
rect -1324 17364 -1320 17396
rect -1360 17316 -1320 17364
rect -1360 17284 -1356 17316
rect -1324 17284 -1320 17316
rect -1360 17236 -1320 17284
rect -1360 17204 -1356 17236
rect -1324 17204 -1320 17236
rect -1360 17156 -1320 17204
rect -1360 17124 -1356 17156
rect -1324 17124 -1320 17156
rect -1360 17076 -1320 17124
rect -1360 17044 -1356 17076
rect -1324 17044 -1320 17076
rect -1360 16996 -1320 17044
rect -1360 16964 -1356 16996
rect -1324 16964 -1320 16996
rect -1360 16916 -1320 16964
rect -1360 16884 -1356 16916
rect -1324 16884 -1320 16916
rect -1360 16836 -1320 16884
rect -1360 16804 -1356 16836
rect -1324 16804 -1320 16836
rect -1360 16756 -1320 16804
rect -1360 16724 -1356 16756
rect -1324 16724 -1320 16756
rect -1360 16636 -1320 16724
rect -1360 16604 -1356 16636
rect -1324 16604 -1320 16636
rect -1360 16556 -1320 16604
rect -1360 16524 -1356 16556
rect -1324 16524 -1320 16556
rect -1520 16445 -1515 16475
rect -1485 16445 -1480 16475
rect -1520 16315 -1480 16445
rect -1520 16285 -1515 16315
rect -1485 16285 -1480 16315
rect -1520 16155 -1480 16285
rect -1520 16125 -1515 16155
rect -1485 16125 -1480 16155
rect -1520 15995 -1480 16125
rect -1520 15965 -1515 15995
rect -1485 15965 -1480 15995
rect -1520 15960 -1480 15965
rect -1440 16475 -1400 16480
rect -1440 16445 -1435 16475
rect -1405 16445 -1400 16475
rect -1440 16315 -1400 16445
rect -1440 16285 -1435 16315
rect -1405 16285 -1400 16315
rect -1440 16155 -1400 16285
rect -1440 16125 -1435 16155
rect -1405 16125 -1400 16155
rect -1440 15995 -1400 16125
rect -1440 15965 -1435 15995
rect -1405 15965 -1400 15995
rect -1440 15960 -1400 15965
rect -1360 16475 -1320 16524
rect -1360 16445 -1355 16475
rect -1325 16445 -1320 16475
rect -1360 16315 -1320 16445
rect -1360 16285 -1355 16315
rect -1325 16285 -1320 16315
rect -1360 16155 -1320 16285
rect -1280 20115 -1240 20120
rect -1280 20085 -1275 20115
rect -1245 20085 -1240 20115
rect -1280 16235 -1240 20085
rect -1200 20035 -1160 20165
rect -1200 20005 -1195 20035
rect -1165 20005 -1160 20035
rect -1200 19955 -1160 20005
rect -1040 20875 -1000 20925
rect -1040 20845 -1035 20875
rect -1005 20845 -1000 20875
rect -1040 20795 -1000 20845
rect -1040 20765 -1035 20795
rect -1005 20765 -1000 20795
rect -1040 20435 -1000 20765
rect -1040 20405 -1035 20435
rect -1005 20405 -1000 20435
rect -1040 20355 -1000 20405
rect -1040 20325 -1035 20355
rect -1005 20325 -1000 20355
rect -1040 20195 -1000 20325
rect -1040 20165 -1035 20195
rect -1005 20165 -1000 20195
rect -1040 20035 -1000 20165
rect -960 20115 -920 21480
rect -960 20085 -955 20115
rect -925 20085 -920 20115
rect -960 20080 -920 20085
rect -880 21435 -840 21480
rect -880 21405 -875 21435
rect -845 21405 -840 21435
rect -880 21275 -840 21405
rect -880 21245 -875 21275
rect -845 21245 -840 21275
rect -880 21115 -840 21245
rect -880 21085 -875 21115
rect -845 21085 -840 21115
rect -880 20955 -840 21085
rect -880 20925 -875 20955
rect -845 20925 -840 20955
rect -880 20875 -840 20925
rect -880 20845 -875 20875
rect -845 20845 -840 20875
rect -880 20795 -840 20845
rect -880 20765 -875 20795
rect -845 20765 -840 20795
rect -880 20435 -840 20765
rect -880 20405 -875 20435
rect -845 20405 -840 20435
rect -880 20355 -840 20405
rect -880 20325 -875 20355
rect -845 20325 -840 20355
rect -880 20195 -840 20325
rect -880 20165 -875 20195
rect -845 20165 -840 20195
rect -1040 20005 -1035 20035
rect -1005 20005 -1000 20035
rect -1200 19925 -1195 19955
rect -1165 19925 -1160 19955
rect -1200 19876 -1160 19925
rect -1200 19844 -1196 19876
rect -1164 19844 -1160 19876
rect -1200 19796 -1160 19844
rect -1200 19764 -1196 19796
rect -1164 19764 -1160 19796
rect -1200 19716 -1160 19764
rect -1200 19684 -1196 19716
rect -1164 19684 -1160 19716
rect -1200 19636 -1160 19684
rect -1200 19604 -1196 19636
rect -1164 19604 -1160 19636
rect -1200 19556 -1160 19604
rect -1200 19524 -1196 19556
rect -1164 19524 -1160 19556
rect -1200 19476 -1160 19524
rect -1200 19444 -1196 19476
rect -1164 19444 -1160 19476
rect -1200 19396 -1160 19444
rect -1200 19364 -1196 19396
rect -1164 19364 -1160 19396
rect -1200 19316 -1160 19364
rect -1200 19284 -1196 19316
rect -1164 19284 -1160 19316
rect -1200 19236 -1160 19284
rect -1200 19204 -1196 19236
rect -1164 19204 -1160 19236
rect -1200 19156 -1160 19204
rect -1200 19124 -1196 19156
rect -1164 19124 -1160 19156
rect -1200 19076 -1160 19124
rect -1200 19044 -1196 19076
rect -1164 19044 -1160 19076
rect -1200 18996 -1160 19044
rect -1200 18964 -1196 18996
rect -1164 18964 -1160 18996
rect -1200 18916 -1160 18964
rect -1200 18884 -1196 18916
rect -1164 18884 -1160 18916
rect -1200 18835 -1160 18884
rect -1200 18805 -1195 18835
rect -1165 18805 -1160 18835
rect -1200 18756 -1160 18805
rect -1200 18724 -1196 18756
rect -1164 18724 -1160 18756
rect -1200 18676 -1160 18724
rect -1200 18644 -1196 18676
rect -1164 18644 -1160 18676
rect -1200 18596 -1160 18644
rect -1200 18564 -1196 18596
rect -1164 18564 -1160 18596
rect -1200 18516 -1160 18564
rect -1200 18484 -1196 18516
rect -1164 18484 -1160 18516
rect -1200 18436 -1160 18484
rect -1200 18404 -1196 18436
rect -1164 18404 -1160 18436
rect -1200 18356 -1160 18404
rect -1200 18324 -1196 18356
rect -1164 18324 -1160 18356
rect -1200 18276 -1160 18324
rect -1200 18244 -1196 18276
rect -1164 18244 -1160 18276
rect -1200 18196 -1160 18244
rect -1200 18164 -1196 18196
rect -1164 18164 -1160 18196
rect -1200 18035 -1160 18164
rect -1200 18005 -1195 18035
rect -1165 18005 -1160 18035
rect -1200 18000 -1160 18005
rect -1120 19955 -1080 19960
rect -1120 19925 -1115 19955
rect -1085 19925 -1080 19955
rect -1280 16205 -1275 16235
rect -1245 16205 -1240 16235
rect -1280 16200 -1240 16205
rect -1200 17876 -1160 17880
rect -1200 17844 -1196 17876
rect -1164 17844 -1160 17876
rect -1200 17796 -1160 17844
rect -1200 17764 -1196 17796
rect -1164 17764 -1160 17796
rect -1200 17716 -1160 17764
rect -1200 17684 -1196 17716
rect -1164 17684 -1160 17716
rect -1200 17636 -1160 17684
rect -1200 17604 -1196 17636
rect -1164 17604 -1160 17636
rect -1200 17556 -1160 17604
rect -1200 17524 -1196 17556
rect -1164 17524 -1160 17556
rect -1200 17476 -1160 17524
rect -1200 17444 -1196 17476
rect -1164 17444 -1160 17476
rect -1200 17396 -1160 17444
rect -1200 17364 -1196 17396
rect -1164 17364 -1160 17396
rect -1200 17316 -1160 17364
rect -1200 17284 -1196 17316
rect -1164 17284 -1160 17316
rect -1200 17236 -1160 17284
rect -1200 17204 -1196 17236
rect -1164 17204 -1160 17236
rect -1200 17156 -1160 17204
rect -1200 17124 -1196 17156
rect -1164 17124 -1160 17156
rect -1200 17076 -1160 17124
rect -1200 17044 -1196 17076
rect -1164 17044 -1160 17076
rect -1200 16996 -1160 17044
rect -1200 16964 -1196 16996
rect -1164 16964 -1160 16996
rect -1200 16916 -1160 16964
rect -1200 16884 -1196 16916
rect -1164 16884 -1160 16916
rect -1200 16836 -1160 16884
rect -1200 16804 -1196 16836
rect -1164 16804 -1160 16836
rect -1200 16756 -1160 16804
rect -1200 16724 -1196 16756
rect -1164 16724 -1160 16756
rect -1200 16636 -1160 16724
rect -1200 16604 -1196 16636
rect -1164 16604 -1160 16636
rect -1200 16556 -1160 16604
rect -1200 16524 -1196 16556
rect -1164 16524 -1160 16556
rect -1200 16475 -1160 16524
rect -1200 16445 -1195 16475
rect -1165 16445 -1160 16475
rect -1200 16315 -1160 16445
rect -1200 16285 -1195 16315
rect -1165 16285 -1160 16315
rect -1360 16125 -1355 16155
rect -1325 16125 -1320 16155
rect -1360 15995 -1320 16125
rect -1360 15965 -1355 15995
rect -1325 15965 -1320 15995
rect -1360 15960 -1320 15965
rect -1200 16155 -1160 16285
rect -1200 16125 -1195 16155
rect -1165 16125 -1160 16155
rect -1200 15995 -1160 16125
rect -1120 16075 -1080 19925
rect -1120 16045 -1115 16075
rect -1085 16045 -1080 16075
rect -1120 16040 -1080 16045
rect -1040 19876 -1000 20005
rect -1040 19844 -1036 19876
rect -1004 19844 -1000 19876
rect -1040 19796 -1000 19844
rect -1040 19764 -1036 19796
rect -1004 19764 -1000 19796
rect -1040 19716 -1000 19764
rect -1040 19684 -1036 19716
rect -1004 19684 -1000 19716
rect -1040 19636 -1000 19684
rect -1040 19604 -1036 19636
rect -1004 19604 -1000 19636
rect -1040 19556 -1000 19604
rect -1040 19524 -1036 19556
rect -1004 19524 -1000 19556
rect -1040 19476 -1000 19524
rect -1040 19444 -1036 19476
rect -1004 19444 -1000 19476
rect -1040 19396 -1000 19444
rect -1040 19364 -1036 19396
rect -1004 19364 -1000 19396
rect -1040 19316 -1000 19364
rect -1040 19284 -1036 19316
rect -1004 19284 -1000 19316
rect -1040 19236 -1000 19284
rect -1040 19204 -1036 19236
rect -1004 19204 -1000 19236
rect -1040 19156 -1000 19204
rect -1040 19124 -1036 19156
rect -1004 19124 -1000 19156
rect -1040 19076 -1000 19124
rect -1040 19044 -1036 19076
rect -1004 19044 -1000 19076
rect -1040 18996 -1000 19044
rect -1040 18964 -1036 18996
rect -1004 18964 -1000 18996
rect -1040 18916 -1000 18964
rect -1040 18884 -1036 18916
rect -1004 18884 -1000 18916
rect -1040 18835 -1000 18884
rect -1040 18805 -1035 18835
rect -1005 18805 -1000 18835
rect -1040 18756 -1000 18805
rect -1040 18724 -1036 18756
rect -1004 18724 -1000 18756
rect -1040 18676 -1000 18724
rect -1040 18644 -1036 18676
rect -1004 18644 -1000 18676
rect -1040 18596 -1000 18644
rect -1040 18564 -1036 18596
rect -1004 18564 -1000 18596
rect -1040 18516 -1000 18564
rect -1040 18484 -1036 18516
rect -1004 18484 -1000 18516
rect -1040 18436 -1000 18484
rect -1040 18404 -1036 18436
rect -1004 18404 -1000 18436
rect -1040 18356 -1000 18404
rect -1040 18324 -1036 18356
rect -1004 18324 -1000 18356
rect -1040 18276 -1000 18324
rect -1040 18244 -1036 18276
rect -1004 18244 -1000 18276
rect -1040 18196 -1000 18244
rect -1040 18164 -1036 18196
rect -1004 18164 -1000 18196
rect -1040 18035 -1000 18164
rect -880 20035 -840 20165
rect -880 20005 -875 20035
rect -845 20005 -840 20035
rect -880 19876 -840 20005
rect -800 19955 -760 21480
rect -800 19925 -795 19955
rect -765 19925 -760 19955
rect -800 19920 -760 19925
rect -720 21435 -680 21480
rect -720 21405 -715 21435
rect -685 21405 -680 21435
rect -720 21275 -680 21405
rect -720 21245 -715 21275
rect -685 21245 -680 21275
rect -720 21115 -680 21245
rect -720 21085 -715 21115
rect -685 21085 -680 21115
rect -720 20955 -680 21085
rect -640 21035 -600 21480
rect -640 21005 -635 21035
rect -605 21005 -600 21035
rect -640 21000 -600 21005
rect -560 21435 -520 21480
rect -560 21405 -555 21435
rect -525 21405 -520 21435
rect -560 21275 -520 21405
rect -560 21245 -555 21275
rect -525 21245 -520 21275
rect -560 21115 -520 21245
rect -560 21085 -555 21115
rect -525 21085 -520 21115
rect -720 20925 -715 20955
rect -685 20925 -680 20955
rect -720 20875 -680 20925
rect -720 20845 -715 20875
rect -685 20845 -680 20875
rect -720 20795 -680 20845
rect -720 20765 -715 20795
rect -685 20765 -680 20795
rect -720 20435 -680 20765
rect -720 20405 -715 20435
rect -685 20405 -680 20435
rect -720 20355 -680 20405
rect -720 20325 -715 20355
rect -685 20325 -680 20355
rect -720 20195 -680 20325
rect -560 20955 -520 21085
rect -560 20925 -555 20955
rect -525 20925 -520 20955
rect -560 20875 -520 20925
rect -560 20845 -555 20875
rect -525 20845 -520 20875
rect -560 20795 -520 20845
rect -560 20765 -555 20795
rect -525 20765 -520 20795
rect -560 20435 -520 20765
rect 20520 20675 20560 20680
rect 20520 20645 20525 20675
rect 20555 20645 20560 20675
rect 20520 20515 20560 20645
rect 20520 20485 20525 20515
rect 20555 20485 20560 20515
rect 20520 20480 20560 20485
rect 20600 20675 20640 20680
rect 20600 20645 20605 20675
rect 20635 20645 20640 20675
rect 20600 20515 20640 20645
rect 20600 20485 20605 20515
rect 20635 20485 20640 20515
rect 20600 20480 20640 20485
rect 20680 20675 20720 20680
rect 20680 20645 20685 20675
rect 20715 20645 20720 20675
rect 20680 20515 20720 20645
rect 20680 20485 20685 20515
rect 20715 20485 20720 20515
rect 20680 20480 20720 20485
rect 20760 20675 20800 20680
rect 20760 20645 20765 20675
rect 20795 20645 20800 20675
rect 20760 20515 20800 20645
rect 20760 20485 20765 20515
rect 20795 20485 20800 20515
rect 20760 20480 20800 20485
rect 20840 20675 20880 20680
rect 20840 20645 20845 20675
rect 20875 20645 20880 20675
rect 20840 20515 20880 20645
rect 20840 20485 20845 20515
rect 20875 20485 20880 20515
rect 20840 20480 20880 20485
rect 20920 20675 20960 20680
rect 20920 20645 20925 20675
rect 20955 20645 20960 20675
rect 20920 20515 20960 20645
rect 20920 20485 20925 20515
rect 20955 20485 20960 20515
rect 20920 20480 20960 20485
rect 21000 20675 21040 20680
rect 21000 20645 21005 20675
rect 21035 20645 21040 20675
rect 21000 20515 21040 20645
rect 21000 20485 21005 20515
rect 21035 20485 21040 20515
rect 21000 20480 21040 20485
rect 21080 20675 21120 20680
rect 21080 20645 21085 20675
rect 21115 20645 21120 20675
rect 21080 20515 21120 20645
rect 21080 20485 21085 20515
rect 21115 20485 21120 20515
rect 21080 20480 21120 20485
rect 21160 20675 21200 20680
rect 21160 20645 21165 20675
rect 21195 20645 21200 20675
rect 21160 20515 21200 20645
rect 21160 20485 21165 20515
rect 21195 20485 21200 20515
rect 21160 20480 21200 20485
rect 21240 20675 21280 20680
rect 21240 20645 21245 20675
rect 21275 20645 21280 20675
rect 21240 20515 21280 20645
rect 21240 20485 21245 20515
rect 21275 20485 21280 20515
rect 21240 20480 21280 20485
rect 21320 20675 21360 20680
rect 21320 20645 21325 20675
rect 21355 20645 21360 20675
rect 21320 20515 21360 20645
rect 21320 20485 21325 20515
rect 21355 20485 21360 20515
rect 21320 20480 21360 20485
rect 21400 20675 21440 20680
rect 21400 20645 21405 20675
rect 21435 20645 21440 20675
rect 21400 20515 21440 20645
rect 21400 20485 21405 20515
rect 21435 20485 21440 20515
rect 21400 20480 21440 20485
rect 21480 20675 21520 20680
rect 21480 20645 21485 20675
rect 21515 20645 21520 20675
rect 21480 20515 21520 20645
rect 21480 20485 21485 20515
rect 21515 20485 21520 20515
rect 21480 20480 21520 20485
rect 21560 20675 21600 20680
rect 21560 20645 21565 20675
rect 21595 20645 21600 20675
rect 21560 20515 21600 20645
rect 21560 20485 21565 20515
rect 21595 20485 21600 20515
rect 21560 20480 21600 20485
rect -560 20405 -555 20435
rect -525 20405 -520 20435
rect -560 20355 -520 20405
rect -560 20325 -555 20355
rect -525 20325 -520 20355
rect -720 20165 -715 20195
rect -685 20165 -680 20195
rect -720 20035 -680 20165
rect -720 20005 -715 20035
rect -685 20005 -680 20035
rect -880 19844 -876 19876
rect -844 19844 -840 19876
rect -880 19796 -840 19844
rect -880 19764 -876 19796
rect -844 19764 -840 19796
rect -880 19716 -840 19764
rect -880 19684 -876 19716
rect -844 19684 -840 19716
rect -880 19636 -840 19684
rect -880 19604 -876 19636
rect -844 19604 -840 19636
rect -880 19556 -840 19604
rect -880 19524 -876 19556
rect -844 19524 -840 19556
rect -880 19476 -840 19524
rect -880 19444 -876 19476
rect -844 19444 -840 19476
rect -880 19396 -840 19444
rect -880 19364 -876 19396
rect -844 19364 -840 19396
rect -880 19316 -840 19364
rect -880 19284 -876 19316
rect -844 19284 -840 19316
rect -880 19236 -840 19284
rect -880 19204 -876 19236
rect -844 19204 -840 19236
rect -880 19156 -840 19204
rect -880 19124 -876 19156
rect -844 19124 -840 19156
rect -880 19076 -840 19124
rect -880 19044 -876 19076
rect -844 19044 -840 19076
rect -880 18996 -840 19044
rect -880 18964 -876 18996
rect -844 18964 -840 18996
rect -880 18916 -840 18964
rect -880 18884 -876 18916
rect -844 18884 -840 18916
rect -880 18835 -840 18884
rect -880 18805 -875 18835
rect -845 18805 -840 18835
rect -880 18756 -840 18805
rect -880 18724 -876 18756
rect -844 18724 -840 18756
rect -880 18676 -840 18724
rect -880 18644 -876 18676
rect -844 18644 -840 18676
rect -880 18596 -840 18644
rect -880 18564 -876 18596
rect -844 18564 -840 18596
rect -880 18516 -840 18564
rect -880 18484 -876 18516
rect -844 18484 -840 18516
rect -880 18436 -840 18484
rect -880 18404 -876 18436
rect -844 18404 -840 18436
rect -880 18356 -840 18404
rect -880 18324 -876 18356
rect -844 18324 -840 18356
rect -880 18276 -840 18324
rect -880 18244 -876 18276
rect -844 18244 -840 18276
rect -880 18196 -840 18244
rect -880 18164 -876 18196
rect -844 18164 -840 18196
rect -1040 18005 -1035 18035
rect -1005 18005 -1000 18035
rect -1040 17876 -1000 18005
rect -1040 17844 -1036 17876
rect -1004 17844 -1000 17876
rect -1040 17796 -1000 17844
rect -1040 17764 -1036 17796
rect -1004 17764 -1000 17796
rect -1040 17716 -1000 17764
rect -1040 17684 -1036 17716
rect -1004 17684 -1000 17716
rect -1040 17636 -1000 17684
rect -1040 17604 -1036 17636
rect -1004 17604 -1000 17636
rect -1040 17556 -1000 17604
rect -1040 17524 -1036 17556
rect -1004 17524 -1000 17556
rect -1040 17476 -1000 17524
rect -1040 17444 -1036 17476
rect -1004 17444 -1000 17476
rect -1040 17396 -1000 17444
rect -1040 17364 -1036 17396
rect -1004 17364 -1000 17396
rect -1040 17316 -1000 17364
rect -1040 17284 -1036 17316
rect -1004 17284 -1000 17316
rect -1040 17236 -1000 17284
rect -1040 17204 -1036 17236
rect -1004 17204 -1000 17236
rect -1040 17156 -1000 17204
rect -1040 17124 -1036 17156
rect -1004 17124 -1000 17156
rect -1040 17076 -1000 17124
rect -1040 17044 -1036 17076
rect -1004 17044 -1000 17076
rect -1040 16996 -1000 17044
rect -1040 16964 -1036 16996
rect -1004 16964 -1000 16996
rect -1040 16916 -1000 16964
rect -1040 16884 -1036 16916
rect -1004 16884 -1000 16916
rect -1040 16836 -1000 16884
rect -1040 16804 -1036 16836
rect -1004 16804 -1000 16836
rect -1040 16756 -1000 16804
rect -1040 16724 -1036 16756
rect -1004 16724 -1000 16756
rect -1040 16636 -1000 16724
rect -1040 16604 -1036 16636
rect -1004 16604 -1000 16636
rect -1040 16556 -1000 16604
rect -1040 16524 -1036 16556
rect -1004 16524 -1000 16556
rect -1040 16475 -1000 16524
rect -1040 16445 -1035 16475
rect -1005 16445 -1000 16475
rect -1040 16315 -1000 16445
rect -1040 16285 -1035 16315
rect -1005 16285 -1000 16315
rect -1040 16155 -1000 16285
rect -1040 16125 -1035 16155
rect -1005 16125 -1000 16155
rect -1200 15965 -1195 15995
rect -1165 15965 -1160 15995
rect -1200 15960 -1160 15965
rect -1040 15995 -1000 16125
rect -1040 15965 -1035 15995
rect -1005 15965 -1000 15995
rect -1040 15920 -1000 15965
rect -960 18115 -920 18120
rect -960 18085 -955 18115
rect -925 18085 -920 18115
rect -960 15920 -920 18085
rect -880 18035 -840 18164
rect -880 18005 -875 18035
rect -845 18005 -840 18035
rect -880 17876 -840 18005
rect -720 19876 -680 20005
rect -720 19844 -716 19876
rect -684 19844 -680 19876
rect -720 19796 -680 19844
rect -720 19764 -716 19796
rect -684 19764 -680 19796
rect -720 19716 -680 19764
rect -720 19684 -716 19716
rect -684 19684 -680 19716
rect -720 19636 -680 19684
rect -720 19604 -716 19636
rect -684 19604 -680 19636
rect -720 19556 -680 19604
rect -720 19524 -716 19556
rect -684 19524 -680 19556
rect -720 19476 -680 19524
rect -720 19444 -716 19476
rect -684 19444 -680 19476
rect -720 19396 -680 19444
rect -720 19364 -716 19396
rect -684 19364 -680 19396
rect -720 19316 -680 19364
rect -720 19284 -716 19316
rect -684 19284 -680 19316
rect -720 19236 -680 19284
rect -720 19204 -716 19236
rect -684 19204 -680 19236
rect -720 19156 -680 19204
rect -720 19124 -716 19156
rect -684 19124 -680 19156
rect -720 19076 -680 19124
rect -720 19044 -716 19076
rect -684 19044 -680 19076
rect -720 18996 -680 19044
rect -720 18964 -716 18996
rect -684 18964 -680 18996
rect -720 18916 -680 18964
rect -720 18884 -716 18916
rect -684 18884 -680 18916
rect -720 18835 -680 18884
rect -720 18805 -715 18835
rect -685 18805 -680 18835
rect -720 18756 -680 18805
rect -640 20275 -600 20280
rect -640 20245 -635 20275
rect -605 20245 -600 20275
rect -640 18835 -600 20245
rect -640 18805 -635 18835
rect -605 18805 -600 18835
rect -640 18800 -600 18805
rect -560 20195 -520 20325
rect -560 20165 -555 20195
rect -525 20165 -520 20195
rect -560 20035 -520 20165
rect -560 20005 -555 20035
rect -525 20005 -520 20035
rect -560 19876 -520 20005
rect -560 19844 -556 19876
rect -524 19844 -520 19876
rect -560 19796 -520 19844
rect 20520 20035 20560 20040
rect 20520 20005 20525 20035
rect 20555 20005 20560 20035
rect 20520 19875 20560 20005
rect 20520 19845 20525 19875
rect 20555 19845 20560 19875
rect 20520 19840 20560 19845
rect 20600 20035 20640 20040
rect 20600 20005 20605 20035
rect 20635 20005 20640 20035
rect 20600 19875 20640 20005
rect 20600 19845 20605 19875
rect 20635 19845 20640 19875
rect 20600 19840 20640 19845
rect 20680 20035 20720 20040
rect 20680 20005 20685 20035
rect 20715 20005 20720 20035
rect 20680 19875 20720 20005
rect 20680 19845 20685 19875
rect 20715 19845 20720 19875
rect 20680 19840 20720 19845
rect 20760 20035 20800 20040
rect 20760 20005 20765 20035
rect 20795 20005 20800 20035
rect 20760 19875 20800 20005
rect 20760 19845 20765 19875
rect 20795 19845 20800 19875
rect 20760 19840 20800 19845
rect 20840 20035 20880 20040
rect 20840 20005 20845 20035
rect 20875 20005 20880 20035
rect 20840 19875 20880 20005
rect 20840 19845 20845 19875
rect 20875 19845 20880 19875
rect 20840 19840 20880 19845
rect 20920 20035 20960 20040
rect 20920 20005 20925 20035
rect 20955 20005 20960 20035
rect 20920 19875 20960 20005
rect 20920 19845 20925 19875
rect 20955 19845 20960 19875
rect 20920 19840 20960 19845
rect 21000 20035 21040 20040
rect 21000 20005 21005 20035
rect 21035 20005 21040 20035
rect 21000 19875 21040 20005
rect 21000 19845 21005 19875
rect 21035 19845 21040 19875
rect 21000 19840 21040 19845
rect 21080 20035 21120 20040
rect 21080 20005 21085 20035
rect 21115 20005 21120 20035
rect 21080 19875 21120 20005
rect 21080 19845 21085 19875
rect 21115 19845 21120 19875
rect 21080 19840 21120 19845
rect 21160 20035 21200 20040
rect 21160 20005 21165 20035
rect 21195 20005 21200 20035
rect 21160 19875 21200 20005
rect 21160 19845 21165 19875
rect 21195 19845 21200 19875
rect 21160 19840 21200 19845
rect 21240 20035 21280 20040
rect 21240 20005 21245 20035
rect 21275 20005 21280 20035
rect 21240 19875 21280 20005
rect 21240 19845 21245 19875
rect 21275 19845 21280 19875
rect 21240 19840 21280 19845
rect 21320 20035 21360 20040
rect 21320 20005 21325 20035
rect 21355 20005 21360 20035
rect 21320 19875 21360 20005
rect 21320 19845 21325 19875
rect 21355 19845 21360 19875
rect 21320 19840 21360 19845
rect 21400 20035 21440 20040
rect 21400 20005 21405 20035
rect 21435 20005 21440 20035
rect 21400 19875 21440 20005
rect 21400 19845 21405 19875
rect 21435 19845 21440 19875
rect 21400 19840 21440 19845
rect 21480 20035 21520 20040
rect 21480 20005 21485 20035
rect 21515 20005 21520 20035
rect 21480 19875 21520 20005
rect 21480 19845 21485 19875
rect 21515 19845 21520 19875
rect 21480 19840 21520 19845
rect 21560 20035 21600 20040
rect 21560 20005 21565 20035
rect 21595 20005 21600 20035
rect 21560 19875 21600 20005
rect 21560 19845 21565 19875
rect 21595 19845 21600 19875
rect 21560 19840 21600 19845
rect -560 19764 -556 19796
rect -524 19764 -520 19796
rect -560 19716 -520 19764
rect -560 19684 -556 19716
rect -524 19684 -520 19716
rect -560 19636 -520 19684
rect -560 19604 -556 19636
rect -524 19604 -520 19636
rect -560 19556 -520 19604
rect -560 19524 -556 19556
rect -524 19524 -520 19556
rect -560 19476 -520 19524
rect -560 19444 -556 19476
rect -524 19444 -520 19476
rect -560 19396 -520 19444
rect -560 19364 -556 19396
rect -524 19364 -520 19396
rect -560 19316 -520 19364
rect -560 19284 -556 19316
rect -524 19284 -520 19316
rect -560 19236 -520 19284
rect -560 19204 -556 19236
rect -524 19204 -520 19236
rect -560 19156 -520 19204
rect -560 19124 -556 19156
rect -524 19124 -520 19156
rect -560 19076 -520 19124
rect -560 19044 -556 19076
rect -524 19044 -520 19076
rect -560 18996 -520 19044
rect -560 18964 -556 18996
rect -524 18964 -520 18996
rect -560 18916 -520 18964
rect -560 18884 -556 18916
rect -524 18884 -520 18916
rect -720 18724 -716 18756
rect -684 18724 -680 18756
rect -720 18676 -680 18724
rect -720 18644 -716 18676
rect -684 18644 -680 18676
rect -720 18596 -680 18644
rect -720 18564 -716 18596
rect -684 18564 -680 18596
rect -720 18516 -680 18564
rect -720 18484 -716 18516
rect -684 18484 -680 18516
rect -720 18436 -680 18484
rect -720 18404 -716 18436
rect -684 18404 -680 18436
rect -720 18356 -680 18404
rect -720 18324 -716 18356
rect -684 18324 -680 18356
rect -720 18276 -680 18324
rect -720 18244 -716 18276
rect -684 18244 -680 18276
rect -720 18196 -680 18244
rect -720 18164 -716 18196
rect -684 18164 -680 18196
rect -720 18035 -680 18164
rect -720 18005 -715 18035
rect -685 18005 -680 18035
rect -880 17844 -876 17876
rect -844 17844 -840 17876
rect -880 17796 -840 17844
rect -880 17764 -876 17796
rect -844 17764 -840 17796
rect -880 17716 -840 17764
rect -880 17684 -876 17716
rect -844 17684 -840 17716
rect -880 17636 -840 17684
rect -880 17604 -876 17636
rect -844 17604 -840 17636
rect -880 17556 -840 17604
rect -880 17524 -876 17556
rect -844 17524 -840 17556
rect -880 17476 -840 17524
rect -880 17444 -876 17476
rect -844 17444 -840 17476
rect -880 17396 -840 17444
rect -880 17364 -876 17396
rect -844 17364 -840 17396
rect -880 17316 -840 17364
rect -880 17284 -876 17316
rect -844 17284 -840 17316
rect -880 17236 -840 17284
rect -880 17204 -876 17236
rect -844 17204 -840 17236
rect -880 17156 -840 17204
rect -880 17124 -876 17156
rect -844 17124 -840 17156
rect -880 17076 -840 17124
rect -880 17044 -876 17076
rect -844 17044 -840 17076
rect -880 16996 -840 17044
rect -880 16964 -876 16996
rect -844 16964 -840 16996
rect -880 16916 -840 16964
rect -880 16884 -876 16916
rect -844 16884 -840 16916
rect -880 16836 -840 16884
rect -880 16804 -876 16836
rect -844 16804 -840 16836
rect -880 16756 -840 16804
rect -880 16724 -876 16756
rect -844 16724 -840 16756
rect -880 16636 -840 16724
rect -880 16604 -876 16636
rect -844 16604 -840 16636
rect -880 16556 -840 16604
rect -880 16524 -876 16556
rect -844 16524 -840 16556
rect -880 16475 -840 16524
rect -880 16445 -875 16475
rect -845 16445 -840 16475
rect -880 16315 -840 16445
rect -880 16285 -875 16315
rect -845 16285 -840 16315
rect -880 16155 -840 16285
rect -880 16125 -875 16155
rect -845 16125 -840 16155
rect -880 15995 -840 16125
rect -880 15965 -875 15995
rect -845 15965 -840 15995
rect -880 15920 -840 15965
rect -800 17955 -760 17960
rect -800 17925 -795 17955
rect -765 17925 -760 17955
rect -800 15920 -760 17925
rect -720 17876 -680 18005
rect -720 17844 -716 17876
rect -684 17844 -680 17876
rect -720 17796 -680 17844
rect -720 17764 -716 17796
rect -684 17764 -680 17796
rect -720 17716 -680 17764
rect -720 17684 -716 17716
rect -684 17684 -680 17716
rect -720 17636 -680 17684
rect -720 17604 -716 17636
rect -684 17604 -680 17636
rect -720 17556 -680 17604
rect -720 17524 -716 17556
rect -684 17524 -680 17556
rect -720 17476 -680 17524
rect -720 17444 -716 17476
rect -684 17444 -680 17476
rect -720 17396 -680 17444
rect -720 17364 -716 17396
rect -684 17364 -680 17396
rect -720 17316 -680 17364
rect -720 17284 -716 17316
rect -684 17284 -680 17316
rect -720 17236 -680 17284
rect -720 17204 -716 17236
rect -684 17204 -680 17236
rect -720 17156 -680 17204
rect -720 17124 -716 17156
rect -684 17124 -680 17156
rect -720 17076 -680 17124
rect -720 17044 -716 17076
rect -684 17044 -680 17076
rect -720 16996 -680 17044
rect -720 16964 -716 16996
rect -684 16964 -680 16996
rect -720 16916 -680 16964
rect -720 16884 -716 16916
rect -684 16884 -680 16916
rect -720 16836 -680 16884
rect -720 16804 -716 16836
rect -684 16804 -680 16836
rect -720 16756 -680 16804
rect -720 16724 -716 16756
rect -684 16724 -680 16756
rect -720 16636 -680 16724
rect -720 16604 -716 16636
rect -684 16604 -680 16636
rect -720 16556 -680 16604
rect -720 16524 -716 16556
rect -684 16524 -680 16556
rect -720 16475 -680 16524
rect -720 16445 -715 16475
rect -685 16445 -680 16475
rect -720 16315 -680 16445
rect -560 18756 -520 18884
rect -560 18724 -556 18756
rect -524 18724 -520 18756
rect -560 18676 -520 18724
rect -560 18644 -556 18676
rect -524 18644 -520 18676
rect -560 18596 -520 18644
rect -560 18564 -556 18596
rect -524 18564 -520 18596
rect -560 18516 -520 18564
rect -560 18484 -556 18516
rect -524 18484 -520 18516
rect -560 18436 -520 18484
rect -560 18404 -556 18436
rect -524 18404 -520 18436
rect -560 18356 -520 18404
rect -560 18324 -556 18356
rect -524 18324 -520 18356
rect -560 18276 -520 18324
rect -560 18244 -556 18276
rect -524 18244 -520 18276
rect -560 18196 -520 18244
rect -560 18164 -556 18196
rect -524 18164 -520 18196
rect -560 18035 -520 18164
rect -560 18005 -555 18035
rect -525 18005 -520 18035
rect -560 17876 -520 18005
rect -560 17844 -556 17876
rect -524 17844 -520 17876
rect -560 17796 -520 17844
rect 20520 18035 20560 18040
rect 20520 18005 20525 18035
rect 20555 18005 20560 18035
rect 20520 17875 20560 18005
rect 20520 17845 20525 17875
rect 20555 17845 20560 17875
rect 20520 17840 20560 17845
rect 20600 18035 20640 18040
rect 20600 18005 20605 18035
rect 20635 18005 20640 18035
rect 20600 17875 20640 18005
rect 20600 17845 20605 17875
rect 20635 17845 20640 17875
rect 20600 17840 20640 17845
rect 20680 18035 20720 18040
rect 20680 18005 20685 18035
rect 20715 18005 20720 18035
rect 20680 17875 20720 18005
rect 20680 17845 20685 17875
rect 20715 17845 20720 17875
rect 20680 17840 20720 17845
rect 20760 18035 20800 18040
rect 20760 18005 20765 18035
rect 20795 18005 20800 18035
rect 20760 17875 20800 18005
rect 20760 17845 20765 17875
rect 20795 17845 20800 17875
rect 20760 17840 20800 17845
rect 20840 18035 20880 18040
rect 20840 18005 20845 18035
rect 20875 18005 20880 18035
rect 20840 17875 20880 18005
rect 20840 17845 20845 17875
rect 20875 17845 20880 17875
rect 20840 17840 20880 17845
rect 20920 18035 20960 18040
rect 20920 18005 20925 18035
rect 20955 18005 20960 18035
rect 20920 17875 20960 18005
rect 20920 17845 20925 17875
rect 20955 17845 20960 17875
rect 20920 17840 20960 17845
rect 21000 18035 21040 18040
rect 21000 18005 21005 18035
rect 21035 18005 21040 18035
rect 21000 17875 21040 18005
rect 21000 17845 21005 17875
rect 21035 17845 21040 17875
rect 21000 17840 21040 17845
rect 21080 18035 21120 18040
rect 21080 18005 21085 18035
rect 21115 18005 21120 18035
rect 21080 17875 21120 18005
rect 21080 17845 21085 17875
rect 21115 17845 21120 17875
rect 21080 17840 21120 17845
rect 21160 18035 21200 18040
rect 21160 18005 21165 18035
rect 21195 18005 21200 18035
rect 21160 17875 21200 18005
rect 21160 17845 21165 17875
rect 21195 17845 21200 17875
rect 21160 17840 21200 17845
rect 21240 18035 21280 18040
rect 21240 18005 21245 18035
rect 21275 18005 21280 18035
rect 21240 17875 21280 18005
rect 21240 17845 21245 17875
rect 21275 17845 21280 17875
rect 21240 17840 21280 17845
rect 21320 18035 21360 18040
rect 21320 18005 21325 18035
rect 21355 18005 21360 18035
rect 21320 17875 21360 18005
rect 21320 17845 21325 17875
rect 21355 17845 21360 17875
rect 21320 17840 21360 17845
rect 21400 18035 21440 18040
rect 21400 18005 21405 18035
rect 21435 18005 21440 18035
rect 21400 17875 21440 18005
rect 21400 17845 21405 17875
rect 21435 17845 21440 17875
rect 21400 17840 21440 17845
rect 21480 18035 21520 18040
rect 21480 18005 21485 18035
rect 21515 18005 21520 18035
rect 21480 17875 21520 18005
rect 21480 17845 21485 17875
rect 21515 17845 21520 17875
rect 21480 17840 21520 17845
rect 21560 18035 21600 18040
rect 21560 18005 21565 18035
rect 21595 18005 21600 18035
rect 21560 17875 21600 18005
rect 21560 17845 21565 17875
rect 21595 17845 21600 17875
rect 21560 17840 21600 17845
rect -560 17764 -556 17796
rect -524 17764 -520 17796
rect -560 17716 -520 17764
rect -560 17684 -556 17716
rect -524 17684 -520 17716
rect -560 17636 -520 17684
rect -560 17604 -556 17636
rect -524 17604 -520 17636
rect -560 17556 -520 17604
rect -560 17524 -556 17556
rect -524 17524 -520 17556
rect -560 17476 -520 17524
rect -560 17444 -556 17476
rect -524 17444 -520 17476
rect -560 17396 -520 17444
rect -560 17364 -556 17396
rect -524 17364 -520 17396
rect -560 17316 -520 17364
rect -560 17284 -556 17316
rect -524 17284 -520 17316
rect -560 17236 -520 17284
rect -560 17204 -556 17236
rect -524 17204 -520 17236
rect -560 17156 -520 17204
rect -560 17124 -556 17156
rect -524 17124 -520 17156
rect -560 17076 -520 17124
rect -560 17044 -556 17076
rect -524 17044 -520 17076
rect -560 16996 -520 17044
rect -560 16964 -556 16996
rect -524 16964 -520 16996
rect -560 16916 -520 16964
rect -560 16884 -556 16916
rect -524 16884 -520 16916
rect -560 16836 -520 16884
rect -560 16804 -556 16836
rect -524 16804 -520 16836
rect -560 16756 -520 16804
rect -560 16724 -556 16756
rect -524 16724 -520 16756
rect -560 16636 -520 16724
rect -560 16604 -556 16636
rect -524 16604 -520 16636
rect -560 16556 -520 16604
rect -560 16524 -556 16556
rect -524 16524 -520 16556
rect -560 16475 -520 16524
rect -560 16445 -555 16475
rect -525 16445 -520 16475
rect -720 16285 -715 16315
rect -685 16285 -680 16315
rect -720 16155 -680 16285
rect -720 16125 -715 16155
rect -685 16125 -680 16155
rect -720 15995 -680 16125
rect -720 15965 -715 15995
rect -685 15965 -680 15995
rect -720 15920 -680 15965
rect -640 16395 -600 16400
rect -640 16365 -635 16395
rect -605 16365 -600 16395
rect -640 15920 -600 16365
rect -560 16315 -520 16445
rect -560 16285 -555 16315
rect -525 16285 -520 16315
rect -560 16155 -520 16285
rect -560 16125 -555 16155
rect -525 16125 -520 16155
rect -560 15995 -520 16125
rect -560 15965 -555 15995
rect -525 15965 -520 15995
rect -560 15920 -520 15965
<< via3 >>
rect -15516 20875 -15484 20876
rect -15516 20845 -15515 20875
rect -15515 20845 -15485 20875
rect -15485 20845 -15484 20875
rect -15516 20844 -15484 20845
rect -15516 20795 -15484 20796
rect -15516 20765 -15515 20795
rect -15515 20765 -15485 20795
rect -15485 20765 -15484 20795
rect -15516 20764 -15484 20765
rect -15516 20395 -15484 20396
rect -15516 20365 -15515 20395
rect -15515 20365 -15485 20395
rect -15485 20365 -15484 20395
rect -15516 20364 -15484 20365
rect -15516 20315 -15484 20316
rect -15516 20285 -15515 20315
rect -15515 20285 -15485 20315
rect -15485 20285 -15484 20315
rect -15516 20284 -15484 20285
rect -15516 20235 -15484 20236
rect -15516 20205 -15515 20235
rect -15515 20205 -15485 20235
rect -15485 20205 -15484 20235
rect -15516 20204 -15484 20205
rect -15516 20155 -15484 20156
rect -15516 20125 -15515 20155
rect -15515 20125 -15485 20155
rect -15485 20125 -15484 20155
rect -15516 20124 -15484 20125
rect -15516 20075 -15484 20076
rect -15516 20045 -15515 20075
rect -15515 20045 -15485 20075
rect -15485 20045 -15484 20075
rect -15516 20044 -15484 20045
rect -15516 19995 -15484 19996
rect -15516 19965 -15515 19995
rect -15515 19965 -15485 19995
rect -15485 19965 -15484 19995
rect -15516 19964 -15484 19965
rect -15516 19915 -15484 19916
rect -15516 19885 -15515 19915
rect -15515 19885 -15485 19915
rect -15485 19885 -15484 19915
rect -15516 19884 -15484 19885
rect -15516 19835 -15484 19836
rect -15516 19805 -15515 19835
rect -15515 19805 -15485 19835
rect -15485 19805 -15484 19835
rect -15516 19804 -15484 19805
rect -15516 19755 -15484 19756
rect -15516 19725 -15515 19755
rect -15515 19725 -15485 19755
rect -15485 19725 -15484 19755
rect -15516 19724 -15484 19725
rect -15516 19675 -15484 19676
rect -15516 19645 -15515 19675
rect -15515 19645 -15485 19675
rect -15485 19645 -15484 19675
rect -15516 19644 -15484 19645
rect -15516 19595 -15484 19596
rect -15516 19565 -15515 19595
rect -15515 19565 -15485 19595
rect -15485 19565 -15484 19595
rect -15516 19564 -15484 19565
rect -15516 19515 -15484 19516
rect -15516 19485 -15515 19515
rect -15515 19485 -15485 19515
rect -15485 19485 -15484 19515
rect -15516 19484 -15484 19485
rect -15516 19435 -15484 19436
rect -15516 19405 -15515 19435
rect -15515 19405 -15485 19435
rect -15485 19405 -15484 19435
rect -15516 19404 -15484 19405
rect -15516 19355 -15484 19356
rect -15516 19325 -15515 19355
rect -15515 19325 -15485 19355
rect -15485 19325 -15484 19355
rect -15516 19324 -15484 19325
rect -15516 19275 -15484 19276
rect -15516 19245 -15515 19275
rect -15515 19245 -15485 19275
rect -15485 19245 -15484 19275
rect -15516 19244 -15484 19245
rect -15516 19195 -15484 19196
rect -15516 19165 -15515 19195
rect -15515 19165 -15485 19195
rect -15485 19165 -15484 19195
rect -15516 19164 -15484 19165
rect -15516 19115 -15484 19116
rect -15516 19085 -15515 19115
rect -15515 19085 -15485 19115
rect -15485 19085 -15484 19115
rect -15516 19084 -15484 19085
rect -15516 19035 -15484 19036
rect -15516 19005 -15515 19035
rect -15515 19005 -15485 19035
rect -15485 19005 -15484 19035
rect -15516 19004 -15484 19005
rect -15516 18955 -15484 18956
rect -15516 18925 -15515 18955
rect -15515 18925 -15485 18955
rect -15485 18925 -15484 18955
rect -15516 18924 -15484 18925
rect -15516 18875 -15484 18876
rect -15516 18845 -15515 18875
rect -15515 18845 -15485 18875
rect -15485 18845 -15484 18875
rect -15516 18844 -15484 18845
rect -15356 20875 -15324 20876
rect -15356 20845 -15355 20875
rect -15355 20845 -15325 20875
rect -15325 20845 -15324 20875
rect -15356 20844 -15324 20845
rect -15356 20795 -15324 20796
rect -15356 20765 -15355 20795
rect -15355 20765 -15325 20795
rect -15325 20765 -15324 20795
rect -15356 20764 -15324 20765
rect -15356 20395 -15324 20396
rect -15356 20365 -15355 20395
rect -15355 20365 -15325 20395
rect -15325 20365 -15324 20395
rect -15356 20364 -15324 20365
rect -15356 20315 -15324 20316
rect -15356 20285 -15355 20315
rect -15355 20285 -15325 20315
rect -15325 20285 -15324 20315
rect -15356 20284 -15324 20285
rect -15356 20235 -15324 20236
rect -15356 20205 -15355 20235
rect -15355 20205 -15325 20235
rect -15325 20205 -15324 20235
rect -15356 20204 -15324 20205
rect -15356 20155 -15324 20156
rect -15356 20125 -15355 20155
rect -15355 20125 -15325 20155
rect -15325 20125 -15324 20155
rect -15356 20124 -15324 20125
rect -15356 20075 -15324 20076
rect -15356 20045 -15355 20075
rect -15355 20045 -15325 20075
rect -15325 20045 -15324 20075
rect -15356 20044 -15324 20045
rect -15356 19995 -15324 19996
rect -15356 19965 -15355 19995
rect -15355 19965 -15325 19995
rect -15325 19965 -15324 19995
rect -15356 19964 -15324 19965
rect -15356 19915 -15324 19916
rect -15356 19885 -15355 19915
rect -15355 19885 -15325 19915
rect -15325 19885 -15324 19915
rect -15356 19884 -15324 19885
rect -15356 19835 -15324 19836
rect -15356 19805 -15355 19835
rect -15355 19805 -15325 19835
rect -15325 19805 -15324 19835
rect -15356 19804 -15324 19805
rect -15356 19755 -15324 19756
rect -15356 19725 -15355 19755
rect -15355 19725 -15325 19755
rect -15325 19725 -15324 19755
rect -15356 19724 -15324 19725
rect -15356 19675 -15324 19676
rect -15356 19645 -15355 19675
rect -15355 19645 -15325 19675
rect -15325 19645 -15324 19675
rect -15356 19644 -15324 19645
rect -15356 19595 -15324 19596
rect -15356 19565 -15355 19595
rect -15355 19565 -15325 19595
rect -15325 19565 -15324 19595
rect -15356 19564 -15324 19565
rect -15356 19515 -15324 19516
rect -15356 19485 -15355 19515
rect -15355 19485 -15325 19515
rect -15325 19485 -15324 19515
rect -15356 19484 -15324 19485
rect -15356 19435 -15324 19436
rect -15356 19405 -15355 19435
rect -15355 19405 -15325 19435
rect -15325 19405 -15324 19435
rect -15356 19404 -15324 19405
rect -15356 19355 -15324 19356
rect -15356 19325 -15355 19355
rect -15355 19325 -15325 19355
rect -15325 19325 -15324 19355
rect -15356 19324 -15324 19325
rect -15356 19275 -15324 19276
rect -15356 19245 -15355 19275
rect -15355 19245 -15325 19275
rect -15325 19245 -15324 19275
rect -15356 19244 -15324 19245
rect -15356 19195 -15324 19196
rect -15356 19165 -15355 19195
rect -15355 19165 -15325 19195
rect -15325 19165 -15324 19195
rect -15356 19164 -15324 19165
rect -15356 19115 -15324 19116
rect -15356 19085 -15355 19115
rect -15355 19085 -15325 19115
rect -15325 19085 -15324 19115
rect -15356 19084 -15324 19085
rect -15356 19035 -15324 19036
rect -15356 19005 -15355 19035
rect -15355 19005 -15325 19035
rect -15325 19005 -15324 19035
rect -15356 19004 -15324 19005
rect -15356 18955 -15324 18956
rect -15356 18925 -15355 18955
rect -15355 18925 -15325 18955
rect -15325 18925 -15324 18955
rect -15356 18924 -15324 18925
rect -15356 18875 -15324 18876
rect -15356 18845 -15355 18875
rect -15355 18845 -15325 18875
rect -15325 18845 -15324 18875
rect -15356 18844 -15324 18845
rect -15196 20875 -15164 20876
rect -15196 20845 -15195 20875
rect -15195 20845 -15165 20875
rect -15165 20845 -15164 20875
rect -15196 20844 -15164 20845
rect -15196 20795 -15164 20796
rect -15196 20765 -15195 20795
rect -15195 20765 -15165 20795
rect -15165 20765 -15164 20795
rect -15196 20764 -15164 20765
rect -15196 20395 -15164 20396
rect -15196 20365 -15195 20395
rect -15195 20365 -15165 20395
rect -15165 20365 -15164 20395
rect -15196 20364 -15164 20365
rect -15196 20315 -15164 20316
rect -15196 20285 -15195 20315
rect -15195 20285 -15165 20315
rect -15165 20285 -15164 20315
rect -15196 20284 -15164 20285
rect -15196 20235 -15164 20236
rect -15196 20205 -15195 20235
rect -15195 20205 -15165 20235
rect -15165 20205 -15164 20235
rect -15196 20204 -15164 20205
rect -15196 20155 -15164 20156
rect -15196 20125 -15195 20155
rect -15195 20125 -15165 20155
rect -15165 20125 -15164 20155
rect -15196 20124 -15164 20125
rect -15196 20075 -15164 20076
rect -15196 20045 -15195 20075
rect -15195 20045 -15165 20075
rect -15165 20045 -15164 20075
rect -15196 20044 -15164 20045
rect -15196 19995 -15164 19996
rect -15196 19965 -15195 19995
rect -15195 19965 -15165 19995
rect -15165 19965 -15164 19995
rect -15196 19964 -15164 19965
rect -15196 19915 -15164 19916
rect -15196 19885 -15195 19915
rect -15195 19885 -15165 19915
rect -15165 19885 -15164 19915
rect -15196 19884 -15164 19885
rect -15196 19835 -15164 19836
rect -15196 19805 -15195 19835
rect -15195 19805 -15165 19835
rect -15165 19805 -15164 19835
rect -15196 19804 -15164 19805
rect -15196 19755 -15164 19756
rect -15196 19725 -15195 19755
rect -15195 19725 -15165 19755
rect -15165 19725 -15164 19755
rect -15196 19724 -15164 19725
rect -15196 19675 -15164 19676
rect -15196 19645 -15195 19675
rect -15195 19645 -15165 19675
rect -15165 19645 -15164 19675
rect -15196 19644 -15164 19645
rect -15196 19595 -15164 19596
rect -15196 19565 -15195 19595
rect -15195 19565 -15165 19595
rect -15165 19565 -15164 19595
rect -15196 19564 -15164 19565
rect -15196 19515 -15164 19516
rect -15196 19485 -15195 19515
rect -15195 19485 -15165 19515
rect -15165 19485 -15164 19515
rect -15196 19484 -15164 19485
rect -15196 19435 -15164 19436
rect -15196 19405 -15195 19435
rect -15195 19405 -15165 19435
rect -15165 19405 -15164 19435
rect -15196 19404 -15164 19405
rect -15196 19355 -15164 19356
rect -15196 19325 -15195 19355
rect -15195 19325 -15165 19355
rect -15165 19325 -15164 19355
rect -15196 19324 -15164 19325
rect -15196 19275 -15164 19276
rect -15196 19245 -15195 19275
rect -15195 19245 -15165 19275
rect -15165 19245 -15164 19275
rect -15196 19244 -15164 19245
rect -15196 19195 -15164 19196
rect -15196 19165 -15195 19195
rect -15195 19165 -15165 19195
rect -15165 19165 -15164 19195
rect -15196 19164 -15164 19165
rect -15196 19115 -15164 19116
rect -15196 19085 -15195 19115
rect -15195 19085 -15165 19115
rect -15165 19085 -15164 19115
rect -15196 19084 -15164 19085
rect -15196 19035 -15164 19036
rect -15196 19005 -15195 19035
rect -15195 19005 -15165 19035
rect -15165 19005 -15164 19035
rect -15196 19004 -15164 19005
rect -15196 18955 -15164 18956
rect -15196 18925 -15195 18955
rect -15195 18925 -15165 18955
rect -15165 18925 -15164 18955
rect -15196 18924 -15164 18925
rect -15196 18875 -15164 18876
rect -15196 18845 -15195 18875
rect -15195 18845 -15165 18875
rect -15165 18845 -15164 18875
rect -15196 18844 -15164 18845
rect -15516 18555 -15484 18556
rect -15516 18525 -15515 18555
rect -15515 18525 -15485 18555
rect -15485 18525 -15484 18555
rect -15516 18524 -15484 18525
rect -15516 18475 -15484 18476
rect -15516 18445 -15515 18475
rect -15515 18445 -15485 18475
rect -15485 18445 -15484 18475
rect -15516 18444 -15484 18445
rect -15516 18395 -15484 18396
rect -15516 18365 -15515 18395
rect -15515 18365 -15485 18395
rect -15485 18365 -15484 18395
rect -15516 18364 -15484 18365
rect -15516 18315 -15484 18316
rect -15516 18285 -15515 18315
rect -15515 18285 -15485 18315
rect -15485 18285 -15484 18315
rect -15516 18284 -15484 18285
rect -15516 18235 -15484 18236
rect -15516 18205 -15515 18235
rect -15515 18205 -15485 18235
rect -15485 18205 -15484 18235
rect -15516 18204 -15484 18205
rect -15516 18155 -15484 18156
rect -15516 18125 -15515 18155
rect -15515 18125 -15485 18155
rect -15485 18125 -15484 18155
rect -15516 18124 -15484 18125
rect -15516 18075 -15484 18076
rect -15516 18045 -15515 18075
rect -15515 18045 -15485 18075
rect -15485 18045 -15484 18075
rect -15516 18044 -15484 18045
rect -15516 17995 -15484 17996
rect -15516 17965 -15515 17995
rect -15515 17965 -15485 17995
rect -15485 17965 -15484 17995
rect -15516 17964 -15484 17965
rect -15516 17915 -15484 17916
rect -15516 17885 -15515 17915
rect -15515 17885 -15485 17915
rect -15485 17885 -15484 17915
rect -15516 17884 -15484 17885
rect -15516 17835 -15484 17836
rect -15516 17805 -15515 17835
rect -15515 17805 -15485 17835
rect -15485 17805 -15484 17835
rect -15516 17804 -15484 17805
rect -15516 17755 -15484 17756
rect -15516 17725 -15515 17755
rect -15515 17725 -15485 17755
rect -15485 17725 -15484 17755
rect -15516 17724 -15484 17725
rect -15516 17675 -15484 17676
rect -15516 17645 -15515 17675
rect -15515 17645 -15485 17675
rect -15485 17645 -15484 17675
rect -15516 17644 -15484 17645
rect -15516 17595 -15484 17596
rect -15516 17565 -15515 17595
rect -15515 17565 -15485 17595
rect -15485 17565 -15484 17595
rect -15516 17564 -15484 17565
rect -15516 17515 -15484 17516
rect -15516 17485 -15515 17515
rect -15515 17485 -15485 17515
rect -15485 17485 -15484 17515
rect -15516 17484 -15484 17485
rect -15516 17435 -15484 17436
rect -15516 17405 -15515 17435
rect -15515 17405 -15485 17435
rect -15485 17405 -15484 17435
rect -15516 17404 -15484 17405
rect -15516 17115 -15484 17116
rect -15516 17085 -15515 17115
rect -15515 17085 -15485 17115
rect -15485 17085 -15484 17115
rect -15516 17084 -15484 17085
rect -15516 17035 -15484 17036
rect -15516 17005 -15515 17035
rect -15515 17005 -15485 17035
rect -15485 17005 -15484 17035
rect -15516 17004 -15484 17005
rect -15516 16955 -15484 16956
rect -15516 16925 -15515 16955
rect -15515 16925 -15485 16955
rect -15485 16925 -15484 16955
rect -15516 16924 -15484 16925
rect -15516 16875 -15484 16876
rect -15516 16845 -15515 16875
rect -15515 16845 -15485 16875
rect -15485 16845 -15484 16875
rect -15516 16844 -15484 16845
rect -15516 16795 -15484 16796
rect -15516 16765 -15515 16795
rect -15515 16765 -15485 16795
rect -15485 16765 -15484 16795
rect -15516 16764 -15484 16765
rect -15516 16715 -15484 16716
rect -15516 16685 -15515 16715
rect -15515 16685 -15485 16715
rect -15485 16685 -15484 16715
rect -15516 16684 -15484 16685
rect -15516 16635 -15484 16636
rect -15516 16605 -15515 16635
rect -15515 16605 -15485 16635
rect -15485 16605 -15484 16635
rect -15516 16604 -15484 16605
rect -15516 16555 -15484 16556
rect -15516 16525 -15515 16555
rect -15515 16525 -15485 16555
rect -15485 16525 -15484 16555
rect -15516 16524 -15484 16525
rect -15516 16475 -15484 16476
rect -15516 16445 -15515 16475
rect -15515 16445 -15485 16475
rect -15485 16445 -15484 16475
rect -15516 16444 -15484 16445
rect -15356 18555 -15324 18556
rect -15356 18525 -15355 18555
rect -15355 18525 -15325 18555
rect -15325 18525 -15324 18555
rect -15356 18524 -15324 18525
rect -15356 18475 -15324 18476
rect -15356 18445 -15355 18475
rect -15355 18445 -15325 18475
rect -15325 18445 -15324 18475
rect -15356 18444 -15324 18445
rect -15356 18395 -15324 18396
rect -15356 18365 -15355 18395
rect -15355 18365 -15325 18395
rect -15325 18365 -15324 18395
rect -15356 18364 -15324 18365
rect -15356 18315 -15324 18316
rect -15356 18285 -15355 18315
rect -15355 18285 -15325 18315
rect -15325 18285 -15324 18315
rect -15356 18284 -15324 18285
rect -15356 18235 -15324 18236
rect -15356 18205 -15355 18235
rect -15355 18205 -15325 18235
rect -15325 18205 -15324 18235
rect -15356 18204 -15324 18205
rect -15356 18155 -15324 18156
rect -15356 18125 -15355 18155
rect -15355 18125 -15325 18155
rect -15325 18125 -15324 18155
rect -15356 18124 -15324 18125
rect -15356 18075 -15324 18076
rect -15356 18045 -15355 18075
rect -15355 18045 -15325 18075
rect -15325 18045 -15324 18075
rect -15356 18044 -15324 18045
rect -15356 17995 -15324 17996
rect -15356 17965 -15355 17995
rect -15355 17965 -15325 17995
rect -15325 17965 -15324 17995
rect -15356 17964 -15324 17965
rect -15356 17915 -15324 17916
rect -15356 17885 -15355 17915
rect -15355 17885 -15325 17915
rect -15325 17885 -15324 17915
rect -15356 17884 -15324 17885
rect -15356 17835 -15324 17836
rect -15356 17805 -15355 17835
rect -15355 17805 -15325 17835
rect -15325 17805 -15324 17835
rect -15356 17804 -15324 17805
rect -15356 17755 -15324 17756
rect -15356 17725 -15355 17755
rect -15355 17725 -15325 17755
rect -15325 17725 -15324 17755
rect -15356 17724 -15324 17725
rect -15356 17675 -15324 17676
rect -15356 17645 -15355 17675
rect -15355 17645 -15325 17675
rect -15325 17645 -15324 17675
rect -15356 17644 -15324 17645
rect -15356 17595 -15324 17596
rect -15356 17565 -15355 17595
rect -15355 17565 -15325 17595
rect -15325 17565 -15324 17595
rect -15356 17564 -15324 17565
rect -15356 17515 -15324 17516
rect -15356 17485 -15355 17515
rect -15355 17485 -15325 17515
rect -15325 17485 -15324 17515
rect -15356 17484 -15324 17485
rect -15356 17435 -15324 17436
rect -15356 17405 -15355 17435
rect -15355 17405 -15325 17435
rect -15325 17405 -15324 17435
rect -15356 17404 -15324 17405
rect -15356 17115 -15324 17116
rect -15356 17085 -15355 17115
rect -15355 17085 -15325 17115
rect -15325 17085 -15324 17115
rect -15356 17084 -15324 17085
rect -15356 17035 -15324 17036
rect -15356 17005 -15355 17035
rect -15355 17005 -15325 17035
rect -15325 17005 -15324 17035
rect -15356 17004 -15324 17005
rect -15356 16955 -15324 16956
rect -15356 16925 -15355 16955
rect -15355 16925 -15325 16955
rect -15325 16925 -15324 16955
rect -15356 16924 -15324 16925
rect -15356 16875 -15324 16876
rect -15356 16845 -15355 16875
rect -15355 16845 -15325 16875
rect -15325 16845 -15324 16875
rect -15356 16844 -15324 16845
rect -15356 16795 -15324 16796
rect -15356 16765 -15355 16795
rect -15355 16765 -15325 16795
rect -15325 16765 -15324 16795
rect -15356 16764 -15324 16765
rect -15356 16715 -15324 16716
rect -15356 16685 -15355 16715
rect -15355 16685 -15325 16715
rect -15325 16685 -15324 16715
rect -15356 16684 -15324 16685
rect -15356 16635 -15324 16636
rect -15356 16605 -15355 16635
rect -15355 16605 -15325 16635
rect -15325 16605 -15324 16635
rect -15356 16604 -15324 16605
rect -15356 16555 -15324 16556
rect -15356 16525 -15355 16555
rect -15355 16525 -15325 16555
rect -15325 16525 -15324 16555
rect -15356 16524 -15324 16525
rect -15356 16475 -15324 16476
rect -15356 16445 -15355 16475
rect -15355 16445 -15325 16475
rect -15325 16445 -15324 16475
rect -15356 16444 -15324 16445
rect -15036 20875 -15004 20876
rect -15036 20845 -15035 20875
rect -15035 20845 -15005 20875
rect -15005 20845 -15004 20875
rect -15036 20844 -15004 20845
rect -15036 20795 -15004 20796
rect -15036 20765 -15035 20795
rect -15035 20765 -15005 20795
rect -15005 20765 -15004 20795
rect -15036 20764 -15004 20765
rect -15036 20395 -15004 20396
rect -15036 20365 -15035 20395
rect -15035 20365 -15005 20395
rect -15005 20365 -15004 20395
rect -15036 20364 -15004 20365
rect -15036 20315 -15004 20316
rect -15036 20285 -15035 20315
rect -15035 20285 -15005 20315
rect -15005 20285 -15004 20315
rect -15036 20284 -15004 20285
rect -15036 20235 -15004 20236
rect -15036 20205 -15035 20235
rect -15035 20205 -15005 20235
rect -15005 20205 -15004 20235
rect -15036 20204 -15004 20205
rect -15036 20155 -15004 20156
rect -15036 20125 -15035 20155
rect -15035 20125 -15005 20155
rect -15005 20125 -15004 20155
rect -15036 20124 -15004 20125
rect -15036 20075 -15004 20076
rect -15036 20045 -15035 20075
rect -15035 20045 -15005 20075
rect -15005 20045 -15004 20075
rect -15036 20044 -15004 20045
rect -15036 19995 -15004 19996
rect -15036 19965 -15035 19995
rect -15035 19965 -15005 19995
rect -15005 19965 -15004 19995
rect -15036 19964 -15004 19965
rect -15036 19915 -15004 19916
rect -15036 19885 -15035 19915
rect -15035 19885 -15005 19915
rect -15005 19885 -15004 19915
rect -15036 19884 -15004 19885
rect -15036 19835 -15004 19836
rect -15036 19805 -15035 19835
rect -15035 19805 -15005 19835
rect -15005 19805 -15004 19835
rect -15036 19804 -15004 19805
rect -15036 19755 -15004 19756
rect -15036 19725 -15035 19755
rect -15035 19725 -15005 19755
rect -15005 19725 -15004 19755
rect -15036 19724 -15004 19725
rect -15036 19675 -15004 19676
rect -15036 19645 -15035 19675
rect -15035 19645 -15005 19675
rect -15005 19645 -15004 19675
rect -15036 19644 -15004 19645
rect -15036 19595 -15004 19596
rect -15036 19565 -15035 19595
rect -15035 19565 -15005 19595
rect -15005 19565 -15004 19595
rect -15036 19564 -15004 19565
rect -15036 19515 -15004 19516
rect -15036 19485 -15035 19515
rect -15035 19485 -15005 19515
rect -15005 19485 -15004 19515
rect -15036 19484 -15004 19485
rect -15036 19435 -15004 19436
rect -15036 19405 -15035 19435
rect -15035 19405 -15005 19435
rect -15005 19405 -15004 19435
rect -15036 19404 -15004 19405
rect -15036 19355 -15004 19356
rect -15036 19325 -15035 19355
rect -15035 19325 -15005 19355
rect -15005 19325 -15004 19355
rect -15036 19324 -15004 19325
rect -15036 19275 -15004 19276
rect -15036 19245 -15035 19275
rect -15035 19245 -15005 19275
rect -15005 19245 -15004 19275
rect -15036 19244 -15004 19245
rect -15036 19195 -15004 19196
rect -15036 19165 -15035 19195
rect -15035 19165 -15005 19195
rect -15005 19165 -15004 19195
rect -15036 19164 -15004 19165
rect -15036 19115 -15004 19116
rect -15036 19085 -15035 19115
rect -15035 19085 -15005 19115
rect -15005 19085 -15004 19115
rect -15036 19084 -15004 19085
rect -15036 19035 -15004 19036
rect -15036 19005 -15035 19035
rect -15035 19005 -15005 19035
rect -15005 19005 -15004 19035
rect -15036 19004 -15004 19005
rect -15036 18955 -15004 18956
rect -15036 18925 -15035 18955
rect -15035 18925 -15005 18955
rect -15005 18925 -15004 18955
rect -15036 18924 -15004 18925
rect -15036 18875 -15004 18876
rect -15036 18845 -15035 18875
rect -15035 18845 -15005 18875
rect -15005 18845 -15004 18875
rect -15036 18844 -15004 18845
rect -15196 18555 -15164 18556
rect -15196 18525 -15195 18555
rect -15195 18525 -15165 18555
rect -15165 18525 -15164 18555
rect -15196 18524 -15164 18525
rect -15196 18475 -15164 18476
rect -15196 18445 -15195 18475
rect -15195 18445 -15165 18475
rect -15165 18445 -15164 18475
rect -15196 18444 -15164 18445
rect -15196 18395 -15164 18396
rect -15196 18365 -15195 18395
rect -15195 18365 -15165 18395
rect -15165 18365 -15164 18395
rect -15196 18364 -15164 18365
rect -15196 18315 -15164 18316
rect -15196 18285 -15195 18315
rect -15195 18285 -15165 18315
rect -15165 18285 -15164 18315
rect -15196 18284 -15164 18285
rect -15196 18235 -15164 18236
rect -15196 18205 -15195 18235
rect -15195 18205 -15165 18235
rect -15165 18205 -15164 18235
rect -15196 18204 -15164 18205
rect -15196 18155 -15164 18156
rect -15196 18125 -15195 18155
rect -15195 18125 -15165 18155
rect -15165 18125 -15164 18155
rect -15196 18124 -15164 18125
rect -15196 18075 -15164 18076
rect -15196 18045 -15195 18075
rect -15195 18045 -15165 18075
rect -15165 18045 -15164 18075
rect -15196 18044 -15164 18045
rect -15196 17995 -15164 17996
rect -15196 17965 -15195 17995
rect -15195 17965 -15165 17995
rect -15165 17965 -15164 17995
rect -15196 17964 -15164 17965
rect -15196 17915 -15164 17916
rect -15196 17885 -15195 17915
rect -15195 17885 -15165 17915
rect -15165 17885 -15164 17915
rect -15196 17884 -15164 17885
rect -15036 18555 -15004 18556
rect -15036 18525 -15035 18555
rect -15035 18525 -15005 18555
rect -15005 18525 -15004 18555
rect -15036 18524 -15004 18525
rect -15036 18475 -15004 18476
rect -15036 18445 -15035 18475
rect -15035 18445 -15005 18475
rect -15005 18445 -15004 18475
rect -15036 18444 -15004 18445
rect -15036 18395 -15004 18396
rect -15036 18365 -15035 18395
rect -15035 18365 -15005 18395
rect -15005 18365 -15004 18395
rect -15036 18364 -15004 18365
rect -15036 18315 -15004 18316
rect -15036 18285 -15035 18315
rect -15035 18285 -15005 18315
rect -15005 18285 -15004 18315
rect -15036 18284 -15004 18285
rect -15036 18235 -15004 18236
rect -15036 18205 -15035 18235
rect -15035 18205 -15005 18235
rect -15005 18205 -15004 18235
rect -15036 18204 -15004 18205
rect -15036 18155 -15004 18156
rect -15036 18125 -15035 18155
rect -15035 18125 -15005 18155
rect -15005 18125 -15004 18155
rect -15036 18124 -15004 18125
rect -15036 18075 -15004 18076
rect -15036 18045 -15035 18075
rect -15035 18045 -15005 18075
rect -15005 18045 -15004 18075
rect -15036 18044 -15004 18045
rect -15036 17995 -15004 17996
rect -15036 17965 -15035 17995
rect -15035 17965 -15005 17995
rect -15005 17965 -15004 17995
rect -15036 17964 -15004 17965
rect -15036 17915 -15004 17916
rect -15036 17885 -15035 17915
rect -15035 17885 -15005 17915
rect -15005 17885 -15004 17915
rect -15036 17884 -15004 17885
rect -15196 17835 -15164 17836
rect -15196 17805 -15195 17835
rect -15195 17805 -15165 17835
rect -15165 17805 -15164 17835
rect -15196 17804 -15164 17805
rect -15196 17755 -15164 17756
rect -15196 17725 -15195 17755
rect -15195 17725 -15165 17755
rect -15165 17725 -15164 17755
rect -15196 17724 -15164 17725
rect -15196 17675 -15164 17676
rect -15196 17645 -15195 17675
rect -15195 17645 -15165 17675
rect -15165 17645 -15164 17675
rect -15196 17644 -15164 17645
rect -15196 17595 -15164 17596
rect -15196 17565 -15195 17595
rect -15195 17565 -15165 17595
rect -15165 17565 -15164 17595
rect -15196 17564 -15164 17565
rect -15196 17515 -15164 17516
rect -15196 17485 -15195 17515
rect -15195 17485 -15165 17515
rect -15165 17485 -15164 17515
rect -15196 17484 -15164 17485
rect -15196 17435 -15164 17436
rect -15196 17405 -15195 17435
rect -15195 17405 -15165 17435
rect -15165 17405 -15164 17435
rect -15196 17404 -15164 17405
rect -15036 17835 -15004 17836
rect -15036 17805 -15035 17835
rect -15035 17805 -15005 17835
rect -15005 17805 -15004 17835
rect -15036 17804 -15004 17805
rect -15036 17755 -15004 17756
rect -15036 17725 -15035 17755
rect -15035 17725 -15005 17755
rect -15005 17725 -15004 17755
rect -15036 17724 -15004 17725
rect -15036 17675 -15004 17676
rect -15036 17645 -15035 17675
rect -15035 17645 -15005 17675
rect -15005 17645 -15004 17675
rect -15036 17644 -15004 17645
rect -15036 17595 -15004 17596
rect -15036 17565 -15035 17595
rect -15035 17565 -15005 17595
rect -15005 17565 -15004 17595
rect -15036 17564 -15004 17565
rect -15036 17515 -15004 17516
rect -15036 17485 -15035 17515
rect -15035 17485 -15005 17515
rect -15005 17485 -15004 17515
rect -15036 17484 -15004 17485
rect -1676 19875 -1644 19876
rect -1676 19845 -1675 19875
rect -1675 19845 -1645 19875
rect -1645 19845 -1644 19875
rect -1676 19844 -1644 19845
rect -1676 19795 -1644 19796
rect -1676 19765 -1675 19795
rect -1675 19765 -1645 19795
rect -1645 19765 -1644 19795
rect -1676 19764 -1644 19765
rect -1676 19715 -1644 19716
rect -1676 19685 -1675 19715
rect -1675 19685 -1645 19715
rect -1645 19685 -1644 19715
rect -1676 19684 -1644 19685
rect -1676 19635 -1644 19636
rect -1676 19605 -1675 19635
rect -1675 19605 -1645 19635
rect -1645 19605 -1644 19635
rect -1676 19604 -1644 19605
rect -1676 19555 -1644 19556
rect -1676 19525 -1675 19555
rect -1675 19525 -1645 19555
rect -1645 19525 -1644 19555
rect -1676 19524 -1644 19525
rect -1676 19475 -1644 19476
rect -1676 19445 -1675 19475
rect -1675 19445 -1645 19475
rect -1645 19445 -1644 19475
rect -1676 19444 -1644 19445
rect -1676 19395 -1644 19396
rect -1676 19365 -1675 19395
rect -1675 19365 -1645 19395
rect -1645 19365 -1644 19395
rect -1676 19364 -1644 19365
rect -1676 19315 -1644 19316
rect -1676 19285 -1675 19315
rect -1675 19285 -1645 19315
rect -1645 19285 -1644 19315
rect -1676 19284 -1644 19285
rect -1676 19235 -1644 19236
rect -1676 19205 -1675 19235
rect -1675 19205 -1645 19235
rect -1645 19205 -1644 19235
rect -1676 19204 -1644 19205
rect -1676 19155 -1644 19156
rect -1676 19125 -1675 19155
rect -1675 19125 -1645 19155
rect -1645 19125 -1644 19155
rect -1676 19124 -1644 19125
rect -1676 19075 -1644 19076
rect -1676 19045 -1675 19075
rect -1675 19045 -1645 19075
rect -1645 19045 -1644 19075
rect -1676 19044 -1644 19045
rect -1676 18995 -1644 18996
rect -1676 18965 -1675 18995
rect -1675 18965 -1645 18995
rect -1645 18965 -1644 18995
rect -1676 18964 -1644 18965
rect -1676 18915 -1644 18916
rect -1676 18885 -1675 18915
rect -1675 18885 -1645 18915
rect -1645 18885 -1644 18915
rect -1676 18884 -1644 18885
rect -1676 18755 -1644 18756
rect -1676 18725 -1675 18755
rect -1675 18725 -1645 18755
rect -1645 18725 -1644 18755
rect -1676 18724 -1644 18725
rect -1676 18675 -1644 18676
rect -1676 18645 -1675 18675
rect -1675 18645 -1645 18675
rect -1645 18645 -1644 18675
rect -1676 18644 -1644 18645
rect -1676 18595 -1644 18596
rect -1676 18565 -1675 18595
rect -1675 18565 -1645 18595
rect -1645 18565 -1644 18595
rect -1676 18564 -1644 18565
rect -1676 18515 -1644 18516
rect -1676 18485 -1675 18515
rect -1675 18485 -1645 18515
rect -1645 18485 -1644 18515
rect -1676 18484 -1644 18485
rect -1676 18435 -1644 18436
rect -1676 18405 -1675 18435
rect -1675 18405 -1645 18435
rect -1645 18405 -1644 18435
rect -1676 18404 -1644 18405
rect -1676 18355 -1644 18356
rect -1676 18325 -1675 18355
rect -1675 18325 -1645 18355
rect -1645 18325 -1644 18355
rect -1676 18324 -1644 18325
rect -1676 18275 -1644 18276
rect -1676 18245 -1675 18275
rect -1675 18245 -1645 18275
rect -1645 18245 -1644 18275
rect -1676 18244 -1644 18245
rect -1676 18195 -1644 18196
rect -1676 18165 -1675 18195
rect -1675 18165 -1645 18195
rect -1645 18165 -1644 18195
rect -1676 18164 -1644 18165
rect -1516 19875 -1484 19876
rect -1516 19845 -1515 19875
rect -1515 19845 -1485 19875
rect -1485 19845 -1484 19875
rect -1516 19844 -1484 19845
rect -1516 19795 -1484 19796
rect -1516 19765 -1515 19795
rect -1515 19765 -1485 19795
rect -1485 19765 -1484 19795
rect -1516 19764 -1484 19765
rect -1516 19715 -1484 19716
rect -1516 19685 -1515 19715
rect -1515 19685 -1485 19715
rect -1485 19685 -1484 19715
rect -1516 19684 -1484 19685
rect -1516 19635 -1484 19636
rect -1516 19605 -1515 19635
rect -1515 19605 -1485 19635
rect -1485 19605 -1484 19635
rect -1516 19604 -1484 19605
rect -1516 19555 -1484 19556
rect -1516 19525 -1515 19555
rect -1515 19525 -1485 19555
rect -1485 19525 -1484 19555
rect -1516 19524 -1484 19525
rect -1516 19475 -1484 19476
rect -1516 19445 -1515 19475
rect -1515 19445 -1485 19475
rect -1485 19445 -1484 19475
rect -1516 19444 -1484 19445
rect -1516 19395 -1484 19396
rect -1516 19365 -1515 19395
rect -1515 19365 -1485 19395
rect -1485 19365 -1484 19395
rect -1516 19364 -1484 19365
rect -1516 19315 -1484 19316
rect -1516 19285 -1515 19315
rect -1515 19285 -1485 19315
rect -1485 19285 -1484 19315
rect -1516 19284 -1484 19285
rect -1516 19235 -1484 19236
rect -1516 19205 -1515 19235
rect -1515 19205 -1485 19235
rect -1485 19205 -1484 19235
rect -1516 19204 -1484 19205
rect -1516 19155 -1484 19156
rect -1516 19125 -1515 19155
rect -1515 19125 -1485 19155
rect -1485 19125 -1484 19155
rect -1516 19124 -1484 19125
rect -1516 19075 -1484 19076
rect -1516 19045 -1515 19075
rect -1515 19045 -1485 19075
rect -1485 19045 -1484 19075
rect -1516 19044 -1484 19045
rect -1516 18995 -1484 18996
rect -1516 18965 -1515 18995
rect -1515 18965 -1485 18995
rect -1485 18965 -1484 18995
rect -1516 18964 -1484 18965
rect -1516 18915 -1484 18916
rect -1516 18885 -1515 18915
rect -1515 18885 -1485 18915
rect -1485 18885 -1484 18915
rect -1516 18884 -1484 18885
rect -1516 18755 -1484 18756
rect -1516 18725 -1515 18755
rect -1515 18725 -1485 18755
rect -1485 18725 -1484 18755
rect -1516 18724 -1484 18725
rect -1516 18675 -1484 18676
rect -1516 18645 -1515 18675
rect -1515 18645 -1485 18675
rect -1485 18645 -1484 18675
rect -1516 18644 -1484 18645
rect -1516 18595 -1484 18596
rect -1516 18565 -1515 18595
rect -1515 18565 -1485 18595
rect -1485 18565 -1484 18595
rect -1516 18564 -1484 18565
rect -1516 18515 -1484 18516
rect -1516 18485 -1515 18515
rect -1515 18485 -1485 18515
rect -1485 18485 -1484 18515
rect -1516 18484 -1484 18485
rect -1516 18435 -1484 18436
rect -1516 18405 -1515 18435
rect -1515 18405 -1485 18435
rect -1485 18405 -1484 18435
rect -1516 18404 -1484 18405
rect -1516 18355 -1484 18356
rect -1516 18325 -1515 18355
rect -1515 18325 -1485 18355
rect -1485 18325 -1484 18355
rect -1516 18324 -1484 18325
rect -1516 18275 -1484 18276
rect -1516 18245 -1515 18275
rect -1515 18245 -1485 18275
rect -1485 18245 -1484 18275
rect -1516 18244 -1484 18245
rect -1516 18195 -1484 18196
rect -1516 18165 -1515 18195
rect -1515 18165 -1485 18195
rect -1485 18165 -1484 18195
rect -1516 18164 -1484 18165
rect -1356 19875 -1324 19876
rect -1356 19845 -1355 19875
rect -1355 19845 -1325 19875
rect -1325 19845 -1324 19875
rect -1356 19844 -1324 19845
rect -1356 19795 -1324 19796
rect -1356 19765 -1355 19795
rect -1355 19765 -1325 19795
rect -1325 19765 -1324 19795
rect -1356 19764 -1324 19765
rect -1356 19715 -1324 19716
rect -1356 19685 -1355 19715
rect -1355 19685 -1325 19715
rect -1325 19685 -1324 19715
rect -1356 19684 -1324 19685
rect -1356 19635 -1324 19636
rect -1356 19605 -1355 19635
rect -1355 19605 -1325 19635
rect -1325 19605 -1324 19635
rect -1356 19604 -1324 19605
rect -1356 19555 -1324 19556
rect -1356 19525 -1355 19555
rect -1355 19525 -1325 19555
rect -1325 19525 -1324 19555
rect -1356 19524 -1324 19525
rect -1356 19475 -1324 19476
rect -1356 19445 -1355 19475
rect -1355 19445 -1325 19475
rect -1325 19445 -1324 19475
rect -1356 19444 -1324 19445
rect -1356 19395 -1324 19396
rect -1356 19365 -1355 19395
rect -1355 19365 -1325 19395
rect -1325 19365 -1324 19395
rect -1356 19364 -1324 19365
rect -1356 19315 -1324 19316
rect -1356 19285 -1355 19315
rect -1355 19285 -1325 19315
rect -1325 19285 -1324 19315
rect -1356 19284 -1324 19285
rect -1356 19235 -1324 19236
rect -1356 19205 -1355 19235
rect -1355 19205 -1325 19235
rect -1325 19205 -1324 19235
rect -1356 19204 -1324 19205
rect -1356 19155 -1324 19156
rect -1356 19125 -1355 19155
rect -1355 19125 -1325 19155
rect -1325 19125 -1324 19155
rect -1356 19124 -1324 19125
rect -1356 19075 -1324 19076
rect -1356 19045 -1355 19075
rect -1355 19045 -1325 19075
rect -1325 19045 -1324 19075
rect -1356 19044 -1324 19045
rect -1356 18995 -1324 18996
rect -1356 18965 -1355 18995
rect -1355 18965 -1325 18995
rect -1325 18965 -1324 18995
rect -1356 18964 -1324 18965
rect -1356 18915 -1324 18916
rect -1356 18885 -1355 18915
rect -1355 18885 -1325 18915
rect -1325 18885 -1324 18915
rect -1356 18884 -1324 18885
rect -1356 18755 -1324 18756
rect -1356 18725 -1355 18755
rect -1355 18725 -1325 18755
rect -1325 18725 -1324 18755
rect -1356 18724 -1324 18725
rect -1356 18675 -1324 18676
rect -1356 18645 -1355 18675
rect -1355 18645 -1325 18675
rect -1325 18645 -1324 18675
rect -1356 18644 -1324 18645
rect -1356 18595 -1324 18596
rect -1356 18565 -1355 18595
rect -1355 18565 -1325 18595
rect -1325 18565 -1324 18595
rect -1356 18564 -1324 18565
rect -1356 18515 -1324 18516
rect -1356 18485 -1355 18515
rect -1355 18485 -1325 18515
rect -1325 18485 -1324 18515
rect -1356 18484 -1324 18485
rect -1356 18435 -1324 18436
rect -1356 18405 -1355 18435
rect -1355 18405 -1325 18435
rect -1325 18405 -1324 18435
rect -1356 18404 -1324 18405
rect -1356 18355 -1324 18356
rect -1356 18325 -1355 18355
rect -1355 18325 -1325 18355
rect -1325 18325 -1324 18355
rect -1356 18324 -1324 18325
rect -1356 18275 -1324 18276
rect -1356 18245 -1355 18275
rect -1355 18245 -1325 18275
rect -1325 18245 -1324 18275
rect -1356 18244 -1324 18245
rect -1356 18195 -1324 18196
rect -1356 18165 -1355 18195
rect -1355 18165 -1325 18195
rect -1325 18165 -1324 18195
rect -1356 18164 -1324 18165
rect -1676 17875 -1644 17876
rect -1676 17845 -1675 17875
rect -1675 17845 -1645 17875
rect -1645 17845 -1644 17875
rect -1676 17844 -1644 17845
rect -1676 17795 -1644 17796
rect -1676 17765 -1675 17795
rect -1675 17765 -1645 17795
rect -1645 17765 -1644 17795
rect -1676 17764 -1644 17765
rect -1676 17715 -1644 17716
rect -1676 17685 -1675 17715
rect -1675 17685 -1645 17715
rect -1645 17685 -1644 17715
rect -1676 17684 -1644 17685
rect -1676 17635 -1644 17636
rect -1676 17605 -1675 17635
rect -1675 17605 -1645 17635
rect -1645 17605 -1644 17635
rect -1676 17604 -1644 17605
rect -1676 17555 -1644 17556
rect -1676 17525 -1675 17555
rect -1675 17525 -1645 17555
rect -1645 17525 -1644 17555
rect -1676 17524 -1644 17525
rect -1676 17475 -1644 17476
rect -1676 17445 -1675 17475
rect -1675 17445 -1645 17475
rect -1645 17445 -1644 17475
rect -1676 17444 -1644 17445
rect -15036 17435 -15004 17436
rect -15036 17405 -15035 17435
rect -15035 17405 -15005 17435
rect -15005 17405 -15004 17435
rect -15036 17404 -15004 17405
rect -15196 17115 -15164 17116
rect -15196 17085 -15195 17115
rect -15195 17085 -15165 17115
rect -15165 17085 -15164 17115
rect -15196 17084 -15164 17085
rect -15196 17035 -15164 17036
rect -15196 17005 -15195 17035
rect -15195 17005 -15165 17035
rect -15165 17005 -15164 17035
rect -15196 17004 -15164 17005
rect -15196 16955 -15164 16956
rect -15196 16925 -15195 16955
rect -15195 16925 -15165 16955
rect -15165 16925 -15164 16955
rect -15196 16924 -15164 16925
rect -15196 16875 -15164 16876
rect -15196 16845 -15195 16875
rect -15195 16845 -15165 16875
rect -15165 16845 -15164 16875
rect -15196 16844 -15164 16845
rect -15196 16795 -15164 16796
rect -15196 16765 -15195 16795
rect -15195 16765 -15165 16795
rect -15165 16765 -15164 16795
rect -15196 16764 -15164 16765
rect -15196 16715 -15164 16716
rect -15196 16685 -15195 16715
rect -15195 16685 -15165 16715
rect -15165 16685 -15164 16715
rect -15196 16684 -15164 16685
rect -15196 16635 -15164 16636
rect -15196 16605 -15195 16635
rect -15195 16605 -15165 16635
rect -15165 16605 -15164 16635
rect -15196 16604 -15164 16605
rect -15196 16555 -15164 16556
rect -15196 16525 -15195 16555
rect -15195 16525 -15165 16555
rect -15165 16525 -15164 16555
rect -15196 16524 -15164 16525
rect -15196 16475 -15164 16476
rect -15196 16445 -15195 16475
rect -15195 16445 -15165 16475
rect -15165 16445 -15164 16475
rect -15196 16444 -15164 16445
rect -15036 17115 -15004 17116
rect -15036 17085 -15035 17115
rect -15035 17085 -15005 17115
rect -15005 17085 -15004 17115
rect -15036 17084 -15004 17085
rect -15036 17035 -15004 17036
rect -15036 17005 -15035 17035
rect -15035 17005 -15005 17035
rect -15005 17005 -15004 17035
rect -15036 17004 -15004 17005
rect -15036 16955 -15004 16956
rect -15036 16925 -15035 16955
rect -15035 16925 -15005 16955
rect -15005 16925 -15004 16955
rect -15036 16924 -15004 16925
rect -15036 16875 -15004 16876
rect -15036 16845 -15035 16875
rect -15035 16845 -15005 16875
rect -15005 16845 -15004 16875
rect -15036 16844 -15004 16845
rect -15036 16795 -15004 16796
rect -15036 16765 -15035 16795
rect -15035 16765 -15005 16795
rect -15005 16765 -15004 16795
rect -15036 16764 -15004 16765
rect -15036 16715 -15004 16716
rect -15036 16685 -15035 16715
rect -15035 16685 -15005 16715
rect -15005 16685 -15004 16715
rect -15036 16684 -15004 16685
rect -15036 16635 -15004 16636
rect -15036 16605 -15035 16635
rect -15035 16605 -15005 16635
rect -15005 16605 -15004 16635
rect -15036 16604 -15004 16605
rect -15036 16555 -15004 16556
rect -15036 16525 -15035 16555
rect -15035 16525 -15005 16555
rect -15005 16525 -15004 16555
rect -15036 16524 -15004 16525
rect -15036 16475 -15004 16476
rect -15036 16445 -15035 16475
rect -15035 16445 -15005 16475
rect -15005 16445 -15004 16475
rect -15036 16444 -15004 16445
rect -1676 17395 -1644 17396
rect -1676 17365 -1675 17395
rect -1675 17365 -1645 17395
rect -1645 17365 -1644 17395
rect -1676 17364 -1644 17365
rect -1676 17315 -1644 17316
rect -1676 17285 -1675 17315
rect -1675 17285 -1645 17315
rect -1645 17285 -1644 17315
rect -1676 17284 -1644 17285
rect -1676 17235 -1644 17236
rect -1676 17205 -1675 17235
rect -1675 17205 -1645 17235
rect -1645 17205 -1644 17235
rect -1676 17204 -1644 17205
rect -1676 17155 -1644 17156
rect -1676 17125 -1675 17155
rect -1675 17125 -1645 17155
rect -1645 17125 -1644 17155
rect -1676 17124 -1644 17125
rect -1676 17075 -1644 17076
rect -1676 17045 -1675 17075
rect -1675 17045 -1645 17075
rect -1645 17045 -1644 17075
rect -1676 17044 -1644 17045
rect -1676 16995 -1644 16996
rect -1676 16965 -1675 16995
rect -1675 16965 -1645 16995
rect -1645 16965 -1644 16995
rect -1676 16964 -1644 16965
rect -1676 16915 -1644 16916
rect -1676 16885 -1675 16915
rect -1675 16885 -1645 16915
rect -1645 16885 -1644 16915
rect -1676 16884 -1644 16885
rect -1676 16835 -1644 16836
rect -1676 16805 -1675 16835
rect -1675 16805 -1645 16835
rect -1645 16805 -1644 16835
rect -1676 16804 -1644 16805
rect -1676 16755 -1644 16756
rect -1676 16725 -1675 16755
rect -1675 16725 -1645 16755
rect -1645 16725 -1644 16755
rect -1676 16724 -1644 16725
rect -1676 16635 -1644 16636
rect -1676 16605 -1675 16635
rect -1675 16605 -1645 16635
rect -1645 16605 -1644 16635
rect -1676 16604 -1644 16605
rect -1676 16555 -1644 16556
rect -1676 16525 -1675 16555
rect -1675 16525 -1645 16555
rect -1645 16525 -1644 16555
rect -1676 16524 -1644 16525
rect -1516 17875 -1484 17876
rect -1516 17845 -1515 17875
rect -1515 17845 -1485 17875
rect -1485 17845 -1484 17875
rect -1516 17844 -1484 17845
rect -1516 17795 -1484 17796
rect -1516 17765 -1515 17795
rect -1515 17765 -1485 17795
rect -1485 17765 -1484 17795
rect -1516 17764 -1484 17765
rect -1516 17715 -1484 17716
rect -1516 17685 -1515 17715
rect -1515 17685 -1485 17715
rect -1485 17685 -1484 17715
rect -1516 17684 -1484 17685
rect -1516 17635 -1484 17636
rect -1516 17605 -1515 17635
rect -1515 17605 -1485 17635
rect -1485 17605 -1484 17635
rect -1516 17604 -1484 17605
rect -1516 17555 -1484 17556
rect -1516 17525 -1515 17555
rect -1515 17525 -1485 17555
rect -1485 17525 -1484 17555
rect -1516 17524 -1484 17525
rect -1516 17475 -1484 17476
rect -1516 17445 -1515 17475
rect -1515 17445 -1485 17475
rect -1485 17445 -1484 17475
rect -1516 17444 -1484 17445
rect -1516 17395 -1484 17396
rect -1516 17365 -1515 17395
rect -1515 17365 -1485 17395
rect -1485 17365 -1484 17395
rect -1516 17364 -1484 17365
rect -1516 17315 -1484 17316
rect -1516 17285 -1515 17315
rect -1515 17285 -1485 17315
rect -1485 17285 -1484 17315
rect -1516 17284 -1484 17285
rect -1516 17235 -1484 17236
rect -1516 17205 -1515 17235
rect -1515 17205 -1485 17235
rect -1485 17205 -1484 17235
rect -1516 17204 -1484 17205
rect -1516 17155 -1484 17156
rect -1516 17125 -1515 17155
rect -1515 17125 -1485 17155
rect -1485 17125 -1484 17155
rect -1516 17124 -1484 17125
rect -1516 17075 -1484 17076
rect -1516 17045 -1515 17075
rect -1515 17045 -1485 17075
rect -1485 17045 -1484 17075
rect -1516 17044 -1484 17045
rect -1516 16995 -1484 16996
rect -1516 16965 -1515 16995
rect -1515 16965 -1485 16995
rect -1485 16965 -1484 16995
rect -1516 16964 -1484 16965
rect -1516 16915 -1484 16916
rect -1516 16885 -1515 16915
rect -1515 16885 -1485 16915
rect -1485 16885 -1484 16915
rect -1516 16884 -1484 16885
rect -1516 16835 -1484 16836
rect -1516 16805 -1515 16835
rect -1515 16805 -1485 16835
rect -1485 16805 -1484 16835
rect -1516 16804 -1484 16805
rect -1516 16755 -1484 16756
rect -1516 16725 -1515 16755
rect -1515 16725 -1485 16755
rect -1485 16725 -1484 16755
rect -1516 16724 -1484 16725
rect -1516 16635 -1484 16636
rect -1516 16605 -1515 16635
rect -1515 16605 -1485 16635
rect -1485 16605 -1484 16635
rect -1516 16604 -1484 16605
rect -1516 16555 -1484 16556
rect -1516 16525 -1515 16555
rect -1515 16525 -1485 16555
rect -1485 16525 -1484 16555
rect -1516 16524 -1484 16525
rect -1356 17875 -1324 17876
rect -1356 17845 -1355 17875
rect -1355 17845 -1325 17875
rect -1325 17845 -1324 17875
rect -1356 17844 -1324 17845
rect -1356 17795 -1324 17796
rect -1356 17765 -1355 17795
rect -1355 17765 -1325 17795
rect -1325 17765 -1324 17795
rect -1356 17764 -1324 17765
rect -1356 17715 -1324 17716
rect -1356 17685 -1355 17715
rect -1355 17685 -1325 17715
rect -1325 17685 -1324 17715
rect -1356 17684 -1324 17685
rect -1356 17635 -1324 17636
rect -1356 17605 -1355 17635
rect -1355 17605 -1325 17635
rect -1325 17605 -1324 17635
rect -1356 17604 -1324 17605
rect -1356 17555 -1324 17556
rect -1356 17525 -1355 17555
rect -1355 17525 -1325 17555
rect -1325 17525 -1324 17555
rect -1356 17524 -1324 17525
rect -1356 17475 -1324 17476
rect -1356 17445 -1355 17475
rect -1355 17445 -1325 17475
rect -1325 17445 -1324 17475
rect -1356 17444 -1324 17445
rect -1356 17395 -1324 17396
rect -1356 17365 -1355 17395
rect -1355 17365 -1325 17395
rect -1325 17365 -1324 17395
rect -1356 17364 -1324 17365
rect -1356 17315 -1324 17316
rect -1356 17285 -1355 17315
rect -1355 17285 -1325 17315
rect -1325 17285 -1324 17315
rect -1356 17284 -1324 17285
rect -1356 17235 -1324 17236
rect -1356 17205 -1355 17235
rect -1355 17205 -1325 17235
rect -1325 17205 -1324 17235
rect -1356 17204 -1324 17205
rect -1356 17155 -1324 17156
rect -1356 17125 -1355 17155
rect -1355 17125 -1325 17155
rect -1325 17125 -1324 17155
rect -1356 17124 -1324 17125
rect -1356 17075 -1324 17076
rect -1356 17045 -1355 17075
rect -1355 17045 -1325 17075
rect -1325 17045 -1324 17075
rect -1356 17044 -1324 17045
rect -1356 16995 -1324 16996
rect -1356 16965 -1355 16995
rect -1355 16965 -1325 16995
rect -1325 16965 -1324 16995
rect -1356 16964 -1324 16965
rect -1356 16915 -1324 16916
rect -1356 16885 -1355 16915
rect -1355 16885 -1325 16915
rect -1325 16885 -1324 16915
rect -1356 16884 -1324 16885
rect -1356 16835 -1324 16836
rect -1356 16805 -1355 16835
rect -1355 16805 -1325 16835
rect -1325 16805 -1324 16835
rect -1356 16804 -1324 16805
rect -1356 16755 -1324 16756
rect -1356 16725 -1355 16755
rect -1355 16725 -1325 16755
rect -1325 16725 -1324 16755
rect -1356 16724 -1324 16725
rect -1356 16635 -1324 16636
rect -1356 16605 -1355 16635
rect -1355 16605 -1325 16635
rect -1325 16605 -1324 16635
rect -1356 16604 -1324 16605
rect -1356 16555 -1324 16556
rect -1356 16525 -1355 16555
rect -1355 16525 -1325 16555
rect -1325 16525 -1324 16555
rect -1356 16524 -1324 16525
rect -1196 19875 -1164 19876
rect -1196 19845 -1195 19875
rect -1195 19845 -1165 19875
rect -1165 19845 -1164 19875
rect -1196 19844 -1164 19845
rect -1196 19795 -1164 19796
rect -1196 19765 -1195 19795
rect -1195 19765 -1165 19795
rect -1165 19765 -1164 19795
rect -1196 19764 -1164 19765
rect -1196 19715 -1164 19716
rect -1196 19685 -1195 19715
rect -1195 19685 -1165 19715
rect -1165 19685 -1164 19715
rect -1196 19684 -1164 19685
rect -1196 19635 -1164 19636
rect -1196 19605 -1195 19635
rect -1195 19605 -1165 19635
rect -1165 19605 -1164 19635
rect -1196 19604 -1164 19605
rect -1196 19555 -1164 19556
rect -1196 19525 -1195 19555
rect -1195 19525 -1165 19555
rect -1165 19525 -1164 19555
rect -1196 19524 -1164 19525
rect -1196 19475 -1164 19476
rect -1196 19445 -1195 19475
rect -1195 19445 -1165 19475
rect -1165 19445 -1164 19475
rect -1196 19444 -1164 19445
rect -1196 19395 -1164 19396
rect -1196 19365 -1195 19395
rect -1195 19365 -1165 19395
rect -1165 19365 -1164 19395
rect -1196 19364 -1164 19365
rect -1196 19315 -1164 19316
rect -1196 19285 -1195 19315
rect -1195 19285 -1165 19315
rect -1165 19285 -1164 19315
rect -1196 19284 -1164 19285
rect -1196 19235 -1164 19236
rect -1196 19205 -1195 19235
rect -1195 19205 -1165 19235
rect -1165 19205 -1164 19235
rect -1196 19204 -1164 19205
rect -1196 19155 -1164 19156
rect -1196 19125 -1195 19155
rect -1195 19125 -1165 19155
rect -1165 19125 -1164 19155
rect -1196 19124 -1164 19125
rect -1196 19075 -1164 19076
rect -1196 19045 -1195 19075
rect -1195 19045 -1165 19075
rect -1165 19045 -1164 19075
rect -1196 19044 -1164 19045
rect -1196 18995 -1164 18996
rect -1196 18965 -1195 18995
rect -1195 18965 -1165 18995
rect -1165 18965 -1164 18995
rect -1196 18964 -1164 18965
rect -1196 18915 -1164 18916
rect -1196 18885 -1195 18915
rect -1195 18885 -1165 18915
rect -1165 18885 -1164 18915
rect -1196 18884 -1164 18885
rect -1196 18755 -1164 18756
rect -1196 18725 -1195 18755
rect -1195 18725 -1165 18755
rect -1165 18725 -1164 18755
rect -1196 18724 -1164 18725
rect -1196 18675 -1164 18676
rect -1196 18645 -1195 18675
rect -1195 18645 -1165 18675
rect -1165 18645 -1164 18675
rect -1196 18644 -1164 18645
rect -1196 18595 -1164 18596
rect -1196 18565 -1195 18595
rect -1195 18565 -1165 18595
rect -1165 18565 -1164 18595
rect -1196 18564 -1164 18565
rect -1196 18515 -1164 18516
rect -1196 18485 -1195 18515
rect -1195 18485 -1165 18515
rect -1165 18485 -1164 18515
rect -1196 18484 -1164 18485
rect -1196 18435 -1164 18436
rect -1196 18405 -1195 18435
rect -1195 18405 -1165 18435
rect -1165 18405 -1164 18435
rect -1196 18404 -1164 18405
rect -1196 18355 -1164 18356
rect -1196 18325 -1195 18355
rect -1195 18325 -1165 18355
rect -1165 18325 -1164 18355
rect -1196 18324 -1164 18325
rect -1196 18275 -1164 18276
rect -1196 18245 -1195 18275
rect -1195 18245 -1165 18275
rect -1165 18245 -1164 18275
rect -1196 18244 -1164 18245
rect -1196 18195 -1164 18196
rect -1196 18165 -1195 18195
rect -1195 18165 -1165 18195
rect -1165 18165 -1164 18195
rect -1196 18164 -1164 18165
rect -1196 17875 -1164 17876
rect -1196 17845 -1195 17875
rect -1195 17845 -1165 17875
rect -1165 17845 -1164 17875
rect -1196 17844 -1164 17845
rect -1196 17795 -1164 17796
rect -1196 17765 -1195 17795
rect -1195 17765 -1165 17795
rect -1165 17765 -1164 17795
rect -1196 17764 -1164 17765
rect -1196 17715 -1164 17716
rect -1196 17685 -1195 17715
rect -1195 17685 -1165 17715
rect -1165 17685 -1164 17715
rect -1196 17684 -1164 17685
rect -1196 17635 -1164 17636
rect -1196 17605 -1195 17635
rect -1195 17605 -1165 17635
rect -1165 17605 -1164 17635
rect -1196 17604 -1164 17605
rect -1196 17555 -1164 17556
rect -1196 17525 -1195 17555
rect -1195 17525 -1165 17555
rect -1165 17525 -1164 17555
rect -1196 17524 -1164 17525
rect -1196 17475 -1164 17476
rect -1196 17445 -1195 17475
rect -1195 17445 -1165 17475
rect -1165 17445 -1164 17475
rect -1196 17444 -1164 17445
rect -1196 17395 -1164 17396
rect -1196 17365 -1195 17395
rect -1195 17365 -1165 17395
rect -1165 17365 -1164 17395
rect -1196 17364 -1164 17365
rect -1196 17315 -1164 17316
rect -1196 17285 -1195 17315
rect -1195 17285 -1165 17315
rect -1165 17285 -1164 17315
rect -1196 17284 -1164 17285
rect -1196 17235 -1164 17236
rect -1196 17205 -1195 17235
rect -1195 17205 -1165 17235
rect -1165 17205 -1164 17235
rect -1196 17204 -1164 17205
rect -1196 17155 -1164 17156
rect -1196 17125 -1195 17155
rect -1195 17125 -1165 17155
rect -1165 17125 -1164 17155
rect -1196 17124 -1164 17125
rect -1196 17075 -1164 17076
rect -1196 17045 -1195 17075
rect -1195 17045 -1165 17075
rect -1165 17045 -1164 17075
rect -1196 17044 -1164 17045
rect -1196 16995 -1164 16996
rect -1196 16965 -1195 16995
rect -1195 16965 -1165 16995
rect -1165 16965 -1164 16995
rect -1196 16964 -1164 16965
rect -1196 16915 -1164 16916
rect -1196 16885 -1195 16915
rect -1195 16885 -1165 16915
rect -1165 16885 -1164 16915
rect -1196 16884 -1164 16885
rect -1196 16835 -1164 16836
rect -1196 16805 -1195 16835
rect -1195 16805 -1165 16835
rect -1165 16805 -1164 16835
rect -1196 16804 -1164 16805
rect -1196 16755 -1164 16756
rect -1196 16725 -1195 16755
rect -1195 16725 -1165 16755
rect -1165 16725 -1164 16755
rect -1196 16724 -1164 16725
rect -1196 16635 -1164 16636
rect -1196 16605 -1195 16635
rect -1195 16605 -1165 16635
rect -1165 16605 -1164 16635
rect -1196 16604 -1164 16605
rect -1196 16555 -1164 16556
rect -1196 16525 -1195 16555
rect -1195 16525 -1165 16555
rect -1165 16525 -1164 16555
rect -1196 16524 -1164 16525
rect -1036 19875 -1004 19876
rect -1036 19845 -1035 19875
rect -1035 19845 -1005 19875
rect -1005 19845 -1004 19875
rect -1036 19844 -1004 19845
rect -1036 19795 -1004 19796
rect -1036 19765 -1035 19795
rect -1035 19765 -1005 19795
rect -1005 19765 -1004 19795
rect -1036 19764 -1004 19765
rect -1036 19715 -1004 19716
rect -1036 19685 -1035 19715
rect -1035 19685 -1005 19715
rect -1005 19685 -1004 19715
rect -1036 19684 -1004 19685
rect -1036 19635 -1004 19636
rect -1036 19605 -1035 19635
rect -1035 19605 -1005 19635
rect -1005 19605 -1004 19635
rect -1036 19604 -1004 19605
rect -1036 19555 -1004 19556
rect -1036 19525 -1035 19555
rect -1035 19525 -1005 19555
rect -1005 19525 -1004 19555
rect -1036 19524 -1004 19525
rect -1036 19475 -1004 19476
rect -1036 19445 -1035 19475
rect -1035 19445 -1005 19475
rect -1005 19445 -1004 19475
rect -1036 19444 -1004 19445
rect -1036 19395 -1004 19396
rect -1036 19365 -1035 19395
rect -1035 19365 -1005 19395
rect -1005 19365 -1004 19395
rect -1036 19364 -1004 19365
rect -1036 19315 -1004 19316
rect -1036 19285 -1035 19315
rect -1035 19285 -1005 19315
rect -1005 19285 -1004 19315
rect -1036 19284 -1004 19285
rect -1036 19235 -1004 19236
rect -1036 19205 -1035 19235
rect -1035 19205 -1005 19235
rect -1005 19205 -1004 19235
rect -1036 19204 -1004 19205
rect -1036 19155 -1004 19156
rect -1036 19125 -1035 19155
rect -1035 19125 -1005 19155
rect -1005 19125 -1004 19155
rect -1036 19124 -1004 19125
rect -1036 19075 -1004 19076
rect -1036 19045 -1035 19075
rect -1035 19045 -1005 19075
rect -1005 19045 -1004 19075
rect -1036 19044 -1004 19045
rect -1036 18995 -1004 18996
rect -1036 18965 -1035 18995
rect -1035 18965 -1005 18995
rect -1005 18965 -1004 18995
rect -1036 18964 -1004 18965
rect -1036 18915 -1004 18916
rect -1036 18885 -1035 18915
rect -1035 18885 -1005 18915
rect -1005 18885 -1004 18915
rect -1036 18884 -1004 18885
rect -1036 18755 -1004 18756
rect -1036 18725 -1035 18755
rect -1035 18725 -1005 18755
rect -1005 18725 -1004 18755
rect -1036 18724 -1004 18725
rect -1036 18675 -1004 18676
rect -1036 18645 -1035 18675
rect -1035 18645 -1005 18675
rect -1005 18645 -1004 18675
rect -1036 18644 -1004 18645
rect -1036 18595 -1004 18596
rect -1036 18565 -1035 18595
rect -1035 18565 -1005 18595
rect -1005 18565 -1004 18595
rect -1036 18564 -1004 18565
rect -1036 18515 -1004 18516
rect -1036 18485 -1035 18515
rect -1035 18485 -1005 18515
rect -1005 18485 -1004 18515
rect -1036 18484 -1004 18485
rect -1036 18435 -1004 18436
rect -1036 18405 -1035 18435
rect -1035 18405 -1005 18435
rect -1005 18405 -1004 18435
rect -1036 18404 -1004 18405
rect -1036 18355 -1004 18356
rect -1036 18325 -1035 18355
rect -1035 18325 -1005 18355
rect -1005 18325 -1004 18355
rect -1036 18324 -1004 18325
rect -1036 18275 -1004 18276
rect -1036 18245 -1035 18275
rect -1035 18245 -1005 18275
rect -1005 18245 -1004 18275
rect -1036 18244 -1004 18245
rect -1036 18195 -1004 18196
rect -1036 18165 -1035 18195
rect -1035 18165 -1005 18195
rect -1005 18165 -1004 18195
rect -1036 18164 -1004 18165
rect -876 19875 -844 19876
rect -876 19845 -875 19875
rect -875 19845 -845 19875
rect -845 19845 -844 19875
rect -876 19844 -844 19845
rect -876 19795 -844 19796
rect -876 19765 -875 19795
rect -875 19765 -845 19795
rect -845 19765 -844 19795
rect -876 19764 -844 19765
rect -876 19715 -844 19716
rect -876 19685 -875 19715
rect -875 19685 -845 19715
rect -845 19685 -844 19715
rect -876 19684 -844 19685
rect -876 19635 -844 19636
rect -876 19605 -875 19635
rect -875 19605 -845 19635
rect -845 19605 -844 19635
rect -876 19604 -844 19605
rect -876 19555 -844 19556
rect -876 19525 -875 19555
rect -875 19525 -845 19555
rect -845 19525 -844 19555
rect -876 19524 -844 19525
rect -876 19475 -844 19476
rect -876 19445 -875 19475
rect -875 19445 -845 19475
rect -845 19445 -844 19475
rect -876 19444 -844 19445
rect -876 19395 -844 19396
rect -876 19365 -875 19395
rect -875 19365 -845 19395
rect -845 19365 -844 19395
rect -876 19364 -844 19365
rect -876 19315 -844 19316
rect -876 19285 -875 19315
rect -875 19285 -845 19315
rect -845 19285 -844 19315
rect -876 19284 -844 19285
rect -876 19235 -844 19236
rect -876 19205 -875 19235
rect -875 19205 -845 19235
rect -845 19205 -844 19235
rect -876 19204 -844 19205
rect -876 19155 -844 19156
rect -876 19125 -875 19155
rect -875 19125 -845 19155
rect -845 19125 -844 19155
rect -876 19124 -844 19125
rect -876 19075 -844 19076
rect -876 19045 -875 19075
rect -875 19045 -845 19075
rect -845 19045 -844 19075
rect -876 19044 -844 19045
rect -876 18995 -844 18996
rect -876 18965 -875 18995
rect -875 18965 -845 18995
rect -845 18965 -844 18995
rect -876 18964 -844 18965
rect -876 18915 -844 18916
rect -876 18885 -875 18915
rect -875 18885 -845 18915
rect -845 18885 -844 18915
rect -876 18884 -844 18885
rect -876 18755 -844 18756
rect -876 18725 -875 18755
rect -875 18725 -845 18755
rect -845 18725 -844 18755
rect -876 18724 -844 18725
rect -876 18675 -844 18676
rect -876 18645 -875 18675
rect -875 18645 -845 18675
rect -845 18645 -844 18675
rect -876 18644 -844 18645
rect -876 18595 -844 18596
rect -876 18565 -875 18595
rect -875 18565 -845 18595
rect -845 18565 -844 18595
rect -876 18564 -844 18565
rect -876 18515 -844 18516
rect -876 18485 -875 18515
rect -875 18485 -845 18515
rect -845 18485 -844 18515
rect -876 18484 -844 18485
rect -876 18435 -844 18436
rect -876 18405 -875 18435
rect -875 18405 -845 18435
rect -845 18405 -844 18435
rect -876 18404 -844 18405
rect -876 18355 -844 18356
rect -876 18325 -875 18355
rect -875 18325 -845 18355
rect -845 18325 -844 18355
rect -876 18324 -844 18325
rect -876 18275 -844 18276
rect -876 18245 -875 18275
rect -875 18245 -845 18275
rect -845 18245 -844 18275
rect -876 18244 -844 18245
rect -876 18195 -844 18196
rect -876 18165 -875 18195
rect -875 18165 -845 18195
rect -845 18165 -844 18195
rect -876 18164 -844 18165
rect -1036 17875 -1004 17876
rect -1036 17845 -1035 17875
rect -1035 17845 -1005 17875
rect -1005 17845 -1004 17875
rect -1036 17844 -1004 17845
rect -1036 17795 -1004 17796
rect -1036 17765 -1035 17795
rect -1035 17765 -1005 17795
rect -1005 17765 -1004 17795
rect -1036 17764 -1004 17765
rect -1036 17715 -1004 17716
rect -1036 17685 -1035 17715
rect -1035 17685 -1005 17715
rect -1005 17685 -1004 17715
rect -1036 17684 -1004 17685
rect -1036 17635 -1004 17636
rect -1036 17605 -1035 17635
rect -1035 17605 -1005 17635
rect -1005 17605 -1004 17635
rect -1036 17604 -1004 17605
rect -1036 17555 -1004 17556
rect -1036 17525 -1035 17555
rect -1035 17525 -1005 17555
rect -1005 17525 -1004 17555
rect -1036 17524 -1004 17525
rect -1036 17475 -1004 17476
rect -1036 17445 -1035 17475
rect -1035 17445 -1005 17475
rect -1005 17445 -1004 17475
rect -1036 17444 -1004 17445
rect -1036 17395 -1004 17396
rect -1036 17365 -1035 17395
rect -1035 17365 -1005 17395
rect -1005 17365 -1004 17395
rect -1036 17364 -1004 17365
rect -1036 17315 -1004 17316
rect -1036 17285 -1035 17315
rect -1035 17285 -1005 17315
rect -1005 17285 -1004 17315
rect -1036 17284 -1004 17285
rect -1036 17235 -1004 17236
rect -1036 17205 -1035 17235
rect -1035 17205 -1005 17235
rect -1005 17205 -1004 17235
rect -1036 17204 -1004 17205
rect -1036 17155 -1004 17156
rect -1036 17125 -1035 17155
rect -1035 17125 -1005 17155
rect -1005 17125 -1004 17155
rect -1036 17124 -1004 17125
rect -1036 17075 -1004 17076
rect -1036 17045 -1035 17075
rect -1035 17045 -1005 17075
rect -1005 17045 -1004 17075
rect -1036 17044 -1004 17045
rect -1036 16995 -1004 16996
rect -1036 16965 -1035 16995
rect -1035 16965 -1005 16995
rect -1005 16965 -1004 16995
rect -1036 16964 -1004 16965
rect -1036 16915 -1004 16916
rect -1036 16885 -1035 16915
rect -1035 16885 -1005 16915
rect -1005 16885 -1004 16915
rect -1036 16884 -1004 16885
rect -1036 16835 -1004 16836
rect -1036 16805 -1035 16835
rect -1035 16805 -1005 16835
rect -1005 16805 -1004 16835
rect -1036 16804 -1004 16805
rect -1036 16755 -1004 16756
rect -1036 16725 -1035 16755
rect -1035 16725 -1005 16755
rect -1005 16725 -1004 16755
rect -1036 16724 -1004 16725
rect -1036 16635 -1004 16636
rect -1036 16605 -1035 16635
rect -1035 16605 -1005 16635
rect -1005 16605 -1004 16635
rect -1036 16604 -1004 16605
rect -1036 16555 -1004 16556
rect -1036 16525 -1035 16555
rect -1035 16525 -1005 16555
rect -1005 16525 -1004 16555
rect -1036 16524 -1004 16525
rect -716 19875 -684 19876
rect -716 19845 -715 19875
rect -715 19845 -685 19875
rect -685 19845 -684 19875
rect -716 19844 -684 19845
rect -716 19795 -684 19796
rect -716 19765 -715 19795
rect -715 19765 -685 19795
rect -685 19765 -684 19795
rect -716 19764 -684 19765
rect -716 19715 -684 19716
rect -716 19685 -715 19715
rect -715 19685 -685 19715
rect -685 19685 -684 19715
rect -716 19684 -684 19685
rect -716 19635 -684 19636
rect -716 19605 -715 19635
rect -715 19605 -685 19635
rect -685 19605 -684 19635
rect -716 19604 -684 19605
rect -716 19555 -684 19556
rect -716 19525 -715 19555
rect -715 19525 -685 19555
rect -685 19525 -684 19555
rect -716 19524 -684 19525
rect -716 19475 -684 19476
rect -716 19445 -715 19475
rect -715 19445 -685 19475
rect -685 19445 -684 19475
rect -716 19444 -684 19445
rect -716 19395 -684 19396
rect -716 19365 -715 19395
rect -715 19365 -685 19395
rect -685 19365 -684 19395
rect -716 19364 -684 19365
rect -716 19315 -684 19316
rect -716 19285 -715 19315
rect -715 19285 -685 19315
rect -685 19285 -684 19315
rect -716 19284 -684 19285
rect -716 19235 -684 19236
rect -716 19205 -715 19235
rect -715 19205 -685 19235
rect -685 19205 -684 19235
rect -716 19204 -684 19205
rect -716 19155 -684 19156
rect -716 19125 -715 19155
rect -715 19125 -685 19155
rect -685 19125 -684 19155
rect -716 19124 -684 19125
rect -716 19075 -684 19076
rect -716 19045 -715 19075
rect -715 19045 -685 19075
rect -685 19045 -684 19075
rect -716 19044 -684 19045
rect -716 18995 -684 18996
rect -716 18965 -715 18995
rect -715 18965 -685 18995
rect -685 18965 -684 18995
rect -716 18964 -684 18965
rect -716 18915 -684 18916
rect -716 18885 -715 18915
rect -715 18885 -685 18915
rect -685 18885 -684 18915
rect -716 18884 -684 18885
rect -556 19875 -524 19876
rect -556 19845 -555 19875
rect -555 19845 -525 19875
rect -525 19845 -524 19875
rect -556 19844 -524 19845
rect -556 19795 -524 19796
rect -556 19765 -555 19795
rect -555 19765 -525 19795
rect -525 19765 -524 19795
rect -556 19764 -524 19765
rect -556 19715 -524 19716
rect -556 19685 -555 19715
rect -555 19685 -525 19715
rect -525 19685 -524 19715
rect -556 19684 -524 19685
rect -556 19635 -524 19636
rect -556 19605 -555 19635
rect -555 19605 -525 19635
rect -525 19605 -524 19635
rect -556 19604 -524 19605
rect -556 19555 -524 19556
rect -556 19525 -555 19555
rect -555 19525 -525 19555
rect -525 19525 -524 19555
rect -556 19524 -524 19525
rect -556 19475 -524 19476
rect -556 19445 -555 19475
rect -555 19445 -525 19475
rect -525 19445 -524 19475
rect -556 19444 -524 19445
rect -556 19395 -524 19396
rect -556 19365 -555 19395
rect -555 19365 -525 19395
rect -525 19365 -524 19395
rect -556 19364 -524 19365
rect -556 19315 -524 19316
rect -556 19285 -555 19315
rect -555 19285 -525 19315
rect -525 19285 -524 19315
rect -556 19284 -524 19285
rect -556 19235 -524 19236
rect -556 19205 -555 19235
rect -555 19205 -525 19235
rect -525 19205 -524 19235
rect -556 19204 -524 19205
rect -556 19155 -524 19156
rect -556 19125 -555 19155
rect -555 19125 -525 19155
rect -525 19125 -524 19155
rect -556 19124 -524 19125
rect -556 19075 -524 19076
rect -556 19045 -555 19075
rect -555 19045 -525 19075
rect -525 19045 -524 19075
rect -556 19044 -524 19045
rect -556 18995 -524 18996
rect -556 18965 -555 18995
rect -555 18965 -525 18995
rect -525 18965 -524 18995
rect -556 18964 -524 18965
rect -556 18915 -524 18916
rect -556 18885 -555 18915
rect -555 18885 -525 18915
rect -525 18885 -524 18915
rect -556 18884 -524 18885
rect -716 18755 -684 18756
rect -716 18725 -715 18755
rect -715 18725 -685 18755
rect -685 18725 -684 18755
rect -716 18724 -684 18725
rect -716 18675 -684 18676
rect -716 18645 -715 18675
rect -715 18645 -685 18675
rect -685 18645 -684 18675
rect -716 18644 -684 18645
rect -716 18595 -684 18596
rect -716 18565 -715 18595
rect -715 18565 -685 18595
rect -685 18565 -684 18595
rect -716 18564 -684 18565
rect -716 18515 -684 18516
rect -716 18485 -715 18515
rect -715 18485 -685 18515
rect -685 18485 -684 18515
rect -716 18484 -684 18485
rect -716 18435 -684 18436
rect -716 18405 -715 18435
rect -715 18405 -685 18435
rect -685 18405 -684 18435
rect -716 18404 -684 18405
rect -716 18355 -684 18356
rect -716 18325 -715 18355
rect -715 18325 -685 18355
rect -685 18325 -684 18355
rect -716 18324 -684 18325
rect -716 18275 -684 18276
rect -716 18245 -715 18275
rect -715 18245 -685 18275
rect -685 18245 -684 18275
rect -716 18244 -684 18245
rect -716 18195 -684 18196
rect -716 18165 -715 18195
rect -715 18165 -685 18195
rect -685 18165 -684 18195
rect -716 18164 -684 18165
rect -876 17875 -844 17876
rect -876 17845 -875 17875
rect -875 17845 -845 17875
rect -845 17845 -844 17875
rect -876 17844 -844 17845
rect -876 17795 -844 17796
rect -876 17765 -875 17795
rect -875 17765 -845 17795
rect -845 17765 -844 17795
rect -876 17764 -844 17765
rect -876 17715 -844 17716
rect -876 17685 -875 17715
rect -875 17685 -845 17715
rect -845 17685 -844 17715
rect -876 17684 -844 17685
rect -876 17635 -844 17636
rect -876 17605 -875 17635
rect -875 17605 -845 17635
rect -845 17605 -844 17635
rect -876 17604 -844 17605
rect -876 17555 -844 17556
rect -876 17525 -875 17555
rect -875 17525 -845 17555
rect -845 17525 -844 17555
rect -876 17524 -844 17525
rect -876 17475 -844 17476
rect -876 17445 -875 17475
rect -875 17445 -845 17475
rect -845 17445 -844 17475
rect -876 17444 -844 17445
rect -876 17395 -844 17396
rect -876 17365 -875 17395
rect -875 17365 -845 17395
rect -845 17365 -844 17395
rect -876 17364 -844 17365
rect -876 17315 -844 17316
rect -876 17285 -875 17315
rect -875 17285 -845 17315
rect -845 17285 -844 17315
rect -876 17284 -844 17285
rect -876 17235 -844 17236
rect -876 17205 -875 17235
rect -875 17205 -845 17235
rect -845 17205 -844 17235
rect -876 17204 -844 17205
rect -876 17155 -844 17156
rect -876 17125 -875 17155
rect -875 17125 -845 17155
rect -845 17125 -844 17155
rect -876 17124 -844 17125
rect -876 17075 -844 17076
rect -876 17045 -875 17075
rect -875 17045 -845 17075
rect -845 17045 -844 17075
rect -876 17044 -844 17045
rect -876 16995 -844 16996
rect -876 16965 -875 16995
rect -875 16965 -845 16995
rect -845 16965 -844 16995
rect -876 16964 -844 16965
rect -876 16915 -844 16916
rect -876 16885 -875 16915
rect -875 16885 -845 16915
rect -845 16885 -844 16915
rect -876 16884 -844 16885
rect -876 16835 -844 16836
rect -876 16805 -875 16835
rect -875 16805 -845 16835
rect -845 16805 -844 16835
rect -876 16804 -844 16805
rect -876 16755 -844 16756
rect -876 16725 -875 16755
rect -875 16725 -845 16755
rect -845 16725 -844 16755
rect -876 16724 -844 16725
rect -876 16635 -844 16636
rect -876 16605 -875 16635
rect -875 16605 -845 16635
rect -845 16605 -844 16635
rect -876 16604 -844 16605
rect -876 16555 -844 16556
rect -876 16525 -875 16555
rect -875 16525 -845 16555
rect -845 16525 -844 16555
rect -876 16524 -844 16525
rect -716 17875 -684 17876
rect -716 17845 -715 17875
rect -715 17845 -685 17875
rect -685 17845 -684 17875
rect -716 17844 -684 17845
rect -716 17795 -684 17796
rect -716 17765 -715 17795
rect -715 17765 -685 17795
rect -685 17765 -684 17795
rect -716 17764 -684 17765
rect -716 17715 -684 17716
rect -716 17685 -715 17715
rect -715 17685 -685 17715
rect -685 17685 -684 17715
rect -716 17684 -684 17685
rect -716 17635 -684 17636
rect -716 17605 -715 17635
rect -715 17605 -685 17635
rect -685 17605 -684 17635
rect -716 17604 -684 17605
rect -716 17555 -684 17556
rect -716 17525 -715 17555
rect -715 17525 -685 17555
rect -685 17525 -684 17555
rect -716 17524 -684 17525
rect -716 17475 -684 17476
rect -716 17445 -715 17475
rect -715 17445 -685 17475
rect -685 17445 -684 17475
rect -716 17444 -684 17445
rect -716 17395 -684 17396
rect -716 17365 -715 17395
rect -715 17365 -685 17395
rect -685 17365 -684 17395
rect -716 17364 -684 17365
rect -716 17315 -684 17316
rect -716 17285 -715 17315
rect -715 17285 -685 17315
rect -685 17285 -684 17315
rect -716 17284 -684 17285
rect -716 17235 -684 17236
rect -716 17205 -715 17235
rect -715 17205 -685 17235
rect -685 17205 -684 17235
rect -716 17204 -684 17205
rect -716 17155 -684 17156
rect -716 17125 -715 17155
rect -715 17125 -685 17155
rect -685 17125 -684 17155
rect -716 17124 -684 17125
rect -716 17075 -684 17076
rect -716 17045 -715 17075
rect -715 17045 -685 17075
rect -685 17045 -684 17075
rect -716 17044 -684 17045
rect -716 16995 -684 16996
rect -716 16965 -715 16995
rect -715 16965 -685 16995
rect -685 16965 -684 16995
rect -716 16964 -684 16965
rect -716 16915 -684 16916
rect -716 16885 -715 16915
rect -715 16885 -685 16915
rect -685 16885 -684 16915
rect -716 16884 -684 16885
rect -716 16835 -684 16836
rect -716 16805 -715 16835
rect -715 16805 -685 16835
rect -685 16805 -684 16835
rect -716 16804 -684 16805
rect -716 16755 -684 16756
rect -716 16725 -715 16755
rect -715 16725 -685 16755
rect -685 16725 -684 16755
rect -716 16724 -684 16725
rect -716 16635 -684 16636
rect -716 16605 -715 16635
rect -715 16605 -685 16635
rect -685 16605 -684 16635
rect -716 16604 -684 16605
rect -716 16555 -684 16556
rect -716 16525 -715 16555
rect -715 16525 -685 16555
rect -685 16525 -684 16555
rect -716 16524 -684 16525
rect -556 18755 -524 18756
rect -556 18725 -555 18755
rect -555 18725 -525 18755
rect -525 18725 -524 18755
rect -556 18724 -524 18725
rect -556 18675 -524 18676
rect -556 18645 -555 18675
rect -555 18645 -525 18675
rect -525 18645 -524 18675
rect -556 18644 -524 18645
rect -556 18595 -524 18596
rect -556 18565 -555 18595
rect -555 18565 -525 18595
rect -525 18565 -524 18595
rect -556 18564 -524 18565
rect -556 18515 -524 18516
rect -556 18485 -555 18515
rect -555 18485 -525 18515
rect -525 18485 -524 18515
rect -556 18484 -524 18485
rect -556 18435 -524 18436
rect -556 18405 -555 18435
rect -555 18405 -525 18435
rect -525 18405 -524 18435
rect -556 18404 -524 18405
rect -556 18355 -524 18356
rect -556 18325 -555 18355
rect -555 18325 -525 18355
rect -525 18325 -524 18355
rect -556 18324 -524 18325
rect -556 18275 -524 18276
rect -556 18245 -555 18275
rect -555 18245 -525 18275
rect -525 18245 -524 18275
rect -556 18244 -524 18245
rect -556 18195 -524 18196
rect -556 18165 -555 18195
rect -555 18165 -525 18195
rect -525 18165 -524 18195
rect -556 18164 -524 18165
rect -556 17875 -524 17876
rect -556 17845 -555 17875
rect -555 17845 -525 17875
rect -525 17845 -524 17875
rect -556 17844 -524 17845
rect -556 17795 -524 17796
rect -556 17765 -555 17795
rect -555 17765 -525 17795
rect -525 17765 -524 17795
rect -556 17764 -524 17765
rect -556 17715 -524 17716
rect -556 17685 -555 17715
rect -555 17685 -525 17715
rect -525 17685 -524 17715
rect -556 17684 -524 17685
rect -556 17635 -524 17636
rect -556 17605 -555 17635
rect -555 17605 -525 17635
rect -525 17605 -524 17635
rect -556 17604 -524 17605
rect -556 17555 -524 17556
rect -556 17525 -555 17555
rect -555 17525 -525 17555
rect -525 17525 -524 17555
rect -556 17524 -524 17525
rect -556 17475 -524 17476
rect -556 17445 -555 17475
rect -555 17445 -525 17475
rect -525 17445 -524 17475
rect -556 17444 -524 17445
rect -556 17395 -524 17396
rect -556 17365 -555 17395
rect -555 17365 -525 17395
rect -525 17365 -524 17395
rect -556 17364 -524 17365
rect -556 17315 -524 17316
rect -556 17285 -555 17315
rect -555 17285 -525 17315
rect -525 17285 -524 17315
rect -556 17284 -524 17285
rect -556 17235 -524 17236
rect -556 17205 -555 17235
rect -555 17205 -525 17235
rect -525 17205 -524 17235
rect -556 17204 -524 17205
rect -556 17155 -524 17156
rect -556 17125 -555 17155
rect -555 17125 -525 17155
rect -525 17125 -524 17155
rect -556 17124 -524 17125
rect -556 17075 -524 17076
rect -556 17045 -555 17075
rect -555 17045 -525 17075
rect -525 17045 -524 17075
rect -556 17044 -524 17045
rect -556 16995 -524 16996
rect -556 16965 -555 16995
rect -555 16965 -525 16995
rect -525 16965 -524 16995
rect -556 16964 -524 16965
rect -556 16915 -524 16916
rect -556 16885 -555 16915
rect -555 16885 -525 16915
rect -525 16885 -524 16915
rect -556 16884 -524 16885
rect -556 16835 -524 16836
rect -556 16805 -555 16835
rect -555 16805 -525 16835
rect -525 16805 -524 16835
rect -556 16804 -524 16805
rect -556 16755 -524 16756
rect -556 16725 -555 16755
rect -555 16725 -525 16755
rect -525 16725 -524 16755
rect -556 16724 -524 16725
rect -556 16635 -524 16636
rect -556 16605 -555 16635
rect -555 16605 -525 16635
rect -525 16605 -524 16635
rect -556 16604 -524 16605
rect -556 16555 -524 16556
rect -556 16525 -555 16555
rect -555 16525 -525 16555
rect -525 16525 -524 16555
rect -556 16524 -524 16525
<< metal4 >>
rect -16560 39480 21600 39520
rect -16560 39360 -16520 39480
rect -16400 39360 21440 39480
rect 21560 39360 21600 39480
rect -16560 39320 21600 39360
rect -16560 39240 21600 39280
rect -16560 39120 -16120 39240
rect -16000 39120 21040 39240
rect 21160 39120 21600 39240
rect -16560 39080 21600 39120
rect -16560 39000 21600 39040
rect -16560 38880 -15720 39000
rect -15600 38880 20640 39000
rect 20760 38880 21600 39000
rect -16560 38840 21600 38880
rect -15760 37400 -15520 37440
rect -15760 37280 -15720 37400
rect -15600 37280 -15520 37400
rect -15760 37240 -15520 37280
rect -520 37240 -480 37440
rect 20480 37400 20800 37440
rect 20480 37280 20640 37400
rect 20760 37280 20800 37400
rect 20480 37240 20800 37280
rect -16160 37160 -15520 37200
rect -16160 37040 -16120 37160
rect -16000 37040 -15520 37160
rect -16160 37000 -15520 37040
rect -520 37000 -480 37200
rect 20480 37160 21200 37200
rect 20480 37040 21040 37160
rect 21160 37040 21200 37160
rect 20480 37000 21200 37040
rect 20480 36680 21600 36720
rect 20480 36560 21440 36680
rect 21560 36560 21600 36680
rect 20480 36520 21600 36560
rect -15520 20876 -15000 20880
rect -15520 20844 -15516 20876
rect -15484 20844 -15356 20876
rect -15324 20844 -15196 20876
rect -15164 20844 -15036 20876
rect -15004 20844 -15000 20876
rect -15520 20840 -15000 20844
rect -15520 20796 -15000 20800
rect -15520 20764 -15516 20796
rect -15484 20764 -15356 20796
rect -15324 20764 -15196 20796
rect -15164 20764 -15036 20796
rect -15004 20764 -15000 20796
rect -15520 20760 -15000 20764
rect -15520 20396 -15000 20400
rect -15520 20364 -15516 20396
rect -15484 20364 -15356 20396
rect -15324 20364 -15196 20396
rect -15164 20364 -15036 20396
rect -15004 20364 -15000 20396
rect -15520 20360 -15000 20364
rect -15520 20316 -15000 20320
rect -15520 20284 -15516 20316
rect -15484 20284 -15356 20316
rect -15324 20284 -15196 20316
rect -15164 20284 -15036 20316
rect -15004 20284 -15000 20316
rect -15520 20280 -15000 20284
rect -15520 20236 -15000 20240
rect -15520 20204 -15516 20236
rect -15484 20204 -15356 20236
rect -15324 20204 -15196 20236
rect -15164 20204 -15036 20236
rect -15004 20204 -15000 20236
rect -15520 20200 -15000 20204
rect -15520 20156 -15000 20160
rect -15520 20124 -15516 20156
rect -15484 20124 -15356 20156
rect -15324 20124 -15196 20156
rect -15164 20124 -15036 20156
rect -15004 20124 -15000 20156
rect -15520 20120 -15000 20124
rect -15520 20076 -15000 20080
rect -15520 20044 -15516 20076
rect -15484 20044 -15356 20076
rect -15324 20044 -15196 20076
rect -15164 20044 -15036 20076
rect -15004 20044 -15000 20076
rect -15520 20040 -15000 20044
rect -15520 19996 -15000 20000
rect -15520 19964 -15516 19996
rect -15484 19964 -15356 19996
rect -15324 19964 -15196 19996
rect -15164 19964 -15036 19996
rect -15004 19964 -15000 19996
rect -15520 19960 -15000 19964
rect -15520 19916 -15000 19920
rect -15520 19884 -15516 19916
rect -15484 19884 -15356 19916
rect -15324 19884 -15196 19916
rect -15164 19884 -15036 19916
rect -15004 19884 -15000 19916
rect -15520 19880 -15000 19884
rect -1680 19876 -520 19880
rect -1680 19844 -1676 19876
rect -1644 19844 -1516 19876
rect -1484 19844 -1356 19876
rect -1324 19844 -1196 19876
rect -1164 19844 -1036 19876
rect -1004 19844 -876 19876
rect -844 19844 -716 19876
rect -684 19844 -556 19876
rect -524 19844 -520 19876
rect -1680 19840 -520 19844
rect -15520 19836 -15000 19840
rect -15520 19804 -15516 19836
rect -15484 19804 -15356 19836
rect -15324 19804 -15196 19836
rect -15164 19804 -15036 19836
rect -15004 19804 -15000 19836
rect -15520 19800 -15000 19804
rect -1680 19796 -520 19800
rect -1680 19764 -1676 19796
rect -1644 19764 -1516 19796
rect -1484 19764 -1356 19796
rect -1324 19764 -1196 19796
rect -1164 19764 -1036 19796
rect -1004 19764 -876 19796
rect -844 19764 -716 19796
rect -684 19764 -556 19796
rect -524 19764 -520 19796
rect -1680 19760 -520 19764
rect -15520 19756 -15000 19760
rect -15520 19724 -15516 19756
rect -15484 19724 -15356 19756
rect -15324 19724 -15196 19756
rect -15164 19724 -15036 19756
rect -15004 19724 -15000 19756
rect -15520 19720 -15000 19724
rect -1680 19716 -520 19720
rect -1680 19684 -1676 19716
rect -1644 19684 -1516 19716
rect -1484 19684 -1356 19716
rect -1324 19684 -1196 19716
rect -1164 19684 -1036 19716
rect -1004 19684 -876 19716
rect -844 19684 -716 19716
rect -684 19684 -556 19716
rect -524 19684 -520 19716
rect -1680 19680 -520 19684
rect -15520 19676 -15000 19680
rect -15520 19644 -15516 19676
rect -15484 19644 -15356 19676
rect -15324 19644 -15196 19676
rect -15164 19644 -15036 19676
rect -15004 19644 -15000 19676
rect -15520 19640 -15000 19644
rect -1680 19636 -520 19640
rect -1680 19604 -1676 19636
rect -1644 19604 -1516 19636
rect -1484 19604 -1356 19636
rect -1324 19604 -1196 19636
rect -1164 19604 -1036 19636
rect -1004 19604 -876 19636
rect -844 19604 -716 19636
rect -684 19604 -556 19636
rect -524 19604 -520 19636
rect -1680 19600 -520 19604
rect -15520 19596 -15000 19600
rect -15520 19564 -15516 19596
rect -15484 19564 -15356 19596
rect -15324 19564 -15196 19596
rect -15164 19564 -15036 19596
rect -15004 19564 -15000 19596
rect -15520 19560 -15000 19564
rect -1680 19556 -520 19560
rect -1680 19524 -1676 19556
rect -1644 19524 -1516 19556
rect -1484 19524 -1356 19556
rect -1324 19524 -1196 19556
rect -1164 19524 -1036 19556
rect -1004 19524 -876 19556
rect -844 19524 -716 19556
rect -684 19524 -556 19556
rect -524 19524 -520 19556
rect -1680 19520 -520 19524
rect -15520 19516 -15000 19520
rect -15520 19484 -15516 19516
rect -15484 19484 -15356 19516
rect -15324 19484 -15196 19516
rect -15164 19484 -15036 19516
rect -15004 19484 -15000 19516
rect -15520 19480 -15000 19484
rect -1680 19476 -520 19480
rect -1680 19444 -1676 19476
rect -1644 19444 -1516 19476
rect -1484 19444 -1356 19476
rect -1324 19444 -1196 19476
rect -1164 19444 -1036 19476
rect -1004 19444 -876 19476
rect -844 19444 -716 19476
rect -684 19444 -556 19476
rect -524 19444 -520 19476
rect -1680 19440 -520 19444
rect -15520 19436 -15000 19440
rect -15520 19404 -15516 19436
rect -15484 19404 -15356 19436
rect -15324 19404 -15196 19436
rect -15164 19404 -15036 19436
rect -15004 19404 -15000 19436
rect -15520 19400 -15000 19404
rect -1680 19396 -520 19400
rect -1680 19364 -1676 19396
rect -1644 19364 -1516 19396
rect -1484 19364 -1356 19396
rect -1324 19364 -1196 19396
rect -1164 19364 -1036 19396
rect -1004 19364 -876 19396
rect -844 19364 -716 19396
rect -684 19364 -556 19396
rect -524 19364 -520 19396
rect -1680 19360 -520 19364
rect -15520 19356 -15000 19360
rect -15520 19324 -15516 19356
rect -15484 19324 -15356 19356
rect -15324 19324 -15196 19356
rect -15164 19324 -15036 19356
rect -15004 19324 -15000 19356
rect -15520 19320 -15000 19324
rect -1680 19316 -520 19320
rect -1680 19284 -1676 19316
rect -1644 19284 -1516 19316
rect -1484 19284 -1356 19316
rect -1324 19284 -1196 19316
rect -1164 19284 -1036 19316
rect -1004 19284 -876 19316
rect -844 19284 -716 19316
rect -684 19284 -556 19316
rect -524 19284 -520 19316
rect -1680 19280 -520 19284
rect -15520 19276 -15000 19280
rect -15520 19244 -15516 19276
rect -15484 19244 -15356 19276
rect -15324 19244 -15196 19276
rect -15164 19244 -15036 19276
rect -15004 19244 -15000 19276
rect -15520 19240 -15000 19244
rect -1680 19236 -520 19240
rect -1680 19204 -1676 19236
rect -1644 19204 -1516 19236
rect -1484 19204 -1356 19236
rect -1324 19204 -1196 19236
rect -1164 19204 -1036 19236
rect -1004 19204 -876 19236
rect -844 19204 -716 19236
rect -684 19204 -556 19236
rect -524 19204 -520 19236
rect -1680 19200 -520 19204
rect -15520 19196 -15000 19200
rect -15520 19164 -15516 19196
rect -15484 19164 -15356 19196
rect -15324 19164 -15196 19196
rect -15164 19164 -15036 19196
rect -15004 19164 -15000 19196
rect -15520 19160 -15000 19164
rect -1680 19156 -520 19160
rect -1680 19124 -1676 19156
rect -1644 19124 -1516 19156
rect -1484 19124 -1356 19156
rect -1324 19124 -1196 19156
rect -1164 19124 -1036 19156
rect -1004 19124 -876 19156
rect -844 19124 -716 19156
rect -684 19124 -556 19156
rect -524 19124 -520 19156
rect -1680 19120 -520 19124
rect -15520 19116 -15000 19120
rect -15520 19084 -15516 19116
rect -15484 19084 -15356 19116
rect -15324 19084 -15196 19116
rect -15164 19084 -15036 19116
rect -15004 19084 -15000 19116
rect -15520 19080 -15000 19084
rect -1680 19076 -520 19080
rect -1680 19044 -1676 19076
rect -1644 19044 -1516 19076
rect -1484 19044 -1356 19076
rect -1324 19044 -1196 19076
rect -1164 19044 -1036 19076
rect -1004 19044 -876 19076
rect -844 19044 -716 19076
rect -684 19044 -556 19076
rect -524 19044 -520 19076
rect -1680 19040 -520 19044
rect -15520 19036 -15000 19040
rect -15520 19004 -15516 19036
rect -15484 19004 -15356 19036
rect -15324 19004 -15196 19036
rect -15164 19004 -15036 19036
rect -15004 19004 -15000 19036
rect -15520 19000 -15000 19004
rect -1680 18996 -520 19000
rect -1680 18964 -1676 18996
rect -1644 18964 -1516 18996
rect -1484 18964 -1356 18996
rect -1324 18964 -1196 18996
rect -1164 18964 -1036 18996
rect -1004 18964 -876 18996
rect -844 18964 -716 18996
rect -684 18964 -556 18996
rect -524 18964 -520 18996
rect -1680 18960 -520 18964
rect -15520 18956 -15000 18960
rect -15520 18924 -15516 18956
rect -15484 18924 -15356 18956
rect -15324 18924 -15196 18956
rect -15164 18924 -15036 18956
rect -15004 18924 -15000 18956
rect -15520 18920 -15000 18924
rect -1680 18916 -520 18920
rect -1680 18884 -1676 18916
rect -1644 18884 -1516 18916
rect -1484 18884 -1356 18916
rect -1324 18884 -1196 18916
rect -1164 18884 -1036 18916
rect -1004 18884 -876 18916
rect -844 18884 -716 18916
rect -684 18884 -556 18916
rect -524 18884 -520 18916
rect -1680 18880 -520 18884
rect -15520 18876 -15000 18880
rect -15520 18844 -15516 18876
rect -15484 18844 -15356 18876
rect -15324 18844 -15196 18876
rect -15164 18844 -15036 18876
rect -15004 18844 -15000 18876
rect -15520 18840 -15000 18844
rect -1680 18756 -520 18760
rect -1680 18724 -1676 18756
rect -1644 18724 -1516 18756
rect -1484 18724 -1356 18756
rect -1324 18724 -1196 18756
rect -1164 18724 -1036 18756
rect -1004 18724 -876 18756
rect -844 18724 -716 18756
rect -684 18724 -556 18756
rect -524 18724 -520 18756
rect -1680 18720 -520 18724
rect -1680 18676 -520 18680
rect -1680 18644 -1676 18676
rect -1644 18644 -1516 18676
rect -1484 18644 -1356 18676
rect -1324 18644 -1196 18676
rect -1164 18644 -1036 18676
rect -1004 18644 -876 18676
rect -844 18644 -716 18676
rect -684 18644 -556 18676
rect -524 18644 -520 18676
rect -1680 18640 -520 18644
rect -1680 18596 -520 18600
rect -1680 18564 -1676 18596
rect -1644 18564 -1516 18596
rect -1484 18564 -1356 18596
rect -1324 18564 -1196 18596
rect -1164 18564 -1036 18596
rect -1004 18564 -876 18596
rect -844 18564 -716 18596
rect -684 18564 -556 18596
rect -524 18564 -520 18596
rect -1680 18560 -520 18564
rect -15520 18556 -15000 18560
rect -15520 18524 -15516 18556
rect -15484 18524 -15356 18556
rect -15324 18524 -15196 18556
rect -15164 18524 -15036 18556
rect -15004 18524 -15000 18556
rect -15520 18520 -15000 18524
rect -1680 18516 -520 18520
rect -1680 18484 -1676 18516
rect -1644 18484 -1516 18516
rect -1484 18484 -1356 18516
rect -1324 18484 -1196 18516
rect -1164 18484 -1036 18516
rect -1004 18484 -876 18516
rect -844 18484 -716 18516
rect -684 18484 -556 18516
rect -524 18484 -520 18516
rect -1680 18480 -520 18484
rect -15520 18476 -15000 18480
rect -15520 18444 -15516 18476
rect -15484 18444 -15356 18476
rect -15324 18444 -15196 18476
rect -15164 18444 -15036 18476
rect -15004 18444 -15000 18476
rect -15520 18440 -15000 18444
rect -1680 18436 -520 18440
rect -1680 18404 -1676 18436
rect -1644 18404 -1516 18436
rect -1484 18404 -1356 18436
rect -1324 18404 -1196 18436
rect -1164 18404 -1036 18436
rect -1004 18404 -876 18436
rect -844 18404 -716 18436
rect -684 18404 -556 18436
rect -524 18404 -520 18436
rect -1680 18400 -520 18404
rect -15520 18396 -15000 18400
rect -15520 18364 -15516 18396
rect -15484 18364 -15356 18396
rect -15324 18364 -15196 18396
rect -15164 18364 -15036 18396
rect -15004 18364 -15000 18396
rect -15520 18360 -15000 18364
rect -1680 18356 -520 18360
rect -1680 18324 -1676 18356
rect -1644 18324 -1516 18356
rect -1484 18324 -1356 18356
rect -1324 18324 -1196 18356
rect -1164 18324 -1036 18356
rect -1004 18324 -876 18356
rect -844 18324 -716 18356
rect -684 18324 -556 18356
rect -524 18324 -520 18356
rect -1680 18320 -520 18324
rect -15520 18316 -15000 18320
rect -15520 18284 -15516 18316
rect -15484 18284 -15356 18316
rect -15324 18284 -15196 18316
rect -15164 18284 -15036 18316
rect -15004 18284 -15000 18316
rect -15520 18280 -15000 18284
rect -1680 18276 -520 18280
rect -1680 18244 -1676 18276
rect -1644 18244 -1516 18276
rect -1484 18244 -1356 18276
rect -1324 18244 -1196 18276
rect -1164 18244 -1036 18276
rect -1004 18244 -876 18276
rect -844 18244 -716 18276
rect -684 18244 -556 18276
rect -524 18244 -520 18276
rect -1680 18240 -520 18244
rect -15520 18236 -15000 18240
rect -15520 18204 -15516 18236
rect -15484 18204 -15356 18236
rect -15324 18204 -15196 18236
rect -15164 18204 -15036 18236
rect -15004 18204 -15000 18236
rect -15520 18200 -15000 18204
rect -1680 18196 -520 18200
rect -1680 18164 -1676 18196
rect -1644 18164 -1516 18196
rect -1484 18164 -1356 18196
rect -1324 18164 -1196 18196
rect -1164 18164 -1036 18196
rect -1004 18164 -876 18196
rect -844 18164 -716 18196
rect -684 18164 -556 18196
rect -524 18164 -520 18196
rect -1680 18160 -520 18164
rect -15520 18156 -15000 18160
rect -15520 18124 -15516 18156
rect -15484 18124 -15356 18156
rect -15324 18124 -15196 18156
rect -15164 18124 -15036 18156
rect -15004 18124 -15000 18156
rect -15520 18120 -15000 18124
rect -15520 18076 -15000 18080
rect -15520 18044 -15516 18076
rect -15484 18044 -15356 18076
rect -15324 18044 -15196 18076
rect -15164 18044 -15036 18076
rect -15004 18044 -15000 18076
rect -15520 18040 -15000 18044
rect -15520 17996 -15000 18000
rect -15520 17964 -15516 17996
rect -15484 17964 -15356 17996
rect -15324 17964 -15196 17996
rect -15164 17964 -15036 17996
rect -15004 17964 -15000 17996
rect -15520 17960 -15000 17964
rect -15520 17916 -15000 17920
rect -15520 17884 -15516 17916
rect -15484 17884 -15356 17916
rect -15324 17884 -15196 17916
rect -15164 17884 -15036 17916
rect -15004 17884 -15000 17916
rect -15520 17880 -15000 17884
rect -1680 17876 -520 17880
rect -1680 17844 -1676 17876
rect -1644 17844 -1516 17876
rect -1484 17844 -1356 17876
rect -1324 17844 -1196 17876
rect -1164 17844 -1036 17876
rect -1004 17844 -876 17876
rect -844 17844 -716 17876
rect -684 17844 -556 17876
rect -524 17844 -520 17876
rect -1680 17840 -520 17844
rect -15520 17836 -15000 17840
rect -15520 17804 -15516 17836
rect -15484 17804 -15356 17836
rect -15324 17804 -15196 17836
rect -15164 17804 -15036 17836
rect -15004 17804 -15000 17836
rect -15520 17800 -15000 17804
rect -1680 17796 -520 17800
rect -1680 17764 -1676 17796
rect -1644 17764 -1516 17796
rect -1484 17764 -1356 17796
rect -1324 17764 -1196 17796
rect -1164 17764 -1036 17796
rect -1004 17764 -876 17796
rect -844 17764 -716 17796
rect -684 17764 -556 17796
rect -524 17764 -520 17796
rect -1680 17760 -520 17764
rect -15520 17756 -15000 17760
rect -15520 17724 -15516 17756
rect -15484 17724 -15356 17756
rect -15324 17724 -15196 17756
rect -15164 17724 -15036 17756
rect -15004 17724 -15000 17756
rect -15520 17720 -15000 17724
rect -1680 17716 -520 17720
rect -1680 17684 -1676 17716
rect -1644 17684 -1516 17716
rect -1484 17684 -1356 17716
rect -1324 17684 -1196 17716
rect -1164 17684 -1036 17716
rect -1004 17684 -876 17716
rect -844 17684 -716 17716
rect -684 17684 -556 17716
rect -524 17684 -520 17716
rect -1680 17680 -520 17684
rect -15520 17676 -15000 17680
rect -15520 17644 -15516 17676
rect -15484 17644 -15356 17676
rect -15324 17644 -15196 17676
rect -15164 17644 -15036 17676
rect -15004 17644 -15000 17676
rect -15520 17640 -15000 17644
rect -1680 17636 -520 17640
rect -1680 17604 -1676 17636
rect -1644 17604 -1516 17636
rect -1484 17604 -1356 17636
rect -1324 17604 -1196 17636
rect -1164 17604 -1036 17636
rect -1004 17604 -876 17636
rect -844 17604 -716 17636
rect -684 17604 -556 17636
rect -524 17604 -520 17636
rect -1680 17600 -520 17604
rect -15520 17596 -15000 17600
rect -15520 17564 -15516 17596
rect -15484 17564 -15356 17596
rect -15324 17564 -15196 17596
rect -15164 17564 -15036 17596
rect -15004 17564 -15000 17596
rect -15520 17560 -15000 17564
rect -1680 17556 -520 17560
rect -1680 17524 -1676 17556
rect -1644 17524 -1516 17556
rect -1484 17524 -1356 17556
rect -1324 17524 -1196 17556
rect -1164 17524 -1036 17556
rect -1004 17524 -876 17556
rect -844 17524 -716 17556
rect -684 17524 -556 17556
rect -524 17524 -520 17556
rect -1680 17520 -520 17524
rect -15520 17516 -15000 17520
rect -15520 17484 -15516 17516
rect -15484 17484 -15356 17516
rect -15324 17484 -15196 17516
rect -15164 17484 -15036 17516
rect -15004 17484 -15000 17516
rect -15520 17480 -15000 17484
rect -1680 17476 -520 17480
rect -1680 17444 -1676 17476
rect -1644 17444 -1516 17476
rect -1484 17444 -1356 17476
rect -1324 17444 -1196 17476
rect -1164 17444 -1036 17476
rect -1004 17444 -876 17476
rect -844 17444 -716 17476
rect -684 17444 -556 17476
rect -524 17444 -520 17476
rect -1680 17440 -520 17444
rect -15520 17436 -15000 17440
rect -15520 17404 -15516 17436
rect -15484 17404 -15356 17436
rect -15324 17404 -15196 17436
rect -15164 17404 -15036 17436
rect -15004 17404 -15000 17436
rect -15520 17400 -15000 17404
rect -1680 17396 -520 17400
rect -1680 17364 -1676 17396
rect -1644 17364 -1516 17396
rect -1484 17364 -1356 17396
rect -1324 17364 -1196 17396
rect -1164 17364 -1036 17396
rect -1004 17364 -876 17396
rect -844 17364 -716 17396
rect -684 17364 -556 17396
rect -524 17364 -520 17396
rect -1680 17360 -520 17364
rect -1680 17316 -520 17320
rect -1680 17284 -1676 17316
rect -1644 17284 -1516 17316
rect -1484 17284 -1356 17316
rect -1324 17284 -1196 17316
rect -1164 17284 -1036 17316
rect -1004 17284 -876 17316
rect -844 17284 -716 17316
rect -684 17284 -556 17316
rect -524 17284 -520 17316
rect -1680 17280 -520 17284
rect -1680 17236 -520 17240
rect -1680 17204 -1676 17236
rect -1644 17204 -1516 17236
rect -1484 17204 -1356 17236
rect -1324 17204 -1196 17236
rect -1164 17204 -1036 17236
rect -1004 17204 -876 17236
rect -844 17204 -716 17236
rect -684 17204 -556 17236
rect -524 17204 -520 17236
rect -1680 17200 -520 17204
rect -1680 17156 -520 17160
rect -1680 17124 -1676 17156
rect -1644 17124 -1516 17156
rect -1484 17124 -1356 17156
rect -1324 17124 -1196 17156
rect -1164 17124 -1036 17156
rect -1004 17124 -876 17156
rect -844 17124 -716 17156
rect -684 17124 -556 17156
rect -524 17124 -520 17156
rect -1680 17120 -520 17124
rect -15520 17116 -15000 17120
rect -15520 17084 -15516 17116
rect -15484 17084 -15356 17116
rect -15324 17084 -15196 17116
rect -15164 17084 -15036 17116
rect -15004 17084 -15000 17116
rect -15520 17080 -15000 17084
rect -1680 17076 -520 17080
rect -1680 17044 -1676 17076
rect -1644 17044 -1516 17076
rect -1484 17044 -1356 17076
rect -1324 17044 -1196 17076
rect -1164 17044 -1036 17076
rect -1004 17044 -876 17076
rect -844 17044 -716 17076
rect -684 17044 -556 17076
rect -524 17044 -520 17076
rect -1680 17040 -520 17044
rect -15520 17036 -15000 17040
rect -15520 17004 -15516 17036
rect -15484 17004 -15356 17036
rect -15324 17004 -15196 17036
rect -15164 17004 -15036 17036
rect -15004 17004 -15000 17036
rect -15520 17000 -15000 17004
rect -1680 16996 -520 17000
rect -1680 16964 -1676 16996
rect -1644 16964 -1516 16996
rect -1484 16964 -1356 16996
rect -1324 16964 -1196 16996
rect -1164 16964 -1036 16996
rect -1004 16964 -876 16996
rect -844 16964 -716 16996
rect -684 16964 -556 16996
rect -524 16964 -520 16996
rect -1680 16960 -520 16964
rect -15520 16956 -15000 16960
rect -15520 16924 -15516 16956
rect -15484 16924 -15356 16956
rect -15324 16924 -15196 16956
rect -15164 16924 -15036 16956
rect -15004 16924 -15000 16956
rect -15520 16920 -15000 16924
rect -1680 16916 -520 16920
rect -1680 16884 -1676 16916
rect -1644 16884 -1516 16916
rect -1484 16884 -1356 16916
rect -1324 16884 -1196 16916
rect -1164 16884 -1036 16916
rect -1004 16884 -876 16916
rect -844 16884 -716 16916
rect -684 16884 -556 16916
rect -524 16884 -520 16916
rect -1680 16880 -520 16884
rect -15520 16876 -15000 16880
rect -15520 16844 -15516 16876
rect -15484 16844 -15356 16876
rect -15324 16844 -15196 16876
rect -15164 16844 -15036 16876
rect -15004 16844 -15000 16876
rect -15520 16840 -15000 16844
rect -1680 16836 -520 16840
rect -1680 16804 -1676 16836
rect -1644 16804 -1516 16836
rect -1484 16804 -1356 16836
rect -1324 16804 -1196 16836
rect -1164 16804 -1036 16836
rect -1004 16804 -876 16836
rect -844 16804 -716 16836
rect -684 16804 -556 16836
rect -524 16804 -520 16836
rect -1680 16800 -520 16804
rect -15520 16796 -15000 16800
rect -15520 16764 -15516 16796
rect -15484 16764 -15356 16796
rect -15324 16764 -15196 16796
rect -15164 16764 -15036 16796
rect -15004 16764 -15000 16796
rect -15520 16760 -15000 16764
rect -1680 16756 -520 16760
rect -1680 16724 -1676 16756
rect -1644 16724 -1516 16756
rect -1484 16724 -1356 16756
rect -1324 16724 -1196 16756
rect -1164 16724 -1036 16756
rect -1004 16724 -876 16756
rect -844 16724 -716 16756
rect -684 16724 -556 16756
rect -524 16724 -520 16756
rect -1680 16720 -520 16724
rect -15520 16716 -15000 16720
rect -15520 16684 -15516 16716
rect -15484 16684 -15356 16716
rect -15324 16684 -15196 16716
rect -15164 16684 -15036 16716
rect -15004 16684 -15000 16716
rect -15520 16680 -15000 16684
rect -15520 16636 -15000 16640
rect -15520 16604 -15516 16636
rect -15484 16604 -15356 16636
rect -15324 16604 -15196 16636
rect -15164 16604 -15036 16636
rect -15004 16604 -15000 16636
rect -15520 16600 -15000 16604
rect -1680 16636 -520 16640
rect -1680 16604 -1676 16636
rect -1644 16604 -1516 16636
rect -1484 16604 -1356 16636
rect -1324 16604 -1196 16636
rect -1164 16604 -1036 16636
rect -1004 16604 -876 16636
rect -844 16604 -716 16636
rect -684 16604 -556 16636
rect -524 16604 -520 16636
rect -1680 16600 -520 16604
rect -15520 16556 -15000 16560
rect -15520 16524 -15516 16556
rect -15484 16524 -15356 16556
rect -15324 16524 -15196 16556
rect -15164 16524 -15036 16556
rect -15004 16524 -15000 16556
rect -15520 16520 -15000 16524
rect -1680 16556 -520 16560
rect -1680 16524 -1676 16556
rect -1644 16524 -1516 16556
rect -1484 16524 -1356 16556
rect -1324 16524 -1196 16556
rect -1164 16524 -1036 16556
rect -1004 16524 -876 16556
rect -844 16524 -716 16556
rect -684 16524 -556 16556
rect -524 16524 -520 16556
rect -1680 16520 -520 16524
rect -15520 16476 -15000 16480
rect -15520 16444 -15516 16476
rect -15484 16444 -15356 16476
rect -15324 16444 -15196 16476
rect -15164 16444 -15036 16476
rect -15004 16444 -15000 16476
rect -15520 16440 -15000 16444
rect -16160 360 -15520 400
rect -16160 240 -16120 360
rect -16000 240 -15520 360
rect -16160 200 -15520 240
rect -520 200 -480 400
rect 20480 360 21200 400
rect 20480 240 21040 360
rect 21160 240 21200 360
rect 20480 200 21200 240
rect -15760 120 -15520 160
rect -15760 0 -15720 120
rect -15600 0 -15520 120
rect -15760 -40 -15520 0
rect -520 -40 -480 160
rect 20480 120 20800 160
rect 20480 0 20640 120
rect 20760 0 20800 120
rect 20480 -40 20800 0
rect -16560 -1480 21600 -1440
rect -16560 -1600 -15720 -1480
rect -15600 -1600 20640 -1480
rect 20760 -1600 21600 -1480
rect -16560 -1640 21600 -1600
rect -16560 -1720 21600 -1680
rect -16560 -1840 -16120 -1720
rect -16000 -1840 21040 -1720
rect 21160 -1840 21600 -1720
rect -16560 -1880 21600 -1840
rect -16560 -1960 21600 -1920
rect -16560 -2080 -16520 -1960
rect -16400 -2080 21440 -1960
rect 21560 -2080 21600 -1960
rect -16560 -2120 21600 -2080
<< via4 >>
rect -16520 39360 -16400 39480
rect 21440 39360 21560 39480
rect -16120 39120 -16000 39240
rect 21040 39120 21160 39240
rect -15720 38880 -15600 39000
rect 20640 38880 20760 39000
rect -15720 37280 -15600 37400
rect 20640 37280 20760 37400
rect -16120 37040 -16000 37160
rect 21040 37040 21160 37160
rect 21440 36560 21560 36680
rect -16120 240 -16000 360
rect 21040 240 21160 360
rect -15720 0 -15600 120
rect 20640 0 20760 120
rect -15720 -1600 -15600 -1480
rect 20640 -1600 20760 -1480
rect -16120 -1840 -16000 -1720
rect 21040 -1840 21160 -1720
rect -16520 -2080 -16400 -1960
rect 21440 -2080 21560 -1960
<< metal5 >>
rect -16560 39480 -16360 39560
rect -16560 39360 -16520 39480
rect -16400 39360 -16360 39480
rect -16560 -1960 -16360 39360
rect -16560 -2080 -16520 -1960
rect -16400 -2080 -16360 -1960
rect -16560 -2120 -16360 -2080
rect -16160 39240 -15960 39560
rect -16160 39120 -16120 39240
rect -16000 39120 -15960 39240
rect -16160 37160 -15960 39120
rect -16160 37040 -16120 37160
rect -16000 37040 -15960 37160
rect -16160 360 -15960 37040
rect -16160 240 -16120 360
rect -16000 240 -15960 360
rect -16160 -1720 -15960 240
rect -16160 -1840 -16120 -1720
rect -16000 -1840 -15960 -1720
rect -16160 -2120 -15960 -1840
rect -15760 39000 -15560 39560
rect -15760 38880 -15720 39000
rect -15600 38880 -15560 39000
rect -15760 37400 -15560 38880
rect 20600 39000 20800 39520
rect 20600 38880 20640 39000
rect 20760 38880 20800 39000
rect -400 37440 -200 37680
rect 3440 37440 3640 37680
rect 5840 37440 6040 37680
rect -15760 37280 -15720 37400
rect -15600 37280 -15560 37400
rect -15760 120 -15560 37280
rect -15760 0 -15720 120
rect -15600 0 -15560 120
rect -15760 -1480 -15560 0
rect -15760 -1600 -15720 -1480
rect -15600 -1600 -15560 -1480
rect -15760 -2120 -15560 -1600
rect 20600 37400 20800 38880
rect 20600 37280 20640 37400
rect 20760 37280 20800 37400
rect 20600 120 20800 37280
rect 20600 0 20640 120
rect 20760 0 20800 120
rect 20600 -1480 20800 0
rect 20600 -1600 20640 -1480
rect 20760 -1600 20800 -1480
rect 20600 -2120 20800 -1600
rect 21000 39240 21200 39520
rect 21000 39120 21040 39240
rect 21160 39120 21200 39240
rect 21000 37160 21200 39120
rect 21000 37040 21040 37160
rect 21160 37040 21200 37160
rect 21000 360 21200 37040
rect 21000 240 21040 360
rect 21160 240 21200 360
rect 21000 -1720 21200 240
rect 21000 -1840 21040 -1720
rect 21160 -1840 21200 -1720
rect 21000 -2120 21200 -1840
rect 21400 39480 21600 39520
rect 21400 39360 21440 39480
rect 21560 39360 21600 39480
rect 21400 36680 21600 39360
rect 21400 36560 21440 36680
rect 21560 36560 21600 36680
rect 21400 -1960 21600 36560
rect 21400 -2080 21440 -1960
rect 21560 -2080 21600 -1960
rect 21400 -2120 21600 -2080
use pseudo  pseudo ../../pseudo/mag
timestamp 1638398147
transform 1 0 -8400 0 1 17800
box -280 -360 6560 2160
use ota  ota ../../ota/mag
timestamp 1638390070
transform 1 0 -480 0 1 2000
box 0 -3400 20960 36800
use cap1_10  cap1 ../../cap1_10/mag
timestamp 1638390070
transform -1 0 -520 0 -1 37440
box 0 0 15000 15960
use cap1_10  cap2
timestamp 1638390070
transform 1 0 -15520 0 1 -40
box 0 0 15000 15960
<< labels >>
rlabel metal2 -640 20240 -600 20280 1 q
rlabel metal2 -640 19920 -600 19960 0 op
rlabel metal2 -640 20080 -600 20120 0 xm
rlabel metal2 -16640 18760 -16600 18800 0 ip
port 0 nsew
rlabel metal2 -16640 18600 -16600 18640 0 im
port 1 nsew
rlabel metal2 21640 19920 21680 19960 1 op
port 2 nsew
rlabel metal2 21640 17920 21680 17960 0 om
port 3 nsew
rlabel metal2 -16640 20560 -16600 20600 0 ib
port 5 nsew
rlabel metal2 -640 17920 -600 17960 0 om
rlabel metal2 -640 18080 -600 18120 0 xp
rlabel metal2 -16640 17240 -16600 17280 1 fsb
port 4 nsew
rlabel metal5 -16560 39520 -16360 39560 1 vdda
port 7 nsew
rlabel metal5 -16160 39520 -15960 39560 0 gnda
port 8 nsew
rlabel metal5 -15760 39520 -15560 39560 0 vssa
port 9 nsew
rlabel metal2 21640 20560 21680 20600 0 ib
port 5 nsew
<< end >>
