magic
tech sky130A
timestamp 1634489271
<< nwell >>
rect -1600 1100 1030 1220
rect -2555 -135 -990 -30
<< poly >>
rect -170 1160 -125 1195
rect -45 1160 0 1195
rect 90 1160 135 1195
<< metal1 >>
rect -2880 -165 -2700 1645
rect -2555 -55 -2375 1640
rect -2270 1195 -2080 1640
rect 810 1540 1070 1650
rect -1690 1230 1280 1540
rect -2270 1180 -1495 1195
rect -2270 1130 -1565 1180
rect -1515 1130 -1495 1180
rect -2270 1110 -1495 1130
rect -2270 905 -1590 1110
rect -1435 820 -1340 1230
rect -1095 1190 -1010 1200
rect -1095 1160 -1075 1190
rect -1080 1155 -1075 1160
rect -1030 1160 -1010 1190
rect -1030 1155 -1025 1160
rect -1080 1150 -1025 1155
rect -860 1150 -710 1230
rect -488 1195 174 1199
rect -488 1165 -420 1195
rect -435 1160 -420 1165
rect -375 1165 -305 1195
rect -375 1160 -350 1165
rect -435 1155 -350 1160
rect -320 1160 -305 1165
rect -260 1165 -170 1195
rect -260 1160 -235 1165
rect -320 1150 -235 1160
rect -180 1160 -170 1165
rect -125 1165 -45 1195
rect -125 1160 -95 1165
rect -180 1150 -95 1160
rect -65 1160 -45 1165
rect 0 1165 90 1195
rect 0 1160 20 1165
rect -65 1150 20 1160
rect 80 1160 90 1165
rect 135 1165 174 1195
rect 135 1160 165 1165
rect 80 1150 165 1160
rect -995 905 -710 1150
rect 230 1090 410 1230
rect 900 1190 980 1195
rect 900 1155 915 1190
rect 960 1155 980 1190
rect 900 1140 980 1155
rect -480 905 410 1090
rect 590 910 895 1115
rect -1495 575 -1340 820
rect -1290 570 -1105 815
rect -350 570 430 820
rect -1290 430 -1160 570
rect -1820 300 -770 430
rect -1820 225 -1670 300
rect -1820 90 -1600 225
rect -900 220 -770 300
rect -1005 90 -770 220
rect 240 125 430 570
rect -485 90 430 125
rect -2555 -115 -2525 -55
rect -2390 -115 -2375 -55
rect -1505 -60 -1330 65
rect -2555 -135 -2375 -115
rect -1600 -165 -1500 -80
rect -2880 -255 -1500 -165
rect -1460 -280 -1330 -60
rect -1785 -410 -1330 -280
rect -1290 -55 -1105 65
rect -485 -30 265 90
rect 380 -30 430 90
rect -1290 -280 -1160 -55
rect -1085 -60 -1005 -45
rect -485 -60 430 -30
rect -1085 -95 -1070 -60
rect -1025 -95 -1005 -60
rect -1085 -110 -1005 -95
rect -350 -265 50 -115
rect -1290 -290 -435 -280
rect -1290 -315 -220 -290
rect -1290 -375 -835 -315
rect -750 -340 -220 -315
rect -750 -375 -705 -340
rect -120 -375 50 -265
rect -1290 -410 -705 -375
rect -1785 -560 -1655 -410
rect -1610 -460 -1330 -410
rect -1610 -540 -1005 -460
rect -940 -560 -810 -410
rect -1785 -645 -1610 -560
rect -1510 -645 -1100 -560
rect -1000 -645 -810 -560
rect -1450 -700 -1185 -645
rect -550 -700 50 -375
rect 240 -445 430 -60
rect 590 410 790 910
rect 1080 815 1280 1230
rect 975 580 1280 815
rect 590 250 1350 410
rect 590 240 1060 250
rect 590 160 790 240
rect 590 -80 900 160
rect 990 -175 1250 -170
rect 985 -420 1250 -175
rect 885 -445 1005 -440
rect 240 -600 1005 -445
rect 1100 -700 1250 -420
rect -1710 -930 1390 -700
<< via1 >>
rect -1565 1130 -1515 1180
rect -1075 1155 -1030 1190
rect -420 1160 -375 1195
rect -305 1160 -260 1195
rect -170 1160 -125 1195
rect -45 1160 0 1195
rect 90 1160 135 1195
rect 915 1155 960 1190
rect -2525 -115 -2390 -55
rect 265 -30 380 90
rect -1070 -95 -1025 -60
rect -835 -375 -750 -315
<< metal2 >>
rect -1600 1195 1030 1220
rect -1600 1190 -420 1195
rect -1600 1180 -1075 1190
rect -1600 1130 -1565 1180
rect -1515 1155 -1075 1180
rect -1030 1160 -420 1190
rect -375 1160 -305 1195
rect -260 1160 -170 1195
rect -125 1160 -45 1195
rect 0 1160 90 1195
rect 135 1190 1030 1195
rect 135 1160 915 1190
rect -1030 1155 915 1160
rect 960 1155 1030 1190
rect -1515 1130 1030 1155
rect -1600 1100 1030 1130
rect 210 90 1435 125
rect 210 -30 265 90
rect 380 -30 1435 90
rect -2555 -55 -990 -30
rect -2555 -115 -2525 -55
rect -2390 -60 -990 -55
rect 210 -60 1435 -30
rect -2390 -95 -1070 -60
rect -1025 -95 -990 -60
rect -2390 -115 -990 -95
rect -2555 -135 -990 -115
rect -855 -315 -715 -280
rect -855 -375 -835 -315
rect -750 -375 -715 -315
rect -855 -1005 -715 -375
rect -1020 -1055 -550 -1005
rect -1020 -1140 -950 -1055
rect -630 -1140 -550 -1055
rect -1020 -1400 -550 -1140
rect 1250 -1295 1435 -60
rect 1250 -1585 1300 -1295
rect 1385 -1585 1435 -1295
rect 1250 -1655 1435 -1585
<< via2 >>
rect -950 -1140 -630 -1055
rect 1300 -1585 1385 -1295
<< metal3 >>
rect -1020 -1055 -550 -1005
rect -1020 -1140 -950 -1055
rect -630 -1140 -550 -1055
rect -1020 -1400 -550 -1140
rect 1250 -1295 1435 -1285
rect 1250 -1585 1300 -1295
rect 1385 -1585 1435 -1295
rect 1250 -1655 1435 -1585
<< via3 >>
rect 1300 -1585 1385 -1295
<< metal4 >>
rect 935 -1295 1435 -1280
rect 935 -1585 1300 -1295
rect 1385 -1585 1435 -1295
rect 935 -1655 1435 -1585
<< labels >>
flabel metal1 -2830 1540 -2730 1640 0 FreeSans 128 0 0 0 in1
port 3 nsew
flabel metal1 -2520 1540 -2420 1640 0 FreeSans 128 0 0 0 in2
port 4 nsew
flabel metal1 -2230 1540 -2130 1640 0 FreeSans 128 0 0 0 ib
port 2 nsew
flabel metal1 890 1550 990 1650 0 FreeSans 128 0 0 0 vd
port 0 nsew
flabel metal1 1250 290 1350 390 0 FreeSans 128 0 0 0 out
port 5 nsew
flabel metal1 1260 -860 1360 -760 0 FreeSans 128 0 0 0 vs
port 1 nsew
<< end >>
