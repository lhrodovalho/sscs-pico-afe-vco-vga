* OpAmp open-loop dc testbench

* Include SkyWater sky130 device models
.lib "/usr/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice" tt
.param mc_mm_switch=0
.include "../mag/opamp_core.spice"

* supply voltages
vdda  vdda 0 1.0
vssa  vssa 0 0.0
egnda gnda vssa vdda vssa 0.5

* input signals
vin in gnda dc 0 ac 1
eip ip gnda in gnda  1.0
eim im gnda in gnda  0.0

* DUT
x0 im ip out ib q vdda bp vddx gnda vssa xn xp x y z opamp_core
ib vdda ib 2n
cl out gnda 10p
ll out gnda 1T

.option gmin=1e-12
.control

	op
	print ib i(vdda)

	ac dec 10 1m 1Meg
	plot vdb(out)
	plot cphase(out)*180/PI
	
*	noise v(out) vin dec 10 1 100
*	print inoise_total onoise_total

.endc

.end
