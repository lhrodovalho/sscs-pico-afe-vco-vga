magic
tech sky130A
magscale 1 2
timestamp 1634487483
<< nwell >>
rect -812 -805 812 805
<< pmos >>
rect -616 -586 -416 586
rect -358 -586 -158 586
rect -100 -586 100 586
rect 158 -586 358 586
rect 416 -586 616 586
<< pdiff >>
rect -674 574 -616 586
rect -674 -574 -662 574
rect -628 -574 -616 574
rect -674 -586 -616 -574
rect -416 574 -358 586
rect -416 -574 -404 574
rect -370 -574 -358 574
rect -416 -586 -358 -574
rect -158 574 -100 586
rect -158 -574 -146 574
rect -112 -574 -100 574
rect -158 -586 -100 -574
rect 100 574 158 586
rect 100 -574 112 574
rect 146 -574 158 574
rect 100 -586 158 -574
rect 358 574 416 586
rect 358 -574 370 574
rect 404 -574 416 574
rect 358 -586 416 -574
rect 616 574 674 586
rect 616 -574 628 574
rect 662 -574 674 574
rect 616 -586 674 -574
<< pdiffc >>
rect -662 -574 -628 574
rect -404 -574 -370 574
rect -146 -574 -112 574
rect 112 -574 146 574
rect 370 -574 404 574
rect 628 -574 662 574
<< nsubdiff >>
rect -776 735 -680 769
rect 680 735 776 769
rect -776 673 -742 735
rect 742 673 776 735
rect -776 -735 -742 -673
rect 742 -735 776 -673
rect -776 -769 -680 -735
rect 680 -769 776 -735
<< nsubdiffcont >>
rect -680 735 680 769
rect -776 -673 -742 673
rect 742 -673 776 673
rect -680 -769 680 -735
<< poly >>
rect -616 667 -416 683
rect -616 633 -600 667
rect -432 633 -416 667
rect -616 586 -416 633
rect -358 667 -158 683
rect -358 633 -342 667
rect -174 633 -158 667
rect -358 586 -158 633
rect -100 667 100 683
rect -100 633 -84 667
rect 84 633 100 667
rect -100 586 100 633
rect 158 667 358 683
rect 158 633 174 667
rect 342 633 358 667
rect 158 586 358 633
rect 416 667 616 683
rect 416 633 432 667
rect 600 633 616 667
rect 416 586 616 633
rect -616 -633 -416 -586
rect -616 -667 -600 -633
rect -432 -667 -416 -633
rect -616 -683 -416 -667
rect -358 -633 -158 -586
rect -358 -667 -342 -633
rect -174 -667 -158 -633
rect -358 -683 -158 -667
rect -100 -633 100 -586
rect -100 -667 -84 -633
rect 84 -667 100 -633
rect -100 -683 100 -667
rect 158 -633 358 -586
rect 158 -667 174 -633
rect 342 -667 358 -633
rect 158 -683 358 -667
rect 416 -633 616 -586
rect 416 -667 432 -633
rect 600 -667 616 -633
rect 416 -683 616 -667
<< polycont >>
rect -600 633 -432 667
rect -342 633 -174 667
rect -84 633 84 667
rect 174 633 342 667
rect 432 633 600 667
rect -600 -667 -432 -633
rect -342 -667 -174 -633
rect -84 -667 84 -633
rect 174 -667 342 -633
rect 432 -667 600 -633
<< locali >>
rect -776 735 -680 769
rect 680 735 776 769
rect -776 673 -742 735
rect 742 673 776 735
rect -616 633 -600 667
rect -432 633 -416 667
rect -358 633 -342 667
rect -174 633 -158 667
rect -100 633 -84 667
rect 84 633 100 667
rect 158 633 174 667
rect 342 633 358 667
rect 416 633 432 667
rect 600 633 616 667
rect -662 574 -628 590
rect -662 -590 -628 -574
rect -404 574 -370 590
rect -404 -590 -370 -574
rect -146 574 -112 590
rect -146 -590 -112 -574
rect 112 574 146 590
rect 112 -590 146 -574
rect 370 574 404 590
rect 370 -590 404 -574
rect 628 574 662 590
rect 628 -590 662 -574
rect -616 -667 -600 -633
rect -432 -667 -416 -633
rect -358 -667 -342 -633
rect -174 -667 -158 -633
rect -100 -667 -84 -633
rect 84 -667 100 -633
rect 158 -667 174 -633
rect 342 -667 358 -633
rect 416 -667 432 -633
rect 600 -667 616 -633
rect -776 -735 -742 -673
rect 742 -735 776 -673
rect -776 -769 -680 -735
rect 680 -769 776 -735
<< viali >>
rect -600 633 -432 667
rect -342 633 -174 667
rect -84 633 84 667
rect 174 633 342 667
rect 432 633 600 667
rect -662 -574 -628 574
rect -404 -574 -370 574
rect -146 -574 -112 574
rect 112 -574 146 574
rect 370 -574 404 574
rect 628 -574 662 574
rect -600 -667 -432 -633
rect -342 -667 -174 -633
rect -84 -667 84 -633
rect 174 -667 342 -633
rect 432 -667 600 -633
<< metal1 >>
rect -612 667 -420 673
rect -612 633 -600 667
rect -432 633 -420 667
rect -612 627 -420 633
rect -354 667 -162 673
rect -354 633 -342 667
rect -174 633 -162 667
rect -354 627 -162 633
rect -96 667 96 673
rect -96 633 -84 667
rect 84 633 96 667
rect -96 627 96 633
rect 162 667 354 673
rect 162 633 174 667
rect 342 633 354 667
rect 162 627 354 633
rect 420 667 612 673
rect 420 633 432 667
rect 600 633 612 667
rect 420 627 612 633
rect -668 574 -622 586
rect -668 -574 -662 574
rect -628 -574 -622 574
rect -668 -586 -622 -574
rect -410 574 -364 586
rect -410 -574 -404 574
rect -370 -574 -364 574
rect -410 -586 -364 -574
rect -152 574 -106 586
rect -152 -574 -146 574
rect -112 -574 -106 574
rect -152 -586 -106 -574
rect 106 574 152 586
rect 106 -574 112 574
rect 146 -574 152 574
rect 106 -586 152 -574
rect 364 574 410 586
rect 364 -574 370 574
rect 404 -574 410 574
rect 364 -586 410 -574
rect 622 574 668 586
rect 622 -574 628 574
rect 662 -574 668 574
rect 622 -586 668 -574
rect -612 -633 -420 -627
rect -612 -667 -600 -633
rect -432 -667 -420 -633
rect -612 -673 -420 -667
rect -354 -633 -162 -627
rect -354 -667 -342 -633
rect -174 -667 -162 -633
rect -354 -673 -162 -667
rect -96 -633 96 -627
rect -96 -667 -84 -633
rect 84 -667 96 -633
rect -96 -673 96 -667
rect 162 -633 354 -627
rect 162 -667 174 -633
rect 342 -667 354 -633
rect 162 -673 354 -667
rect 420 -633 612 -627
rect 420 -667 432 -633
rect 600 -667 612 -633
rect 420 -673 612 -667
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -759 -752 759 752
string parameters w 5.86 l 1.0 m 1 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagt 0 viagr 0 viagl 0
string library sky130
<< end >>
