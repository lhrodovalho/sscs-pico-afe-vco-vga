* NGSPICE file created from opamp_pair.ext - technology: sky130A

.subckt invt in out xpb xn xpa vddx bp gnda vssa
X0 xpa bp pa1 xpa sky130_fd_pr__pfet_01v8_lvt ad=2.4e+12p pd=4.6e+06u as=2.4e+12p ps=4.6e+06u w=3e+06u l=8e+06u
X1 vddx bp xpa xpa sky130_fd_pr__pfet_01v8_lvt ad=2.85e+12p pd=7.15e+06u as=2.4e+12p ps=4.6e+06u w=3e+06u l=8e+06u
X2 n2 in xn vssa sky130_fd_pr__nfet_01v8 ad=8e+11p pd=2.6e+06u as=8e+11p ps=2.6e+06u w=1e+06u l=8e+06u
X3 xn in n1 vssa sky130_fd_pr__nfet_01v8 ad=8e+11p pd=2.6e+06u as=8e+11p ps=2.6e+06u w=1e+06u l=8e+06u
X4 pa2 bp xpa xpa sky130_fd_pr__pfet_01v8_lvt ad=2.4e+12p pd=4.6e+06u as=2.4e+12p ps=4.6e+06u w=3e+06u l=8e+06u
X5 pb1 in vddx vddx sky130_fd_pr__pfet_01v8_lvt ad=2.4e+12p pd=4.6e+06u as=2.85e+12p ps=7.15e+06u w=3e+06u l=8e+06u
X6 xn in out vssa sky130_fd_pr__nfet_01v8 ad=8e+11p pd=2.6e+06u as=9e+11p ps=3.3e+06u w=1e+06u l=8e+06u
X7 vddx bp pa2 xpa sky130_fd_pr__pfet_01v8_lvt ad=2.85e+12p pd=7.15e+06u as=2.4e+12p ps=4.6e+06u w=3e+06u l=8e+06u
X8 xpb in out vddx sky130_fd_pr__pfet_01v8_lvt ad=2.4e+12p pd=4.6e+06u as=2.7e+12p ps=6.3e+06u w=3e+06u l=8e+06u
X9 xpb in pb1 vddx sky130_fd_pr__pfet_01v8_lvt ad=2.4e+12p pd=4.6e+06u as=2.4e+12p ps=4.6e+06u w=3e+06u l=8e+06u
X10 out in xpb vddx sky130_fd_pr__pfet_01v8_lvt ad=2.7e+12p pd=6.3e+06u as=2.4e+12p ps=4.6e+06u w=3e+06u l=8e+06u
X11 n1 in vssa vssa sky130_fd_pr__nfet_01v8 ad=8e+11p pd=2.6e+06u as=1e+12p ps=4e+06u w=1e+06u l=8e+06u
X12 pb2 in xpb vddx sky130_fd_pr__pfet_01v8_lvt ad=2.4e+12p pd=4.6e+06u as=2.4e+12p ps=4.6e+06u w=3e+06u l=8e+06u
X13 xpb in out vddx sky130_fd_pr__pfet_01v8_lvt ad=2.4e+12p pd=4.6e+06u as=2.7e+12p ps=6.3e+06u w=3e+06u l=8e+06u
X14 xpa bp vddx xpa sky130_fd_pr__pfet_01v8_lvt ad=2.4e+12p pd=4.6e+06u as=2.85e+12p ps=7.15e+06u w=3e+06u l=8e+06u
X15 vddx in pb2 vddx sky130_fd_pr__pfet_01v8_lvt ad=2.85e+12p pd=7.15e+06u as=2.4e+12p ps=4.6e+06u w=3e+06u l=8e+06u
X16 out in xpb vddx sky130_fd_pr__pfet_01v8_lvt ad=2.7e+12p pd=6.3e+06u as=2.4e+12p ps=4.6e+06u w=3e+06u l=8e+06u
X17 out in xn vssa sky130_fd_pr__nfet_01v8 ad=9e+11p pd=3.3e+06u as=8e+11p ps=2.6e+06u w=1e+06u l=8e+06u
X18 vddx bp xpa xpa sky130_fd_pr__pfet_01v8_lvt ad=2.85e+12p pd=7.15e+06u as=2.4e+12p ps=4.6e+06u w=3e+06u l=8e+06u
X19 xn in out vssa sky130_fd_pr__nfet_01v8 ad=8e+11p pd=2.6e+06u as=9e+11p ps=3.3e+06u w=1e+06u l=8e+06u
X20 pa1 bp vddx xpa sky130_fd_pr__pfet_01v8_lvt ad=2.4e+12p pd=4.6e+06u as=2.85e+12p ps=7.15e+06u w=3e+06u l=8e+06u
X21 xpa bp vddx xpa sky130_fd_pr__pfet_01v8_lvt ad=2.4e+12p pd=4.6e+06u as=2.85e+12p ps=7.15e+06u w=3e+06u l=8e+06u
X22 vssa in n2 vssa sky130_fd_pr__nfet_01v8 ad=1e+12p pd=4e+06u as=8e+11p ps=2.6e+06u w=1e+06u l=8e+06u
X23 out in xn vssa sky130_fd_pr__nfet_01v8 ad=9e+11p pd=3.3e+06u as=8e+11p ps=2.6e+06u w=1e+06u l=8e+06u
.ends

.subckt inv_2_2 in out vdda bp vddx gnda vssa
X0 pb1 in vddx vddx sky130_fd_pr__pfet_01v8_lvt ad=2.4e+12p pd=4.6e+06u as=3e+12p ps=8e+06u w=3e+06u l=8e+06u
X1 n2 in out vssa sky130_fd_pr__nfet_01v8 ad=8e+11p pd=2.6e+06u as=8e+11p ps=2.6e+06u w=1e+06u l=8e+06u
X2 out in pb1 vddx sky130_fd_pr__pfet_01v8_lvt ad=2.4e+12p pd=4.6e+06u as=2.4e+12p ps=4.6e+06u w=3e+06u l=8e+06u
X3 out in n1 vssa sky130_fd_pr__nfet_01v8 ad=8e+11p pd=2.6e+06u as=8e+11p ps=2.6e+06u w=1e+06u l=8e+06u
X4 pa1 bp vddx vdda sky130_fd_pr__pfet_01v8_lvt ad=2.4e+12p pd=4.6e+06u as=3e+12p ps=8e+06u w=3e+06u l=8e+06u
X5 vdda bp pa1 vdda sky130_fd_pr__pfet_01v8_lvt ad=2.4e+12p pd=4.6e+06u as=2.4e+12p ps=4.6e+06u w=3e+06u l=8e+06u
X6 pb2 in out vddx sky130_fd_pr__pfet_01v8_lvt ad=2.4e+12p pd=4.6e+06u as=2.4e+12p ps=4.6e+06u w=3e+06u l=8e+06u
X7 vddx in pb2 vddx sky130_fd_pr__pfet_01v8_lvt ad=3e+12p pd=8e+06u as=2.4e+12p ps=4.6e+06u w=3e+06u l=8e+06u
X8 pa2 bp vdda vdda sky130_fd_pr__pfet_01v8_lvt ad=2.4e+12p pd=4.6e+06u as=2.4e+12p ps=4.6e+06u w=3e+06u l=8e+06u
X9 n1 in vssa vssa sky130_fd_pr__nfet_01v8 ad=8e+11p pd=2.6e+06u as=1e+12p ps=4e+06u w=1e+06u l=8e+06u
X10 vddx bp pa2 vdda sky130_fd_pr__pfet_01v8_lvt ad=3e+12p pd=8e+06u as=2.4e+12p ps=4.6e+06u w=3e+06u l=8e+06u
X11 vssa in n2 vssa sky130_fd_pr__nfet_01v8 ad=1e+12p pd=4e+06u as=8e+11p ps=2.6e+06u w=1e+06u l=8e+06u
.ends

.subckt inv_bias bpa bpb gnda na nb qa qb vdda vddx vssa xa xb
X0 qa6 qa vddx vddx sky130_fd_pr__pfet_01v8_lvt ad=2.4e+12p pd=4.6e+06u as=3e+12p ps=8e+06u w=3e+06u l=8e+06u
X1 qa3 qa qa2 vssa sky130_fd_pr__nfet_01v8 ad=8e+11p pd=2.6e+06u as=8e+11p ps=2.6e+06u w=1e+06u l=8e+06u
X2 qb2 qb qb1 vssa sky130_fd_pr__nfet_01v8 ad=8e+11p pd=2.6e+06u as=8e+11p ps=2.6e+06u w=1e+06u l=8e+06u
X3 qb1 qb vssa vssa sky130_fd_pr__nfet_01v8 ad=8e+11p pd=2.6e+06u as=1e+12p ps=4e+06u w=1e+06u l=8e+06u
X4 qa5 qa qa6 vddx sky130_fd_pr__pfet_01v8_lvt ad=2.4e+12p pd=4.6e+06u as=2.4e+12p ps=4.6e+06u w=3e+06u l=8e+06u
X5 qa2 qa qa1 vssa sky130_fd_pr__nfet_01v8 ad=8e+11p pd=2.6e+06u as=8e+11p ps=2.6e+06u w=1e+06u l=8e+06u
X6 bpa3 bpa vddx vdda sky130_fd_pr__pfet_01v8_lvt ad=2.4e+12p pd=4.6e+06u as=3e+12p ps=8e+06u w=3e+06u l=8e+06u
X7 nb2 nb nb1 vssa sky130_fd_pr__nfet_01v8 ad=8e+11p pd=2.6e+06u as=8e+11p ps=2.6e+06u w=1e+06u l=8e+06u
X8 na2 na na1 vssa sky130_fd_pr__nfet_01v8 ad=8e+11p pd=2.6e+06u as=8e+11p ps=2.6e+06u w=1e+06u l=8e+06u
X9 xb1 xb vdda vdda sky130_fd_pr__pfet_01v8_lvt ad=2.4e+12p pd=4.6e+06u as=3e+12p ps=8e+06u w=3e+06u l=8e+06u
X10 nb1 nb vssa vssa sky130_fd_pr__nfet_01v8 ad=8e+11p pd=2.6e+06u as=1e+12p ps=4e+06u w=1e+06u l=8e+06u
X11 na1 na vssa vssa sky130_fd_pr__nfet_01v8 ad=8e+11p pd=2.6e+06u as=1e+12p ps=4e+06u w=1e+06u l=8e+06u
X12 bpa2 bpa bpa3 vdda sky130_fd_pr__pfet_01v8_lvt ad=2.4e+12p pd=4.6e+06u as=2.4e+12p ps=4.6e+06u w=3e+06u l=8e+06u
X13 qa4 qa qa5 vddx sky130_fd_pr__pfet_01v8_lvt ad=2.4e+12p pd=4.6e+06u as=2.4e+12p ps=4.6e+06u w=3e+06u l=8e+06u
X14 xb2 xb xb1 vdda sky130_fd_pr__pfet_01v8_lvt ad=2.4e+12p pd=4.6e+06u as=2.4e+12p ps=4.6e+06u w=3e+06u l=8e+06u
X15 xb qb qb3 vssa sky130_fd_pr__nfet_01v8 ad=1e+12p pd=4e+06u as=8e+11p ps=2.6e+06u w=1e+06u l=8e+06u
X16 qa qa qa4 vddx sky130_fd_pr__pfet_01v8_lvt ad=3e+12p pd=8e+06u as=2.4e+12p ps=4.6e+06u w=3e+06u l=8e+06u
X17 bpa1 bpa bpa2 vdda sky130_fd_pr__pfet_01v8_lvt ad=2.4e+12p pd=4.6e+06u as=2.4e+12p ps=4.6e+06u w=3e+06u l=8e+06u
X18 qa1 qa vssa vssa sky130_fd_pr__nfet_01v8 ad=8e+11p pd=2.6e+06u as=1e+12p ps=4e+06u w=1e+06u l=8e+06u
X19 bpb nb nb3 vssa sky130_fd_pr__nfet_01v8 ad=1e+12p pd=4e+06u as=8e+11p ps=2.6e+06u w=1e+06u l=8e+06u
X20 xa1 xa vdda vdda sky130_fd_pr__pfet_01v8_lvt ad=2.4e+12p pd=4.6e+06u as=3e+12p ps=8e+06u w=3e+06u l=8e+06u
X21 na na na3 vssa sky130_fd_pr__nfet_01v8 ad=1e+12p pd=4e+06u as=8e+11p ps=2.6e+06u w=1e+06u l=8e+06u
X22 xb3 xb xb2 vdda sky130_fd_pr__pfet_01v8_lvt ad=2.4e+12p pd=4.6e+06u as=2.4e+12p ps=4.6e+06u w=3e+06u l=8e+06u
X23 vdda bpa bpa1 vdda sky130_fd_pr__pfet_01v8_lvt ad=3e+12p pd=8e+06u as=2.4e+12p ps=4.6e+06u w=3e+06u l=8e+06u
X24 xa2 xa xa1 vdda sky130_fd_pr__pfet_01v8_lvt ad=2.4e+12p pd=4.6e+06u as=2.4e+12p ps=4.6e+06u w=3e+06u l=8e+06u
X25 xb xb xb3 vdda sky130_fd_pr__pfet_01v8_lvt ad=3e+12p pd=8e+06u as=2.4e+12p ps=4.6e+06u w=3e+06u l=8e+06u
X26 qb3 qb qb2 vssa sky130_fd_pr__nfet_01v8 ad=8e+11p pd=2.6e+06u as=8e+11p ps=2.6e+06u w=1e+06u l=8e+06u
X27 xa3 xa xa2 vdda sky130_fd_pr__pfet_01v8_lvt ad=2.4e+12p pd=4.6e+06u as=2.4e+12p ps=4.6e+06u w=3e+06u l=8e+06u
X28 nb3 nb nb2 vssa sky130_fd_pr__nfet_01v8 ad=8e+11p pd=2.6e+06u as=8e+11p ps=2.6e+06u w=1e+06u l=8e+06u
X29 na3 na na2 vssa sky130_fd_pr__nfet_01v8 ad=8e+11p pd=2.6e+06u as=8e+11p ps=2.6e+06u w=1e+06u l=8e+06u
X30 bpb xa xa3 vdda sky130_fd_pr__pfet_01v8_lvt ad=3e+12p pd=8e+06u as=2.4e+12p ps=4.6e+06u w=3e+06u l=8e+06u
X31 qa qa qa3 vssa sky130_fd_pr__nfet_01v8 ad=1e+12p pd=4e+06u as=8e+11p ps=2.6e+06u w=1e+06u l=8e+06u
.ends

.subckt opamp_core im ip out ib q vdda bp vddx gnda vssa xn xp x y z
Xbl x y xp xn vdda vddx bp gnda vssa invt
Xcl y out vdda bp vddx gnda vssa inv_2_2
Xal im x vdda bp vddx gnda vssa inv_2_2
Xcr y out vdda bp vddx gnda vssa inv_2_2
Xbr ip y xp xn vdda vddx bp gnda vssa invt
Xar x x vdda bp vddx gnda vssa inv_2_2
Xbiasl bp bp gnda ib ib q q vdda vddx vssa z z inv_bias
Xbiasr bp bp gnda ib ib q q vdda vddx vssa z z inv_bias
X0 vddx bp sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=9.2e+06u
X1 out xn sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=9.2e+06u
X2 vddx bp sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=9.2e+06u
X3 out xn sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=9.2e+06u
X4 vddx bp sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=9.2e+06u
X5 vddx bp sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=9.2e+06u
X6 vddx bp sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=9.2e+06u
X7 vddx bp sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=9.2e+06u
X8 out xn sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=9.2e+06u
X9 out xn sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=9.2e+06u
X10 vddx bp sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=9.2e+06u
X11 vddx bp sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=9.2e+06u
X12 out xp sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=9.2e+06u
X13 out xp sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=9.2e+06u
X14 out xp sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=9.2e+06u
X15 out xp sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=9.2e+06u
.ends

.subckt opamp_pair ima ipa outa imb ipb outb ib vdda gnda vssa
Xb1 imb ipb outb ib q vdda bp vddx gnda vssa xpb xpb xb yb z opamp_core
Xa1 ima ipa outa ib q vdda bp vddx gnda vssa xpa xpa xa ya z opamp_core
Xb2 imb ipb outb ib q vdda bp vddx gnda vssa xpb xpb xb yb z opamp_core
Xa2 ima ipa outa ib q vdda bp vddx gnda vssa xpa xpa xa ya z opamp_core
.ends

