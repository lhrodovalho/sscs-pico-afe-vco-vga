magic
tech sky130A
timestamp 1634487483
<< pwell >>
rect -148 -148 148 148
<< nmos >>
rect -50 -43 50 43
<< ndiff >>
rect -79 37 -50 43
rect -79 -37 -73 37
rect -56 -37 -50 37
rect -79 -43 -50 -37
rect 50 37 79 43
rect 50 -37 56 37
rect 73 -37 79 37
rect 50 -43 79 -37
<< ndiffc >>
rect -73 -37 -56 37
rect 56 -37 73 37
<< psubdiff >>
rect -130 113 -82 130
rect 82 113 130 130
rect -130 82 -113 113
rect 113 82 130 113
rect -130 -113 -113 -82
rect 113 -113 130 -82
rect -130 -130 -82 -113
rect 82 -130 130 -113
<< psubdiffcont >>
rect -82 113 82 130
rect -130 -82 -113 82
rect 113 -82 130 82
rect -82 -130 82 -113
<< poly >>
rect -50 79 50 87
rect -50 62 -42 79
rect 42 62 50 79
rect -50 43 50 62
rect -50 -62 50 -43
rect -50 -79 -42 -62
rect 42 -79 50 -62
rect -50 -87 50 -79
<< polycont >>
rect -42 62 42 79
rect -42 -79 42 -62
<< locali >>
rect -130 113 -82 130
rect 82 113 130 130
rect -130 82 -113 113
rect 113 82 130 113
rect -50 62 -42 79
rect 42 62 50 79
rect -73 37 -56 45
rect -73 -45 -56 -37
rect 56 37 73 45
rect 56 -45 73 -37
rect -50 -79 -42 -62
rect 42 -79 50 -62
rect -130 -113 -113 -82
rect 113 -113 130 -82
rect -130 -130 -82 -113
rect 82 -130 130 -113
<< viali >>
rect -42 62 42 79
rect -73 -37 -56 37
rect 56 -37 73 37
rect -42 -79 42 -62
<< metal1 >>
rect -48 79 48 82
rect -48 62 -42 79
rect 42 62 48 79
rect -48 59 48 62
rect -76 37 -53 43
rect -76 -37 -73 37
rect -56 -37 -53 37
rect -76 -43 -53 -37
rect 53 37 76 43
rect 53 -37 56 37
rect 73 -37 76 37
rect 53 -43 76 -37
rect -48 -62 48 -59
rect -48 -79 -42 -62
rect 42 -79 48 -62
rect -48 -82 48 -79
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string FIXED_BBOX -121 -121 121 121
string parameters w 0.861 l 1.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
