* NGSPICE file created from cap1_10_core.ext - technology: sky130A

.subckt cap1_10_core a b1 b2 c1 c2 gnda vssa
X0 a c1 sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=9.2e+06u
X1 a c1 sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=9.2e+06u
X2 gnda gnda sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1.2e+06u
X3 a c2 sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=9.2e+06u
X4 a c2 sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=9.2e+06u
X5 gnda gnda sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1.2e+06u
X6 a c2 sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=9.2e+06u
X7 a c1 sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=9.2e+06u
X8 a c1 sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=9.2e+06u
X9 a b2 sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=9.2e+06u
X10 a c2 sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=9.2e+06u
X11 a c1 sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=9.2e+06u
X12 a c2 sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=9.2e+06u
X13 a c1 sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=9.2e+06u
X14 a b1 sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=9.2e+06u
X15 a c1 sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=9.2e+06u
X16 gnda gnda sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1.2e+06u
X17 a c2 sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=9.2e+06u
X18 gnda gnda sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1.2e+06u
X19 a c1 sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=9.2e+06u
X20 a c2 sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=9.2e+06u
X21 a c2 sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=9.2e+06u
X22 a c1 sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=9.2e+06u
X23 a c2 sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=9.2e+06u
X24 a c1 sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=9.2e+06u
X25 a c2 sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=9.2e+06u
.ends

