magic
tech sky130A
timestamp 1638207559
<< psubdiff >>
rect 560 480 600 520
<< locali >>
rect 560 510 600 15960
rect 560 490 570 510
rect 590 490 600 510
rect 560 480 600 490
rect 14400 510 14440 15960
rect 14400 490 14410 510
rect 14430 490 14440 510
rect 14400 480 14440 490
<< viali >>
rect 570 490 590 510
rect 14410 490 14430 510
<< metal1 >>
rect 560 515 600 520
rect 560 485 565 515
rect 595 485 600 515
rect 560 480 600 485
rect 14400 515 14440 520
rect 14400 485 14405 515
rect 14435 485 14440 515
rect 14400 480 14440 485
<< via1 >>
rect 565 510 595 515
rect 565 490 570 510
rect 570 490 590 510
rect 590 490 595 510
rect 565 485 595 490
rect 14405 510 14435 515
rect 14405 490 14410 510
rect 14410 490 14430 510
rect 14430 490 14435 510
rect 14405 485 14435 490
<< metal2 >>
rect 0 15955 520 15960
rect 0 15925 5 15955
rect 35 15925 165 15955
rect 195 15925 325 15955
rect 355 15925 485 15955
rect 515 15925 520 15955
rect 0 15920 520 15925
rect 14480 15955 15000 15960
rect 14480 15925 14485 15955
rect 14515 15925 14645 15955
rect 14675 15925 14805 15955
rect 14835 15925 14965 15955
rect 14995 15925 15000 15955
rect 14480 15920 15000 15925
rect 0 15875 520 15880
rect 0 15845 5 15875
rect 35 15845 165 15875
rect 195 15845 325 15875
rect 355 15845 485 15875
rect 515 15845 520 15875
rect 0 15840 520 15845
rect 14480 15875 15000 15880
rect 14480 15845 14485 15875
rect 14515 15845 14645 15875
rect 14675 15845 14805 15875
rect 14835 15845 14965 15875
rect 14995 15845 15000 15875
rect 14480 15840 15000 15845
rect 0 15795 520 15800
rect 0 15765 5 15795
rect 35 15765 165 15795
rect 195 15765 325 15795
rect 355 15765 485 15795
rect 515 15765 520 15795
rect 0 15760 520 15765
rect 14480 15795 15000 15800
rect 14480 15765 14485 15795
rect 14515 15765 14645 15795
rect 14675 15765 14805 15795
rect 14835 15765 14965 15795
rect 14995 15765 15000 15795
rect 14480 15760 15000 15765
rect 0 15715 520 15720
rect 0 15685 5 15715
rect 35 15685 165 15715
rect 195 15685 325 15715
rect 355 15685 485 15715
rect 515 15685 520 15715
rect 0 15680 520 15685
rect 14480 15715 15000 15720
rect 14480 15685 14485 15715
rect 14515 15685 14645 15715
rect 14675 15685 14805 15715
rect 14835 15685 14965 15715
rect 14995 15685 15000 15715
rect 14480 15680 15000 15685
rect 0 15635 520 15640
rect 0 15605 5 15635
rect 35 15605 165 15635
rect 195 15605 325 15635
rect 355 15605 485 15635
rect 515 15605 520 15635
rect 0 15600 520 15605
rect 14480 15635 15000 15640
rect 14480 15605 14485 15635
rect 14515 15605 14645 15635
rect 14675 15605 14805 15635
rect 14835 15605 14965 15635
rect 14995 15605 15000 15635
rect 14480 15600 15000 15605
rect 0 15555 520 15560
rect 0 15525 5 15555
rect 35 15525 165 15555
rect 195 15525 325 15555
rect 355 15525 485 15555
rect 515 15525 520 15555
rect 0 15520 520 15525
rect 14480 15555 15000 15560
rect 14480 15525 14485 15555
rect 14515 15525 14645 15555
rect 14675 15525 14805 15555
rect 14835 15525 14965 15555
rect 14995 15525 15000 15555
rect 14480 15520 15000 15525
rect 0 15475 520 15480
rect 0 15445 5 15475
rect 35 15445 165 15475
rect 195 15445 325 15475
rect 355 15445 485 15475
rect 515 15445 520 15475
rect 0 15440 520 15445
rect 14480 15475 15000 15480
rect 14480 15445 14485 15475
rect 14515 15445 14645 15475
rect 14675 15445 14805 15475
rect 14835 15445 14965 15475
rect 14995 15445 15000 15475
rect 14480 15440 15000 15445
rect 0 15395 520 15400
rect 0 15365 5 15395
rect 35 15365 165 15395
rect 195 15365 325 15395
rect 355 15365 485 15395
rect 515 15365 520 15395
rect 0 15360 520 15365
rect 14480 15395 15000 15400
rect 14480 15365 14485 15395
rect 14515 15365 14645 15395
rect 14675 15365 14805 15395
rect 14835 15365 14965 15395
rect 14995 15365 15000 15395
rect 14480 15360 15000 15365
rect 0 15315 520 15320
rect 0 15285 5 15315
rect 35 15285 165 15315
rect 195 15285 325 15315
rect 355 15285 485 15315
rect 515 15285 520 15315
rect 0 15280 520 15285
rect 14480 15315 15000 15320
rect 14480 15285 14485 15315
rect 14515 15285 14645 15315
rect 14675 15285 14805 15315
rect 14835 15285 14965 15315
rect 14995 15285 15000 15315
rect 14480 15280 15000 15285
rect 0 15235 520 15240
rect 0 15205 5 15235
rect 35 15205 165 15235
rect 195 15205 325 15235
rect 355 15205 485 15235
rect 515 15205 520 15235
rect 0 15200 520 15205
rect 14480 15235 15000 15240
rect 14480 15205 14485 15235
rect 14515 15205 14645 15235
rect 14675 15205 14805 15235
rect 14835 15205 14965 15235
rect 14995 15205 15000 15235
rect 14480 15200 15000 15205
rect 0 15155 520 15160
rect 0 15125 5 15155
rect 35 15125 165 15155
rect 195 15125 325 15155
rect 355 15125 485 15155
rect 515 15125 520 15155
rect 0 15120 520 15125
rect 14480 15155 15000 15160
rect 14480 15125 14485 15155
rect 14515 15125 14645 15155
rect 14675 15125 14805 15155
rect 14835 15125 14965 15155
rect 14995 15125 15000 15155
rect 14480 15120 15000 15125
rect 0 15075 520 15080
rect 0 15045 5 15075
rect 35 15045 165 15075
rect 195 15045 325 15075
rect 355 15045 485 15075
rect 515 15045 520 15075
rect 0 15040 520 15045
rect 14480 15075 15000 15080
rect 14480 15045 14485 15075
rect 14515 15045 14645 15075
rect 14675 15045 14805 15075
rect 14835 15045 14965 15075
rect 14995 15045 15000 15075
rect 14480 15040 15000 15045
rect 0 14995 520 15000
rect 0 14965 5 14995
rect 35 14965 165 14995
rect 195 14965 325 14995
rect 355 14965 485 14995
rect 515 14965 520 14995
rect 0 14960 520 14965
rect 14480 14995 15000 15000
rect 14480 14965 14485 14995
rect 14515 14965 14645 14995
rect 14675 14965 14805 14995
rect 14835 14965 14965 14995
rect 14995 14965 15000 14995
rect 14480 14960 15000 14965
rect 0 14915 520 14920
rect 0 14885 5 14915
rect 35 14885 165 14915
rect 195 14885 325 14915
rect 355 14885 485 14915
rect 515 14885 520 14915
rect 0 14880 520 14885
rect 14480 14915 15000 14920
rect 14480 14885 14485 14915
rect 14515 14885 14645 14915
rect 14675 14885 14805 14915
rect 14835 14885 14965 14915
rect 14995 14885 15000 14915
rect 14480 14880 15000 14885
rect 0 14835 520 14840
rect 0 14805 5 14835
rect 35 14805 165 14835
rect 195 14805 325 14835
rect 355 14805 485 14835
rect 515 14805 520 14835
rect 0 14800 520 14805
rect 14480 14835 15000 14840
rect 14480 14805 14485 14835
rect 14515 14805 14645 14835
rect 14675 14805 14805 14835
rect 14835 14805 14965 14835
rect 14995 14805 15000 14835
rect 14480 14800 15000 14805
rect 0 14755 520 14760
rect 0 14725 5 14755
rect 35 14725 165 14755
rect 195 14725 325 14755
rect 355 14725 485 14755
rect 515 14725 520 14755
rect 0 14720 520 14725
rect 14480 14755 15000 14760
rect 14480 14725 14485 14755
rect 14515 14725 14645 14755
rect 14675 14725 14805 14755
rect 14835 14725 14965 14755
rect 14995 14725 15000 14755
rect 14480 14720 15000 14725
rect 0 14675 520 14680
rect 0 14645 5 14675
rect 35 14645 165 14675
rect 195 14645 325 14675
rect 355 14645 485 14675
rect 515 14645 520 14675
rect 0 14640 520 14645
rect 14480 14675 15000 14680
rect 14480 14645 14485 14675
rect 14515 14645 14645 14675
rect 14675 14645 14805 14675
rect 14835 14645 14965 14675
rect 14995 14645 15000 14675
rect 14480 14640 15000 14645
rect 0 14595 520 14600
rect 0 14565 5 14595
rect 35 14565 165 14595
rect 195 14565 325 14595
rect 355 14565 485 14595
rect 515 14565 520 14595
rect 0 14560 520 14565
rect 0 14515 520 14520
rect 0 14485 5 14515
rect 35 14485 165 14515
rect 195 14485 325 14515
rect 355 14485 485 14515
rect 515 14485 520 14515
rect 0 14480 520 14485
rect 14480 14515 15000 14520
rect 14480 14485 14485 14515
rect 14515 14485 14645 14515
rect 14675 14485 14805 14515
rect 14835 14485 14965 14515
rect 14995 14485 15000 14515
rect 14480 14480 15000 14485
rect 0 14435 520 14440
rect 0 14405 5 14435
rect 35 14405 165 14435
rect 195 14405 325 14435
rect 355 14405 485 14435
rect 515 14405 520 14435
rect 0 14400 520 14405
rect 14800 14435 15000 14440
rect 14800 14405 14805 14435
rect 14835 14405 14965 14435
rect 14995 14405 15000 14435
rect 14800 14400 15000 14405
rect 0 14355 520 14360
rect 0 14325 5 14355
rect 35 14325 165 14355
rect 195 14325 325 14355
rect 355 14325 485 14355
rect 515 14325 520 14355
rect 0 14320 520 14325
rect 14480 14355 15000 14360
rect 14480 14325 14485 14355
rect 14515 14325 14645 14355
rect 14675 14325 14805 14355
rect 14835 14325 14965 14355
rect 14995 14325 15000 14355
rect 14480 14320 15000 14325
rect 0 14275 520 14280
rect 0 14245 5 14275
rect 35 14245 165 14275
rect 195 14245 325 14275
rect 355 14245 485 14275
rect 515 14245 520 14275
rect 0 14240 520 14245
rect 14480 14275 15000 14280
rect 14480 14245 14485 14275
rect 14515 14245 14645 14275
rect 14675 14245 14805 14275
rect 14835 14245 14965 14275
rect 14995 14245 15000 14275
rect 14480 14240 15000 14245
rect 0 14195 520 14200
rect 0 14165 5 14195
rect 35 14165 165 14195
rect 195 14165 325 14195
rect 355 14165 485 14195
rect 515 14165 520 14195
rect 0 14160 520 14165
rect 14480 14195 15000 14200
rect 14480 14165 14485 14195
rect 14515 14165 14645 14195
rect 14675 14165 14805 14195
rect 14835 14165 14965 14195
rect 14995 14165 15000 14195
rect 14480 14160 15000 14165
rect 0 14115 520 14120
rect 0 14085 5 14115
rect 35 14085 165 14115
rect 195 14085 325 14115
rect 355 14085 485 14115
rect 515 14085 520 14115
rect 0 14080 520 14085
rect 14480 14115 15000 14120
rect 14480 14085 14485 14115
rect 14515 14085 14645 14115
rect 14675 14085 14805 14115
rect 14835 14085 14965 14115
rect 14995 14085 15000 14115
rect 14480 14080 15000 14085
rect 0 14035 520 14040
rect 0 14005 5 14035
rect 35 14005 165 14035
rect 195 14005 325 14035
rect 355 14005 485 14035
rect 515 14005 520 14035
rect 0 14000 520 14005
rect 14480 14035 15000 14040
rect 14480 14005 14485 14035
rect 14515 14005 14645 14035
rect 14675 14005 14805 14035
rect 14835 14005 14965 14035
rect 14995 14005 15000 14035
rect 14480 14000 15000 14005
rect 0 13955 520 13960
rect 0 13925 5 13955
rect 35 13925 165 13955
rect 195 13925 325 13955
rect 355 13925 485 13955
rect 515 13925 520 13955
rect 0 13920 520 13925
rect 14480 13955 15000 13960
rect 14480 13925 14485 13955
rect 14515 13925 14645 13955
rect 14675 13925 14805 13955
rect 14835 13925 14965 13955
rect 14995 13925 15000 13955
rect 14480 13920 15000 13925
rect 0 13875 520 13880
rect 0 13845 5 13875
rect 35 13845 165 13875
rect 195 13845 325 13875
rect 355 13845 485 13875
rect 515 13845 520 13875
rect 0 13840 520 13845
rect 14480 13875 15000 13880
rect 14480 13845 14485 13875
rect 14515 13845 14645 13875
rect 14675 13845 14805 13875
rect 14835 13845 14965 13875
rect 14995 13845 15000 13875
rect 14480 13840 15000 13845
rect 0 13795 520 13800
rect 0 13765 5 13795
rect 35 13765 165 13795
rect 195 13765 325 13795
rect 355 13765 485 13795
rect 515 13765 520 13795
rect 0 13760 520 13765
rect 14480 13795 15000 13800
rect 14480 13765 14485 13795
rect 14515 13765 14645 13795
rect 14675 13765 14805 13795
rect 14835 13765 14965 13795
rect 14995 13765 15000 13795
rect 14480 13760 15000 13765
rect 0 13715 520 13720
rect 0 13685 5 13715
rect 35 13685 165 13715
rect 195 13685 325 13715
rect 355 13685 485 13715
rect 515 13685 520 13715
rect 0 13680 520 13685
rect 14480 13715 15000 13720
rect 14480 13685 14485 13715
rect 14515 13685 14645 13715
rect 14675 13685 14805 13715
rect 14835 13685 14965 13715
rect 14995 13685 15000 13715
rect 14480 13680 15000 13685
rect 0 13635 520 13640
rect 0 13605 5 13635
rect 35 13605 165 13635
rect 195 13605 325 13635
rect 355 13605 485 13635
rect 515 13605 520 13635
rect 0 13600 520 13605
rect 14480 13635 15000 13640
rect 14480 13605 14485 13635
rect 14515 13605 14645 13635
rect 14675 13605 14805 13635
rect 14835 13605 14965 13635
rect 14995 13605 15000 13635
rect 14480 13600 15000 13605
rect 0 13555 520 13560
rect 0 13525 5 13555
rect 35 13525 165 13555
rect 195 13525 325 13555
rect 355 13525 485 13555
rect 515 13525 520 13555
rect 0 13520 520 13525
rect 14480 13555 15000 13560
rect 14480 13525 14485 13555
rect 14515 13525 14645 13555
rect 14675 13525 14805 13555
rect 14835 13525 14965 13555
rect 14995 13525 15000 13555
rect 14480 13520 15000 13525
rect 0 13475 520 13480
rect 0 13445 5 13475
rect 35 13445 165 13475
rect 195 13445 325 13475
rect 355 13445 485 13475
rect 515 13445 520 13475
rect 0 13440 520 13445
rect 14480 13475 15000 13480
rect 14480 13445 14485 13475
rect 14515 13445 14645 13475
rect 14675 13445 14805 13475
rect 14835 13445 14965 13475
rect 14995 13445 15000 13475
rect 14480 13440 15000 13445
rect 0 13395 520 13400
rect 0 13365 5 13395
rect 35 13365 165 13395
rect 195 13365 325 13395
rect 355 13365 485 13395
rect 515 13365 520 13395
rect 0 13360 520 13365
rect 14480 13395 15000 13400
rect 14480 13365 14485 13395
rect 14515 13365 14645 13395
rect 14675 13365 14805 13395
rect 14835 13365 14965 13395
rect 14995 13365 15000 13395
rect 14480 13360 15000 13365
rect 0 13315 520 13320
rect 0 13285 5 13315
rect 35 13285 165 13315
rect 195 13285 325 13315
rect 355 13285 485 13315
rect 515 13285 520 13315
rect 0 13280 520 13285
rect 14480 13315 15000 13320
rect 14480 13285 14485 13315
rect 14515 13285 14645 13315
rect 14675 13285 14805 13315
rect 14835 13285 14965 13315
rect 14995 13285 15000 13315
rect 14480 13280 15000 13285
rect 0 13235 520 13240
rect 0 13205 5 13235
rect 35 13205 165 13235
rect 195 13205 325 13235
rect 355 13205 485 13235
rect 515 13205 520 13235
rect 0 13200 520 13205
rect 14480 13235 15000 13240
rect 14480 13205 14485 13235
rect 14515 13205 14645 13235
rect 14675 13205 14805 13235
rect 14835 13205 14965 13235
rect 14995 13205 15000 13235
rect 14480 13200 15000 13205
rect 0 13155 520 13160
rect 0 13125 5 13155
rect 35 13125 165 13155
rect 195 13125 325 13155
rect 355 13125 485 13155
rect 515 13125 520 13155
rect 0 13120 520 13125
rect 14640 13155 15000 13160
rect 14640 13125 14645 13155
rect 14675 13125 14805 13155
rect 14835 13125 14965 13155
rect 14995 13125 15000 13155
rect 14640 13120 15000 13125
rect 0 13075 520 13080
rect 0 13045 5 13075
rect 35 13045 165 13075
rect 195 13045 325 13075
rect 355 13045 485 13075
rect 515 13045 520 13075
rect 0 13040 520 13045
rect 14480 13075 15000 13080
rect 14480 13045 14485 13075
rect 14515 13045 14645 13075
rect 14675 13045 14805 13075
rect 14835 13045 14965 13075
rect 14995 13045 15000 13075
rect 14480 13040 15000 13045
rect 0 12995 520 13000
rect 0 12965 5 12995
rect 35 12965 165 12995
rect 195 12965 325 12995
rect 355 12965 485 12995
rect 515 12965 520 12995
rect 0 12960 520 12965
rect 14480 12995 15000 13000
rect 14480 12965 14485 12995
rect 14515 12965 14645 12995
rect 14675 12965 14805 12995
rect 14835 12965 14965 12995
rect 14995 12965 15000 12995
rect 14480 12960 15000 12965
rect 0 12915 520 12920
rect 0 12885 5 12915
rect 35 12885 165 12915
rect 195 12885 325 12915
rect 355 12885 485 12915
rect 515 12885 520 12915
rect 0 12880 520 12885
rect 14480 12915 15000 12920
rect 14480 12885 14485 12915
rect 14515 12885 14645 12915
rect 14675 12885 14805 12915
rect 14835 12885 14965 12915
rect 14995 12885 15000 12915
rect 14480 12880 15000 12885
rect 0 12835 520 12840
rect 0 12805 5 12835
rect 35 12805 165 12835
rect 195 12805 325 12835
rect 355 12805 485 12835
rect 515 12805 520 12835
rect 0 12800 520 12805
rect 14480 12835 15000 12840
rect 14480 12805 14485 12835
rect 14515 12805 14645 12835
rect 14675 12805 14805 12835
rect 14835 12805 14965 12835
rect 14995 12805 15000 12835
rect 14480 12800 15000 12805
rect 0 12755 520 12760
rect 0 12725 5 12755
rect 35 12725 165 12755
rect 195 12725 325 12755
rect 355 12725 485 12755
rect 515 12725 520 12755
rect 0 12720 520 12725
rect 14480 12755 15000 12760
rect 14480 12725 14485 12755
rect 14515 12725 14645 12755
rect 14675 12725 14805 12755
rect 14835 12725 14965 12755
rect 14995 12725 15000 12755
rect 14480 12720 15000 12725
rect 0 12675 520 12680
rect 0 12645 5 12675
rect 35 12645 165 12675
rect 195 12645 325 12675
rect 355 12645 485 12675
rect 515 12645 520 12675
rect 0 12640 520 12645
rect 14480 12675 15000 12680
rect 14480 12645 14485 12675
rect 14515 12645 14645 12675
rect 14675 12645 14805 12675
rect 14835 12645 14965 12675
rect 14995 12645 15000 12675
rect 14480 12640 15000 12645
rect 0 12595 520 12600
rect 0 12565 5 12595
rect 35 12565 165 12595
rect 195 12565 325 12595
rect 355 12565 485 12595
rect 515 12565 520 12595
rect 0 12560 520 12565
rect 14480 12595 15000 12600
rect 14480 12565 14485 12595
rect 14515 12565 14645 12595
rect 14675 12565 14805 12595
rect 14835 12565 14965 12595
rect 14995 12565 15000 12595
rect 14480 12560 15000 12565
rect 0 12515 520 12520
rect 0 12485 5 12515
rect 35 12485 165 12515
rect 195 12485 325 12515
rect 355 12485 485 12515
rect 515 12485 520 12515
rect 0 12480 520 12485
rect 14480 12515 15000 12520
rect 14480 12485 14485 12515
rect 14515 12485 14645 12515
rect 14675 12485 14805 12515
rect 14835 12485 14965 12515
rect 14995 12485 15000 12515
rect 14480 12480 15000 12485
rect 0 12435 520 12440
rect 0 12405 5 12435
rect 35 12405 165 12435
rect 195 12405 325 12435
rect 355 12405 485 12435
rect 515 12405 520 12435
rect 0 12400 520 12405
rect 14480 12435 15000 12440
rect 14480 12405 14485 12435
rect 14515 12405 14645 12435
rect 14675 12405 14805 12435
rect 14835 12405 14965 12435
rect 14995 12405 15000 12435
rect 14480 12400 15000 12405
rect 0 12355 520 12360
rect 0 12325 5 12355
rect 35 12325 165 12355
rect 195 12325 325 12355
rect 355 12325 485 12355
rect 515 12325 520 12355
rect 0 12320 520 12325
rect 14480 12355 15000 12360
rect 14480 12325 14485 12355
rect 14515 12325 14645 12355
rect 14675 12325 14805 12355
rect 14835 12325 14965 12355
rect 14995 12325 15000 12355
rect 14480 12320 15000 12325
rect 0 12275 520 12280
rect 0 12245 5 12275
rect 35 12245 165 12275
rect 195 12245 325 12275
rect 355 12245 485 12275
rect 515 12245 520 12275
rect 0 12240 520 12245
rect 14480 12275 15000 12280
rect 14480 12245 14485 12275
rect 14515 12245 14645 12275
rect 14675 12245 14805 12275
rect 14835 12245 14965 12275
rect 14995 12245 15000 12275
rect 14480 12240 15000 12245
rect 0 12195 520 12200
rect 0 12165 5 12195
rect 35 12165 165 12195
rect 195 12165 325 12195
rect 355 12165 485 12195
rect 515 12165 520 12195
rect 0 12160 520 12165
rect 14480 12195 15000 12200
rect 14480 12165 14485 12195
rect 14515 12165 14645 12195
rect 14675 12165 14805 12195
rect 14835 12165 14965 12195
rect 14995 12165 15000 12195
rect 14480 12160 15000 12165
rect 0 12115 520 12120
rect 0 12085 5 12115
rect 35 12085 165 12115
rect 195 12085 325 12115
rect 355 12085 485 12115
rect 515 12085 520 12115
rect 0 12080 520 12085
rect 14480 12115 15000 12120
rect 14480 12085 14485 12115
rect 14515 12085 14645 12115
rect 14675 12085 14805 12115
rect 14835 12085 14965 12115
rect 14995 12085 15000 12115
rect 14480 12080 15000 12085
rect 0 12035 520 12040
rect 0 12005 5 12035
rect 35 12005 165 12035
rect 195 12005 325 12035
rect 355 12005 485 12035
rect 515 12005 520 12035
rect 0 12000 520 12005
rect 14480 12035 15000 12040
rect 14480 12005 14485 12035
rect 14515 12005 14645 12035
rect 14675 12005 14805 12035
rect 14835 12005 14965 12035
rect 14995 12005 15000 12035
rect 14480 12000 15000 12005
rect 0 11955 520 11960
rect 0 11925 5 11955
rect 35 11925 165 11955
rect 195 11925 325 11955
rect 355 11925 485 11955
rect 515 11925 520 11955
rect 0 11920 520 11925
rect 14480 11955 15000 11960
rect 14480 11925 14485 11955
rect 14515 11925 14645 11955
rect 14675 11925 14805 11955
rect 14835 11925 14965 11955
rect 14995 11925 15000 11955
rect 14480 11920 15000 11925
rect 0 11875 520 11880
rect 0 11845 5 11875
rect 35 11845 165 11875
rect 195 11845 325 11875
rect 355 11845 485 11875
rect 515 11845 520 11875
rect 0 11840 520 11845
rect 14800 11875 15000 11880
rect 14800 11845 14805 11875
rect 14835 11845 14965 11875
rect 14995 11845 15000 11875
rect 14800 11840 15000 11845
rect 0 11795 520 11800
rect 0 11765 5 11795
rect 35 11765 165 11795
rect 195 11765 325 11795
rect 355 11765 485 11795
rect 515 11765 520 11795
rect 0 11760 520 11765
rect 14480 11795 15000 11800
rect 14480 11765 14485 11795
rect 14515 11765 14645 11795
rect 14675 11765 14805 11795
rect 14835 11765 14965 11795
rect 14995 11765 15000 11795
rect 14480 11760 15000 11765
rect 0 11715 520 11720
rect 0 11685 5 11715
rect 35 11685 165 11715
rect 195 11685 325 11715
rect 355 11685 485 11715
rect 515 11685 520 11715
rect 0 11680 520 11685
rect 0 11635 520 11640
rect 0 11605 5 11635
rect 35 11605 165 11635
rect 195 11605 325 11635
rect 355 11605 485 11635
rect 515 11605 520 11635
rect 0 11600 520 11605
rect 14480 11635 15000 11640
rect 14480 11605 14485 11635
rect 14515 11605 14645 11635
rect 14675 11605 14805 11635
rect 14835 11605 14965 11635
rect 14995 11605 15000 11635
rect 14480 11600 15000 11605
rect 0 11555 520 11560
rect 0 11525 5 11555
rect 35 11525 165 11555
rect 195 11525 325 11555
rect 355 11525 485 11555
rect 515 11525 520 11555
rect 0 11520 520 11525
rect 14480 11555 15000 11560
rect 14480 11525 14485 11555
rect 14515 11525 14645 11555
rect 14675 11525 14805 11555
rect 14835 11525 14965 11555
rect 14995 11525 15000 11555
rect 14480 11520 15000 11525
rect 0 11475 520 11480
rect 0 11445 5 11475
rect 35 11445 165 11475
rect 195 11445 325 11475
rect 355 11445 485 11475
rect 515 11445 520 11475
rect 0 11440 520 11445
rect 14480 11475 15000 11480
rect 14480 11445 14485 11475
rect 14515 11445 14645 11475
rect 14675 11445 14805 11475
rect 14835 11445 14965 11475
rect 14995 11445 15000 11475
rect 14480 11440 15000 11445
rect 0 11395 520 11400
rect 0 11365 5 11395
rect 35 11365 165 11395
rect 195 11365 325 11395
rect 355 11365 485 11395
rect 515 11365 520 11395
rect 0 11360 520 11365
rect 14480 11395 15000 11400
rect 14480 11365 14485 11395
rect 14515 11365 14645 11395
rect 14675 11365 14805 11395
rect 14835 11365 14965 11395
rect 14995 11365 15000 11395
rect 14480 11360 15000 11365
rect 14480 11315 15000 11320
rect 14480 11285 14485 11315
rect 14515 11285 14645 11315
rect 14675 11285 14805 11315
rect 14835 11285 14965 11315
rect 14995 11285 15000 11315
rect 14480 11280 15000 11285
rect 0 11235 520 11240
rect 0 11205 5 11235
rect 35 11205 165 11235
rect 195 11205 325 11235
rect 355 11205 485 11235
rect 515 11205 520 11235
rect 0 11200 520 11205
rect 14480 11235 15000 11240
rect 14480 11205 14485 11235
rect 14515 11205 14645 11235
rect 14675 11205 14805 11235
rect 14835 11205 14965 11235
rect 14995 11205 15000 11235
rect 14480 11200 15000 11205
rect 0 11155 200 11160
rect 0 11125 5 11155
rect 35 11125 165 11155
rect 195 11125 200 11155
rect 0 11120 200 11125
rect 14480 11155 15000 11160
rect 14480 11125 14485 11155
rect 14515 11125 14645 11155
rect 14675 11125 14805 11155
rect 14835 11125 14965 11155
rect 14995 11125 15000 11155
rect 14480 11120 15000 11125
rect 0 11075 520 11080
rect 0 11045 5 11075
rect 35 11045 165 11075
rect 195 11045 325 11075
rect 355 11045 485 11075
rect 515 11045 520 11075
rect 0 11040 520 11045
rect 14480 11075 15000 11080
rect 14480 11045 14485 11075
rect 14515 11045 14645 11075
rect 14675 11045 14805 11075
rect 14835 11045 14965 11075
rect 14995 11045 15000 11075
rect 14480 11040 15000 11045
rect 0 10995 520 11000
rect 0 10965 5 10995
rect 35 10965 165 10995
rect 195 10965 325 10995
rect 355 10965 485 10995
rect 515 10965 520 10995
rect 0 10960 520 10965
rect 14480 10995 15000 11000
rect 14480 10965 14485 10995
rect 14515 10965 14645 10995
rect 14675 10965 14805 10995
rect 14835 10965 14965 10995
rect 14995 10965 15000 10995
rect 14480 10960 15000 10965
rect 0 10915 520 10920
rect 0 10885 5 10915
rect 35 10885 165 10915
rect 195 10885 325 10915
rect 355 10885 485 10915
rect 515 10885 520 10915
rect 0 10880 520 10885
rect 14480 10915 15000 10920
rect 14480 10885 14485 10915
rect 14515 10885 14645 10915
rect 14675 10885 14805 10915
rect 14835 10885 14965 10915
rect 14995 10885 15000 10915
rect 14480 10880 15000 10885
rect 0 10835 520 10840
rect 0 10805 5 10835
rect 35 10805 165 10835
rect 195 10805 325 10835
rect 355 10805 485 10835
rect 515 10805 520 10835
rect 0 10800 520 10805
rect 14480 10835 15000 10840
rect 14480 10805 14485 10835
rect 14515 10805 14645 10835
rect 14675 10805 14805 10835
rect 14835 10805 14965 10835
rect 14995 10805 15000 10835
rect 14480 10800 15000 10805
rect 0 10755 520 10760
rect 0 10725 5 10755
rect 35 10725 165 10755
rect 195 10725 325 10755
rect 355 10725 485 10755
rect 515 10725 520 10755
rect 0 10720 520 10725
rect 14480 10755 15000 10760
rect 14480 10725 14485 10755
rect 14515 10725 14645 10755
rect 14675 10725 14805 10755
rect 14835 10725 14965 10755
rect 14995 10725 15000 10755
rect 14480 10720 15000 10725
rect 0 10675 520 10680
rect 0 10645 5 10675
rect 35 10645 165 10675
rect 195 10645 325 10675
rect 355 10645 485 10675
rect 515 10645 520 10675
rect 0 10640 520 10645
rect 14480 10675 15000 10680
rect 14480 10645 14485 10675
rect 14515 10645 14645 10675
rect 14675 10645 14805 10675
rect 14835 10645 14965 10675
rect 14995 10645 15000 10675
rect 14480 10640 15000 10645
rect 0 10595 520 10600
rect 0 10565 5 10595
rect 35 10565 165 10595
rect 195 10565 325 10595
rect 355 10565 485 10595
rect 515 10565 520 10595
rect 0 10560 520 10565
rect 14480 10595 15000 10600
rect 14480 10565 14485 10595
rect 14515 10565 14645 10595
rect 14675 10565 14805 10595
rect 14835 10565 14965 10595
rect 14995 10565 15000 10595
rect 14480 10560 15000 10565
rect 0 10515 520 10520
rect 0 10485 5 10515
rect 35 10485 165 10515
rect 195 10485 325 10515
rect 355 10485 485 10515
rect 515 10485 520 10515
rect 0 10480 520 10485
rect 14480 10515 15000 10520
rect 14480 10485 14485 10515
rect 14515 10485 14645 10515
rect 14675 10485 14805 10515
rect 14835 10485 14965 10515
rect 14995 10485 15000 10515
rect 14480 10480 15000 10485
rect 0 10435 520 10440
rect 0 10405 5 10435
rect 35 10405 165 10435
rect 195 10405 325 10435
rect 355 10405 485 10435
rect 515 10405 520 10435
rect 0 10400 520 10405
rect 14480 10435 15000 10440
rect 14480 10405 14485 10435
rect 14515 10405 14645 10435
rect 14675 10405 14805 10435
rect 14835 10405 14965 10435
rect 14995 10405 15000 10435
rect 14480 10400 15000 10405
rect 0 10355 520 10360
rect 0 10325 5 10355
rect 35 10325 165 10355
rect 195 10325 325 10355
rect 355 10325 485 10355
rect 515 10325 520 10355
rect 0 10320 520 10325
rect 14480 10355 15000 10360
rect 14480 10325 14485 10355
rect 14515 10325 14645 10355
rect 14675 10325 14805 10355
rect 14835 10325 14965 10355
rect 14995 10325 15000 10355
rect 14480 10320 15000 10325
rect 0 10275 520 10280
rect 0 10245 5 10275
rect 35 10245 165 10275
rect 195 10245 325 10275
rect 355 10245 485 10275
rect 515 10245 520 10275
rect 0 10240 520 10245
rect 14480 10275 15000 10280
rect 14480 10245 14485 10275
rect 14515 10245 14645 10275
rect 14675 10245 14805 10275
rect 14835 10245 14965 10275
rect 14995 10245 15000 10275
rect 14480 10240 15000 10245
rect 0 10195 520 10200
rect 0 10165 5 10195
rect 35 10165 165 10195
rect 195 10165 325 10195
rect 355 10165 485 10195
rect 515 10165 520 10195
rect 0 10160 520 10165
rect 14480 10195 15000 10200
rect 14480 10165 14485 10195
rect 14515 10165 14645 10195
rect 14675 10165 14805 10195
rect 14835 10165 14965 10195
rect 14995 10165 15000 10195
rect 14480 10160 15000 10165
rect 0 10115 520 10120
rect 0 10085 5 10115
rect 35 10085 165 10115
rect 195 10085 325 10115
rect 355 10085 485 10115
rect 515 10085 520 10115
rect 0 10080 520 10085
rect 14480 10115 15000 10120
rect 14480 10085 14485 10115
rect 14515 10085 14645 10115
rect 14675 10085 14805 10115
rect 14835 10085 14965 10115
rect 14995 10085 15000 10115
rect 14480 10080 15000 10085
rect 0 10035 520 10040
rect 0 10005 5 10035
rect 35 10005 165 10035
rect 195 10005 325 10035
rect 355 10005 485 10035
rect 515 10005 520 10035
rect 0 10000 520 10005
rect 14480 10035 15000 10040
rect 14480 10005 14485 10035
rect 14515 10005 14645 10035
rect 14675 10005 14805 10035
rect 14835 10005 14965 10035
rect 14995 10005 15000 10035
rect 14480 10000 15000 10005
rect 0 9955 520 9960
rect 0 9925 5 9955
rect 35 9925 165 9955
rect 195 9925 325 9955
rect 355 9925 485 9955
rect 515 9925 520 9955
rect 0 9920 520 9925
rect 14480 9955 15000 9960
rect 14480 9925 14485 9955
rect 14515 9925 14645 9955
rect 14675 9925 14805 9955
rect 14835 9925 14965 9955
rect 14995 9925 15000 9955
rect 14480 9920 15000 9925
rect 0 9875 360 9880
rect 0 9845 5 9875
rect 35 9845 165 9875
rect 195 9845 325 9875
rect 355 9845 360 9875
rect 0 9840 360 9845
rect 14480 9875 15000 9880
rect 14480 9845 14485 9875
rect 14515 9845 14645 9875
rect 14675 9845 14805 9875
rect 14835 9845 14965 9875
rect 14995 9845 15000 9875
rect 14480 9840 15000 9845
rect 0 9795 520 9800
rect 0 9765 5 9795
rect 35 9765 165 9795
rect 195 9765 325 9795
rect 355 9765 485 9795
rect 515 9765 520 9795
rect 0 9760 520 9765
rect 14480 9795 15000 9800
rect 14480 9765 14485 9795
rect 14515 9765 14645 9795
rect 14675 9765 14805 9795
rect 14835 9765 14965 9795
rect 14995 9765 15000 9795
rect 14480 9760 15000 9765
rect 0 9715 520 9720
rect 0 9685 5 9715
rect 35 9685 165 9715
rect 195 9685 325 9715
rect 355 9685 485 9715
rect 515 9685 520 9715
rect 0 9680 520 9685
rect 14480 9715 15000 9720
rect 14480 9685 14485 9715
rect 14515 9685 14645 9715
rect 14675 9685 14805 9715
rect 14835 9685 14965 9715
rect 14995 9685 15000 9715
rect 14480 9680 15000 9685
rect 0 9635 520 9640
rect 0 9605 5 9635
rect 35 9605 165 9635
rect 195 9605 325 9635
rect 355 9605 485 9635
rect 515 9605 520 9635
rect 0 9600 520 9605
rect 14480 9635 15000 9640
rect 14480 9605 14485 9635
rect 14515 9605 14645 9635
rect 14675 9605 14805 9635
rect 14835 9605 14965 9635
rect 14995 9605 15000 9635
rect 14480 9600 15000 9605
rect 0 9555 520 9560
rect 0 9525 5 9555
rect 35 9525 165 9555
rect 195 9525 325 9555
rect 355 9525 485 9555
rect 515 9525 520 9555
rect 0 9520 520 9525
rect 14480 9555 15000 9560
rect 14480 9525 14485 9555
rect 14515 9525 14645 9555
rect 14675 9525 14805 9555
rect 14835 9525 14965 9555
rect 14995 9525 15000 9555
rect 14480 9520 15000 9525
rect 0 9475 520 9480
rect 0 9445 5 9475
rect 35 9445 165 9475
rect 195 9445 325 9475
rect 355 9445 485 9475
rect 515 9445 520 9475
rect 0 9440 520 9445
rect 14480 9475 15000 9480
rect 14480 9445 14485 9475
rect 14515 9445 14645 9475
rect 14675 9445 14805 9475
rect 14835 9445 14965 9475
rect 14995 9445 15000 9475
rect 14480 9440 15000 9445
rect 0 9395 520 9400
rect 0 9365 5 9395
rect 35 9365 165 9395
rect 195 9365 325 9395
rect 355 9365 485 9395
rect 515 9365 520 9395
rect 0 9360 520 9365
rect 14480 9395 15000 9400
rect 14480 9365 14485 9395
rect 14515 9365 14645 9395
rect 14675 9365 14805 9395
rect 14835 9365 14965 9395
rect 14995 9365 15000 9395
rect 14480 9360 15000 9365
rect 0 9315 520 9320
rect 0 9285 5 9315
rect 35 9285 165 9315
rect 195 9285 325 9315
rect 355 9285 485 9315
rect 515 9285 520 9315
rect 0 9280 520 9285
rect 14480 9315 15000 9320
rect 14480 9285 14485 9315
rect 14515 9285 14645 9315
rect 14675 9285 14805 9315
rect 14835 9285 14965 9315
rect 14995 9285 15000 9315
rect 14480 9280 15000 9285
rect 0 9235 520 9240
rect 0 9205 5 9235
rect 35 9205 165 9235
rect 195 9205 325 9235
rect 355 9205 485 9235
rect 515 9205 520 9235
rect 0 9200 520 9205
rect 14480 9235 15000 9240
rect 14480 9205 14485 9235
rect 14515 9205 14645 9235
rect 14675 9205 14805 9235
rect 14835 9205 14965 9235
rect 14995 9205 15000 9235
rect 14480 9200 15000 9205
rect 0 9155 520 9160
rect 0 9125 5 9155
rect 35 9125 165 9155
rect 195 9125 325 9155
rect 355 9125 485 9155
rect 515 9125 520 9155
rect 0 9120 520 9125
rect 14480 9155 15000 9160
rect 14480 9125 14485 9155
rect 14515 9125 14645 9155
rect 14675 9125 14805 9155
rect 14835 9125 14965 9155
rect 14995 9125 15000 9155
rect 14480 9120 15000 9125
rect 0 9075 520 9080
rect 0 9045 5 9075
rect 35 9045 165 9075
rect 195 9045 325 9075
rect 355 9045 485 9075
rect 515 9045 520 9075
rect 0 9040 520 9045
rect 14480 9075 15000 9080
rect 14480 9045 14485 9075
rect 14515 9045 14645 9075
rect 14675 9045 14805 9075
rect 14835 9045 14965 9075
rect 14995 9045 15000 9075
rect 14480 9040 15000 9045
rect 0 8995 520 9000
rect 0 8965 5 8995
rect 35 8965 165 8995
rect 195 8965 325 8995
rect 355 8965 485 8995
rect 515 8965 520 8995
rect 0 8960 520 8965
rect 14480 8995 15000 9000
rect 14480 8965 14485 8995
rect 14515 8965 14645 8995
rect 14675 8965 14805 8995
rect 14835 8965 14965 8995
rect 14995 8965 15000 8995
rect 14480 8960 15000 8965
rect 0 8915 520 8920
rect 0 8885 5 8915
rect 35 8885 165 8915
rect 195 8885 325 8915
rect 355 8885 485 8915
rect 515 8885 520 8915
rect 0 8880 520 8885
rect 14480 8915 15000 8920
rect 14480 8885 14485 8915
rect 14515 8885 14645 8915
rect 14675 8885 14805 8915
rect 14835 8885 14965 8915
rect 14995 8885 15000 8915
rect 14480 8880 15000 8885
rect 0 8835 520 8840
rect 0 8805 5 8835
rect 35 8805 165 8835
rect 195 8805 325 8835
rect 355 8805 485 8835
rect 515 8805 520 8835
rect 0 8800 520 8805
rect 14480 8835 15000 8840
rect 14480 8805 14485 8835
rect 14515 8805 14645 8835
rect 14675 8805 14805 8835
rect 14835 8805 14965 8835
rect 14995 8805 15000 8835
rect 14480 8800 15000 8805
rect 0 8755 520 8760
rect 0 8725 5 8755
rect 35 8725 165 8755
rect 195 8725 325 8755
rect 355 8725 485 8755
rect 515 8725 520 8755
rect 0 8720 520 8725
rect 14480 8755 15000 8760
rect 14480 8725 14485 8755
rect 14515 8725 14645 8755
rect 14675 8725 14805 8755
rect 14835 8725 14965 8755
rect 14995 8725 15000 8755
rect 14480 8720 15000 8725
rect 0 8675 520 8680
rect 0 8645 5 8675
rect 35 8645 165 8675
rect 195 8645 325 8675
rect 355 8645 485 8675
rect 515 8645 520 8675
rect 0 8640 520 8645
rect 14480 8675 15000 8680
rect 14480 8645 14485 8675
rect 14515 8645 14645 8675
rect 14675 8645 14805 8675
rect 14835 8645 14965 8675
rect 14995 8645 15000 8675
rect 14480 8640 15000 8645
rect 0 8595 200 8600
rect 0 8565 5 8595
rect 35 8565 165 8595
rect 195 8565 200 8595
rect 0 8560 200 8565
rect 14480 8595 15000 8600
rect 14480 8565 14485 8595
rect 14515 8565 14645 8595
rect 14675 8565 14805 8595
rect 14835 8565 14965 8595
rect 14995 8565 15000 8595
rect 14480 8560 15000 8565
rect 0 8515 520 8520
rect 0 8485 5 8515
rect 35 8485 165 8515
rect 195 8485 325 8515
rect 355 8485 485 8515
rect 515 8485 520 8515
rect 0 8480 520 8485
rect 14480 8515 15000 8520
rect 14480 8485 14485 8515
rect 14515 8485 14645 8515
rect 14675 8485 14805 8515
rect 14835 8485 14965 8515
rect 14995 8485 15000 8515
rect 14480 8480 15000 8485
rect 14480 8435 15000 8440
rect 14480 8405 14485 8435
rect 14515 8405 14645 8435
rect 14675 8405 14805 8435
rect 14835 8405 14965 8435
rect 14995 8405 15000 8435
rect 14480 8400 15000 8405
rect 0 8355 520 8360
rect 0 8325 5 8355
rect 35 8325 165 8355
rect 195 8325 325 8355
rect 355 8325 485 8355
rect 515 8325 520 8355
rect 0 8320 520 8325
rect 14480 8355 15000 8360
rect 14480 8325 14485 8355
rect 14515 8325 14645 8355
rect 14675 8325 14805 8355
rect 14835 8325 14965 8355
rect 14995 8325 15000 8355
rect 14480 8320 15000 8325
rect 0 8275 520 8280
rect 0 8245 5 8275
rect 35 8245 165 8275
rect 195 8245 325 8275
rect 355 8245 485 8275
rect 515 8245 520 8275
rect 0 8240 520 8245
rect 14480 8275 15000 8280
rect 14480 8245 14485 8275
rect 14515 8245 14645 8275
rect 14675 8245 14805 8275
rect 14835 8245 14965 8275
rect 14995 8245 15000 8275
rect 14480 8240 15000 8245
rect 0 8195 520 8200
rect 0 8165 5 8195
rect 35 8165 165 8195
rect 195 8165 325 8195
rect 355 8165 485 8195
rect 515 8165 520 8195
rect 0 8160 520 8165
rect 14480 8195 15000 8200
rect 14480 8165 14485 8195
rect 14515 8165 14645 8195
rect 14675 8165 14805 8195
rect 14835 8165 14965 8195
rect 14995 8165 15000 8195
rect 14480 8160 15000 8165
rect 0 8115 520 8120
rect 0 8085 5 8115
rect 35 8085 165 8115
rect 195 8085 325 8115
rect 355 8085 485 8115
rect 515 8085 520 8115
rect 0 8080 520 8085
rect 14480 8115 15000 8120
rect 14480 8085 14485 8115
rect 14515 8085 14645 8115
rect 14675 8085 14805 8115
rect 14835 8085 14965 8115
rect 14995 8085 15000 8115
rect 14480 8080 15000 8085
rect 14480 8035 15000 8040
rect 14480 8005 14485 8035
rect 14515 8005 14645 8035
rect 14675 8005 14805 8035
rect 14835 8005 14965 8035
rect 14995 8005 15000 8035
rect 14480 8000 15000 8005
rect 0 7955 520 7960
rect 0 7925 5 7955
rect 35 7925 165 7955
rect 195 7925 325 7955
rect 355 7925 485 7955
rect 515 7925 520 7955
rect 0 7920 520 7925
rect 14480 7955 15000 7960
rect 14480 7925 14485 7955
rect 14515 7925 14645 7955
rect 14675 7925 14805 7955
rect 14835 7925 14965 7955
rect 14995 7925 15000 7955
rect 14480 7920 15000 7925
rect 0 7875 200 7880
rect 0 7845 5 7875
rect 35 7845 165 7875
rect 195 7845 200 7875
rect 0 7840 200 7845
rect 14480 7875 15000 7880
rect 14480 7845 14485 7875
rect 14515 7845 14645 7875
rect 14675 7845 14805 7875
rect 14835 7845 14965 7875
rect 14995 7845 15000 7875
rect 14480 7840 15000 7845
rect 0 7795 520 7800
rect 0 7765 5 7795
rect 35 7765 165 7795
rect 195 7765 325 7795
rect 355 7765 485 7795
rect 515 7765 520 7795
rect 0 7760 520 7765
rect 14480 7795 15000 7800
rect 14480 7765 14485 7795
rect 14515 7765 14645 7795
rect 14675 7765 14805 7795
rect 14835 7765 14965 7795
rect 14995 7765 15000 7795
rect 14480 7760 15000 7765
rect 0 7715 520 7720
rect 0 7685 5 7715
rect 35 7685 165 7715
rect 195 7685 325 7715
rect 355 7685 485 7715
rect 515 7685 520 7715
rect 0 7680 520 7685
rect 14480 7715 15000 7720
rect 14480 7685 14485 7715
rect 14515 7685 14645 7715
rect 14675 7685 14805 7715
rect 14835 7685 14965 7715
rect 14995 7685 15000 7715
rect 14480 7680 15000 7685
rect 0 7635 520 7640
rect 0 7605 5 7635
rect 35 7605 165 7635
rect 195 7605 325 7635
rect 355 7605 485 7635
rect 515 7605 520 7635
rect 0 7600 520 7605
rect 14480 7635 15000 7640
rect 14480 7605 14485 7635
rect 14515 7605 14645 7635
rect 14675 7605 14805 7635
rect 14835 7605 14965 7635
rect 14995 7605 15000 7635
rect 14480 7600 15000 7605
rect 0 7555 520 7560
rect 0 7525 5 7555
rect 35 7525 165 7555
rect 195 7525 325 7555
rect 355 7525 485 7555
rect 515 7525 520 7555
rect 0 7520 520 7525
rect 14480 7555 15000 7560
rect 14480 7525 14485 7555
rect 14515 7525 14645 7555
rect 14675 7525 14805 7555
rect 14835 7525 14965 7555
rect 14995 7525 15000 7555
rect 14480 7520 15000 7525
rect 0 7475 520 7480
rect 0 7445 5 7475
rect 35 7445 165 7475
rect 195 7445 325 7475
rect 355 7445 485 7475
rect 515 7445 520 7475
rect 0 7440 520 7445
rect 14480 7475 15000 7480
rect 14480 7445 14485 7475
rect 14515 7445 14645 7475
rect 14675 7445 14805 7475
rect 14835 7445 14965 7475
rect 14995 7445 15000 7475
rect 14480 7440 15000 7445
rect 0 7395 520 7400
rect 0 7365 5 7395
rect 35 7365 165 7395
rect 195 7365 325 7395
rect 355 7365 485 7395
rect 515 7365 520 7395
rect 0 7360 520 7365
rect 14480 7395 15000 7400
rect 14480 7365 14485 7395
rect 14515 7365 14645 7395
rect 14675 7365 14805 7395
rect 14835 7365 14965 7395
rect 14995 7365 15000 7395
rect 14480 7360 15000 7365
rect 0 7315 520 7320
rect 0 7285 5 7315
rect 35 7285 165 7315
rect 195 7285 325 7315
rect 355 7285 485 7315
rect 515 7285 520 7315
rect 0 7280 520 7285
rect 14480 7315 15000 7320
rect 14480 7285 14485 7315
rect 14515 7285 14645 7315
rect 14675 7285 14805 7315
rect 14835 7285 14965 7315
rect 14995 7285 15000 7315
rect 14480 7280 15000 7285
rect 0 7235 520 7240
rect 0 7205 5 7235
rect 35 7205 165 7235
rect 195 7205 325 7235
rect 355 7205 485 7235
rect 515 7205 520 7235
rect 0 7200 520 7205
rect 14480 7235 15000 7240
rect 14480 7205 14485 7235
rect 14515 7205 14645 7235
rect 14675 7205 14805 7235
rect 14835 7205 14965 7235
rect 14995 7205 15000 7235
rect 14480 7200 15000 7205
rect 0 7155 520 7160
rect 0 7125 5 7155
rect 35 7125 165 7155
rect 195 7125 325 7155
rect 355 7125 485 7155
rect 515 7125 520 7155
rect 0 7120 520 7125
rect 14480 7155 15000 7160
rect 14480 7125 14485 7155
rect 14515 7125 14645 7155
rect 14675 7125 14805 7155
rect 14835 7125 14965 7155
rect 14995 7125 15000 7155
rect 14480 7120 15000 7125
rect 0 7075 520 7080
rect 0 7045 5 7075
rect 35 7045 165 7075
rect 195 7045 325 7075
rect 355 7045 485 7075
rect 515 7045 520 7075
rect 0 7040 520 7045
rect 14480 7075 15000 7080
rect 14480 7045 14485 7075
rect 14515 7045 14645 7075
rect 14675 7045 14805 7075
rect 14835 7045 14965 7075
rect 14995 7045 15000 7075
rect 14480 7040 15000 7045
rect 0 6995 520 7000
rect 0 6965 5 6995
rect 35 6965 165 6995
rect 195 6965 325 6995
rect 355 6965 485 6995
rect 515 6965 520 6995
rect 0 6960 520 6965
rect 14480 6995 15000 7000
rect 14480 6965 14485 6995
rect 14515 6965 14645 6995
rect 14675 6965 14805 6995
rect 14835 6965 14965 6995
rect 14995 6965 15000 6995
rect 14480 6960 15000 6965
rect 0 6915 520 6920
rect 0 6885 5 6915
rect 35 6885 165 6915
rect 195 6885 325 6915
rect 355 6885 485 6915
rect 515 6885 520 6915
rect 0 6880 520 6885
rect 14480 6915 15000 6920
rect 14480 6885 14485 6915
rect 14515 6885 14645 6915
rect 14675 6885 14805 6915
rect 14835 6885 14965 6915
rect 14995 6885 15000 6915
rect 14480 6880 15000 6885
rect 0 6835 520 6840
rect 0 6805 5 6835
rect 35 6805 165 6835
rect 195 6805 325 6835
rect 355 6805 485 6835
rect 515 6805 520 6835
rect 0 6800 520 6805
rect 14480 6835 15000 6840
rect 14480 6805 14485 6835
rect 14515 6805 14645 6835
rect 14675 6805 14805 6835
rect 14835 6805 14965 6835
rect 14995 6805 15000 6835
rect 14480 6800 15000 6805
rect 0 6755 520 6760
rect 0 6725 5 6755
rect 35 6725 165 6755
rect 195 6725 325 6755
rect 355 6725 485 6755
rect 515 6725 520 6755
rect 0 6720 520 6725
rect 14480 6755 15000 6760
rect 14480 6725 14485 6755
rect 14515 6725 14645 6755
rect 14675 6725 14805 6755
rect 14835 6725 14965 6755
rect 14995 6725 15000 6755
rect 14480 6720 15000 6725
rect 0 6675 520 6680
rect 0 6645 5 6675
rect 35 6645 165 6675
rect 195 6645 325 6675
rect 355 6645 485 6675
rect 515 6645 520 6675
rect 0 6640 520 6645
rect 14480 6675 15000 6680
rect 14480 6645 14485 6675
rect 14515 6645 14645 6675
rect 14675 6645 14805 6675
rect 14835 6645 14965 6675
rect 14995 6645 15000 6675
rect 14480 6640 15000 6645
rect 0 6595 360 6600
rect 0 6565 5 6595
rect 35 6565 165 6595
rect 195 6565 325 6595
rect 355 6565 360 6595
rect 0 6560 360 6565
rect 14480 6595 15000 6600
rect 14480 6565 14485 6595
rect 14515 6565 14645 6595
rect 14675 6565 14805 6595
rect 14835 6565 14965 6595
rect 14995 6565 15000 6595
rect 14480 6560 15000 6565
rect 0 6515 520 6520
rect 0 6485 5 6515
rect 35 6485 165 6515
rect 195 6485 325 6515
rect 355 6485 485 6515
rect 515 6485 520 6515
rect 0 6480 520 6485
rect 14480 6515 15000 6520
rect 14480 6485 14485 6515
rect 14515 6485 14645 6515
rect 14675 6485 14805 6515
rect 14835 6485 14965 6515
rect 14995 6485 15000 6515
rect 14480 6480 15000 6485
rect 0 6435 520 6440
rect 0 6405 5 6435
rect 35 6405 165 6435
rect 195 6405 325 6435
rect 355 6405 485 6435
rect 515 6405 520 6435
rect 0 6400 520 6405
rect 14480 6435 15000 6440
rect 14480 6405 14485 6435
rect 14515 6405 14645 6435
rect 14675 6405 14805 6435
rect 14835 6405 14965 6435
rect 14995 6405 15000 6435
rect 14480 6400 15000 6405
rect 0 6355 520 6360
rect 0 6325 5 6355
rect 35 6325 165 6355
rect 195 6325 325 6355
rect 355 6325 485 6355
rect 515 6325 520 6355
rect 0 6320 520 6325
rect 14480 6355 15000 6360
rect 14480 6325 14485 6355
rect 14515 6325 14645 6355
rect 14675 6325 14805 6355
rect 14835 6325 14965 6355
rect 14995 6325 15000 6355
rect 14480 6320 15000 6325
rect 0 6275 520 6280
rect 0 6245 5 6275
rect 35 6245 165 6275
rect 195 6245 325 6275
rect 355 6245 485 6275
rect 515 6245 520 6275
rect 0 6240 520 6245
rect 14480 6275 15000 6280
rect 14480 6245 14485 6275
rect 14515 6245 14645 6275
rect 14675 6245 14805 6275
rect 14835 6245 14965 6275
rect 14995 6245 15000 6275
rect 14480 6240 15000 6245
rect 0 6195 520 6200
rect 0 6165 5 6195
rect 35 6165 165 6195
rect 195 6165 325 6195
rect 355 6165 485 6195
rect 515 6165 520 6195
rect 0 6160 520 6165
rect 14480 6195 15000 6200
rect 14480 6165 14485 6195
rect 14515 6165 14645 6195
rect 14675 6165 14805 6195
rect 14835 6165 14965 6195
rect 14995 6165 15000 6195
rect 14480 6160 15000 6165
rect 0 6115 520 6120
rect 0 6085 5 6115
rect 35 6085 165 6115
rect 195 6085 325 6115
rect 355 6085 485 6115
rect 515 6085 520 6115
rect 0 6080 520 6085
rect 14480 6115 15000 6120
rect 14480 6085 14485 6115
rect 14515 6085 14645 6115
rect 14675 6085 14805 6115
rect 14835 6085 14965 6115
rect 14995 6085 15000 6115
rect 14480 6080 15000 6085
rect 0 6035 520 6040
rect 0 6005 5 6035
rect 35 6005 165 6035
rect 195 6005 325 6035
rect 355 6005 485 6035
rect 515 6005 520 6035
rect 0 6000 520 6005
rect 14480 6035 15000 6040
rect 14480 6005 14485 6035
rect 14515 6005 14645 6035
rect 14675 6005 14805 6035
rect 14835 6005 14965 6035
rect 14995 6005 15000 6035
rect 14480 6000 15000 6005
rect 0 5955 520 5960
rect 0 5925 5 5955
rect 35 5925 165 5955
rect 195 5925 325 5955
rect 355 5925 485 5955
rect 515 5925 520 5955
rect 0 5920 520 5925
rect 14480 5955 15000 5960
rect 14480 5925 14485 5955
rect 14515 5925 14645 5955
rect 14675 5925 14805 5955
rect 14835 5925 14965 5955
rect 14995 5925 15000 5955
rect 14480 5920 15000 5925
rect 0 5875 520 5880
rect 0 5845 5 5875
rect 35 5845 165 5875
rect 195 5845 325 5875
rect 355 5845 485 5875
rect 515 5845 520 5875
rect 0 5840 520 5845
rect 14480 5875 15000 5880
rect 14480 5845 14485 5875
rect 14515 5845 14645 5875
rect 14675 5845 14805 5875
rect 14835 5845 14965 5875
rect 14995 5845 15000 5875
rect 14480 5840 15000 5845
rect 0 5795 520 5800
rect 0 5765 5 5795
rect 35 5765 165 5795
rect 195 5765 325 5795
rect 355 5765 485 5795
rect 515 5765 520 5795
rect 0 5760 520 5765
rect 14480 5795 15000 5800
rect 14480 5765 14485 5795
rect 14515 5765 14645 5795
rect 14675 5765 14805 5795
rect 14835 5765 14965 5795
rect 14995 5765 15000 5795
rect 14480 5760 15000 5765
rect 0 5715 520 5720
rect 0 5685 5 5715
rect 35 5685 165 5715
rect 195 5685 325 5715
rect 355 5685 485 5715
rect 515 5685 520 5715
rect 0 5680 520 5685
rect 14480 5715 15000 5720
rect 14480 5685 14485 5715
rect 14515 5685 14645 5715
rect 14675 5685 14805 5715
rect 14835 5685 14965 5715
rect 14995 5685 15000 5715
rect 14480 5680 15000 5685
rect 0 5635 520 5640
rect 0 5605 5 5635
rect 35 5605 165 5635
rect 195 5605 325 5635
rect 355 5605 485 5635
rect 515 5605 520 5635
rect 0 5600 520 5605
rect 14480 5635 15000 5640
rect 14480 5605 14485 5635
rect 14515 5605 14645 5635
rect 14675 5605 14805 5635
rect 14835 5605 14965 5635
rect 14995 5605 15000 5635
rect 14480 5600 15000 5605
rect 0 5555 520 5560
rect 0 5525 5 5555
rect 35 5525 165 5555
rect 195 5525 325 5555
rect 355 5525 485 5555
rect 515 5525 520 5555
rect 0 5520 520 5525
rect 14480 5555 15000 5560
rect 14480 5525 14485 5555
rect 14515 5525 14645 5555
rect 14675 5525 14805 5555
rect 14835 5525 14965 5555
rect 14995 5525 15000 5555
rect 14480 5520 15000 5525
rect 0 5475 520 5480
rect 0 5445 5 5475
rect 35 5445 165 5475
rect 195 5445 325 5475
rect 355 5445 485 5475
rect 515 5445 520 5475
rect 0 5440 520 5445
rect 14480 5475 15000 5480
rect 14480 5445 14485 5475
rect 14515 5445 14645 5475
rect 14675 5445 14805 5475
rect 14835 5445 14965 5475
rect 14995 5445 15000 5475
rect 14480 5440 15000 5445
rect 0 5395 520 5400
rect 0 5365 5 5395
rect 35 5365 165 5395
rect 195 5365 325 5395
rect 355 5365 485 5395
rect 515 5365 520 5395
rect 0 5360 520 5365
rect 14480 5395 15000 5400
rect 14480 5365 14485 5395
rect 14515 5365 14645 5395
rect 14675 5365 14805 5395
rect 14835 5365 14965 5395
rect 14995 5365 15000 5395
rect 14480 5360 15000 5365
rect 0 5315 200 5320
rect 0 5285 5 5315
rect 35 5285 165 5315
rect 195 5285 200 5315
rect 0 5280 200 5285
rect 14480 5315 15000 5320
rect 14480 5285 14485 5315
rect 14515 5285 14645 5315
rect 14675 5285 14805 5315
rect 14835 5285 14965 5315
rect 14995 5285 15000 5315
rect 14480 5280 15000 5285
rect 0 5235 520 5240
rect 0 5205 5 5235
rect 35 5205 165 5235
rect 195 5205 325 5235
rect 355 5205 485 5235
rect 515 5205 520 5235
rect 0 5200 520 5205
rect 14480 5235 15000 5240
rect 14480 5205 14485 5235
rect 14515 5205 14645 5235
rect 14675 5205 14805 5235
rect 14835 5205 14965 5235
rect 14995 5205 15000 5235
rect 14480 5200 15000 5205
rect 14480 5155 15000 5160
rect 14480 5125 14485 5155
rect 14515 5125 14645 5155
rect 14675 5125 14805 5155
rect 14835 5125 14965 5155
rect 14995 5125 15000 5155
rect 14480 5120 15000 5125
rect 0 5075 520 5080
rect 0 5045 5 5075
rect 35 5045 165 5075
rect 195 5045 325 5075
rect 355 5045 485 5075
rect 515 5045 520 5075
rect 0 5040 520 5045
rect 14480 5075 15000 5080
rect 14480 5045 14485 5075
rect 14515 5045 14645 5075
rect 14675 5045 14805 5075
rect 14835 5045 14965 5075
rect 14995 5045 15000 5075
rect 14480 5040 15000 5045
rect 0 4995 520 5000
rect 0 4965 5 4995
rect 35 4965 165 4995
rect 195 4965 325 4995
rect 355 4965 485 4995
rect 515 4965 520 4995
rect 0 4960 520 4965
rect 14480 4995 15000 5000
rect 14480 4965 14485 4995
rect 14515 4965 14645 4995
rect 14675 4965 14805 4995
rect 14835 4965 14965 4995
rect 14995 4965 15000 4995
rect 14480 4960 15000 4965
rect 0 4915 520 4920
rect 0 4885 5 4915
rect 35 4885 165 4915
rect 195 4885 325 4915
rect 355 4885 485 4915
rect 515 4885 520 4915
rect 0 4880 520 4885
rect 14480 4915 15000 4920
rect 14480 4885 14485 4915
rect 14515 4885 14645 4915
rect 14675 4885 14805 4915
rect 14835 4885 14965 4915
rect 14995 4885 15000 4915
rect 14480 4880 15000 4885
rect 0 4835 520 4840
rect 0 4805 5 4835
rect 35 4805 165 4835
rect 195 4805 325 4835
rect 355 4805 485 4835
rect 515 4805 520 4835
rect 0 4800 520 4805
rect 14480 4835 15000 4840
rect 14480 4805 14485 4835
rect 14515 4805 14645 4835
rect 14675 4805 14805 4835
rect 14835 4805 14965 4835
rect 14995 4805 15000 4835
rect 14480 4800 15000 4805
rect 0 4755 520 4760
rect 0 4725 5 4755
rect 35 4725 165 4755
rect 195 4725 325 4755
rect 355 4725 485 4755
rect 515 4725 520 4755
rect 0 4720 520 4725
rect 0 4675 520 4680
rect 0 4645 5 4675
rect 35 4645 165 4675
rect 195 4645 325 4675
rect 355 4645 485 4675
rect 515 4645 520 4675
rect 0 4640 520 4645
rect 14480 4675 15000 4680
rect 14480 4645 14485 4675
rect 14515 4645 14645 4675
rect 14675 4645 14805 4675
rect 14835 4645 14965 4675
rect 14995 4645 15000 4675
rect 14480 4640 15000 4645
rect 0 4595 520 4600
rect 0 4565 5 4595
rect 35 4565 165 4595
rect 195 4565 325 4595
rect 355 4565 485 4595
rect 515 4565 520 4595
rect 0 4560 520 4565
rect 14800 4595 15000 4600
rect 14800 4565 14805 4595
rect 14835 4565 14965 4595
rect 14995 4565 15000 4595
rect 14800 4560 15000 4565
rect 0 4515 520 4520
rect 0 4485 5 4515
rect 35 4485 165 4515
rect 195 4485 325 4515
rect 355 4485 485 4515
rect 515 4485 520 4515
rect 0 4480 520 4485
rect 14480 4515 15000 4520
rect 14480 4485 14485 4515
rect 14515 4485 14645 4515
rect 14675 4485 14805 4515
rect 14835 4485 14965 4515
rect 14995 4485 15000 4515
rect 14480 4480 15000 4485
rect 0 4435 520 4440
rect 0 4405 5 4435
rect 35 4405 165 4435
rect 195 4405 325 4435
rect 355 4405 485 4435
rect 515 4405 520 4435
rect 0 4400 520 4405
rect 14480 4435 15000 4440
rect 14480 4405 14485 4435
rect 14515 4405 14645 4435
rect 14675 4405 14805 4435
rect 14835 4405 14965 4435
rect 14995 4405 15000 4435
rect 14480 4400 15000 4405
rect 0 4355 520 4360
rect 0 4325 5 4355
rect 35 4325 165 4355
rect 195 4325 325 4355
rect 355 4325 485 4355
rect 515 4325 520 4355
rect 0 4320 520 4325
rect 14480 4355 15000 4360
rect 14480 4325 14485 4355
rect 14515 4325 14645 4355
rect 14675 4325 14805 4355
rect 14835 4325 14965 4355
rect 14995 4325 15000 4355
rect 14480 4320 15000 4325
rect 0 4275 520 4280
rect 0 4245 5 4275
rect 35 4245 165 4275
rect 195 4245 325 4275
rect 355 4245 485 4275
rect 515 4245 520 4275
rect 0 4240 520 4245
rect 14480 4275 15000 4280
rect 14480 4245 14485 4275
rect 14515 4245 14645 4275
rect 14675 4245 14805 4275
rect 14835 4245 14965 4275
rect 14995 4245 15000 4275
rect 14480 4240 15000 4245
rect 0 4195 520 4200
rect 0 4165 5 4195
rect 35 4165 165 4195
rect 195 4165 325 4195
rect 355 4165 485 4195
rect 515 4165 520 4195
rect 0 4160 520 4165
rect 14480 4195 15000 4200
rect 14480 4165 14485 4195
rect 14515 4165 14645 4195
rect 14675 4165 14805 4195
rect 14835 4165 14965 4195
rect 14995 4165 15000 4195
rect 14480 4160 15000 4165
rect 0 4115 520 4120
rect 0 4085 5 4115
rect 35 4085 165 4115
rect 195 4085 325 4115
rect 355 4085 485 4115
rect 515 4085 520 4115
rect 0 4080 520 4085
rect 14480 4115 15000 4120
rect 14480 4085 14485 4115
rect 14515 4085 14645 4115
rect 14675 4085 14805 4115
rect 14835 4085 14965 4115
rect 14995 4085 15000 4115
rect 14480 4080 15000 4085
rect 0 4035 520 4040
rect 0 4005 5 4035
rect 35 4005 165 4035
rect 195 4005 325 4035
rect 355 4005 485 4035
rect 515 4005 520 4035
rect 0 4000 520 4005
rect 14480 4035 15000 4040
rect 14480 4005 14485 4035
rect 14515 4005 14645 4035
rect 14675 4005 14805 4035
rect 14835 4005 14965 4035
rect 14995 4005 15000 4035
rect 14480 4000 15000 4005
rect 0 3955 520 3960
rect 0 3925 5 3955
rect 35 3925 165 3955
rect 195 3925 325 3955
rect 355 3925 485 3955
rect 515 3925 520 3955
rect 0 3920 520 3925
rect 14480 3955 15000 3960
rect 14480 3925 14485 3955
rect 14515 3925 14645 3955
rect 14675 3925 14805 3955
rect 14835 3925 14965 3955
rect 14995 3925 15000 3955
rect 14480 3920 15000 3925
rect 0 3875 520 3880
rect 0 3845 5 3875
rect 35 3845 165 3875
rect 195 3845 325 3875
rect 355 3845 485 3875
rect 515 3845 520 3875
rect 0 3840 520 3845
rect 14480 3875 15000 3880
rect 14480 3845 14485 3875
rect 14515 3845 14645 3875
rect 14675 3845 14805 3875
rect 14835 3845 14965 3875
rect 14995 3845 15000 3875
rect 14480 3840 15000 3845
rect 0 3795 520 3800
rect 0 3765 5 3795
rect 35 3765 165 3795
rect 195 3765 325 3795
rect 355 3765 485 3795
rect 515 3765 520 3795
rect 0 3760 520 3765
rect 14480 3795 15000 3800
rect 14480 3765 14485 3795
rect 14515 3765 14645 3795
rect 14675 3765 14805 3795
rect 14835 3765 14965 3795
rect 14995 3765 15000 3795
rect 14480 3760 15000 3765
rect 0 3715 520 3720
rect 0 3685 5 3715
rect 35 3685 165 3715
rect 195 3685 325 3715
rect 355 3685 485 3715
rect 515 3685 520 3715
rect 0 3680 520 3685
rect 14480 3715 15000 3720
rect 14480 3685 14485 3715
rect 14515 3685 14645 3715
rect 14675 3685 14805 3715
rect 14835 3685 14965 3715
rect 14995 3685 15000 3715
rect 14480 3680 15000 3685
rect 0 3635 520 3640
rect 0 3605 5 3635
rect 35 3605 165 3635
rect 195 3605 325 3635
rect 355 3605 485 3635
rect 515 3605 520 3635
rect 0 3600 520 3605
rect 14480 3635 15000 3640
rect 14480 3605 14485 3635
rect 14515 3605 14645 3635
rect 14675 3605 14805 3635
rect 14835 3605 14965 3635
rect 14995 3605 15000 3635
rect 14480 3600 15000 3605
rect 0 3555 520 3560
rect 0 3525 5 3555
rect 35 3525 165 3555
rect 195 3525 325 3555
rect 355 3525 485 3555
rect 515 3525 520 3555
rect 0 3520 520 3525
rect 14480 3555 15000 3560
rect 14480 3525 14485 3555
rect 14515 3525 14645 3555
rect 14675 3525 14805 3555
rect 14835 3525 14965 3555
rect 14995 3525 15000 3555
rect 14480 3520 15000 3525
rect 0 3475 520 3480
rect 0 3445 5 3475
rect 35 3445 165 3475
rect 195 3445 325 3475
rect 355 3445 485 3475
rect 515 3445 520 3475
rect 0 3440 520 3445
rect 14480 3475 15000 3480
rect 14480 3445 14485 3475
rect 14515 3445 14645 3475
rect 14675 3445 14805 3475
rect 14835 3445 14965 3475
rect 14995 3445 15000 3475
rect 14480 3440 15000 3445
rect 0 3395 520 3400
rect 0 3365 5 3395
rect 35 3365 165 3395
rect 195 3365 325 3395
rect 355 3365 485 3395
rect 515 3365 520 3395
rect 0 3360 520 3365
rect 14480 3395 15000 3400
rect 14480 3365 14485 3395
rect 14515 3365 14645 3395
rect 14675 3365 14805 3395
rect 14835 3365 14965 3395
rect 14995 3365 15000 3395
rect 14480 3360 15000 3365
rect 0 3315 520 3320
rect 0 3285 5 3315
rect 35 3285 165 3315
rect 195 3285 325 3315
rect 355 3285 485 3315
rect 515 3285 520 3315
rect 0 3280 520 3285
rect 14640 3315 15000 3320
rect 14640 3285 14645 3315
rect 14675 3285 14805 3315
rect 14835 3285 14965 3315
rect 14995 3285 15000 3315
rect 14640 3280 15000 3285
rect 0 3235 520 3240
rect 0 3205 5 3235
rect 35 3205 165 3235
rect 195 3205 325 3235
rect 355 3205 485 3235
rect 515 3205 520 3235
rect 0 3200 520 3205
rect 14480 3235 15000 3240
rect 14480 3205 14485 3235
rect 14515 3205 14645 3235
rect 14675 3205 14805 3235
rect 14835 3205 14965 3235
rect 14995 3205 15000 3235
rect 14480 3200 15000 3205
rect 0 3155 520 3160
rect 0 3125 5 3155
rect 35 3125 165 3155
rect 195 3125 325 3155
rect 355 3125 485 3155
rect 515 3125 520 3155
rect 0 3120 520 3125
rect 14480 3155 15000 3160
rect 14480 3125 14485 3155
rect 14515 3125 14645 3155
rect 14675 3125 14805 3155
rect 14835 3125 14965 3155
rect 14995 3125 15000 3155
rect 14480 3120 15000 3125
rect 0 3075 520 3080
rect 0 3045 5 3075
rect 35 3045 165 3075
rect 195 3045 325 3075
rect 355 3045 485 3075
rect 515 3045 520 3075
rect 0 3040 520 3045
rect 14480 3075 15000 3080
rect 14480 3045 14485 3075
rect 14515 3045 14645 3075
rect 14675 3045 14805 3075
rect 14835 3045 14965 3075
rect 14995 3045 15000 3075
rect 14480 3040 15000 3045
rect 0 2995 520 3000
rect 0 2965 5 2995
rect 35 2965 165 2995
rect 195 2965 325 2995
rect 355 2965 485 2995
rect 515 2965 520 2995
rect 0 2960 520 2965
rect 14480 2995 15000 3000
rect 14480 2965 14485 2995
rect 14515 2965 14645 2995
rect 14675 2965 14805 2995
rect 14835 2965 14965 2995
rect 14995 2965 15000 2995
rect 14480 2960 15000 2965
rect 0 2915 520 2920
rect 0 2885 5 2915
rect 35 2885 165 2915
rect 195 2885 325 2915
rect 355 2885 485 2915
rect 515 2885 520 2915
rect 0 2880 520 2885
rect 14480 2915 15000 2920
rect 14480 2885 14485 2915
rect 14515 2885 14645 2915
rect 14675 2885 14805 2915
rect 14835 2885 14965 2915
rect 14995 2885 15000 2915
rect 14480 2880 15000 2885
rect 0 2835 520 2840
rect 0 2805 5 2835
rect 35 2805 165 2835
rect 195 2805 325 2835
rect 355 2805 485 2835
rect 515 2805 520 2835
rect 0 2800 520 2805
rect 14480 2835 15000 2840
rect 14480 2805 14485 2835
rect 14515 2805 14645 2835
rect 14675 2805 14805 2835
rect 14835 2805 14965 2835
rect 14995 2805 15000 2835
rect 14480 2800 15000 2805
rect 0 2755 520 2760
rect 0 2725 5 2755
rect 35 2725 165 2755
rect 195 2725 325 2755
rect 355 2725 485 2755
rect 515 2725 520 2755
rect 0 2720 520 2725
rect 14480 2755 15000 2760
rect 14480 2725 14485 2755
rect 14515 2725 14645 2755
rect 14675 2725 14805 2755
rect 14835 2725 14965 2755
rect 14995 2725 15000 2755
rect 14480 2720 15000 2725
rect 0 2675 520 2680
rect 0 2645 5 2675
rect 35 2645 165 2675
rect 195 2645 325 2675
rect 355 2645 485 2675
rect 515 2645 520 2675
rect 0 2640 520 2645
rect 14480 2675 15000 2680
rect 14480 2645 14485 2675
rect 14515 2645 14645 2675
rect 14675 2645 14805 2675
rect 14835 2645 14965 2675
rect 14995 2645 15000 2675
rect 14480 2640 15000 2645
rect 0 2595 520 2600
rect 0 2565 5 2595
rect 35 2565 165 2595
rect 195 2565 325 2595
rect 355 2565 485 2595
rect 515 2565 520 2595
rect 0 2560 520 2565
rect 14480 2595 15000 2600
rect 14480 2565 14485 2595
rect 14515 2565 14645 2595
rect 14675 2565 14805 2595
rect 14835 2565 14965 2595
rect 14995 2565 15000 2595
rect 14480 2560 15000 2565
rect 0 2515 520 2520
rect 0 2485 5 2515
rect 35 2485 165 2515
rect 195 2485 325 2515
rect 355 2485 485 2515
rect 515 2485 520 2515
rect 0 2480 520 2485
rect 14480 2515 15000 2520
rect 14480 2485 14485 2515
rect 14515 2485 14645 2515
rect 14675 2485 14805 2515
rect 14835 2485 14965 2515
rect 14995 2485 15000 2515
rect 14480 2480 15000 2485
rect 0 2435 520 2440
rect 0 2405 5 2435
rect 35 2405 165 2435
rect 195 2405 325 2435
rect 355 2405 485 2435
rect 515 2405 520 2435
rect 0 2400 520 2405
rect 14480 2435 15000 2440
rect 14480 2405 14485 2435
rect 14515 2405 14645 2435
rect 14675 2405 14805 2435
rect 14835 2405 14965 2435
rect 14995 2405 15000 2435
rect 14480 2400 15000 2405
rect 0 2355 520 2360
rect 0 2325 5 2355
rect 35 2325 165 2355
rect 195 2325 325 2355
rect 355 2325 485 2355
rect 515 2325 520 2355
rect 0 2320 520 2325
rect 14480 2355 15000 2360
rect 14480 2325 14485 2355
rect 14515 2325 14645 2355
rect 14675 2325 14805 2355
rect 14835 2325 14965 2355
rect 14995 2325 15000 2355
rect 14480 2320 15000 2325
rect 0 2275 520 2280
rect 0 2245 5 2275
rect 35 2245 165 2275
rect 195 2245 325 2275
rect 355 2245 485 2275
rect 515 2245 520 2275
rect 0 2240 520 2245
rect 14480 2275 15000 2280
rect 14480 2245 14485 2275
rect 14515 2245 14645 2275
rect 14675 2245 14805 2275
rect 14835 2245 14965 2275
rect 14995 2245 15000 2275
rect 14480 2240 15000 2245
rect 0 2195 520 2200
rect 0 2165 5 2195
rect 35 2165 165 2195
rect 195 2165 325 2195
rect 355 2165 485 2195
rect 515 2165 520 2195
rect 0 2160 520 2165
rect 14480 2195 15000 2200
rect 14480 2165 14485 2195
rect 14515 2165 14645 2195
rect 14675 2165 14805 2195
rect 14835 2165 14965 2195
rect 14995 2165 15000 2195
rect 14480 2160 15000 2165
rect 0 2115 520 2120
rect 0 2085 5 2115
rect 35 2085 165 2115
rect 195 2085 325 2115
rect 355 2085 485 2115
rect 515 2085 520 2115
rect 0 2080 520 2085
rect 14480 2115 15000 2120
rect 14480 2085 14485 2115
rect 14515 2085 14645 2115
rect 14675 2085 14805 2115
rect 14835 2085 14965 2115
rect 14995 2085 15000 2115
rect 14480 2080 15000 2085
rect 0 2035 520 2040
rect 0 2005 5 2035
rect 35 2005 165 2035
rect 195 2005 325 2035
rect 355 2005 485 2035
rect 515 2005 520 2035
rect 0 2000 520 2005
rect 14800 2035 15000 2040
rect 14800 2005 14805 2035
rect 14835 2005 14965 2035
rect 14995 2005 15000 2035
rect 14800 2000 15000 2005
rect 0 1955 520 1960
rect 0 1925 5 1955
rect 35 1925 165 1955
rect 195 1925 325 1955
rect 355 1925 485 1955
rect 515 1925 520 1955
rect 0 1920 520 1925
rect 14480 1955 15000 1960
rect 14480 1925 14485 1955
rect 14515 1925 14645 1955
rect 14675 1925 14805 1955
rect 14835 1925 14965 1955
rect 14995 1925 15000 1955
rect 14480 1920 15000 1925
rect 0 1875 520 1880
rect 0 1845 5 1875
rect 35 1845 165 1875
rect 195 1845 325 1875
rect 355 1845 485 1875
rect 515 1845 520 1875
rect 0 1840 520 1845
rect 0 1795 520 1800
rect 0 1765 5 1795
rect 35 1765 165 1795
rect 195 1765 325 1795
rect 355 1765 485 1795
rect 515 1765 520 1795
rect 0 1760 520 1765
rect 14480 1795 15000 1800
rect 14480 1765 14485 1795
rect 14515 1765 14645 1795
rect 14675 1765 14805 1795
rect 14835 1765 14965 1795
rect 14995 1765 15000 1795
rect 14480 1760 15000 1765
rect 0 1715 520 1720
rect 0 1685 5 1715
rect 35 1685 165 1715
rect 195 1685 325 1715
rect 355 1685 485 1715
rect 515 1685 520 1715
rect 0 1680 520 1685
rect 14480 1715 15000 1720
rect 14480 1685 14485 1715
rect 14515 1685 14645 1715
rect 14675 1685 14805 1715
rect 14835 1685 14965 1715
rect 14995 1685 15000 1715
rect 14480 1680 15000 1685
rect 0 1635 520 1640
rect 0 1605 5 1635
rect 35 1605 165 1635
rect 195 1605 325 1635
rect 355 1605 485 1635
rect 515 1605 520 1635
rect 0 1600 520 1605
rect 14480 1635 15000 1640
rect 14480 1605 14485 1635
rect 14515 1605 14645 1635
rect 14675 1605 14805 1635
rect 14835 1605 14965 1635
rect 14995 1605 15000 1635
rect 14480 1600 15000 1605
rect 0 1555 520 1560
rect 0 1525 5 1555
rect 35 1525 165 1555
rect 195 1525 325 1555
rect 355 1525 485 1555
rect 515 1525 520 1555
rect 0 1520 520 1525
rect 14480 1555 15000 1560
rect 14480 1525 14485 1555
rect 14515 1525 14645 1555
rect 14675 1525 14805 1555
rect 14835 1525 14965 1555
rect 14995 1525 15000 1555
rect 14480 1520 15000 1525
rect 0 1475 520 1480
rect 0 1445 5 1475
rect 35 1445 165 1475
rect 195 1445 325 1475
rect 355 1445 485 1475
rect 515 1445 520 1475
rect 0 1440 520 1445
rect 14480 1475 15000 1480
rect 14480 1445 14485 1475
rect 14515 1445 14645 1475
rect 14675 1445 14805 1475
rect 14835 1445 14965 1475
rect 14995 1445 15000 1475
rect 14480 1440 15000 1445
rect 0 1395 520 1400
rect 0 1365 5 1395
rect 35 1365 165 1395
rect 195 1365 325 1395
rect 355 1365 485 1395
rect 515 1365 520 1395
rect 0 1360 520 1365
rect 14480 1395 15000 1400
rect 14480 1365 14485 1395
rect 14515 1365 14645 1395
rect 14675 1365 14805 1395
rect 14835 1365 14965 1395
rect 14995 1365 15000 1395
rect 14480 1360 15000 1365
rect 0 1315 520 1320
rect 0 1285 5 1315
rect 35 1285 165 1315
rect 195 1285 325 1315
rect 355 1285 485 1315
rect 515 1285 520 1315
rect 0 1280 520 1285
rect 14480 1315 15000 1320
rect 14480 1285 14485 1315
rect 14515 1285 14645 1315
rect 14675 1285 14805 1315
rect 14835 1285 14965 1315
rect 14995 1285 15000 1315
rect 14480 1280 15000 1285
rect 0 1235 520 1240
rect 0 1205 5 1235
rect 35 1205 165 1235
rect 195 1205 325 1235
rect 355 1205 485 1235
rect 515 1205 520 1235
rect 0 1200 520 1205
rect 14480 1235 15000 1240
rect 14480 1205 14485 1235
rect 14515 1205 14645 1235
rect 14675 1205 14805 1235
rect 14835 1205 14965 1235
rect 14995 1205 15000 1235
rect 14480 1200 15000 1205
rect 0 1155 520 1160
rect 0 1125 5 1155
rect 35 1125 165 1155
rect 195 1125 325 1155
rect 355 1125 485 1155
rect 515 1125 520 1155
rect 0 1120 520 1125
rect 14480 1155 15000 1160
rect 14480 1125 14485 1155
rect 14515 1125 14645 1155
rect 14675 1125 14805 1155
rect 14835 1125 14965 1155
rect 14995 1125 15000 1155
rect 14480 1120 15000 1125
rect 0 1075 520 1080
rect 0 1045 5 1075
rect 35 1045 165 1075
rect 195 1045 325 1075
rect 355 1045 485 1075
rect 515 1045 520 1075
rect 0 1040 520 1045
rect 14480 1075 15000 1080
rect 14480 1045 14485 1075
rect 14515 1045 14645 1075
rect 14675 1045 14805 1075
rect 14835 1045 14965 1075
rect 14995 1045 15000 1075
rect 14480 1040 15000 1045
rect 0 995 520 1000
rect 0 965 5 995
rect 35 965 165 995
rect 195 965 325 995
rect 355 965 485 995
rect 515 965 520 995
rect 0 960 520 965
rect 14480 995 15000 1000
rect 14480 965 14485 995
rect 14515 965 14645 995
rect 14675 965 14805 995
rect 14835 965 14965 995
rect 14995 965 15000 995
rect 14480 960 15000 965
rect 0 915 520 920
rect 0 885 5 915
rect 35 885 165 915
rect 195 885 325 915
rect 355 885 485 915
rect 515 885 520 915
rect 0 880 520 885
rect 14480 915 15000 920
rect 14480 885 14485 915
rect 14515 885 14645 915
rect 14675 885 14805 915
rect 14835 885 14965 915
rect 14995 885 15000 915
rect 14480 880 15000 885
rect 0 835 520 840
rect 0 805 5 835
rect 35 805 165 835
rect 195 805 325 835
rect 355 805 485 835
rect 515 805 520 835
rect 0 800 520 805
rect 14480 835 15000 840
rect 14480 805 14485 835
rect 14515 805 14645 835
rect 14675 805 14805 835
rect 14835 805 14965 835
rect 14995 805 15000 835
rect 14480 800 15000 805
rect 0 755 520 760
rect 0 725 5 755
rect 35 725 165 755
rect 195 725 325 755
rect 355 725 485 755
rect 515 725 520 755
rect 0 720 520 725
rect 14480 755 15000 760
rect 14480 725 14485 755
rect 14515 725 14645 755
rect 14675 725 14805 755
rect 14835 725 14965 755
rect 14995 725 15000 755
rect 14480 720 15000 725
rect 0 675 520 680
rect 0 645 5 675
rect 35 645 165 675
rect 195 645 325 675
rect 355 645 485 675
rect 515 645 520 675
rect 0 640 520 645
rect 14480 675 15000 680
rect 14480 645 14485 675
rect 14515 645 14645 675
rect 14675 645 14805 675
rect 14835 645 14965 675
rect 14995 645 15000 675
rect 14480 640 15000 645
rect 0 595 520 600
rect 0 565 5 595
rect 35 565 165 595
rect 195 565 325 595
rect 355 565 485 595
rect 515 565 520 595
rect 0 560 520 565
rect 14480 595 15000 600
rect 14480 565 14485 595
rect 14515 565 14645 595
rect 14675 565 14805 595
rect 14835 565 14965 595
rect 14995 565 15000 595
rect 14480 560 15000 565
rect 0 515 520 520
rect 0 485 5 515
rect 35 485 165 515
rect 195 485 325 515
rect 355 485 485 515
rect 515 485 520 515
rect 0 480 520 485
rect 560 515 600 520
rect 560 485 565 515
rect 595 485 600 515
rect 560 480 600 485
rect 14400 515 14440 520
rect 14400 485 14405 515
rect 14435 485 14440 515
rect 14400 480 14440 485
rect 14480 515 15000 520
rect 14480 485 14485 515
rect 14515 485 14645 515
rect 14675 485 14805 515
rect 14835 485 14965 515
rect 14995 485 15000 515
rect 14480 480 15000 485
<< via2 >>
rect 5 15925 35 15955
rect 165 15925 195 15955
rect 325 15925 355 15955
rect 485 15925 515 15955
rect 14485 15925 14515 15955
rect 14645 15925 14675 15955
rect 14805 15925 14835 15955
rect 14965 15925 14995 15955
rect 5 15845 35 15875
rect 165 15845 195 15875
rect 325 15845 355 15875
rect 485 15845 515 15875
rect 14485 15845 14515 15875
rect 14645 15845 14675 15875
rect 14805 15845 14835 15875
rect 14965 15845 14995 15875
rect 5 15765 35 15795
rect 165 15765 195 15795
rect 325 15765 355 15795
rect 485 15765 515 15795
rect 14485 15765 14515 15795
rect 14645 15765 14675 15795
rect 14805 15765 14835 15795
rect 14965 15765 14995 15795
rect 5 15685 35 15715
rect 165 15685 195 15715
rect 325 15685 355 15715
rect 485 15685 515 15715
rect 14485 15685 14515 15715
rect 14645 15685 14675 15715
rect 14805 15685 14835 15715
rect 14965 15685 14995 15715
rect 5 15605 35 15635
rect 165 15605 195 15635
rect 325 15605 355 15635
rect 485 15605 515 15635
rect 14485 15605 14515 15635
rect 14645 15605 14675 15635
rect 14805 15605 14835 15635
rect 14965 15605 14995 15635
rect 5 15525 35 15555
rect 165 15525 195 15555
rect 325 15525 355 15555
rect 485 15525 515 15555
rect 14485 15525 14515 15555
rect 14645 15525 14675 15555
rect 14805 15525 14835 15555
rect 14965 15525 14995 15555
rect 5 15445 35 15475
rect 165 15445 195 15475
rect 325 15445 355 15475
rect 485 15445 515 15475
rect 14485 15445 14515 15475
rect 14645 15445 14675 15475
rect 14805 15445 14835 15475
rect 14965 15445 14995 15475
rect 5 15365 35 15395
rect 165 15365 195 15395
rect 325 15365 355 15395
rect 485 15365 515 15395
rect 14485 15365 14515 15395
rect 14645 15365 14675 15395
rect 14805 15365 14835 15395
rect 14965 15365 14995 15395
rect 5 15285 35 15315
rect 165 15285 195 15315
rect 325 15285 355 15315
rect 485 15285 515 15315
rect 14485 15285 14515 15315
rect 14645 15285 14675 15315
rect 14805 15285 14835 15315
rect 14965 15285 14995 15315
rect 5 15205 35 15235
rect 165 15205 195 15235
rect 325 15205 355 15235
rect 485 15205 515 15235
rect 14485 15205 14515 15235
rect 14645 15205 14675 15235
rect 14805 15205 14835 15235
rect 14965 15205 14995 15235
rect 5 15125 35 15155
rect 165 15125 195 15155
rect 325 15125 355 15155
rect 485 15125 515 15155
rect 14485 15125 14515 15155
rect 14645 15125 14675 15155
rect 14805 15125 14835 15155
rect 14965 15125 14995 15155
rect 5 15045 35 15075
rect 165 15045 195 15075
rect 325 15045 355 15075
rect 485 15045 515 15075
rect 14485 15045 14515 15075
rect 14645 15045 14675 15075
rect 14805 15045 14835 15075
rect 14965 15045 14995 15075
rect 5 14965 35 14995
rect 165 14965 195 14995
rect 325 14965 355 14995
rect 485 14965 515 14995
rect 14485 14965 14515 14995
rect 14645 14965 14675 14995
rect 14805 14965 14835 14995
rect 14965 14965 14995 14995
rect 5 14885 35 14915
rect 165 14885 195 14915
rect 325 14885 355 14915
rect 485 14885 515 14915
rect 14485 14885 14515 14915
rect 14645 14885 14675 14915
rect 14805 14885 14835 14915
rect 14965 14885 14995 14915
rect 5 14805 35 14835
rect 165 14805 195 14835
rect 325 14805 355 14835
rect 485 14805 515 14835
rect 14485 14805 14515 14835
rect 14645 14805 14675 14835
rect 14805 14805 14835 14835
rect 14965 14805 14995 14835
rect 5 14725 35 14755
rect 165 14725 195 14755
rect 325 14725 355 14755
rect 485 14725 515 14755
rect 14485 14725 14515 14755
rect 14645 14725 14675 14755
rect 14805 14725 14835 14755
rect 14965 14725 14995 14755
rect 5 14645 35 14675
rect 165 14645 195 14675
rect 325 14645 355 14675
rect 485 14645 515 14675
rect 14485 14645 14515 14675
rect 14645 14645 14675 14675
rect 14805 14645 14835 14675
rect 14965 14645 14995 14675
rect 5 14565 35 14595
rect 165 14565 195 14595
rect 325 14565 355 14595
rect 485 14565 515 14595
rect 5 14485 35 14515
rect 165 14485 195 14515
rect 325 14485 355 14515
rect 485 14485 515 14515
rect 14485 14485 14515 14515
rect 14645 14485 14675 14515
rect 14805 14485 14835 14515
rect 14965 14485 14995 14515
rect 5 14405 35 14435
rect 165 14405 195 14435
rect 325 14405 355 14435
rect 485 14405 515 14435
rect 14805 14405 14835 14435
rect 14965 14405 14995 14435
rect 5 14325 35 14355
rect 165 14325 195 14355
rect 325 14325 355 14355
rect 485 14325 515 14355
rect 14485 14325 14515 14355
rect 14645 14325 14675 14355
rect 14805 14325 14835 14355
rect 14965 14325 14995 14355
rect 5 14245 35 14275
rect 165 14245 195 14275
rect 325 14245 355 14275
rect 485 14245 515 14275
rect 14485 14245 14515 14275
rect 14645 14245 14675 14275
rect 14805 14245 14835 14275
rect 14965 14245 14995 14275
rect 5 14165 35 14195
rect 165 14165 195 14195
rect 325 14165 355 14195
rect 485 14165 515 14195
rect 14485 14165 14515 14195
rect 14645 14165 14675 14195
rect 14805 14165 14835 14195
rect 14965 14165 14995 14195
rect 5 14085 35 14115
rect 165 14085 195 14115
rect 325 14085 355 14115
rect 485 14085 515 14115
rect 14485 14085 14515 14115
rect 14645 14085 14675 14115
rect 14805 14085 14835 14115
rect 14965 14085 14995 14115
rect 5 14005 35 14035
rect 165 14005 195 14035
rect 325 14005 355 14035
rect 485 14005 515 14035
rect 14485 14005 14515 14035
rect 14645 14005 14675 14035
rect 14805 14005 14835 14035
rect 14965 14005 14995 14035
rect 5 13925 35 13955
rect 165 13925 195 13955
rect 325 13925 355 13955
rect 485 13925 515 13955
rect 14485 13925 14515 13955
rect 14645 13925 14675 13955
rect 14805 13925 14835 13955
rect 14965 13925 14995 13955
rect 5 13845 35 13875
rect 165 13845 195 13875
rect 325 13845 355 13875
rect 485 13845 515 13875
rect 14485 13845 14515 13875
rect 14645 13845 14675 13875
rect 14805 13845 14835 13875
rect 14965 13845 14995 13875
rect 5 13765 35 13795
rect 165 13765 195 13795
rect 325 13765 355 13795
rect 485 13765 515 13795
rect 14485 13765 14515 13795
rect 14645 13765 14675 13795
rect 14805 13765 14835 13795
rect 14965 13765 14995 13795
rect 5 13685 35 13715
rect 165 13685 195 13715
rect 325 13685 355 13715
rect 485 13685 515 13715
rect 14485 13685 14515 13715
rect 14645 13685 14675 13715
rect 14805 13685 14835 13715
rect 14965 13685 14995 13715
rect 5 13605 35 13635
rect 165 13605 195 13635
rect 325 13605 355 13635
rect 485 13605 515 13635
rect 14485 13605 14515 13635
rect 14645 13605 14675 13635
rect 14805 13605 14835 13635
rect 14965 13605 14995 13635
rect 5 13525 35 13555
rect 165 13525 195 13555
rect 325 13525 355 13555
rect 485 13525 515 13555
rect 14485 13525 14515 13555
rect 14645 13525 14675 13555
rect 14805 13525 14835 13555
rect 14965 13525 14995 13555
rect 5 13445 35 13475
rect 165 13445 195 13475
rect 325 13445 355 13475
rect 485 13445 515 13475
rect 14485 13445 14515 13475
rect 14645 13445 14675 13475
rect 14805 13445 14835 13475
rect 14965 13445 14995 13475
rect 5 13365 35 13395
rect 165 13365 195 13395
rect 325 13365 355 13395
rect 485 13365 515 13395
rect 14485 13365 14515 13395
rect 14645 13365 14675 13395
rect 14805 13365 14835 13395
rect 14965 13365 14995 13395
rect 5 13285 35 13315
rect 165 13285 195 13315
rect 325 13285 355 13315
rect 485 13285 515 13315
rect 14485 13285 14515 13315
rect 14645 13285 14675 13315
rect 14805 13285 14835 13315
rect 14965 13285 14995 13315
rect 5 13205 35 13235
rect 165 13205 195 13235
rect 325 13205 355 13235
rect 485 13205 515 13235
rect 14485 13205 14515 13235
rect 14645 13205 14675 13235
rect 14805 13205 14835 13235
rect 14965 13205 14995 13235
rect 5 13125 35 13155
rect 165 13125 195 13155
rect 325 13125 355 13155
rect 485 13125 515 13155
rect 14645 13125 14675 13155
rect 14805 13125 14835 13155
rect 14965 13125 14995 13155
rect 5 13045 35 13075
rect 165 13045 195 13075
rect 325 13045 355 13075
rect 485 13045 515 13075
rect 14485 13045 14515 13075
rect 14645 13045 14675 13075
rect 14805 13045 14835 13075
rect 14965 13045 14995 13075
rect 5 12965 35 12995
rect 165 12965 195 12995
rect 325 12965 355 12995
rect 485 12965 515 12995
rect 14485 12965 14515 12995
rect 14645 12965 14675 12995
rect 14805 12965 14835 12995
rect 14965 12965 14995 12995
rect 5 12885 35 12915
rect 165 12885 195 12915
rect 325 12885 355 12915
rect 485 12885 515 12915
rect 14485 12885 14515 12915
rect 14645 12885 14675 12915
rect 14805 12885 14835 12915
rect 14965 12885 14995 12915
rect 5 12805 35 12835
rect 165 12805 195 12835
rect 325 12805 355 12835
rect 485 12805 515 12835
rect 14485 12805 14515 12835
rect 14645 12805 14675 12835
rect 14805 12805 14835 12835
rect 14965 12805 14995 12835
rect 5 12725 35 12755
rect 165 12725 195 12755
rect 325 12725 355 12755
rect 485 12725 515 12755
rect 14485 12725 14515 12755
rect 14645 12725 14675 12755
rect 14805 12725 14835 12755
rect 14965 12725 14995 12755
rect 5 12645 35 12675
rect 165 12645 195 12675
rect 325 12645 355 12675
rect 485 12645 515 12675
rect 14485 12645 14515 12675
rect 14645 12645 14675 12675
rect 14805 12645 14835 12675
rect 14965 12645 14995 12675
rect 5 12565 35 12595
rect 165 12565 195 12595
rect 325 12565 355 12595
rect 485 12565 515 12595
rect 14485 12565 14515 12595
rect 14645 12565 14675 12595
rect 14805 12565 14835 12595
rect 14965 12565 14995 12595
rect 5 12485 35 12515
rect 165 12485 195 12515
rect 325 12485 355 12515
rect 485 12485 515 12515
rect 14485 12485 14515 12515
rect 14645 12485 14675 12515
rect 14805 12485 14835 12515
rect 14965 12485 14995 12515
rect 5 12405 35 12435
rect 165 12405 195 12435
rect 325 12405 355 12435
rect 485 12405 515 12435
rect 14485 12405 14515 12435
rect 14645 12405 14675 12435
rect 14805 12405 14835 12435
rect 14965 12405 14995 12435
rect 5 12325 35 12355
rect 165 12325 195 12355
rect 325 12325 355 12355
rect 485 12325 515 12355
rect 14485 12325 14515 12355
rect 14645 12325 14675 12355
rect 14805 12325 14835 12355
rect 14965 12325 14995 12355
rect 5 12245 35 12275
rect 165 12245 195 12275
rect 325 12245 355 12275
rect 485 12245 515 12275
rect 14485 12245 14515 12275
rect 14645 12245 14675 12275
rect 14805 12245 14835 12275
rect 14965 12245 14995 12275
rect 5 12165 35 12195
rect 165 12165 195 12195
rect 325 12165 355 12195
rect 485 12165 515 12195
rect 14485 12165 14515 12195
rect 14645 12165 14675 12195
rect 14805 12165 14835 12195
rect 14965 12165 14995 12195
rect 5 12085 35 12115
rect 165 12085 195 12115
rect 325 12085 355 12115
rect 485 12085 515 12115
rect 14485 12085 14515 12115
rect 14645 12085 14675 12115
rect 14805 12085 14835 12115
rect 14965 12085 14995 12115
rect 5 12005 35 12035
rect 165 12005 195 12035
rect 325 12005 355 12035
rect 485 12005 515 12035
rect 14485 12005 14515 12035
rect 14645 12005 14675 12035
rect 14805 12005 14835 12035
rect 14965 12005 14995 12035
rect 5 11925 35 11955
rect 165 11925 195 11955
rect 325 11925 355 11955
rect 485 11925 515 11955
rect 14485 11925 14515 11955
rect 14645 11925 14675 11955
rect 14805 11925 14835 11955
rect 14965 11925 14995 11955
rect 5 11845 35 11875
rect 165 11845 195 11875
rect 325 11845 355 11875
rect 485 11845 515 11875
rect 14805 11845 14835 11875
rect 14965 11845 14995 11875
rect 5 11765 35 11795
rect 165 11765 195 11795
rect 325 11765 355 11795
rect 485 11765 515 11795
rect 14485 11765 14515 11795
rect 14645 11765 14675 11795
rect 14805 11765 14835 11795
rect 14965 11765 14995 11795
rect 5 11685 35 11715
rect 165 11685 195 11715
rect 325 11685 355 11715
rect 485 11685 515 11715
rect 5 11605 35 11635
rect 165 11605 195 11635
rect 325 11605 355 11635
rect 485 11605 515 11635
rect 14485 11605 14515 11635
rect 14645 11605 14675 11635
rect 14805 11605 14835 11635
rect 14965 11605 14995 11635
rect 5 11525 35 11555
rect 165 11525 195 11555
rect 325 11525 355 11555
rect 485 11525 515 11555
rect 14485 11525 14515 11555
rect 14645 11525 14675 11555
rect 14805 11525 14835 11555
rect 14965 11525 14995 11555
rect 5 11445 35 11475
rect 165 11445 195 11475
rect 325 11445 355 11475
rect 485 11445 515 11475
rect 14485 11445 14515 11475
rect 14645 11445 14675 11475
rect 14805 11445 14835 11475
rect 14965 11445 14995 11475
rect 5 11365 35 11395
rect 165 11365 195 11395
rect 325 11365 355 11395
rect 485 11365 515 11395
rect 14485 11365 14515 11395
rect 14645 11365 14675 11395
rect 14805 11365 14835 11395
rect 14965 11365 14995 11395
rect 14485 11285 14515 11315
rect 14645 11285 14675 11315
rect 14805 11285 14835 11315
rect 14965 11285 14995 11315
rect 5 11205 35 11235
rect 165 11205 195 11235
rect 325 11205 355 11235
rect 485 11205 515 11235
rect 14485 11205 14515 11235
rect 14645 11205 14675 11235
rect 14805 11205 14835 11235
rect 14965 11205 14995 11235
rect 5 11125 35 11155
rect 165 11125 195 11155
rect 14485 11125 14515 11155
rect 14645 11125 14675 11155
rect 14805 11125 14835 11155
rect 14965 11125 14995 11155
rect 5 11045 35 11075
rect 165 11045 195 11075
rect 325 11045 355 11075
rect 485 11045 515 11075
rect 14485 11045 14515 11075
rect 14645 11045 14675 11075
rect 14805 11045 14835 11075
rect 14965 11045 14995 11075
rect 5 10965 35 10995
rect 165 10965 195 10995
rect 325 10965 355 10995
rect 485 10965 515 10995
rect 14485 10965 14515 10995
rect 14645 10965 14675 10995
rect 14805 10965 14835 10995
rect 14965 10965 14995 10995
rect 5 10885 35 10915
rect 165 10885 195 10915
rect 325 10885 355 10915
rect 485 10885 515 10915
rect 14485 10885 14515 10915
rect 14645 10885 14675 10915
rect 14805 10885 14835 10915
rect 14965 10885 14995 10915
rect 5 10805 35 10835
rect 165 10805 195 10835
rect 325 10805 355 10835
rect 485 10805 515 10835
rect 14485 10805 14515 10835
rect 14645 10805 14675 10835
rect 14805 10805 14835 10835
rect 14965 10805 14995 10835
rect 5 10725 35 10755
rect 165 10725 195 10755
rect 325 10725 355 10755
rect 485 10725 515 10755
rect 14485 10725 14515 10755
rect 14645 10725 14675 10755
rect 14805 10725 14835 10755
rect 14965 10725 14995 10755
rect 5 10645 35 10675
rect 165 10645 195 10675
rect 325 10645 355 10675
rect 485 10645 515 10675
rect 14485 10645 14515 10675
rect 14645 10645 14675 10675
rect 14805 10645 14835 10675
rect 14965 10645 14995 10675
rect 5 10565 35 10595
rect 165 10565 195 10595
rect 325 10565 355 10595
rect 485 10565 515 10595
rect 14485 10565 14515 10595
rect 14645 10565 14675 10595
rect 14805 10565 14835 10595
rect 14965 10565 14995 10595
rect 5 10485 35 10515
rect 165 10485 195 10515
rect 325 10485 355 10515
rect 485 10485 515 10515
rect 14485 10485 14515 10515
rect 14645 10485 14675 10515
rect 14805 10485 14835 10515
rect 14965 10485 14995 10515
rect 5 10405 35 10435
rect 165 10405 195 10435
rect 325 10405 355 10435
rect 485 10405 515 10435
rect 14485 10405 14515 10435
rect 14645 10405 14675 10435
rect 14805 10405 14835 10435
rect 14965 10405 14995 10435
rect 5 10325 35 10355
rect 165 10325 195 10355
rect 325 10325 355 10355
rect 485 10325 515 10355
rect 14485 10325 14515 10355
rect 14645 10325 14675 10355
rect 14805 10325 14835 10355
rect 14965 10325 14995 10355
rect 5 10245 35 10275
rect 165 10245 195 10275
rect 325 10245 355 10275
rect 485 10245 515 10275
rect 14485 10245 14515 10275
rect 14645 10245 14675 10275
rect 14805 10245 14835 10275
rect 14965 10245 14995 10275
rect 5 10165 35 10195
rect 165 10165 195 10195
rect 325 10165 355 10195
rect 485 10165 515 10195
rect 14485 10165 14515 10195
rect 14645 10165 14675 10195
rect 14805 10165 14835 10195
rect 14965 10165 14995 10195
rect 5 10085 35 10115
rect 165 10085 195 10115
rect 325 10085 355 10115
rect 485 10085 515 10115
rect 14485 10085 14515 10115
rect 14645 10085 14675 10115
rect 14805 10085 14835 10115
rect 14965 10085 14995 10115
rect 5 10005 35 10035
rect 165 10005 195 10035
rect 325 10005 355 10035
rect 485 10005 515 10035
rect 14485 10005 14515 10035
rect 14645 10005 14675 10035
rect 14805 10005 14835 10035
rect 14965 10005 14995 10035
rect 5 9925 35 9955
rect 165 9925 195 9955
rect 325 9925 355 9955
rect 485 9925 515 9955
rect 14485 9925 14515 9955
rect 14645 9925 14675 9955
rect 14805 9925 14835 9955
rect 14965 9925 14995 9955
rect 5 9845 35 9875
rect 165 9845 195 9875
rect 325 9845 355 9875
rect 14485 9845 14515 9875
rect 14645 9845 14675 9875
rect 14805 9845 14835 9875
rect 14965 9845 14995 9875
rect 5 9765 35 9795
rect 165 9765 195 9795
rect 325 9765 355 9795
rect 485 9765 515 9795
rect 14485 9765 14515 9795
rect 14645 9765 14675 9795
rect 14805 9765 14835 9795
rect 14965 9765 14995 9795
rect 5 9685 35 9715
rect 165 9685 195 9715
rect 325 9685 355 9715
rect 485 9685 515 9715
rect 14485 9685 14515 9715
rect 14645 9685 14675 9715
rect 14805 9685 14835 9715
rect 14965 9685 14995 9715
rect 5 9605 35 9635
rect 165 9605 195 9635
rect 325 9605 355 9635
rect 485 9605 515 9635
rect 14485 9605 14515 9635
rect 14645 9605 14675 9635
rect 14805 9605 14835 9635
rect 14965 9605 14995 9635
rect 5 9525 35 9555
rect 165 9525 195 9555
rect 325 9525 355 9555
rect 485 9525 515 9555
rect 14485 9525 14515 9555
rect 14645 9525 14675 9555
rect 14805 9525 14835 9555
rect 14965 9525 14995 9555
rect 5 9445 35 9475
rect 165 9445 195 9475
rect 325 9445 355 9475
rect 485 9445 515 9475
rect 14485 9445 14515 9475
rect 14645 9445 14675 9475
rect 14805 9445 14835 9475
rect 14965 9445 14995 9475
rect 5 9365 35 9395
rect 165 9365 195 9395
rect 325 9365 355 9395
rect 485 9365 515 9395
rect 14485 9365 14515 9395
rect 14645 9365 14675 9395
rect 14805 9365 14835 9395
rect 14965 9365 14995 9395
rect 5 9285 35 9315
rect 165 9285 195 9315
rect 325 9285 355 9315
rect 485 9285 515 9315
rect 14485 9285 14515 9315
rect 14645 9285 14675 9315
rect 14805 9285 14835 9315
rect 14965 9285 14995 9315
rect 5 9205 35 9235
rect 165 9205 195 9235
rect 325 9205 355 9235
rect 485 9205 515 9235
rect 14485 9205 14515 9235
rect 14645 9205 14675 9235
rect 14805 9205 14835 9235
rect 14965 9205 14995 9235
rect 5 9125 35 9155
rect 165 9125 195 9155
rect 325 9125 355 9155
rect 485 9125 515 9155
rect 14485 9125 14515 9155
rect 14645 9125 14675 9155
rect 14805 9125 14835 9155
rect 14965 9125 14995 9155
rect 5 9045 35 9075
rect 165 9045 195 9075
rect 325 9045 355 9075
rect 485 9045 515 9075
rect 14485 9045 14515 9075
rect 14645 9045 14675 9075
rect 14805 9045 14835 9075
rect 14965 9045 14995 9075
rect 5 8965 35 8995
rect 165 8965 195 8995
rect 325 8965 355 8995
rect 485 8965 515 8995
rect 14485 8965 14515 8995
rect 14645 8965 14675 8995
rect 14805 8965 14835 8995
rect 14965 8965 14995 8995
rect 5 8885 35 8915
rect 165 8885 195 8915
rect 325 8885 355 8915
rect 485 8885 515 8915
rect 14485 8885 14515 8915
rect 14645 8885 14675 8915
rect 14805 8885 14835 8915
rect 14965 8885 14995 8915
rect 5 8805 35 8835
rect 165 8805 195 8835
rect 325 8805 355 8835
rect 485 8805 515 8835
rect 14485 8805 14515 8835
rect 14645 8805 14675 8835
rect 14805 8805 14835 8835
rect 14965 8805 14995 8835
rect 5 8725 35 8755
rect 165 8725 195 8755
rect 325 8725 355 8755
rect 485 8725 515 8755
rect 14485 8725 14515 8755
rect 14645 8725 14675 8755
rect 14805 8725 14835 8755
rect 14965 8725 14995 8755
rect 5 8645 35 8675
rect 165 8645 195 8675
rect 325 8645 355 8675
rect 485 8645 515 8675
rect 14485 8645 14515 8675
rect 14645 8645 14675 8675
rect 14805 8645 14835 8675
rect 14965 8645 14995 8675
rect 5 8565 35 8595
rect 165 8565 195 8595
rect 14485 8565 14515 8595
rect 14645 8565 14675 8595
rect 14805 8565 14835 8595
rect 14965 8565 14995 8595
rect 5 8485 35 8515
rect 165 8485 195 8515
rect 325 8485 355 8515
rect 485 8485 515 8515
rect 14485 8485 14515 8515
rect 14645 8485 14675 8515
rect 14805 8485 14835 8515
rect 14965 8485 14995 8515
rect 14485 8405 14515 8435
rect 14645 8405 14675 8435
rect 14805 8405 14835 8435
rect 14965 8405 14995 8435
rect 5 8325 35 8355
rect 165 8325 195 8355
rect 325 8325 355 8355
rect 485 8325 515 8355
rect 14485 8325 14515 8355
rect 14645 8325 14675 8355
rect 14805 8325 14835 8355
rect 14965 8325 14995 8355
rect 5 8245 35 8275
rect 165 8245 195 8275
rect 325 8245 355 8275
rect 485 8245 515 8275
rect 14485 8245 14515 8275
rect 14645 8245 14675 8275
rect 14805 8245 14835 8275
rect 14965 8245 14995 8275
rect 5 8165 35 8195
rect 165 8165 195 8195
rect 325 8165 355 8195
rect 485 8165 515 8195
rect 14485 8165 14515 8195
rect 14645 8165 14675 8195
rect 14805 8165 14835 8195
rect 14965 8165 14995 8195
rect 5 8085 35 8115
rect 165 8085 195 8115
rect 325 8085 355 8115
rect 485 8085 515 8115
rect 14485 8085 14515 8115
rect 14645 8085 14675 8115
rect 14805 8085 14835 8115
rect 14965 8085 14995 8115
rect 14485 8005 14515 8035
rect 14645 8005 14675 8035
rect 14805 8005 14835 8035
rect 14965 8005 14995 8035
rect 5 7925 35 7955
rect 165 7925 195 7955
rect 325 7925 355 7955
rect 485 7925 515 7955
rect 14485 7925 14515 7955
rect 14645 7925 14675 7955
rect 14805 7925 14835 7955
rect 14965 7925 14995 7955
rect 5 7845 35 7875
rect 165 7845 195 7875
rect 14485 7845 14515 7875
rect 14645 7845 14675 7875
rect 14805 7845 14835 7875
rect 14965 7845 14995 7875
rect 5 7765 35 7795
rect 165 7765 195 7795
rect 325 7765 355 7795
rect 485 7765 515 7795
rect 14485 7765 14515 7795
rect 14645 7765 14675 7795
rect 14805 7765 14835 7795
rect 14965 7765 14995 7795
rect 5 7685 35 7715
rect 165 7685 195 7715
rect 325 7685 355 7715
rect 485 7685 515 7715
rect 14485 7685 14515 7715
rect 14645 7685 14675 7715
rect 14805 7685 14835 7715
rect 14965 7685 14995 7715
rect 5 7605 35 7635
rect 165 7605 195 7635
rect 325 7605 355 7635
rect 485 7605 515 7635
rect 14485 7605 14515 7635
rect 14645 7605 14675 7635
rect 14805 7605 14835 7635
rect 14965 7605 14995 7635
rect 5 7525 35 7555
rect 165 7525 195 7555
rect 325 7525 355 7555
rect 485 7525 515 7555
rect 14485 7525 14515 7555
rect 14645 7525 14675 7555
rect 14805 7525 14835 7555
rect 14965 7525 14995 7555
rect 5 7445 35 7475
rect 165 7445 195 7475
rect 325 7445 355 7475
rect 485 7445 515 7475
rect 14485 7445 14515 7475
rect 14645 7445 14675 7475
rect 14805 7445 14835 7475
rect 14965 7445 14995 7475
rect 5 7365 35 7395
rect 165 7365 195 7395
rect 325 7365 355 7395
rect 485 7365 515 7395
rect 14485 7365 14515 7395
rect 14645 7365 14675 7395
rect 14805 7365 14835 7395
rect 14965 7365 14995 7395
rect 5 7285 35 7315
rect 165 7285 195 7315
rect 325 7285 355 7315
rect 485 7285 515 7315
rect 14485 7285 14515 7315
rect 14645 7285 14675 7315
rect 14805 7285 14835 7315
rect 14965 7285 14995 7315
rect 5 7205 35 7235
rect 165 7205 195 7235
rect 325 7205 355 7235
rect 485 7205 515 7235
rect 14485 7205 14515 7235
rect 14645 7205 14675 7235
rect 14805 7205 14835 7235
rect 14965 7205 14995 7235
rect 5 7125 35 7155
rect 165 7125 195 7155
rect 325 7125 355 7155
rect 485 7125 515 7155
rect 14485 7125 14515 7155
rect 14645 7125 14675 7155
rect 14805 7125 14835 7155
rect 14965 7125 14995 7155
rect 5 7045 35 7075
rect 165 7045 195 7075
rect 325 7045 355 7075
rect 485 7045 515 7075
rect 14485 7045 14515 7075
rect 14645 7045 14675 7075
rect 14805 7045 14835 7075
rect 14965 7045 14995 7075
rect 5 6965 35 6995
rect 165 6965 195 6995
rect 325 6965 355 6995
rect 485 6965 515 6995
rect 14485 6965 14515 6995
rect 14645 6965 14675 6995
rect 14805 6965 14835 6995
rect 14965 6965 14995 6995
rect 5 6885 35 6915
rect 165 6885 195 6915
rect 325 6885 355 6915
rect 485 6885 515 6915
rect 14485 6885 14515 6915
rect 14645 6885 14675 6915
rect 14805 6885 14835 6915
rect 14965 6885 14995 6915
rect 5 6805 35 6835
rect 165 6805 195 6835
rect 325 6805 355 6835
rect 485 6805 515 6835
rect 14485 6805 14515 6835
rect 14645 6805 14675 6835
rect 14805 6805 14835 6835
rect 14965 6805 14995 6835
rect 5 6725 35 6755
rect 165 6725 195 6755
rect 325 6725 355 6755
rect 485 6725 515 6755
rect 14485 6725 14515 6755
rect 14645 6725 14675 6755
rect 14805 6725 14835 6755
rect 14965 6725 14995 6755
rect 5 6645 35 6675
rect 165 6645 195 6675
rect 325 6645 355 6675
rect 485 6645 515 6675
rect 14485 6645 14515 6675
rect 14645 6645 14675 6675
rect 14805 6645 14835 6675
rect 14965 6645 14995 6675
rect 5 6565 35 6595
rect 165 6565 195 6595
rect 325 6565 355 6595
rect 14485 6565 14515 6595
rect 14645 6565 14675 6595
rect 14805 6565 14835 6595
rect 14965 6565 14995 6595
rect 5 6485 35 6515
rect 165 6485 195 6515
rect 325 6485 355 6515
rect 485 6485 515 6515
rect 14485 6485 14515 6515
rect 14645 6485 14675 6515
rect 14805 6485 14835 6515
rect 14965 6485 14995 6515
rect 5 6405 35 6435
rect 165 6405 195 6435
rect 325 6405 355 6435
rect 485 6405 515 6435
rect 14485 6405 14515 6435
rect 14645 6405 14675 6435
rect 14805 6405 14835 6435
rect 14965 6405 14995 6435
rect 5 6325 35 6355
rect 165 6325 195 6355
rect 325 6325 355 6355
rect 485 6325 515 6355
rect 14485 6325 14515 6355
rect 14645 6325 14675 6355
rect 14805 6325 14835 6355
rect 14965 6325 14995 6355
rect 5 6245 35 6275
rect 165 6245 195 6275
rect 325 6245 355 6275
rect 485 6245 515 6275
rect 14485 6245 14515 6275
rect 14645 6245 14675 6275
rect 14805 6245 14835 6275
rect 14965 6245 14995 6275
rect 5 6165 35 6195
rect 165 6165 195 6195
rect 325 6165 355 6195
rect 485 6165 515 6195
rect 14485 6165 14515 6195
rect 14645 6165 14675 6195
rect 14805 6165 14835 6195
rect 14965 6165 14995 6195
rect 5 6085 35 6115
rect 165 6085 195 6115
rect 325 6085 355 6115
rect 485 6085 515 6115
rect 14485 6085 14515 6115
rect 14645 6085 14675 6115
rect 14805 6085 14835 6115
rect 14965 6085 14995 6115
rect 5 6005 35 6035
rect 165 6005 195 6035
rect 325 6005 355 6035
rect 485 6005 515 6035
rect 14485 6005 14515 6035
rect 14645 6005 14675 6035
rect 14805 6005 14835 6035
rect 14965 6005 14995 6035
rect 5 5925 35 5955
rect 165 5925 195 5955
rect 325 5925 355 5955
rect 485 5925 515 5955
rect 14485 5925 14515 5955
rect 14645 5925 14675 5955
rect 14805 5925 14835 5955
rect 14965 5925 14995 5955
rect 5 5845 35 5875
rect 165 5845 195 5875
rect 325 5845 355 5875
rect 485 5845 515 5875
rect 14485 5845 14515 5875
rect 14645 5845 14675 5875
rect 14805 5845 14835 5875
rect 14965 5845 14995 5875
rect 5 5765 35 5795
rect 165 5765 195 5795
rect 325 5765 355 5795
rect 485 5765 515 5795
rect 14485 5765 14515 5795
rect 14645 5765 14675 5795
rect 14805 5765 14835 5795
rect 14965 5765 14995 5795
rect 5 5685 35 5715
rect 165 5685 195 5715
rect 325 5685 355 5715
rect 485 5685 515 5715
rect 14485 5685 14515 5715
rect 14645 5685 14675 5715
rect 14805 5685 14835 5715
rect 14965 5685 14995 5715
rect 5 5605 35 5635
rect 165 5605 195 5635
rect 325 5605 355 5635
rect 485 5605 515 5635
rect 14485 5605 14515 5635
rect 14645 5605 14675 5635
rect 14805 5605 14835 5635
rect 14965 5605 14995 5635
rect 5 5525 35 5555
rect 165 5525 195 5555
rect 325 5525 355 5555
rect 485 5525 515 5555
rect 14485 5525 14515 5555
rect 14645 5525 14675 5555
rect 14805 5525 14835 5555
rect 14965 5525 14995 5555
rect 5 5445 35 5475
rect 165 5445 195 5475
rect 325 5445 355 5475
rect 485 5445 515 5475
rect 14485 5445 14515 5475
rect 14645 5445 14675 5475
rect 14805 5445 14835 5475
rect 14965 5445 14995 5475
rect 5 5365 35 5395
rect 165 5365 195 5395
rect 325 5365 355 5395
rect 485 5365 515 5395
rect 14485 5365 14515 5395
rect 14645 5365 14675 5395
rect 14805 5365 14835 5395
rect 14965 5365 14995 5395
rect 5 5285 35 5315
rect 165 5285 195 5315
rect 14485 5285 14515 5315
rect 14645 5285 14675 5315
rect 14805 5285 14835 5315
rect 14965 5285 14995 5315
rect 5 5205 35 5235
rect 165 5205 195 5235
rect 325 5205 355 5235
rect 485 5205 515 5235
rect 14485 5205 14515 5235
rect 14645 5205 14675 5235
rect 14805 5205 14835 5235
rect 14965 5205 14995 5235
rect 14485 5125 14515 5155
rect 14645 5125 14675 5155
rect 14805 5125 14835 5155
rect 14965 5125 14995 5155
rect 5 5045 35 5075
rect 165 5045 195 5075
rect 325 5045 355 5075
rect 485 5045 515 5075
rect 14485 5045 14515 5075
rect 14645 5045 14675 5075
rect 14805 5045 14835 5075
rect 14965 5045 14995 5075
rect 5 4965 35 4995
rect 165 4965 195 4995
rect 325 4965 355 4995
rect 485 4965 515 4995
rect 14485 4965 14515 4995
rect 14645 4965 14675 4995
rect 14805 4965 14835 4995
rect 14965 4965 14995 4995
rect 5 4885 35 4915
rect 165 4885 195 4915
rect 325 4885 355 4915
rect 485 4885 515 4915
rect 14485 4885 14515 4915
rect 14645 4885 14675 4915
rect 14805 4885 14835 4915
rect 14965 4885 14995 4915
rect 5 4805 35 4835
rect 165 4805 195 4835
rect 325 4805 355 4835
rect 485 4805 515 4835
rect 14485 4805 14515 4835
rect 14645 4805 14675 4835
rect 14805 4805 14835 4835
rect 14965 4805 14995 4835
rect 5 4725 35 4755
rect 165 4725 195 4755
rect 325 4725 355 4755
rect 485 4725 515 4755
rect 5 4645 35 4675
rect 165 4645 195 4675
rect 325 4645 355 4675
rect 485 4645 515 4675
rect 14485 4645 14515 4675
rect 14645 4645 14675 4675
rect 14805 4645 14835 4675
rect 14965 4645 14995 4675
rect 5 4565 35 4595
rect 165 4565 195 4595
rect 325 4565 355 4595
rect 485 4565 515 4595
rect 14805 4565 14835 4595
rect 14965 4565 14995 4595
rect 5 4485 35 4515
rect 165 4485 195 4515
rect 325 4485 355 4515
rect 485 4485 515 4515
rect 14485 4485 14515 4515
rect 14645 4485 14675 4515
rect 14805 4485 14835 4515
rect 14965 4485 14995 4515
rect 5 4405 35 4435
rect 165 4405 195 4435
rect 325 4405 355 4435
rect 485 4405 515 4435
rect 14485 4405 14515 4435
rect 14645 4405 14675 4435
rect 14805 4405 14835 4435
rect 14965 4405 14995 4435
rect 5 4325 35 4355
rect 165 4325 195 4355
rect 325 4325 355 4355
rect 485 4325 515 4355
rect 14485 4325 14515 4355
rect 14645 4325 14675 4355
rect 14805 4325 14835 4355
rect 14965 4325 14995 4355
rect 5 4245 35 4275
rect 165 4245 195 4275
rect 325 4245 355 4275
rect 485 4245 515 4275
rect 14485 4245 14515 4275
rect 14645 4245 14675 4275
rect 14805 4245 14835 4275
rect 14965 4245 14995 4275
rect 5 4165 35 4195
rect 165 4165 195 4195
rect 325 4165 355 4195
rect 485 4165 515 4195
rect 14485 4165 14515 4195
rect 14645 4165 14675 4195
rect 14805 4165 14835 4195
rect 14965 4165 14995 4195
rect 5 4085 35 4115
rect 165 4085 195 4115
rect 325 4085 355 4115
rect 485 4085 515 4115
rect 14485 4085 14515 4115
rect 14645 4085 14675 4115
rect 14805 4085 14835 4115
rect 14965 4085 14995 4115
rect 5 4005 35 4035
rect 165 4005 195 4035
rect 325 4005 355 4035
rect 485 4005 515 4035
rect 14485 4005 14515 4035
rect 14645 4005 14675 4035
rect 14805 4005 14835 4035
rect 14965 4005 14995 4035
rect 5 3925 35 3955
rect 165 3925 195 3955
rect 325 3925 355 3955
rect 485 3925 515 3955
rect 14485 3925 14515 3955
rect 14645 3925 14675 3955
rect 14805 3925 14835 3955
rect 14965 3925 14995 3955
rect 5 3845 35 3875
rect 165 3845 195 3875
rect 325 3845 355 3875
rect 485 3845 515 3875
rect 14485 3845 14515 3875
rect 14645 3845 14675 3875
rect 14805 3845 14835 3875
rect 14965 3845 14995 3875
rect 5 3765 35 3795
rect 165 3765 195 3795
rect 325 3765 355 3795
rect 485 3765 515 3795
rect 14485 3765 14515 3795
rect 14645 3765 14675 3795
rect 14805 3765 14835 3795
rect 14965 3765 14995 3795
rect 5 3685 35 3715
rect 165 3685 195 3715
rect 325 3685 355 3715
rect 485 3685 515 3715
rect 14485 3685 14515 3715
rect 14645 3685 14675 3715
rect 14805 3685 14835 3715
rect 14965 3685 14995 3715
rect 5 3605 35 3635
rect 165 3605 195 3635
rect 325 3605 355 3635
rect 485 3605 515 3635
rect 14485 3605 14515 3635
rect 14645 3605 14675 3635
rect 14805 3605 14835 3635
rect 14965 3605 14995 3635
rect 5 3525 35 3555
rect 165 3525 195 3555
rect 325 3525 355 3555
rect 485 3525 515 3555
rect 14485 3525 14515 3555
rect 14645 3525 14675 3555
rect 14805 3525 14835 3555
rect 14965 3525 14995 3555
rect 5 3445 35 3475
rect 165 3445 195 3475
rect 325 3445 355 3475
rect 485 3445 515 3475
rect 14485 3445 14515 3475
rect 14645 3445 14675 3475
rect 14805 3445 14835 3475
rect 14965 3445 14995 3475
rect 5 3365 35 3395
rect 165 3365 195 3395
rect 325 3365 355 3395
rect 485 3365 515 3395
rect 14485 3365 14515 3395
rect 14645 3365 14675 3395
rect 14805 3365 14835 3395
rect 14965 3365 14995 3395
rect 5 3285 35 3315
rect 165 3285 195 3315
rect 325 3285 355 3315
rect 485 3285 515 3315
rect 14645 3285 14675 3315
rect 14805 3285 14835 3315
rect 14965 3285 14995 3315
rect 5 3205 35 3235
rect 165 3205 195 3235
rect 325 3205 355 3235
rect 485 3205 515 3235
rect 14485 3205 14515 3235
rect 14645 3205 14675 3235
rect 14805 3205 14835 3235
rect 14965 3205 14995 3235
rect 5 3125 35 3155
rect 165 3125 195 3155
rect 325 3125 355 3155
rect 485 3125 515 3155
rect 14485 3125 14515 3155
rect 14645 3125 14675 3155
rect 14805 3125 14835 3155
rect 14965 3125 14995 3155
rect 5 3045 35 3075
rect 165 3045 195 3075
rect 325 3045 355 3075
rect 485 3045 515 3075
rect 14485 3045 14515 3075
rect 14645 3045 14675 3075
rect 14805 3045 14835 3075
rect 14965 3045 14995 3075
rect 5 2965 35 2995
rect 165 2965 195 2995
rect 325 2965 355 2995
rect 485 2965 515 2995
rect 14485 2965 14515 2995
rect 14645 2965 14675 2995
rect 14805 2965 14835 2995
rect 14965 2965 14995 2995
rect 5 2885 35 2915
rect 165 2885 195 2915
rect 325 2885 355 2915
rect 485 2885 515 2915
rect 14485 2885 14515 2915
rect 14645 2885 14675 2915
rect 14805 2885 14835 2915
rect 14965 2885 14995 2915
rect 5 2805 35 2835
rect 165 2805 195 2835
rect 325 2805 355 2835
rect 485 2805 515 2835
rect 14485 2805 14515 2835
rect 14645 2805 14675 2835
rect 14805 2805 14835 2835
rect 14965 2805 14995 2835
rect 5 2725 35 2755
rect 165 2725 195 2755
rect 325 2725 355 2755
rect 485 2725 515 2755
rect 14485 2725 14515 2755
rect 14645 2725 14675 2755
rect 14805 2725 14835 2755
rect 14965 2725 14995 2755
rect 5 2645 35 2675
rect 165 2645 195 2675
rect 325 2645 355 2675
rect 485 2645 515 2675
rect 14485 2645 14515 2675
rect 14645 2645 14675 2675
rect 14805 2645 14835 2675
rect 14965 2645 14995 2675
rect 5 2565 35 2595
rect 165 2565 195 2595
rect 325 2565 355 2595
rect 485 2565 515 2595
rect 14485 2565 14515 2595
rect 14645 2565 14675 2595
rect 14805 2565 14835 2595
rect 14965 2565 14995 2595
rect 5 2485 35 2515
rect 165 2485 195 2515
rect 325 2485 355 2515
rect 485 2485 515 2515
rect 14485 2485 14515 2515
rect 14645 2485 14675 2515
rect 14805 2485 14835 2515
rect 14965 2485 14995 2515
rect 5 2405 35 2435
rect 165 2405 195 2435
rect 325 2405 355 2435
rect 485 2405 515 2435
rect 14485 2405 14515 2435
rect 14645 2405 14675 2435
rect 14805 2405 14835 2435
rect 14965 2405 14995 2435
rect 5 2325 35 2355
rect 165 2325 195 2355
rect 325 2325 355 2355
rect 485 2325 515 2355
rect 14485 2325 14515 2355
rect 14645 2325 14675 2355
rect 14805 2325 14835 2355
rect 14965 2325 14995 2355
rect 5 2245 35 2275
rect 165 2245 195 2275
rect 325 2245 355 2275
rect 485 2245 515 2275
rect 14485 2245 14515 2275
rect 14645 2245 14675 2275
rect 14805 2245 14835 2275
rect 14965 2245 14995 2275
rect 5 2165 35 2195
rect 165 2165 195 2195
rect 325 2165 355 2195
rect 485 2165 515 2195
rect 14485 2165 14515 2195
rect 14645 2165 14675 2195
rect 14805 2165 14835 2195
rect 14965 2165 14995 2195
rect 5 2085 35 2115
rect 165 2085 195 2115
rect 325 2085 355 2115
rect 485 2085 515 2115
rect 14485 2085 14515 2115
rect 14645 2085 14675 2115
rect 14805 2085 14835 2115
rect 14965 2085 14995 2115
rect 5 2005 35 2035
rect 165 2005 195 2035
rect 325 2005 355 2035
rect 485 2005 515 2035
rect 14805 2005 14835 2035
rect 14965 2005 14995 2035
rect 5 1925 35 1955
rect 165 1925 195 1955
rect 325 1925 355 1955
rect 485 1925 515 1955
rect 14485 1925 14515 1955
rect 14645 1925 14675 1955
rect 14805 1925 14835 1955
rect 14965 1925 14995 1955
rect 5 1845 35 1875
rect 165 1845 195 1875
rect 325 1845 355 1875
rect 485 1845 515 1875
rect 5 1765 35 1795
rect 165 1765 195 1795
rect 325 1765 355 1795
rect 485 1765 515 1795
rect 14485 1765 14515 1795
rect 14645 1765 14675 1795
rect 14805 1765 14835 1795
rect 14965 1765 14995 1795
rect 5 1685 35 1715
rect 165 1685 195 1715
rect 325 1685 355 1715
rect 485 1685 515 1715
rect 14485 1685 14515 1715
rect 14645 1685 14675 1715
rect 14805 1685 14835 1715
rect 14965 1685 14995 1715
rect 5 1605 35 1635
rect 165 1605 195 1635
rect 325 1605 355 1635
rect 485 1605 515 1635
rect 14485 1605 14515 1635
rect 14645 1605 14675 1635
rect 14805 1605 14835 1635
rect 14965 1605 14995 1635
rect 5 1525 35 1555
rect 165 1525 195 1555
rect 325 1525 355 1555
rect 485 1525 515 1555
rect 14485 1525 14515 1555
rect 14645 1525 14675 1555
rect 14805 1525 14835 1555
rect 14965 1525 14995 1555
rect 5 1445 35 1475
rect 165 1445 195 1475
rect 325 1445 355 1475
rect 485 1445 515 1475
rect 14485 1445 14515 1475
rect 14645 1445 14675 1475
rect 14805 1445 14835 1475
rect 14965 1445 14995 1475
rect 5 1365 35 1395
rect 165 1365 195 1395
rect 325 1365 355 1395
rect 485 1365 515 1395
rect 14485 1365 14515 1395
rect 14645 1365 14675 1395
rect 14805 1365 14835 1395
rect 14965 1365 14995 1395
rect 5 1285 35 1315
rect 165 1285 195 1315
rect 325 1285 355 1315
rect 485 1285 515 1315
rect 14485 1285 14515 1315
rect 14645 1285 14675 1315
rect 14805 1285 14835 1315
rect 14965 1285 14995 1315
rect 5 1205 35 1235
rect 165 1205 195 1235
rect 325 1205 355 1235
rect 485 1205 515 1235
rect 14485 1205 14515 1235
rect 14645 1205 14675 1235
rect 14805 1205 14835 1235
rect 14965 1205 14995 1235
rect 5 1125 35 1155
rect 165 1125 195 1155
rect 325 1125 355 1155
rect 485 1125 515 1155
rect 14485 1125 14515 1155
rect 14645 1125 14675 1155
rect 14805 1125 14835 1155
rect 14965 1125 14995 1155
rect 5 1045 35 1075
rect 165 1045 195 1075
rect 325 1045 355 1075
rect 485 1045 515 1075
rect 14485 1045 14515 1075
rect 14645 1045 14675 1075
rect 14805 1045 14835 1075
rect 14965 1045 14995 1075
rect 5 965 35 995
rect 165 965 195 995
rect 325 965 355 995
rect 485 965 515 995
rect 14485 965 14515 995
rect 14645 965 14675 995
rect 14805 965 14835 995
rect 14965 965 14995 995
rect 5 885 35 915
rect 165 885 195 915
rect 325 885 355 915
rect 485 885 515 915
rect 14485 885 14515 915
rect 14645 885 14675 915
rect 14805 885 14835 915
rect 14965 885 14995 915
rect 5 805 35 835
rect 165 805 195 835
rect 325 805 355 835
rect 485 805 515 835
rect 14485 805 14515 835
rect 14645 805 14675 835
rect 14805 805 14835 835
rect 14965 805 14995 835
rect 5 725 35 755
rect 165 725 195 755
rect 325 725 355 755
rect 485 725 515 755
rect 14485 725 14515 755
rect 14645 725 14675 755
rect 14805 725 14835 755
rect 14965 725 14995 755
rect 5 645 35 675
rect 165 645 195 675
rect 325 645 355 675
rect 485 645 515 675
rect 14485 645 14515 675
rect 14645 645 14675 675
rect 14805 645 14835 675
rect 14965 645 14995 675
rect 5 565 35 595
rect 165 565 195 595
rect 325 565 355 595
rect 485 565 515 595
rect 14485 565 14515 595
rect 14645 565 14675 595
rect 14805 565 14835 595
rect 14965 565 14995 595
rect 5 485 35 515
rect 165 485 195 515
rect 325 485 355 515
rect 485 485 515 515
rect 565 485 595 515
rect 14405 485 14435 515
rect 14485 485 14515 515
rect 14645 485 14675 515
rect 14805 485 14835 515
rect 14965 485 14995 515
<< metal3 >>
rect 0 15956 40 15960
rect 0 15924 4 15956
rect 36 15924 40 15956
rect 0 15876 40 15924
rect 0 15844 4 15876
rect 36 15844 40 15876
rect 0 15796 40 15844
rect 0 15764 4 15796
rect 36 15764 40 15796
rect 0 15716 40 15764
rect 0 15684 4 15716
rect 36 15684 40 15716
rect 0 15636 40 15684
rect 0 15604 4 15636
rect 36 15604 40 15636
rect 0 15556 40 15604
rect 0 15524 4 15556
rect 36 15524 40 15556
rect 0 15476 40 15524
rect 0 15444 4 15476
rect 36 15444 40 15476
rect 0 15396 40 15444
rect 0 15364 4 15396
rect 36 15364 40 15396
rect 0 15316 40 15364
rect 0 15284 4 15316
rect 36 15284 40 15316
rect 0 15236 40 15284
rect 0 15204 4 15236
rect 36 15204 40 15236
rect 0 15156 40 15204
rect 0 15124 4 15156
rect 36 15124 40 15156
rect 0 15076 40 15124
rect 0 15044 4 15076
rect 36 15044 40 15076
rect 0 14996 40 15044
rect 0 14964 4 14996
rect 36 14964 40 14996
rect 0 14916 40 14964
rect 0 14884 4 14916
rect 36 14884 40 14916
rect 0 14836 40 14884
rect 0 14804 4 14836
rect 36 14804 40 14836
rect 0 14756 40 14804
rect 0 14724 4 14756
rect 36 14724 40 14756
rect 0 14676 40 14724
rect 0 14644 4 14676
rect 36 14644 40 14676
rect 0 14596 40 14644
rect 0 14564 4 14596
rect 36 14564 40 14596
rect 0 14516 40 14564
rect 0 14484 4 14516
rect 36 14484 40 14516
rect 0 14436 40 14484
rect 0 14404 4 14436
rect 36 14404 40 14436
rect 0 14356 40 14404
rect 0 14324 4 14356
rect 36 14324 40 14356
rect 0 14276 40 14324
rect 0 14244 4 14276
rect 36 14244 40 14276
rect 0 14196 40 14244
rect 0 14164 4 14196
rect 36 14164 40 14196
rect 0 14116 40 14164
rect 0 14084 4 14116
rect 36 14084 40 14116
rect 0 14036 40 14084
rect 0 14004 4 14036
rect 36 14004 40 14036
rect 0 13956 40 14004
rect 0 13924 4 13956
rect 36 13924 40 13956
rect 0 13876 40 13924
rect 0 13844 4 13876
rect 36 13844 40 13876
rect 0 13796 40 13844
rect 0 13764 4 13796
rect 36 13764 40 13796
rect 0 13716 40 13764
rect 0 13684 4 13716
rect 36 13684 40 13716
rect 0 13636 40 13684
rect 0 13604 4 13636
rect 36 13604 40 13636
rect 0 13556 40 13604
rect 0 13524 4 13556
rect 36 13524 40 13556
rect 0 13476 40 13524
rect 0 13444 4 13476
rect 36 13444 40 13476
rect 0 13396 40 13444
rect 0 13364 4 13396
rect 36 13364 40 13396
rect 0 13316 40 13364
rect 0 13284 4 13316
rect 36 13284 40 13316
rect 0 13236 40 13284
rect 0 13204 4 13236
rect 36 13204 40 13236
rect 0 13156 40 13204
rect 0 13124 4 13156
rect 36 13124 40 13156
rect 0 13076 40 13124
rect 0 13044 4 13076
rect 36 13044 40 13076
rect 0 12996 40 13044
rect 0 12964 4 12996
rect 36 12964 40 12996
rect 0 12916 40 12964
rect 0 12884 4 12916
rect 36 12884 40 12916
rect 0 12836 40 12884
rect 0 12804 4 12836
rect 36 12804 40 12836
rect 0 12756 40 12804
rect 0 12724 4 12756
rect 36 12724 40 12756
rect 0 12676 40 12724
rect 0 12644 4 12676
rect 36 12644 40 12676
rect 0 12596 40 12644
rect 0 12564 4 12596
rect 36 12564 40 12596
rect 0 12516 40 12564
rect 0 12484 4 12516
rect 36 12484 40 12516
rect 0 12436 40 12484
rect 0 12404 4 12436
rect 36 12404 40 12436
rect 0 12356 40 12404
rect 0 12324 4 12356
rect 36 12324 40 12356
rect 0 12276 40 12324
rect 0 12244 4 12276
rect 36 12244 40 12276
rect 0 12196 40 12244
rect 0 12164 4 12196
rect 36 12164 40 12196
rect 0 12116 40 12164
rect 0 12084 4 12116
rect 36 12084 40 12116
rect 0 12036 40 12084
rect 0 12004 4 12036
rect 36 12004 40 12036
rect 0 11956 40 12004
rect 0 11924 4 11956
rect 36 11924 40 11956
rect 0 11876 40 11924
rect 0 11844 4 11876
rect 36 11844 40 11876
rect 0 11796 40 11844
rect 0 11764 4 11796
rect 36 11764 40 11796
rect 0 11716 40 11764
rect 0 11684 4 11716
rect 36 11684 40 11716
rect 0 11636 40 11684
rect 0 11604 4 11636
rect 36 11604 40 11636
rect 0 11556 40 11604
rect 0 11524 4 11556
rect 36 11524 40 11556
rect 0 11476 40 11524
rect 0 11444 4 11476
rect 36 11444 40 11476
rect 0 11396 40 11444
rect 0 11364 4 11396
rect 36 11364 40 11396
rect 0 11236 40 11364
rect 0 11204 4 11236
rect 36 11204 40 11236
rect 0 11156 40 11204
rect 0 11124 4 11156
rect 36 11124 40 11156
rect 0 11076 40 11124
rect 0 11044 4 11076
rect 36 11044 40 11076
rect 0 10996 40 11044
rect 0 10964 4 10996
rect 36 10964 40 10996
rect 0 10916 40 10964
rect 0 10884 4 10916
rect 36 10884 40 10916
rect 0 10836 40 10884
rect 0 10804 4 10836
rect 36 10804 40 10836
rect 0 10756 40 10804
rect 0 10724 4 10756
rect 36 10724 40 10756
rect 0 10676 40 10724
rect 0 10644 4 10676
rect 36 10644 40 10676
rect 0 10596 40 10644
rect 0 10564 4 10596
rect 36 10564 40 10596
rect 0 10516 40 10564
rect 0 10484 4 10516
rect 36 10484 40 10516
rect 0 10436 40 10484
rect 0 10404 4 10436
rect 36 10404 40 10436
rect 0 10356 40 10404
rect 0 10324 4 10356
rect 36 10324 40 10356
rect 0 10276 40 10324
rect 0 10244 4 10276
rect 36 10244 40 10276
rect 0 10196 40 10244
rect 0 10164 4 10196
rect 36 10164 40 10196
rect 0 10116 40 10164
rect 0 10084 4 10116
rect 36 10084 40 10116
rect 0 10036 40 10084
rect 0 10004 4 10036
rect 36 10004 40 10036
rect 0 9956 40 10004
rect 0 9924 4 9956
rect 36 9924 40 9956
rect 0 9876 40 9924
rect 0 9844 4 9876
rect 36 9844 40 9876
rect 0 9796 40 9844
rect 0 9764 4 9796
rect 36 9764 40 9796
rect 0 9716 40 9764
rect 0 9684 4 9716
rect 36 9684 40 9716
rect 0 9636 40 9684
rect 0 9604 4 9636
rect 36 9604 40 9636
rect 0 9556 40 9604
rect 0 9524 4 9556
rect 36 9524 40 9556
rect 0 9476 40 9524
rect 0 9444 4 9476
rect 36 9444 40 9476
rect 0 9396 40 9444
rect 0 9364 4 9396
rect 36 9364 40 9396
rect 0 9316 40 9364
rect 0 9284 4 9316
rect 36 9284 40 9316
rect 0 9236 40 9284
rect 0 9204 4 9236
rect 36 9204 40 9236
rect 0 9156 40 9204
rect 0 9124 4 9156
rect 36 9124 40 9156
rect 0 9076 40 9124
rect 0 9044 4 9076
rect 36 9044 40 9076
rect 0 8996 40 9044
rect 0 8964 4 8996
rect 36 8964 40 8996
rect 0 8916 40 8964
rect 0 8884 4 8916
rect 36 8884 40 8916
rect 0 8836 40 8884
rect 0 8804 4 8836
rect 36 8804 40 8836
rect 0 8756 40 8804
rect 0 8724 4 8756
rect 36 8724 40 8756
rect 0 8676 40 8724
rect 0 8644 4 8676
rect 36 8644 40 8676
rect 0 8596 40 8644
rect 0 8564 4 8596
rect 36 8564 40 8596
rect 0 8516 40 8564
rect 0 8484 4 8516
rect 36 8484 40 8516
rect 0 8356 40 8484
rect 0 8324 4 8356
rect 36 8324 40 8356
rect 0 8276 40 8324
rect 0 8244 4 8276
rect 36 8244 40 8276
rect 0 8196 40 8244
rect 0 8164 4 8196
rect 36 8164 40 8196
rect 0 8116 40 8164
rect 0 8084 4 8116
rect 36 8084 40 8116
rect 0 7956 40 8084
rect 0 7924 4 7956
rect 36 7924 40 7956
rect 0 7876 40 7924
rect 0 7844 4 7876
rect 36 7844 40 7876
rect 0 7796 40 7844
rect 0 7764 4 7796
rect 36 7764 40 7796
rect 0 7716 40 7764
rect 0 7684 4 7716
rect 36 7684 40 7716
rect 0 7636 40 7684
rect 0 7604 4 7636
rect 36 7604 40 7636
rect 0 7556 40 7604
rect 0 7524 4 7556
rect 36 7524 40 7556
rect 0 7476 40 7524
rect 0 7444 4 7476
rect 36 7444 40 7476
rect 0 7396 40 7444
rect 0 7364 4 7396
rect 36 7364 40 7396
rect 0 7316 40 7364
rect 0 7284 4 7316
rect 36 7284 40 7316
rect 0 7236 40 7284
rect 0 7204 4 7236
rect 36 7204 40 7236
rect 0 7156 40 7204
rect 0 7124 4 7156
rect 36 7124 40 7156
rect 0 7076 40 7124
rect 0 7044 4 7076
rect 36 7044 40 7076
rect 0 6996 40 7044
rect 0 6964 4 6996
rect 36 6964 40 6996
rect 0 6916 40 6964
rect 0 6884 4 6916
rect 36 6884 40 6916
rect 0 6836 40 6884
rect 0 6804 4 6836
rect 36 6804 40 6836
rect 0 6756 40 6804
rect 0 6724 4 6756
rect 36 6724 40 6756
rect 0 6676 40 6724
rect 0 6644 4 6676
rect 36 6644 40 6676
rect 0 6596 40 6644
rect 0 6564 4 6596
rect 36 6564 40 6596
rect 0 6516 40 6564
rect 0 6484 4 6516
rect 36 6484 40 6516
rect 0 6436 40 6484
rect 0 6404 4 6436
rect 36 6404 40 6436
rect 0 6356 40 6404
rect 0 6324 4 6356
rect 36 6324 40 6356
rect 0 6276 40 6324
rect 0 6244 4 6276
rect 36 6244 40 6276
rect 0 6196 40 6244
rect 0 6164 4 6196
rect 36 6164 40 6196
rect 0 6116 40 6164
rect 0 6084 4 6116
rect 36 6084 40 6116
rect 0 6036 40 6084
rect 0 6004 4 6036
rect 36 6004 40 6036
rect 0 5956 40 6004
rect 0 5924 4 5956
rect 36 5924 40 5956
rect 0 5876 40 5924
rect 0 5844 4 5876
rect 36 5844 40 5876
rect 0 5796 40 5844
rect 0 5764 4 5796
rect 36 5764 40 5796
rect 0 5716 40 5764
rect 0 5684 4 5716
rect 36 5684 40 5716
rect 0 5636 40 5684
rect 0 5604 4 5636
rect 36 5604 40 5636
rect 0 5556 40 5604
rect 0 5524 4 5556
rect 36 5524 40 5556
rect 0 5476 40 5524
rect 0 5444 4 5476
rect 36 5444 40 5476
rect 0 5396 40 5444
rect 0 5364 4 5396
rect 36 5364 40 5396
rect 0 5316 40 5364
rect 0 5284 4 5316
rect 36 5284 40 5316
rect 0 5236 40 5284
rect 0 5204 4 5236
rect 36 5204 40 5236
rect 0 5076 40 5204
rect 0 5044 4 5076
rect 36 5044 40 5076
rect 0 4996 40 5044
rect 0 4964 4 4996
rect 36 4964 40 4996
rect 0 4916 40 4964
rect 0 4884 4 4916
rect 36 4884 40 4916
rect 0 4836 40 4884
rect 0 4804 4 4836
rect 36 4804 40 4836
rect 0 4756 40 4804
rect 0 4724 4 4756
rect 36 4724 40 4756
rect 0 4676 40 4724
rect 0 4644 4 4676
rect 36 4644 40 4676
rect 0 4596 40 4644
rect 0 4564 4 4596
rect 36 4564 40 4596
rect 0 4516 40 4564
rect 0 4484 4 4516
rect 36 4484 40 4516
rect 0 4436 40 4484
rect 0 4404 4 4436
rect 36 4404 40 4436
rect 0 4356 40 4404
rect 0 4324 4 4356
rect 36 4324 40 4356
rect 0 4276 40 4324
rect 0 4244 4 4276
rect 36 4244 40 4276
rect 0 4196 40 4244
rect 0 4164 4 4196
rect 36 4164 40 4196
rect 0 4116 40 4164
rect 0 4084 4 4116
rect 36 4084 40 4116
rect 0 4036 40 4084
rect 0 4004 4 4036
rect 36 4004 40 4036
rect 0 3956 40 4004
rect 0 3924 4 3956
rect 36 3924 40 3956
rect 0 3876 40 3924
rect 0 3844 4 3876
rect 36 3844 40 3876
rect 0 3796 40 3844
rect 0 3764 4 3796
rect 36 3764 40 3796
rect 0 3716 40 3764
rect 0 3684 4 3716
rect 36 3684 40 3716
rect 0 3636 40 3684
rect 0 3604 4 3636
rect 36 3604 40 3636
rect 0 3556 40 3604
rect 0 3524 4 3556
rect 36 3524 40 3556
rect 0 3476 40 3524
rect 0 3444 4 3476
rect 36 3444 40 3476
rect 0 3396 40 3444
rect 0 3364 4 3396
rect 36 3364 40 3396
rect 0 3316 40 3364
rect 0 3284 4 3316
rect 36 3284 40 3316
rect 0 3236 40 3284
rect 0 3204 4 3236
rect 36 3204 40 3236
rect 0 3156 40 3204
rect 0 3124 4 3156
rect 36 3124 40 3156
rect 0 3076 40 3124
rect 0 3044 4 3076
rect 36 3044 40 3076
rect 0 2996 40 3044
rect 0 2964 4 2996
rect 36 2964 40 2996
rect 0 2916 40 2964
rect 0 2884 4 2916
rect 36 2884 40 2916
rect 0 2836 40 2884
rect 0 2804 4 2836
rect 36 2804 40 2836
rect 0 2756 40 2804
rect 0 2724 4 2756
rect 36 2724 40 2756
rect 0 2676 40 2724
rect 0 2644 4 2676
rect 36 2644 40 2676
rect 0 2596 40 2644
rect 0 2564 4 2596
rect 36 2564 40 2596
rect 0 2516 40 2564
rect 0 2484 4 2516
rect 36 2484 40 2516
rect 0 2436 40 2484
rect 0 2404 4 2436
rect 36 2404 40 2436
rect 0 2356 40 2404
rect 0 2324 4 2356
rect 36 2324 40 2356
rect 0 2276 40 2324
rect 0 2244 4 2276
rect 36 2244 40 2276
rect 0 2196 40 2244
rect 0 2164 4 2196
rect 36 2164 40 2196
rect 0 2116 40 2164
rect 0 2084 4 2116
rect 36 2084 40 2116
rect 0 2036 40 2084
rect 0 2004 4 2036
rect 36 2004 40 2036
rect 0 1956 40 2004
rect 0 1924 4 1956
rect 36 1924 40 1956
rect 0 1876 40 1924
rect 0 1844 4 1876
rect 36 1844 40 1876
rect 0 1796 40 1844
rect 0 1764 4 1796
rect 36 1764 40 1796
rect 0 1716 40 1764
rect 0 1684 4 1716
rect 36 1684 40 1716
rect 0 1636 40 1684
rect 0 1604 4 1636
rect 36 1604 40 1636
rect 0 1556 40 1604
rect 0 1524 4 1556
rect 36 1524 40 1556
rect 0 1476 40 1524
rect 0 1444 4 1476
rect 36 1444 40 1476
rect 0 1396 40 1444
rect 0 1364 4 1396
rect 36 1364 40 1396
rect 0 1316 40 1364
rect 0 1284 4 1316
rect 36 1284 40 1316
rect 0 1236 40 1284
rect 0 1204 4 1236
rect 36 1204 40 1236
rect 0 1156 40 1204
rect 0 1124 4 1156
rect 36 1124 40 1156
rect 0 1076 40 1124
rect 0 1044 4 1076
rect 36 1044 40 1076
rect 0 996 40 1044
rect 0 964 4 996
rect 36 964 40 996
rect 0 916 40 964
rect 0 884 4 916
rect 36 884 40 916
rect 0 836 40 884
rect 0 804 4 836
rect 36 804 40 836
rect 0 756 40 804
rect 0 724 4 756
rect 36 724 40 756
rect 0 676 40 724
rect 0 644 4 676
rect 36 644 40 676
rect 0 596 40 644
rect 0 564 4 596
rect 36 564 40 596
rect 0 516 40 564
rect 0 484 4 516
rect 36 484 40 516
rect 0 436 40 484
rect 80 11316 120 15960
rect 80 11284 84 11316
rect 116 11284 120 11316
rect 80 8436 120 11284
rect 80 8404 84 8436
rect 116 8404 120 8436
rect 80 8036 120 8404
rect 80 8004 84 8036
rect 116 8004 120 8036
rect 80 5156 120 8004
rect 80 5124 84 5156
rect 116 5124 120 5156
rect 80 480 120 5124
rect 160 15956 200 15960
rect 160 15924 164 15956
rect 196 15924 200 15956
rect 160 15876 200 15924
rect 160 15844 164 15876
rect 196 15844 200 15876
rect 160 15796 200 15844
rect 160 15764 164 15796
rect 196 15764 200 15796
rect 160 15716 200 15764
rect 160 15684 164 15716
rect 196 15684 200 15716
rect 160 15636 200 15684
rect 160 15604 164 15636
rect 196 15604 200 15636
rect 160 15556 200 15604
rect 160 15524 164 15556
rect 196 15524 200 15556
rect 160 15476 200 15524
rect 160 15444 164 15476
rect 196 15444 200 15476
rect 160 15396 200 15444
rect 160 15364 164 15396
rect 196 15364 200 15396
rect 160 15316 200 15364
rect 160 15284 164 15316
rect 196 15284 200 15316
rect 160 15236 200 15284
rect 160 15204 164 15236
rect 196 15204 200 15236
rect 160 15156 200 15204
rect 160 15124 164 15156
rect 196 15124 200 15156
rect 160 15076 200 15124
rect 160 15044 164 15076
rect 196 15044 200 15076
rect 160 14996 200 15044
rect 160 14964 164 14996
rect 196 14964 200 14996
rect 160 14916 200 14964
rect 160 14884 164 14916
rect 196 14884 200 14916
rect 160 14836 200 14884
rect 160 14804 164 14836
rect 196 14804 200 14836
rect 160 14756 200 14804
rect 160 14724 164 14756
rect 196 14724 200 14756
rect 160 14676 200 14724
rect 160 14644 164 14676
rect 196 14644 200 14676
rect 160 14596 200 14644
rect 160 14564 164 14596
rect 196 14564 200 14596
rect 160 14516 200 14564
rect 160 14484 164 14516
rect 196 14484 200 14516
rect 160 14436 200 14484
rect 160 14404 164 14436
rect 196 14404 200 14436
rect 160 14356 200 14404
rect 160 14324 164 14356
rect 196 14324 200 14356
rect 160 14276 200 14324
rect 160 14244 164 14276
rect 196 14244 200 14276
rect 160 14196 200 14244
rect 160 14164 164 14196
rect 196 14164 200 14196
rect 160 14116 200 14164
rect 160 14084 164 14116
rect 196 14084 200 14116
rect 160 14036 200 14084
rect 160 14004 164 14036
rect 196 14004 200 14036
rect 160 13956 200 14004
rect 160 13924 164 13956
rect 196 13924 200 13956
rect 160 13876 200 13924
rect 160 13844 164 13876
rect 196 13844 200 13876
rect 160 13796 200 13844
rect 160 13764 164 13796
rect 196 13764 200 13796
rect 160 13716 200 13764
rect 160 13684 164 13716
rect 196 13684 200 13716
rect 160 13636 200 13684
rect 160 13604 164 13636
rect 196 13604 200 13636
rect 160 13556 200 13604
rect 160 13524 164 13556
rect 196 13524 200 13556
rect 160 13476 200 13524
rect 160 13444 164 13476
rect 196 13444 200 13476
rect 160 13396 200 13444
rect 160 13364 164 13396
rect 196 13364 200 13396
rect 160 13316 200 13364
rect 160 13284 164 13316
rect 196 13284 200 13316
rect 160 13236 200 13284
rect 160 13204 164 13236
rect 196 13204 200 13236
rect 160 13156 200 13204
rect 160 13124 164 13156
rect 196 13124 200 13156
rect 160 13076 200 13124
rect 160 13044 164 13076
rect 196 13044 200 13076
rect 160 12996 200 13044
rect 160 12964 164 12996
rect 196 12964 200 12996
rect 160 12916 200 12964
rect 160 12884 164 12916
rect 196 12884 200 12916
rect 160 12836 200 12884
rect 160 12804 164 12836
rect 196 12804 200 12836
rect 160 12756 200 12804
rect 160 12724 164 12756
rect 196 12724 200 12756
rect 160 12676 200 12724
rect 160 12644 164 12676
rect 196 12644 200 12676
rect 160 12596 200 12644
rect 160 12564 164 12596
rect 196 12564 200 12596
rect 160 12516 200 12564
rect 160 12484 164 12516
rect 196 12484 200 12516
rect 160 12436 200 12484
rect 160 12404 164 12436
rect 196 12404 200 12436
rect 160 12356 200 12404
rect 160 12324 164 12356
rect 196 12324 200 12356
rect 160 12276 200 12324
rect 160 12244 164 12276
rect 196 12244 200 12276
rect 160 12196 200 12244
rect 160 12164 164 12196
rect 196 12164 200 12196
rect 160 12116 200 12164
rect 160 12084 164 12116
rect 196 12084 200 12116
rect 160 12036 200 12084
rect 160 12004 164 12036
rect 196 12004 200 12036
rect 160 11956 200 12004
rect 160 11924 164 11956
rect 196 11924 200 11956
rect 160 11876 200 11924
rect 160 11844 164 11876
rect 196 11844 200 11876
rect 160 11796 200 11844
rect 160 11764 164 11796
rect 196 11764 200 11796
rect 160 11716 200 11764
rect 160 11684 164 11716
rect 196 11684 200 11716
rect 160 11636 200 11684
rect 160 11604 164 11636
rect 196 11604 200 11636
rect 160 11556 200 11604
rect 160 11524 164 11556
rect 196 11524 200 11556
rect 160 11476 200 11524
rect 160 11444 164 11476
rect 196 11444 200 11476
rect 160 11396 200 11444
rect 160 11364 164 11396
rect 196 11364 200 11396
rect 160 11236 200 11364
rect 160 11204 164 11236
rect 196 11204 200 11236
rect 160 11156 200 11204
rect 160 11124 164 11156
rect 196 11124 200 11156
rect 160 11076 200 11124
rect 160 11044 164 11076
rect 196 11044 200 11076
rect 160 10996 200 11044
rect 160 10964 164 10996
rect 196 10964 200 10996
rect 160 10916 200 10964
rect 160 10884 164 10916
rect 196 10884 200 10916
rect 160 10836 200 10884
rect 160 10804 164 10836
rect 196 10804 200 10836
rect 160 10756 200 10804
rect 160 10724 164 10756
rect 196 10724 200 10756
rect 160 10676 200 10724
rect 160 10644 164 10676
rect 196 10644 200 10676
rect 160 10596 200 10644
rect 160 10564 164 10596
rect 196 10564 200 10596
rect 160 10516 200 10564
rect 160 10484 164 10516
rect 196 10484 200 10516
rect 160 10436 200 10484
rect 160 10404 164 10436
rect 196 10404 200 10436
rect 160 10356 200 10404
rect 160 10324 164 10356
rect 196 10324 200 10356
rect 160 10276 200 10324
rect 160 10244 164 10276
rect 196 10244 200 10276
rect 160 10196 200 10244
rect 160 10164 164 10196
rect 196 10164 200 10196
rect 160 10116 200 10164
rect 160 10084 164 10116
rect 196 10084 200 10116
rect 160 10036 200 10084
rect 160 10004 164 10036
rect 196 10004 200 10036
rect 160 9956 200 10004
rect 160 9924 164 9956
rect 196 9924 200 9956
rect 160 9876 200 9924
rect 160 9844 164 9876
rect 196 9844 200 9876
rect 160 9796 200 9844
rect 160 9764 164 9796
rect 196 9764 200 9796
rect 160 9716 200 9764
rect 160 9684 164 9716
rect 196 9684 200 9716
rect 160 9636 200 9684
rect 160 9604 164 9636
rect 196 9604 200 9636
rect 160 9556 200 9604
rect 160 9524 164 9556
rect 196 9524 200 9556
rect 160 9476 200 9524
rect 160 9444 164 9476
rect 196 9444 200 9476
rect 160 9396 200 9444
rect 160 9364 164 9396
rect 196 9364 200 9396
rect 160 9316 200 9364
rect 160 9284 164 9316
rect 196 9284 200 9316
rect 160 9236 200 9284
rect 160 9204 164 9236
rect 196 9204 200 9236
rect 160 9156 200 9204
rect 160 9124 164 9156
rect 196 9124 200 9156
rect 160 9076 200 9124
rect 160 9044 164 9076
rect 196 9044 200 9076
rect 160 8996 200 9044
rect 160 8964 164 8996
rect 196 8964 200 8996
rect 160 8916 200 8964
rect 160 8884 164 8916
rect 196 8884 200 8916
rect 160 8836 200 8884
rect 160 8804 164 8836
rect 196 8804 200 8836
rect 160 8756 200 8804
rect 160 8724 164 8756
rect 196 8724 200 8756
rect 160 8676 200 8724
rect 160 8644 164 8676
rect 196 8644 200 8676
rect 160 8596 200 8644
rect 160 8564 164 8596
rect 196 8564 200 8596
rect 160 8516 200 8564
rect 160 8484 164 8516
rect 196 8484 200 8516
rect 160 8356 200 8484
rect 160 8324 164 8356
rect 196 8324 200 8356
rect 160 8276 200 8324
rect 160 8244 164 8276
rect 196 8244 200 8276
rect 160 8196 200 8244
rect 160 8164 164 8196
rect 196 8164 200 8196
rect 160 8116 200 8164
rect 160 8084 164 8116
rect 196 8084 200 8116
rect 160 7956 200 8084
rect 160 7924 164 7956
rect 196 7924 200 7956
rect 160 7876 200 7924
rect 160 7844 164 7876
rect 196 7844 200 7876
rect 160 7796 200 7844
rect 160 7764 164 7796
rect 196 7764 200 7796
rect 160 7716 200 7764
rect 160 7684 164 7716
rect 196 7684 200 7716
rect 160 7636 200 7684
rect 160 7604 164 7636
rect 196 7604 200 7636
rect 160 7556 200 7604
rect 160 7524 164 7556
rect 196 7524 200 7556
rect 160 7476 200 7524
rect 160 7444 164 7476
rect 196 7444 200 7476
rect 160 7396 200 7444
rect 160 7364 164 7396
rect 196 7364 200 7396
rect 160 7316 200 7364
rect 160 7284 164 7316
rect 196 7284 200 7316
rect 160 7236 200 7284
rect 160 7204 164 7236
rect 196 7204 200 7236
rect 160 7156 200 7204
rect 160 7124 164 7156
rect 196 7124 200 7156
rect 160 7076 200 7124
rect 160 7044 164 7076
rect 196 7044 200 7076
rect 160 6996 200 7044
rect 160 6964 164 6996
rect 196 6964 200 6996
rect 160 6916 200 6964
rect 160 6884 164 6916
rect 196 6884 200 6916
rect 160 6836 200 6884
rect 160 6804 164 6836
rect 196 6804 200 6836
rect 160 6756 200 6804
rect 160 6724 164 6756
rect 196 6724 200 6756
rect 160 6676 200 6724
rect 160 6644 164 6676
rect 196 6644 200 6676
rect 160 6596 200 6644
rect 160 6564 164 6596
rect 196 6564 200 6596
rect 160 6516 200 6564
rect 160 6484 164 6516
rect 196 6484 200 6516
rect 160 6436 200 6484
rect 160 6404 164 6436
rect 196 6404 200 6436
rect 160 6356 200 6404
rect 160 6324 164 6356
rect 196 6324 200 6356
rect 160 6276 200 6324
rect 160 6244 164 6276
rect 196 6244 200 6276
rect 160 6196 200 6244
rect 160 6164 164 6196
rect 196 6164 200 6196
rect 160 6116 200 6164
rect 160 6084 164 6116
rect 196 6084 200 6116
rect 160 6036 200 6084
rect 160 6004 164 6036
rect 196 6004 200 6036
rect 160 5956 200 6004
rect 160 5924 164 5956
rect 196 5924 200 5956
rect 160 5876 200 5924
rect 160 5844 164 5876
rect 196 5844 200 5876
rect 160 5796 200 5844
rect 160 5764 164 5796
rect 196 5764 200 5796
rect 160 5716 200 5764
rect 160 5684 164 5716
rect 196 5684 200 5716
rect 160 5636 200 5684
rect 160 5604 164 5636
rect 196 5604 200 5636
rect 160 5556 200 5604
rect 160 5524 164 5556
rect 196 5524 200 5556
rect 160 5476 200 5524
rect 160 5444 164 5476
rect 196 5444 200 5476
rect 160 5396 200 5444
rect 160 5364 164 5396
rect 196 5364 200 5396
rect 160 5316 200 5364
rect 160 5284 164 5316
rect 196 5284 200 5316
rect 160 5236 200 5284
rect 160 5204 164 5236
rect 196 5204 200 5236
rect 160 5076 200 5204
rect 160 5044 164 5076
rect 196 5044 200 5076
rect 160 4996 200 5044
rect 160 4964 164 4996
rect 196 4964 200 4996
rect 160 4916 200 4964
rect 160 4884 164 4916
rect 196 4884 200 4916
rect 160 4836 200 4884
rect 160 4804 164 4836
rect 196 4804 200 4836
rect 160 4756 200 4804
rect 160 4724 164 4756
rect 196 4724 200 4756
rect 160 4676 200 4724
rect 160 4644 164 4676
rect 196 4644 200 4676
rect 160 4596 200 4644
rect 160 4564 164 4596
rect 196 4564 200 4596
rect 160 4516 200 4564
rect 160 4484 164 4516
rect 196 4484 200 4516
rect 160 4436 200 4484
rect 160 4404 164 4436
rect 196 4404 200 4436
rect 160 4356 200 4404
rect 160 4324 164 4356
rect 196 4324 200 4356
rect 160 4276 200 4324
rect 160 4244 164 4276
rect 196 4244 200 4276
rect 160 4196 200 4244
rect 160 4164 164 4196
rect 196 4164 200 4196
rect 160 4116 200 4164
rect 160 4084 164 4116
rect 196 4084 200 4116
rect 160 4036 200 4084
rect 160 4004 164 4036
rect 196 4004 200 4036
rect 160 3956 200 4004
rect 160 3924 164 3956
rect 196 3924 200 3956
rect 160 3876 200 3924
rect 160 3844 164 3876
rect 196 3844 200 3876
rect 160 3796 200 3844
rect 160 3764 164 3796
rect 196 3764 200 3796
rect 160 3716 200 3764
rect 160 3684 164 3716
rect 196 3684 200 3716
rect 160 3636 200 3684
rect 160 3604 164 3636
rect 196 3604 200 3636
rect 160 3556 200 3604
rect 160 3524 164 3556
rect 196 3524 200 3556
rect 160 3476 200 3524
rect 160 3444 164 3476
rect 196 3444 200 3476
rect 160 3396 200 3444
rect 160 3364 164 3396
rect 196 3364 200 3396
rect 160 3316 200 3364
rect 160 3284 164 3316
rect 196 3284 200 3316
rect 160 3236 200 3284
rect 160 3204 164 3236
rect 196 3204 200 3236
rect 160 3156 200 3204
rect 160 3124 164 3156
rect 196 3124 200 3156
rect 160 3076 200 3124
rect 160 3044 164 3076
rect 196 3044 200 3076
rect 160 2996 200 3044
rect 160 2964 164 2996
rect 196 2964 200 2996
rect 160 2916 200 2964
rect 160 2884 164 2916
rect 196 2884 200 2916
rect 160 2836 200 2884
rect 160 2804 164 2836
rect 196 2804 200 2836
rect 160 2756 200 2804
rect 160 2724 164 2756
rect 196 2724 200 2756
rect 160 2676 200 2724
rect 160 2644 164 2676
rect 196 2644 200 2676
rect 160 2596 200 2644
rect 160 2564 164 2596
rect 196 2564 200 2596
rect 160 2516 200 2564
rect 160 2484 164 2516
rect 196 2484 200 2516
rect 160 2436 200 2484
rect 160 2404 164 2436
rect 196 2404 200 2436
rect 160 2356 200 2404
rect 160 2324 164 2356
rect 196 2324 200 2356
rect 160 2276 200 2324
rect 160 2244 164 2276
rect 196 2244 200 2276
rect 160 2196 200 2244
rect 160 2164 164 2196
rect 196 2164 200 2196
rect 160 2116 200 2164
rect 160 2084 164 2116
rect 196 2084 200 2116
rect 160 2036 200 2084
rect 160 2004 164 2036
rect 196 2004 200 2036
rect 160 1956 200 2004
rect 160 1924 164 1956
rect 196 1924 200 1956
rect 160 1876 200 1924
rect 160 1844 164 1876
rect 196 1844 200 1876
rect 160 1796 200 1844
rect 160 1764 164 1796
rect 196 1764 200 1796
rect 160 1716 200 1764
rect 160 1684 164 1716
rect 196 1684 200 1716
rect 160 1636 200 1684
rect 160 1604 164 1636
rect 196 1604 200 1636
rect 160 1556 200 1604
rect 160 1524 164 1556
rect 196 1524 200 1556
rect 160 1476 200 1524
rect 160 1444 164 1476
rect 196 1444 200 1476
rect 160 1396 200 1444
rect 160 1364 164 1396
rect 196 1364 200 1396
rect 160 1316 200 1364
rect 160 1284 164 1316
rect 196 1284 200 1316
rect 160 1236 200 1284
rect 160 1204 164 1236
rect 196 1204 200 1236
rect 160 1156 200 1204
rect 160 1124 164 1156
rect 196 1124 200 1156
rect 160 1076 200 1124
rect 160 1044 164 1076
rect 196 1044 200 1076
rect 160 996 200 1044
rect 160 964 164 996
rect 196 964 200 996
rect 160 916 200 964
rect 160 884 164 916
rect 196 884 200 916
rect 160 836 200 884
rect 160 804 164 836
rect 196 804 200 836
rect 160 756 200 804
rect 160 724 164 756
rect 196 724 200 756
rect 160 676 200 724
rect 160 644 164 676
rect 196 644 200 676
rect 160 596 200 644
rect 160 564 164 596
rect 196 564 200 596
rect 160 516 200 564
rect 160 484 164 516
rect 196 484 200 516
rect 0 244 4 436
rect 36 244 40 436
rect 0 240 40 244
rect 160 436 200 484
rect 240 11156 280 15960
rect 240 11124 244 11156
rect 276 11124 280 11156
rect 240 8596 280 11124
rect 240 8564 244 8596
rect 276 8564 280 8596
rect 240 7876 280 8564
rect 240 7844 244 7876
rect 276 7844 280 7876
rect 240 5316 280 7844
rect 240 5284 244 5316
rect 276 5284 280 5316
rect 240 480 280 5284
rect 320 15956 360 15960
rect 320 15924 324 15956
rect 356 15924 360 15956
rect 320 15876 360 15924
rect 320 15844 324 15876
rect 356 15844 360 15876
rect 320 15796 360 15844
rect 320 15764 324 15796
rect 356 15764 360 15796
rect 320 15716 360 15764
rect 320 15684 324 15716
rect 356 15684 360 15716
rect 320 15636 360 15684
rect 320 15604 324 15636
rect 356 15604 360 15636
rect 320 15556 360 15604
rect 320 15524 324 15556
rect 356 15524 360 15556
rect 320 15476 360 15524
rect 320 15444 324 15476
rect 356 15444 360 15476
rect 320 15396 360 15444
rect 320 15364 324 15396
rect 356 15364 360 15396
rect 320 15316 360 15364
rect 320 15284 324 15316
rect 356 15284 360 15316
rect 320 15236 360 15284
rect 320 15204 324 15236
rect 356 15204 360 15236
rect 320 15156 360 15204
rect 320 15124 324 15156
rect 356 15124 360 15156
rect 320 15076 360 15124
rect 320 15044 324 15076
rect 356 15044 360 15076
rect 320 14996 360 15044
rect 320 14964 324 14996
rect 356 14964 360 14996
rect 320 14916 360 14964
rect 320 14884 324 14916
rect 356 14884 360 14916
rect 320 14836 360 14884
rect 320 14804 324 14836
rect 356 14804 360 14836
rect 320 14756 360 14804
rect 320 14724 324 14756
rect 356 14724 360 14756
rect 320 14676 360 14724
rect 320 14644 324 14676
rect 356 14644 360 14676
rect 320 14596 360 14644
rect 320 14564 324 14596
rect 356 14564 360 14596
rect 320 14516 360 14564
rect 320 14484 324 14516
rect 356 14484 360 14516
rect 320 14436 360 14484
rect 320 14404 324 14436
rect 356 14404 360 14436
rect 320 14356 360 14404
rect 320 14324 324 14356
rect 356 14324 360 14356
rect 320 14276 360 14324
rect 320 14244 324 14276
rect 356 14244 360 14276
rect 320 14196 360 14244
rect 320 14164 324 14196
rect 356 14164 360 14196
rect 320 14116 360 14164
rect 320 14084 324 14116
rect 356 14084 360 14116
rect 320 14036 360 14084
rect 320 14004 324 14036
rect 356 14004 360 14036
rect 320 13956 360 14004
rect 320 13924 324 13956
rect 356 13924 360 13956
rect 320 13876 360 13924
rect 320 13844 324 13876
rect 356 13844 360 13876
rect 320 13796 360 13844
rect 320 13764 324 13796
rect 356 13764 360 13796
rect 320 13716 360 13764
rect 320 13684 324 13716
rect 356 13684 360 13716
rect 320 13636 360 13684
rect 320 13604 324 13636
rect 356 13604 360 13636
rect 320 13556 360 13604
rect 320 13524 324 13556
rect 356 13524 360 13556
rect 320 13476 360 13524
rect 320 13444 324 13476
rect 356 13444 360 13476
rect 320 13396 360 13444
rect 320 13364 324 13396
rect 356 13364 360 13396
rect 320 13316 360 13364
rect 320 13284 324 13316
rect 356 13284 360 13316
rect 320 13236 360 13284
rect 320 13204 324 13236
rect 356 13204 360 13236
rect 320 13156 360 13204
rect 320 13124 324 13156
rect 356 13124 360 13156
rect 320 13076 360 13124
rect 320 13044 324 13076
rect 356 13044 360 13076
rect 320 12996 360 13044
rect 320 12964 324 12996
rect 356 12964 360 12996
rect 320 12916 360 12964
rect 320 12884 324 12916
rect 356 12884 360 12916
rect 320 12836 360 12884
rect 320 12804 324 12836
rect 356 12804 360 12836
rect 320 12756 360 12804
rect 320 12724 324 12756
rect 356 12724 360 12756
rect 320 12676 360 12724
rect 320 12644 324 12676
rect 356 12644 360 12676
rect 320 12596 360 12644
rect 320 12564 324 12596
rect 356 12564 360 12596
rect 320 12516 360 12564
rect 320 12484 324 12516
rect 356 12484 360 12516
rect 320 12436 360 12484
rect 320 12404 324 12436
rect 356 12404 360 12436
rect 320 12356 360 12404
rect 320 12324 324 12356
rect 356 12324 360 12356
rect 320 12276 360 12324
rect 320 12244 324 12276
rect 356 12244 360 12276
rect 320 12196 360 12244
rect 320 12164 324 12196
rect 356 12164 360 12196
rect 320 12116 360 12164
rect 320 12084 324 12116
rect 356 12084 360 12116
rect 320 12036 360 12084
rect 320 12004 324 12036
rect 356 12004 360 12036
rect 320 11956 360 12004
rect 320 11924 324 11956
rect 356 11924 360 11956
rect 320 11876 360 11924
rect 320 11844 324 11876
rect 356 11844 360 11876
rect 320 11796 360 11844
rect 320 11764 324 11796
rect 356 11764 360 11796
rect 320 11716 360 11764
rect 320 11684 324 11716
rect 356 11684 360 11716
rect 320 11636 360 11684
rect 320 11604 324 11636
rect 356 11604 360 11636
rect 320 11556 360 11604
rect 320 11524 324 11556
rect 356 11524 360 11556
rect 320 11476 360 11524
rect 320 11444 324 11476
rect 356 11444 360 11476
rect 320 11396 360 11444
rect 320 11364 324 11396
rect 356 11364 360 11396
rect 320 11236 360 11364
rect 320 11204 324 11236
rect 356 11204 360 11236
rect 320 11076 360 11204
rect 320 11044 324 11076
rect 356 11044 360 11076
rect 320 10996 360 11044
rect 320 10964 324 10996
rect 356 10964 360 10996
rect 320 10916 360 10964
rect 320 10884 324 10916
rect 356 10884 360 10916
rect 320 10836 360 10884
rect 320 10804 324 10836
rect 356 10804 360 10836
rect 320 10756 360 10804
rect 320 10724 324 10756
rect 356 10724 360 10756
rect 320 10676 360 10724
rect 320 10644 324 10676
rect 356 10644 360 10676
rect 320 10596 360 10644
rect 320 10564 324 10596
rect 356 10564 360 10596
rect 320 10516 360 10564
rect 320 10484 324 10516
rect 356 10484 360 10516
rect 320 10436 360 10484
rect 320 10404 324 10436
rect 356 10404 360 10436
rect 320 10356 360 10404
rect 320 10324 324 10356
rect 356 10324 360 10356
rect 320 10276 360 10324
rect 320 10244 324 10276
rect 356 10244 360 10276
rect 320 10196 360 10244
rect 320 10164 324 10196
rect 356 10164 360 10196
rect 320 10116 360 10164
rect 320 10084 324 10116
rect 356 10084 360 10116
rect 320 10036 360 10084
rect 320 10004 324 10036
rect 356 10004 360 10036
rect 320 9956 360 10004
rect 320 9924 324 9956
rect 356 9924 360 9956
rect 320 9876 360 9924
rect 320 9844 324 9876
rect 356 9844 360 9876
rect 320 9796 360 9844
rect 320 9764 324 9796
rect 356 9764 360 9796
rect 320 9716 360 9764
rect 320 9684 324 9716
rect 356 9684 360 9716
rect 320 9636 360 9684
rect 320 9604 324 9636
rect 356 9604 360 9636
rect 320 9556 360 9604
rect 320 9524 324 9556
rect 356 9524 360 9556
rect 320 9476 360 9524
rect 320 9444 324 9476
rect 356 9444 360 9476
rect 320 9396 360 9444
rect 320 9364 324 9396
rect 356 9364 360 9396
rect 320 9316 360 9364
rect 320 9284 324 9316
rect 356 9284 360 9316
rect 320 9236 360 9284
rect 320 9204 324 9236
rect 356 9204 360 9236
rect 320 9156 360 9204
rect 320 9124 324 9156
rect 356 9124 360 9156
rect 320 9076 360 9124
rect 320 9044 324 9076
rect 356 9044 360 9076
rect 320 8996 360 9044
rect 320 8964 324 8996
rect 356 8964 360 8996
rect 320 8916 360 8964
rect 320 8884 324 8916
rect 356 8884 360 8916
rect 320 8836 360 8884
rect 320 8804 324 8836
rect 356 8804 360 8836
rect 320 8756 360 8804
rect 320 8724 324 8756
rect 356 8724 360 8756
rect 320 8676 360 8724
rect 320 8644 324 8676
rect 356 8644 360 8676
rect 320 8516 360 8644
rect 320 8484 324 8516
rect 356 8484 360 8516
rect 320 8356 360 8484
rect 320 8324 324 8356
rect 356 8324 360 8356
rect 320 8276 360 8324
rect 320 8244 324 8276
rect 356 8244 360 8276
rect 320 8196 360 8244
rect 320 8164 324 8196
rect 356 8164 360 8196
rect 320 8116 360 8164
rect 320 8084 324 8116
rect 356 8084 360 8116
rect 320 7956 360 8084
rect 320 7924 324 7956
rect 356 7924 360 7956
rect 320 7796 360 7924
rect 320 7764 324 7796
rect 356 7764 360 7796
rect 320 7716 360 7764
rect 320 7684 324 7716
rect 356 7684 360 7716
rect 320 7636 360 7684
rect 320 7604 324 7636
rect 356 7604 360 7636
rect 320 7556 360 7604
rect 320 7524 324 7556
rect 356 7524 360 7556
rect 320 7476 360 7524
rect 320 7444 324 7476
rect 356 7444 360 7476
rect 320 7396 360 7444
rect 320 7364 324 7396
rect 356 7364 360 7396
rect 320 7316 360 7364
rect 320 7284 324 7316
rect 356 7284 360 7316
rect 320 7236 360 7284
rect 320 7204 324 7236
rect 356 7204 360 7236
rect 320 7156 360 7204
rect 320 7124 324 7156
rect 356 7124 360 7156
rect 320 7076 360 7124
rect 320 7044 324 7076
rect 356 7044 360 7076
rect 320 6996 360 7044
rect 320 6964 324 6996
rect 356 6964 360 6996
rect 320 6916 360 6964
rect 320 6884 324 6916
rect 356 6884 360 6916
rect 320 6836 360 6884
rect 320 6804 324 6836
rect 356 6804 360 6836
rect 320 6756 360 6804
rect 320 6724 324 6756
rect 356 6724 360 6756
rect 320 6676 360 6724
rect 320 6644 324 6676
rect 356 6644 360 6676
rect 320 6596 360 6644
rect 320 6564 324 6596
rect 356 6564 360 6596
rect 320 6516 360 6564
rect 320 6484 324 6516
rect 356 6484 360 6516
rect 320 6436 360 6484
rect 320 6404 324 6436
rect 356 6404 360 6436
rect 320 6356 360 6404
rect 320 6324 324 6356
rect 356 6324 360 6356
rect 320 6276 360 6324
rect 320 6244 324 6276
rect 356 6244 360 6276
rect 320 6196 360 6244
rect 320 6164 324 6196
rect 356 6164 360 6196
rect 320 6116 360 6164
rect 320 6084 324 6116
rect 356 6084 360 6116
rect 320 6036 360 6084
rect 320 6004 324 6036
rect 356 6004 360 6036
rect 320 5956 360 6004
rect 320 5924 324 5956
rect 356 5924 360 5956
rect 320 5876 360 5924
rect 320 5844 324 5876
rect 356 5844 360 5876
rect 320 5796 360 5844
rect 320 5764 324 5796
rect 356 5764 360 5796
rect 320 5716 360 5764
rect 320 5684 324 5716
rect 356 5684 360 5716
rect 320 5636 360 5684
rect 320 5604 324 5636
rect 356 5604 360 5636
rect 320 5556 360 5604
rect 320 5524 324 5556
rect 356 5524 360 5556
rect 320 5476 360 5524
rect 320 5444 324 5476
rect 356 5444 360 5476
rect 320 5396 360 5444
rect 320 5364 324 5396
rect 356 5364 360 5396
rect 320 5236 360 5364
rect 320 5204 324 5236
rect 356 5204 360 5236
rect 320 5076 360 5204
rect 320 5044 324 5076
rect 356 5044 360 5076
rect 320 4996 360 5044
rect 320 4964 324 4996
rect 356 4964 360 4996
rect 320 4916 360 4964
rect 320 4884 324 4916
rect 356 4884 360 4916
rect 320 4836 360 4884
rect 320 4804 324 4836
rect 356 4804 360 4836
rect 320 4756 360 4804
rect 320 4724 324 4756
rect 356 4724 360 4756
rect 320 4676 360 4724
rect 320 4644 324 4676
rect 356 4644 360 4676
rect 320 4596 360 4644
rect 320 4564 324 4596
rect 356 4564 360 4596
rect 320 4516 360 4564
rect 320 4484 324 4516
rect 356 4484 360 4516
rect 320 4436 360 4484
rect 320 4404 324 4436
rect 356 4404 360 4436
rect 320 4356 360 4404
rect 320 4324 324 4356
rect 356 4324 360 4356
rect 320 4276 360 4324
rect 320 4244 324 4276
rect 356 4244 360 4276
rect 320 4196 360 4244
rect 320 4164 324 4196
rect 356 4164 360 4196
rect 320 4116 360 4164
rect 320 4084 324 4116
rect 356 4084 360 4116
rect 320 4036 360 4084
rect 320 4004 324 4036
rect 356 4004 360 4036
rect 320 3956 360 4004
rect 320 3924 324 3956
rect 356 3924 360 3956
rect 320 3876 360 3924
rect 320 3844 324 3876
rect 356 3844 360 3876
rect 320 3796 360 3844
rect 320 3764 324 3796
rect 356 3764 360 3796
rect 320 3716 360 3764
rect 320 3684 324 3716
rect 356 3684 360 3716
rect 320 3636 360 3684
rect 320 3604 324 3636
rect 356 3604 360 3636
rect 320 3556 360 3604
rect 320 3524 324 3556
rect 356 3524 360 3556
rect 320 3476 360 3524
rect 320 3444 324 3476
rect 356 3444 360 3476
rect 320 3396 360 3444
rect 320 3364 324 3396
rect 356 3364 360 3396
rect 320 3316 360 3364
rect 320 3284 324 3316
rect 356 3284 360 3316
rect 320 3236 360 3284
rect 320 3204 324 3236
rect 356 3204 360 3236
rect 320 3156 360 3204
rect 320 3124 324 3156
rect 356 3124 360 3156
rect 320 3076 360 3124
rect 320 3044 324 3076
rect 356 3044 360 3076
rect 320 2996 360 3044
rect 320 2964 324 2996
rect 356 2964 360 2996
rect 320 2916 360 2964
rect 320 2884 324 2916
rect 356 2884 360 2916
rect 320 2836 360 2884
rect 320 2804 324 2836
rect 356 2804 360 2836
rect 320 2756 360 2804
rect 320 2724 324 2756
rect 356 2724 360 2756
rect 320 2676 360 2724
rect 320 2644 324 2676
rect 356 2644 360 2676
rect 320 2596 360 2644
rect 320 2564 324 2596
rect 356 2564 360 2596
rect 320 2516 360 2564
rect 320 2484 324 2516
rect 356 2484 360 2516
rect 320 2436 360 2484
rect 320 2404 324 2436
rect 356 2404 360 2436
rect 320 2356 360 2404
rect 320 2324 324 2356
rect 356 2324 360 2356
rect 320 2276 360 2324
rect 320 2244 324 2276
rect 356 2244 360 2276
rect 320 2196 360 2244
rect 320 2164 324 2196
rect 356 2164 360 2196
rect 320 2116 360 2164
rect 320 2084 324 2116
rect 356 2084 360 2116
rect 320 2036 360 2084
rect 320 2004 324 2036
rect 356 2004 360 2036
rect 320 1956 360 2004
rect 320 1924 324 1956
rect 356 1924 360 1956
rect 320 1876 360 1924
rect 320 1844 324 1876
rect 356 1844 360 1876
rect 320 1796 360 1844
rect 320 1764 324 1796
rect 356 1764 360 1796
rect 320 1716 360 1764
rect 320 1684 324 1716
rect 356 1684 360 1716
rect 320 1636 360 1684
rect 320 1604 324 1636
rect 356 1604 360 1636
rect 320 1556 360 1604
rect 320 1524 324 1556
rect 356 1524 360 1556
rect 320 1476 360 1524
rect 320 1444 324 1476
rect 356 1444 360 1476
rect 320 1396 360 1444
rect 320 1364 324 1396
rect 356 1364 360 1396
rect 320 1316 360 1364
rect 320 1284 324 1316
rect 356 1284 360 1316
rect 320 1236 360 1284
rect 320 1204 324 1236
rect 356 1204 360 1236
rect 320 1156 360 1204
rect 320 1124 324 1156
rect 356 1124 360 1156
rect 320 1076 360 1124
rect 320 1044 324 1076
rect 356 1044 360 1076
rect 320 996 360 1044
rect 320 964 324 996
rect 356 964 360 996
rect 320 916 360 964
rect 320 884 324 916
rect 356 884 360 916
rect 320 836 360 884
rect 320 804 324 836
rect 356 804 360 836
rect 320 756 360 804
rect 320 724 324 756
rect 356 724 360 756
rect 320 676 360 724
rect 320 644 324 676
rect 356 644 360 676
rect 320 596 360 644
rect 320 564 324 596
rect 356 564 360 596
rect 320 516 360 564
rect 320 484 324 516
rect 356 484 360 516
rect 160 244 164 436
rect 196 244 200 436
rect 160 240 200 244
rect 320 436 360 484
rect 400 9876 440 15960
rect 400 9844 404 9876
rect 436 9844 440 9876
rect 400 6596 440 9844
rect 400 6564 404 6596
rect 436 6564 440 6596
rect 400 480 440 6564
rect 480 15956 520 15960
rect 480 15924 484 15956
rect 516 15924 520 15956
rect 480 15876 520 15924
rect 480 15844 484 15876
rect 516 15844 520 15876
rect 480 15796 520 15844
rect 480 15764 484 15796
rect 516 15764 520 15796
rect 480 15716 520 15764
rect 480 15684 484 15716
rect 516 15684 520 15716
rect 480 15636 520 15684
rect 480 15604 484 15636
rect 516 15604 520 15636
rect 480 15556 520 15604
rect 480 15524 484 15556
rect 516 15524 520 15556
rect 480 15476 520 15524
rect 480 15444 484 15476
rect 516 15444 520 15476
rect 480 15396 520 15444
rect 480 15364 484 15396
rect 516 15364 520 15396
rect 480 15316 520 15364
rect 480 15284 484 15316
rect 516 15284 520 15316
rect 480 15236 520 15284
rect 480 15204 484 15236
rect 516 15204 520 15236
rect 480 15156 520 15204
rect 480 15124 484 15156
rect 516 15124 520 15156
rect 480 15076 520 15124
rect 480 15044 484 15076
rect 516 15044 520 15076
rect 480 14996 520 15044
rect 480 14964 484 14996
rect 516 14964 520 14996
rect 480 14916 520 14964
rect 480 14884 484 14916
rect 516 14884 520 14916
rect 480 14836 520 14884
rect 480 14804 484 14836
rect 516 14804 520 14836
rect 480 14756 520 14804
rect 480 14724 484 14756
rect 516 14724 520 14756
rect 480 14676 520 14724
rect 480 14644 484 14676
rect 516 14644 520 14676
rect 480 14596 520 14644
rect 480 14564 484 14596
rect 516 14564 520 14596
rect 480 14516 520 14564
rect 480 14484 484 14516
rect 516 14484 520 14516
rect 480 14436 520 14484
rect 480 14404 484 14436
rect 516 14404 520 14436
rect 480 14356 520 14404
rect 480 14324 484 14356
rect 516 14324 520 14356
rect 480 14276 520 14324
rect 480 14244 484 14276
rect 516 14244 520 14276
rect 480 14196 520 14244
rect 480 14164 484 14196
rect 516 14164 520 14196
rect 480 14116 520 14164
rect 480 14084 484 14116
rect 516 14084 520 14116
rect 480 14036 520 14084
rect 480 14004 484 14036
rect 516 14004 520 14036
rect 480 13956 520 14004
rect 480 13924 484 13956
rect 516 13924 520 13956
rect 480 13876 520 13924
rect 480 13844 484 13876
rect 516 13844 520 13876
rect 480 13796 520 13844
rect 480 13764 484 13796
rect 516 13764 520 13796
rect 480 13716 520 13764
rect 480 13684 484 13716
rect 516 13684 520 13716
rect 480 13636 520 13684
rect 480 13604 484 13636
rect 516 13604 520 13636
rect 480 13556 520 13604
rect 480 13524 484 13556
rect 516 13524 520 13556
rect 480 13476 520 13524
rect 480 13444 484 13476
rect 516 13444 520 13476
rect 480 13396 520 13444
rect 480 13364 484 13396
rect 516 13364 520 13396
rect 480 13316 520 13364
rect 480 13284 484 13316
rect 516 13284 520 13316
rect 480 13236 520 13284
rect 480 13204 484 13236
rect 516 13204 520 13236
rect 480 13156 520 13204
rect 480 13124 484 13156
rect 516 13124 520 13156
rect 480 13076 520 13124
rect 480 13044 484 13076
rect 516 13044 520 13076
rect 480 12996 520 13044
rect 480 12964 484 12996
rect 516 12964 520 12996
rect 480 12916 520 12964
rect 480 12884 484 12916
rect 516 12884 520 12916
rect 480 12836 520 12884
rect 480 12804 484 12836
rect 516 12804 520 12836
rect 480 12756 520 12804
rect 480 12724 484 12756
rect 516 12724 520 12756
rect 480 12676 520 12724
rect 480 12644 484 12676
rect 516 12644 520 12676
rect 480 12596 520 12644
rect 480 12564 484 12596
rect 516 12564 520 12596
rect 480 12516 520 12564
rect 480 12484 484 12516
rect 516 12484 520 12516
rect 480 12436 520 12484
rect 480 12404 484 12436
rect 516 12404 520 12436
rect 480 12356 520 12404
rect 480 12324 484 12356
rect 516 12324 520 12356
rect 480 12276 520 12324
rect 480 12244 484 12276
rect 516 12244 520 12276
rect 480 12196 520 12244
rect 480 12164 484 12196
rect 516 12164 520 12196
rect 480 12116 520 12164
rect 480 12084 484 12116
rect 516 12084 520 12116
rect 480 12036 520 12084
rect 480 12004 484 12036
rect 516 12004 520 12036
rect 480 11956 520 12004
rect 480 11924 484 11956
rect 516 11924 520 11956
rect 480 11876 520 11924
rect 480 11844 484 11876
rect 516 11844 520 11876
rect 480 11796 520 11844
rect 480 11764 484 11796
rect 516 11764 520 11796
rect 480 11716 520 11764
rect 480 11684 484 11716
rect 516 11684 520 11716
rect 480 11636 520 11684
rect 480 11604 484 11636
rect 516 11604 520 11636
rect 480 11556 520 11604
rect 480 11524 484 11556
rect 516 11524 520 11556
rect 480 11476 520 11524
rect 480 11444 484 11476
rect 516 11444 520 11476
rect 480 11396 520 11444
rect 480 11364 484 11396
rect 516 11364 520 11396
rect 480 11236 520 11364
rect 480 11204 484 11236
rect 516 11204 520 11236
rect 480 11076 520 11204
rect 480 11044 484 11076
rect 516 11044 520 11076
rect 480 10996 520 11044
rect 480 10964 484 10996
rect 516 10964 520 10996
rect 480 10916 520 10964
rect 480 10884 484 10916
rect 516 10884 520 10916
rect 480 10836 520 10884
rect 480 10804 484 10836
rect 516 10804 520 10836
rect 480 10756 520 10804
rect 480 10724 484 10756
rect 516 10724 520 10756
rect 480 10676 520 10724
rect 480 10644 484 10676
rect 516 10644 520 10676
rect 480 10596 520 10644
rect 480 10564 484 10596
rect 516 10564 520 10596
rect 480 10516 520 10564
rect 480 10484 484 10516
rect 516 10484 520 10516
rect 480 10436 520 10484
rect 480 10404 484 10436
rect 516 10404 520 10436
rect 480 10356 520 10404
rect 480 10324 484 10356
rect 516 10324 520 10356
rect 480 10276 520 10324
rect 480 10244 484 10276
rect 516 10244 520 10276
rect 480 10196 520 10244
rect 480 10164 484 10196
rect 516 10164 520 10196
rect 480 10116 520 10164
rect 480 10084 484 10116
rect 516 10084 520 10116
rect 480 10036 520 10084
rect 480 10004 484 10036
rect 516 10004 520 10036
rect 480 9956 520 10004
rect 480 9924 484 9956
rect 516 9924 520 9956
rect 480 9796 520 9924
rect 480 9764 484 9796
rect 516 9764 520 9796
rect 480 9716 520 9764
rect 480 9684 484 9716
rect 516 9684 520 9716
rect 480 9636 520 9684
rect 480 9604 484 9636
rect 516 9604 520 9636
rect 480 9556 520 9604
rect 480 9524 484 9556
rect 516 9524 520 9556
rect 480 9476 520 9524
rect 480 9444 484 9476
rect 516 9444 520 9476
rect 480 9396 520 9444
rect 480 9364 484 9396
rect 516 9364 520 9396
rect 480 9316 520 9364
rect 480 9284 484 9316
rect 516 9284 520 9316
rect 480 9236 520 9284
rect 480 9204 484 9236
rect 516 9204 520 9236
rect 480 9156 520 9204
rect 480 9124 484 9156
rect 516 9124 520 9156
rect 480 9076 520 9124
rect 480 9044 484 9076
rect 516 9044 520 9076
rect 480 8996 520 9044
rect 480 8964 484 8996
rect 516 8964 520 8996
rect 480 8916 520 8964
rect 480 8884 484 8916
rect 516 8884 520 8916
rect 480 8836 520 8884
rect 480 8804 484 8836
rect 516 8804 520 8836
rect 480 8756 520 8804
rect 480 8724 484 8756
rect 516 8724 520 8756
rect 480 8676 520 8724
rect 480 8644 484 8676
rect 516 8644 520 8676
rect 480 8516 520 8644
rect 480 8484 484 8516
rect 516 8484 520 8516
rect 480 8356 520 8484
rect 480 8324 484 8356
rect 516 8324 520 8356
rect 480 8276 520 8324
rect 480 8244 484 8276
rect 516 8244 520 8276
rect 480 8196 520 8244
rect 480 8164 484 8196
rect 516 8164 520 8196
rect 480 8116 520 8164
rect 480 8084 484 8116
rect 516 8084 520 8116
rect 480 7956 520 8084
rect 480 7924 484 7956
rect 516 7924 520 7956
rect 480 7796 520 7924
rect 480 7764 484 7796
rect 516 7764 520 7796
rect 480 7716 520 7764
rect 480 7684 484 7716
rect 516 7684 520 7716
rect 480 7636 520 7684
rect 480 7604 484 7636
rect 516 7604 520 7636
rect 480 7556 520 7604
rect 480 7524 484 7556
rect 516 7524 520 7556
rect 480 7476 520 7524
rect 480 7444 484 7476
rect 516 7444 520 7476
rect 480 7396 520 7444
rect 480 7364 484 7396
rect 516 7364 520 7396
rect 480 7316 520 7364
rect 480 7284 484 7316
rect 516 7284 520 7316
rect 480 7236 520 7284
rect 480 7204 484 7236
rect 516 7204 520 7236
rect 480 7156 520 7204
rect 480 7124 484 7156
rect 516 7124 520 7156
rect 480 7076 520 7124
rect 480 7044 484 7076
rect 516 7044 520 7076
rect 480 6996 520 7044
rect 480 6964 484 6996
rect 516 6964 520 6996
rect 480 6916 520 6964
rect 480 6884 484 6916
rect 516 6884 520 6916
rect 480 6836 520 6884
rect 480 6804 484 6836
rect 516 6804 520 6836
rect 480 6756 520 6804
rect 480 6724 484 6756
rect 516 6724 520 6756
rect 480 6676 520 6724
rect 480 6644 484 6676
rect 516 6644 520 6676
rect 480 6516 520 6644
rect 480 6484 484 6516
rect 516 6484 520 6516
rect 480 6436 520 6484
rect 480 6404 484 6436
rect 516 6404 520 6436
rect 480 6356 520 6404
rect 480 6324 484 6356
rect 516 6324 520 6356
rect 480 6276 520 6324
rect 480 6244 484 6276
rect 516 6244 520 6276
rect 480 6196 520 6244
rect 480 6164 484 6196
rect 516 6164 520 6196
rect 480 6116 520 6164
rect 480 6084 484 6116
rect 516 6084 520 6116
rect 480 6036 520 6084
rect 480 6004 484 6036
rect 516 6004 520 6036
rect 480 5956 520 6004
rect 480 5924 484 5956
rect 516 5924 520 5956
rect 480 5876 520 5924
rect 480 5844 484 5876
rect 516 5844 520 5876
rect 480 5796 520 5844
rect 480 5764 484 5796
rect 516 5764 520 5796
rect 480 5716 520 5764
rect 480 5684 484 5716
rect 516 5684 520 5716
rect 480 5636 520 5684
rect 480 5604 484 5636
rect 516 5604 520 5636
rect 480 5556 520 5604
rect 480 5524 484 5556
rect 516 5524 520 5556
rect 480 5476 520 5524
rect 480 5444 484 5476
rect 516 5444 520 5476
rect 480 5396 520 5444
rect 480 5364 484 5396
rect 516 5364 520 5396
rect 480 5236 520 5364
rect 480 5204 484 5236
rect 516 5204 520 5236
rect 480 5076 520 5204
rect 480 5044 484 5076
rect 516 5044 520 5076
rect 480 4996 520 5044
rect 480 4964 484 4996
rect 516 4964 520 4996
rect 480 4916 520 4964
rect 480 4884 484 4916
rect 516 4884 520 4916
rect 480 4836 520 4884
rect 480 4804 484 4836
rect 516 4804 520 4836
rect 480 4756 520 4804
rect 480 4724 484 4756
rect 516 4724 520 4756
rect 480 4676 520 4724
rect 480 4644 484 4676
rect 516 4644 520 4676
rect 480 4596 520 4644
rect 480 4564 484 4596
rect 516 4564 520 4596
rect 480 4516 520 4564
rect 480 4484 484 4516
rect 516 4484 520 4516
rect 480 4436 520 4484
rect 480 4404 484 4436
rect 516 4404 520 4436
rect 480 4356 520 4404
rect 480 4324 484 4356
rect 516 4324 520 4356
rect 480 4276 520 4324
rect 480 4244 484 4276
rect 516 4244 520 4276
rect 480 4196 520 4244
rect 480 4164 484 4196
rect 516 4164 520 4196
rect 480 4116 520 4164
rect 480 4084 484 4116
rect 516 4084 520 4116
rect 480 4036 520 4084
rect 480 4004 484 4036
rect 516 4004 520 4036
rect 480 3956 520 4004
rect 480 3924 484 3956
rect 516 3924 520 3956
rect 480 3876 520 3924
rect 480 3844 484 3876
rect 516 3844 520 3876
rect 480 3796 520 3844
rect 480 3764 484 3796
rect 516 3764 520 3796
rect 480 3716 520 3764
rect 480 3684 484 3716
rect 516 3684 520 3716
rect 480 3636 520 3684
rect 480 3604 484 3636
rect 516 3604 520 3636
rect 480 3556 520 3604
rect 480 3524 484 3556
rect 516 3524 520 3556
rect 480 3476 520 3524
rect 480 3444 484 3476
rect 516 3444 520 3476
rect 480 3396 520 3444
rect 480 3364 484 3396
rect 516 3364 520 3396
rect 480 3316 520 3364
rect 480 3284 484 3316
rect 516 3284 520 3316
rect 480 3236 520 3284
rect 480 3204 484 3236
rect 516 3204 520 3236
rect 480 3156 520 3204
rect 480 3124 484 3156
rect 516 3124 520 3156
rect 480 3076 520 3124
rect 480 3044 484 3076
rect 516 3044 520 3076
rect 480 2996 520 3044
rect 480 2964 484 2996
rect 516 2964 520 2996
rect 480 2916 520 2964
rect 480 2884 484 2916
rect 516 2884 520 2916
rect 480 2836 520 2884
rect 480 2804 484 2836
rect 516 2804 520 2836
rect 480 2756 520 2804
rect 480 2724 484 2756
rect 516 2724 520 2756
rect 480 2676 520 2724
rect 480 2644 484 2676
rect 516 2644 520 2676
rect 480 2596 520 2644
rect 480 2564 484 2596
rect 516 2564 520 2596
rect 480 2516 520 2564
rect 480 2484 484 2516
rect 516 2484 520 2516
rect 480 2436 520 2484
rect 480 2404 484 2436
rect 516 2404 520 2436
rect 480 2356 520 2404
rect 480 2324 484 2356
rect 516 2324 520 2356
rect 480 2276 520 2324
rect 480 2244 484 2276
rect 516 2244 520 2276
rect 480 2196 520 2244
rect 480 2164 484 2196
rect 516 2164 520 2196
rect 480 2116 520 2164
rect 480 2084 484 2116
rect 516 2084 520 2116
rect 480 2036 520 2084
rect 480 2004 484 2036
rect 516 2004 520 2036
rect 480 1956 520 2004
rect 480 1924 484 1956
rect 516 1924 520 1956
rect 480 1876 520 1924
rect 480 1844 484 1876
rect 516 1844 520 1876
rect 480 1796 520 1844
rect 480 1764 484 1796
rect 516 1764 520 1796
rect 480 1716 520 1764
rect 480 1684 484 1716
rect 516 1684 520 1716
rect 480 1636 520 1684
rect 480 1604 484 1636
rect 516 1604 520 1636
rect 480 1556 520 1604
rect 480 1524 484 1556
rect 516 1524 520 1556
rect 480 1476 520 1524
rect 480 1444 484 1476
rect 516 1444 520 1476
rect 480 1396 520 1444
rect 480 1364 484 1396
rect 516 1364 520 1396
rect 480 1316 520 1364
rect 480 1284 484 1316
rect 516 1284 520 1316
rect 480 1236 520 1284
rect 480 1204 484 1236
rect 516 1204 520 1236
rect 480 1156 520 1204
rect 480 1124 484 1156
rect 516 1124 520 1156
rect 480 1076 520 1124
rect 480 1044 484 1076
rect 516 1044 520 1076
rect 480 996 520 1044
rect 480 964 484 996
rect 516 964 520 996
rect 480 916 520 964
rect 480 884 484 916
rect 516 884 520 916
rect 480 836 520 884
rect 480 804 484 836
rect 516 804 520 836
rect 480 756 520 804
rect 480 724 484 756
rect 516 724 520 756
rect 480 676 520 724
rect 480 644 484 676
rect 516 644 520 676
rect 480 596 520 644
rect 480 564 484 596
rect 516 564 520 596
rect 480 516 520 564
rect 14480 15956 14520 15960
rect 14480 15924 14484 15956
rect 14516 15924 14520 15956
rect 14480 15876 14520 15924
rect 14480 15844 14484 15876
rect 14516 15844 14520 15876
rect 14480 15796 14520 15844
rect 14480 15764 14484 15796
rect 14516 15764 14520 15796
rect 14480 15716 14520 15764
rect 14480 15684 14484 15716
rect 14516 15684 14520 15716
rect 14480 15636 14520 15684
rect 14480 15604 14484 15636
rect 14516 15604 14520 15636
rect 14480 15556 14520 15604
rect 14480 15524 14484 15556
rect 14516 15524 14520 15556
rect 14480 15476 14520 15524
rect 14480 15444 14484 15476
rect 14516 15444 14520 15476
rect 14480 15396 14520 15444
rect 14480 15364 14484 15396
rect 14516 15364 14520 15396
rect 14480 15316 14520 15364
rect 14480 15284 14484 15316
rect 14516 15284 14520 15316
rect 14480 15236 14520 15284
rect 14480 15204 14484 15236
rect 14516 15204 14520 15236
rect 14480 15156 14520 15204
rect 14480 15124 14484 15156
rect 14516 15124 14520 15156
rect 14480 15076 14520 15124
rect 14480 15044 14484 15076
rect 14516 15044 14520 15076
rect 14480 14996 14520 15044
rect 14480 14964 14484 14996
rect 14516 14964 14520 14996
rect 14480 14916 14520 14964
rect 14480 14884 14484 14916
rect 14516 14884 14520 14916
rect 14480 14836 14520 14884
rect 14480 14804 14484 14836
rect 14516 14804 14520 14836
rect 14480 14756 14520 14804
rect 14480 14724 14484 14756
rect 14516 14724 14520 14756
rect 14480 14676 14520 14724
rect 14480 14644 14484 14676
rect 14516 14644 14520 14676
rect 14480 14516 14520 14644
rect 14480 14484 14484 14516
rect 14516 14484 14520 14516
rect 14480 14356 14520 14484
rect 14480 14324 14484 14356
rect 14516 14324 14520 14356
rect 14480 14276 14520 14324
rect 14480 14244 14484 14276
rect 14516 14244 14520 14276
rect 14480 14196 14520 14244
rect 14480 14164 14484 14196
rect 14516 14164 14520 14196
rect 14480 14116 14520 14164
rect 14480 14084 14484 14116
rect 14516 14084 14520 14116
rect 14480 14036 14520 14084
rect 14480 14004 14484 14036
rect 14516 14004 14520 14036
rect 14480 13956 14520 14004
rect 14480 13924 14484 13956
rect 14516 13924 14520 13956
rect 14480 13876 14520 13924
rect 14480 13844 14484 13876
rect 14516 13844 14520 13876
rect 14480 13796 14520 13844
rect 14480 13764 14484 13796
rect 14516 13764 14520 13796
rect 14480 13716 14520 13764
rect 14480 13684 14484 13716
rect 14516 13684 14520 13716
rect 14480 13636 14520 13684
rect 14480 13604 14484 13636
rect 14516 13604 14520 13636
rect 14480 13556 14520 13604
rect 14480 13524 14484 13556
rect 14516 13524 14520 13556
rect 14480 13476 14520 13524
rect 14480 13444 14484 13476
rect 14516 13444 14520 13476
rect 14480 13396 14520 13444
rect 14480 13364 14484 13396
rect 14516 13364 14520 13396
rect 14480 13316 14520 13364
rect 14480 13284 14484 13316
rect 14516 13284 14520 13316
rect 14480 13236 14520 13284
rect 14480 13204 14484 13236
rect 14516 13204 14520 13236
rect 14480 13076 14520 13204
rect 14480 13044 14484 13076
rect 14516 13044 14520 13076
rect 14480 12996 14520 13044
rect 14480 12964 14484 12996
rect 14516 12964 14520 12996
rect 14480 12916 14520 12964
rect 14480 12884 14484 12916
rect 14516 12884 14520 12916
rect 14480 12836 14520 12884
rect 14480 12804 14484 12836
rect 14516 12804 14520 12836
rect 14480 12756 14520 12804
rect 14480 12724 14484 12756
rect 14516 12724 14520 12756
rect 14480 12676 14520 12724
rect 14480 12644 14484 12676
rect 14516 12644 14520 12676
rect 14480 12596 14520 12644
rect 14480 12564 14484 12596
rect 14516 12564 14520 12596
rect 14480 12516 14520 12564
rect 14480 12484 14484 12516
rect 14516 12484 14520 12516
rect 14480 12436 14520 12484
rect 14480 12404 14484 12436
rect 14516 12404 14520 12436
rect 14480 12356 14520 12404
rect 14480 12324 14484 12356
rect 14516 12324 14520 12356
rect 14480 12276 14520 12324
rect 14480 12244 14484 12276
rect 14516 12244 14520 12276
rect 14480 12196 14520 12244
rect 14480 12164 14484 12196
rect 14516 12164 14520 12196
rect 14480 12116 14520 12164
rect 14480 12084 14484 12116
rect 14516 12084 14520 12116
rect 14480 12036 14520 12084
rect 14480 12004 14484 12036
rect 14516 12004 14520 12036
rect 14480 11956 14520 12004
rect 14480 11924 14484 11956
rect 14516 11924 14520 11956
rect 14480 11796 14520 11924
rect 14480 11764 14484 11796
rect 14516 11764 14520 11796
rect 14480 11636 14520 11764
rect 14480 11604 14484 11636
rect 14516 11604 14520 11636
rect 14480 11556 14520 11604
rect 14480 11524 14484 11556
rect 14516 11524 14520 11556
rect 14480 11476 14520 11524
rect 14480 11444 14484 11476
rect 14516 11444 14520 11476
rect 14480 11396 14520 11444
rect 14480 11364 14484 11396
rect 14516 11364 14520 11396
rect 14480 11316 14520 11364
rect 14480 11284 14484 11316
rect 14516 11284 14520 11316
rect 14480 11236 14520 11284
rect 14480 11204 14484 11236
rect 14516 11204 14520 11236
rect 14480 11156 14520 11204
rect 14480 11124 14484 11156
rect 14516 11124 14520 11156
rect 14480 11076 14520 11124
rect 14480 11044 14484 11076
rect 14516 11044 14520 11076
rect 14480 10996 14520 11044
rect 14480 10964 14484 10996
rect 14516 10964 14520 10996
rect 14480 10916 14520 10964
rect 14480 10884 14484 10916
rect 14516 10884 14520 10916
rect 14480 10836 14520 10884
rect 14480 10804 14484 10836
rect 14516 10804 14520 10836
rect 14480 10756 14520 10804
rect 14480 10724 14484 10756
rect 14516 10724 14520 10756
rect 14480 10676 14520 10724
rect 14480 10644 14484 10676
rect 14516 10644 14520 10676
rect 14480 10596 14520 10644
rect 14480 10564 14484 10596
rect 14516 10564 14520 10596
rect 14480 10516 14520 10564
rect 14480 10484 14484 10516
rect 14516 10484 14520 10516
rect 14480 10436 14520 10484
rect 14480 10404 14484 10436
rect 14516 10404 14520 10436
rect 14480 10356 14520 10404
rect 14480 10324 14484 10356
rect 14516 10324 14520 10356
rect 14480 10276 14520 10324
rect 14480 10244 14484 10276
rect 14516 10244 14520 10276
rect 14480 10196 14520 10244
rect 14480 10164 14484 10196
rect 14516 10164 14520 10196
rect 14480 10116 14520 10164
rect 14480 10084 14484 10116
rect 14516 10084 14520 10116
rect 14480 10036 14520 10084
rect 14480 10004 14484 10036
rect 14516 10004 14520 10036
rect 14480 9956 14520 10004
rect 14480 9924 14484 9956
rect 14516 9924 14520 9956
rect 14480 9876 14520 9924
rect 14480 9844 14484 9876
rect 14516 9844 14520 9876
rect 14480 9796 14520 9844
rect 14480 9764 14484 9796
rect 14516 9764 14520 9796
rect 14480 9716 14520 9764
rect 14480 9684 14484 9716
rect 14516 9684 14520 9716
rect 14480 9636 14520 9684
rect 14480 9604 14484 9636
rect 14516 9604 14520 9636
rect 14480 9556 14520 9604
rect 14480 9524 14484 9556
rect 14516 9524 14520 9556
rect 14480 9476 14520 9524
rect 14480 9444 14484 9476
rect 14516 9444 14520 9476
rect 14480 9396 14520 9444
rect 14480 9364 14484 9396
rect 14516 9364 14520 9396
rect 14480 9316 14520 9364
rect 14480 9284 14484 9316
rect 14516 9284 14520 9316
rect 14480 9236 14520 9284
rect 14480 9204 14484 9236
rect 14516 9204 14520 9236
rect 14480 9156 14520 9204
rect 14480 9124 14484 9156
rect 14516 9124 14520 9156
rect 14480 9076 14520 9124
rect 14480 9044 14484 9076
rect 14516 9044 14520 9076
rect 14480 8996 14520 9044
rect 14480 8964 14484 8996
rect 14516 8964 14520 8996
rect 14480 8916 14520 8964
rect 14480 8884 14484 8916
rect 14516 8884 14520 8916
rect 14480 8836 14520 8884
rect 14480 8804 14484 8836
rect 14516 8804 14520 8836
rect 14480 8756 14520 8804
rect 14480 8724 14484 8756
rect 14516 8724 14520 8756
rect 14480 8676 14520 8724
rect 14480 8644 14484 8676
rect 14516 8644 14520 8676
rect 14480 8596 14520 8644
rect 14480 8564 14484 8596
rect 14516 8564 14520 8596
rect 14480 8516 14520 8564
rect 14480 8484 14484 8516
rect 14516 8484 14520 8516
rect 14480 8436 14520 8484
rect 14480 8404 14484 8436
rect 14516 8404 14520 8436
rect 14480 8356 14520 8404
rect 14480 8324 14484 8356
rect 14516 8324 14520 8356
rect 14480 8276 14520 8324
rect 14480 8244 14484 8276
rect 14516 8244 14520 8276
rect 14480 8196 14520 8244
rect 14480 8164 14484 8196
rect 14516 8164 14520 8196
rect 14480 8116 14520 8164
rect 14480 8084 14484 8116
rect 14516 8084 14520 8116
rect 14480 8036 14520 8084
rect 14480 8004 14484 8036
rect 14516 8004 14520 8036
rect 14480 7956 14520 8004
rect 14480 7924 14484 7956
rect 14516 7924 14520 7956
rect 14480 7876 14520 7924
rect 14480 7844 14484 7876
rect 14516 7844 14520 7876
rect 14480 7796 14520 7844
rect 14480 7764 14484 7796
rect 14516 7764 14520 7796
rect 14480 7716 14520 7764
rect 14480 7684 14484 7716
rect 14516 7684 14520 7716
rect 14480 7636 14520 7684
rect 14480 7604 14484 7636
rect 14516 7604 14520 7636
rect 14480 7556 14520 7604
rect 14480 7524 14484 7556
rect 14516 7524 14520 7556
rect 14480 7476 14520 7524
rect 14480 7444 14484 7476
rect 14516 7444 14520 7476
rect 14480 7396 14520 7444
rect 14480 7364 14484 7396
rect 14516 7364 14520 7396
rect 14480 7316 14520 7364
rect 14480 7284 14484 7316
rect 14516 7284 14520 7316
rect 14480 7236 14520 7284
rect 14480 7204 14484 7236
rect 14516 7204 14520 7236
rect 14480 7156 14520 7204
rect 14480 7124 14484 7156
rect 14516 7124 14520 7156
rect 14480 7076 14520 7124
rect 14480 7044 14484 7076
rect 14516 7044 14520 7076
rect 14480 6996 14520 7044
rect 14480 6964 14484 6996
rect 14516 6964 14520 6996
rect 14480 6916 14520 6964
rect 14480 6884 14484 6916
rect 14516 6884 14520 6916
rect 14480 6836 14520 6884
rect 14480 6804 14484 6836
rect 14516 6804 14520 6836
rect 14480 6756 14520 6804
rect 14480 6724 14484 6756
rect 14516 6724 14520 6756
rect 14480 6676 14520 6724
rect 14480 6644 14484 6676
rect 14516 6644 14520 6676
rect 14480 6596 14520 6644
rect 14480 6564 14484 6596
rect 14516 6564 14520 6596
rect 14480 6516 14520 6564
rect 14480 6484 14484 6516
rect 14516 6484 14520 6516
rect 14480 6436 14520 6484
rect 14480 6404 14484 6436
rect 14516 6404 14520 6436
rect 14480 6356 14520 6404
rect 14480 6324 14484 6356
rect 14516 6324 14520 6356
rect 14480 6276 14520 6324
rect 14480 6244 14484 6276
rect 14516 6244 14520 6276
rect 14480 6196 14520 6244
rect 14480 6164 14484 6196
rect 14516 6164 14520 6196
rect 14480 6116 14520 6164
rect 14480 6084 14484 6116
rect 14516 6084 14520 6116
rect 14480 6036 14520 6084
rect 14480 6004 14484 6036
rect 14516 6004 14520 6036
rect 14480 5956 14520 6004
rect 14480 5924 14484 5956
rect 14516 5924 14520 5956
rect 14480 5876 14520 5924
rect 14480 5844 14484 5876
rect 14516 5844 14520 5876
rect 14480 5796 14520 5844
rect 14480 5764 14484 5796
rect 14516 5764 14520 5796
rect 14480 5716 14520 5764
rect 14480 5684 14484 5716
rect 14516 5684 14520 5716
rect 14480 5636 14520 5684
rect 14480 5604 14484 5636
rect 14516 5604 14520 5636
rect 14480 5556 14520 5604
rect 14480 5524 14484 5556
rect 14516 5524 14520 5556
rect 14480 5476 14520 5524
rect 14480 5444 14484 5476
rect 14516 5444 14520 5476
rect 14480 5396 14520 5444
rect 14480 5364 14484 5396
rect 14516 5364 14520 5396
rect 14480 5316 14520 5364
rect 14480 5284 14484 5316
rect 14516 5284 14520 5316
rect 14480 5236 14520 5284
rect 14480 5204 14484 5236
rect 14516 5204 14520 5236
rect 14480 5156 14520 5204
rect 14480 5124 14484 5156
rect 14516 5124 14520 5156
rect 14480 5076 14520 5124
rect 14480 5044 14484 5076
rect 14516 5044 14520 5076
rect 14480 4996 14520 5044
rect 14480 4964 14484 4996
rect 14516 4964 14520 4996
rect 14480 4916 14520 4964
rect 14480 4884 14484 4916
rect 14516 4884 14520 4916
rect 14480 4836 14520 4884
rect 14480 4804 14484 4836
rect 14516 4804 14520 4836
rect 14480 4676 14520 4804
rect 14480 4644 14484 4676
rect 14516 4644 14520 4676
rect 14480 4516 14520 4644
rect 14480 4484 14484 4516
rect 14516 4484 14520 4516
rect 14480 4436 14520 4484
rect 14480 4404 14484 4436
rect 14516 4404 14520 4436
rect 14480 4356 14520 4404
rect 14480 4324 14484 4356
rect 14516 4324 14520 4356
rect 14480 4276 14520 4324
rect 14480 4244 14484 4276
rect 14516 4244 14520 4276
rect 14480 4196 14520 4244
rect 14480 4164 14484 4196
rect 14516 4164 14520 4196
rect 14480 4116 14520 4164
rect 14480 4084 14484 4116
rect 14516 4084 14520 4116
rect 14480 4036 14520 4084
rect 14480 4004 14484 4036
rect 14516 4004 14520 4036
rect 14480 3956 14520 4004
rect 14480 3924 14484 3956
rect 14516 3924 14520 3956
rect 14480 3876 14520 3924
rect 14480 3844 14484 3876
rect 14516 3844 14520 3876
rect 14480 3796 14520 3844
rect 14480 3764 14484 3796
rect 14516 3764 14520 3796
rect 14480 3716 14520 3764
rect 14480 3684 14484 3716
rect 14516 3684 14520 3716
rect 14480 3636 14520 3684
rect 14480 3604 14484 3636
rect 14516 3604 14520 3636
rect 14480 3556 14520 3604
rect 14480 3524 14484 3556
rect 14516 3524 14520 3556
rect 14480 3476 14520 3524
rect 14480 3444 14484 3476
rect 14516 3444 14520 3476
rect 14480 3396 14520 3444
rect 14480 3364 14484 3396
rect 14516 3364 14520 3396
rect 14480 3236 14520 3364
rect 14480 3204 14484 3236
rect 14516 3204 14520 3236
rect 14480 3156 14520 3204
rect 14480 3124 14484 3156
rect 14516 3124 14520 3156
rect 14480 3076 14520 3124
rect 14480 3044 14484 3076
rect 14516 3044 14520 3076
rect 14480 2996 14520 3044
rect 14480 2964 14484 2996
rect 14516 2964 14520 2996
rect 14480 2916 14520 2964
rect 14480 2884 14484 2916
rect 14516 2884 14520 2916
rect 14480 2836 14520 2884
rect 14480 2804 14484 2836
rect 14516 2804 14520 2836
rect 14480 2756 14520 2804
rect 14480 2724 14484 2756
rect 14516 2724 14520 2756
rect 14480 2676 14520 2724
rect 14480 2644 14484 2676
rect 14516 2644 14520 2676
rect 14480 2596 14520 2644
rect 14480 2564 14484 2596
rect 14516 2564 14520 2596
rect 14480 2516 14520 2564
rect 14480 2484 14484 2516
rect 14516 2484 14520 2516
rect 14480 2436 14520 2484
rect 14480 2404 14484 2436
rect 14516 2404 14520 2436
rect 14480 2356 14520 2404
rect 14480 2324 14484 2356
rect 14516 2324 14520 2356
rect 14480 2276 14520 2324
rect 14480 2244 14484 2276
rect 14516 2244 14520 2276
rect 14480 2196 14520 2244
rect 14480 2164 14484 2196
rect 14516 2164 14520 2196
rect 14480 2116 14520 2164
rect 14480 2084 14484 2116
rect 14516 2084 14520 2116
rect 14480 1956 14520 2084
rect 14480 1924 14484 1956
rect 14516 1924 14520 1956
rect 14480 1796 14520 1924
rect 14480 1764 14484 1796
rect 14516 1764 14520 1796
rect 14480 1716 14520 1764
rect 14480 1684 14484 1716
rect 14516 1684 14520 1716
rect 14480 1636 14520 1684
rect 14480 1604 14484 1636
rect 14516 1604 14520 1636
rect 14480 1556 14520 1604
rect 14480 1524 14484 1556
rect 14516 1524 14520 1556
rect 14480 1476 14520 1524
rect 14480 1444 14484 1476
rect 14516 1444 14520 1476
rect 14480 1396 14520 1444
rect 14480 1364 14484 1396
rect 14516 1364 14520 1396
rect 14480 1316 14520 1364
rect 14480 1284 14484 1316
rect 14516 1284 14520 1316
rect 14480 1236 14520 1284
rect 14480 1204 14484 1236
rect 14516 1204 14520 1236
rect 14480 1156 14520 1204
rect 14480 1124 14484 1156
rect 14516 1124 14520 1156
rect 14480 1076 14520 1124
rect 14480 1044 14484 1076
rect 14516 1044 14520 1076
rect 14480 996 14520 1044
rect 14480 964 14484 996
rect 14516 964 14520 996
rect 14480 916 14520 964
rect 14480 884 14484 916
rect 14516 884 14520 916
rect 14480 836 14520 884
rect 14480 804 14484 836
rect 14516 804 14520 836
rect 14480 756 14520 804
rect 14480 724 14484 756
rect 14516 724 14520 756
rect 14480 676 14520 724
rect 14480 644 14484 676
rect 14516 644 14520 676
rect 14480 596 14520 644
rect 14480 564 14484 596
rect 14516 564 14520 596
rect 480 484 484 516
rect 516 484 520 516
rect 320 244 324 436
rect 356 244 360 436
rect 320 240 360 244
rect 480 436 520 484
rect 480 244 484 436
rect 516 244 520 436
rect 480 240 520 244
rect 560 515 600 520
rect 560 485 565 515
rect 595 485 600 515
rect 560 196 600 485
rect 560 4 564 196
rect 596 4 600 196
rect 560 0 600 4
rect 14400 515 14440 520
rect 14400 485 14405 515
rect 14435 485 14440 515
rect 14400 196 14440 485
rect 14480 516 14520 564
rect 14480 484 14484 516
rect 14516 484 14520 516
rect 14480 436 14520 484
rect 14560 13156 14600 15960
rect 14560 13124 14564 13156
rect 14596 13124 14600 13156
rect 14560 3316 14600 13124
rect 14560 3284 14564 3316
rect 14596 3284 14600 3316
rect 14560 480 14600 3284
rect 14640 15956 14680 15960
rect 14640 15924 14644 15956
rect 14676 15924 14680 15956
rect 14640 15876 14680 15924
rect 14640 15844 14644 15876
rect 14676 15844 14680 15876
rect 14640 15796 14680 15844
rect 14640 15764 14644 15796
rect 14676 15764 14680 15796
rect 14640 15716 14680 15764
rect 14640 15684 14644 15716
rect 14676 15684 14680 15716
rect 14640 15636 14680 15684
rect 14640 15604 14644 15636
rect 14676 15604 14680 15636
rect 14640 15556 14680 15604
rect 14640 15524 14644 15556
rect 14676 15524 14680 15556
rect 14640 15476 14680 15524
rect 14640 15444 14644 15476
rect 14676 15444 14680 15476
rect 14640 15396 14680 15444
rect 14640 15364 14644 15396
rect 14676 15364 14680 15396
rect 14640 15316 14680 15364
rect 14640 15284 14644 15316
rect 14676 15284 14680 15316
rect 14640 15236 14680 15284
rect 14640 15204 14644 15236
rect 14676 15204 14680 15236
rect 14640 15156 14680 15204
rect 14640 15124 14644 15156
rect 14676 15124 14680 15156
rect 14640 15076 14680 15124
rect 14640 15044 14644 15076
rect 14676 15044 14680 15076
rect 14640 14996 14680 15044
rect 14640 14964 14644 14996
rect 14676 14964 14680 14996
rect 14640 14916 14680 14964
rect 14640 14884 14644 14916
rect 14676 14884 14680 14916
rect 14640 14836 14680 14884
rect 14640 14804 14644 14836
rect 14676 14804 14680 14836
rect 14640 14756 14680 14804
rect 14640 14724 14644 14756
rect 14676 14724 14680 14756
rect 14640 14676 14680 14724
rect 14640 14644 14644 14676
rect 14676 14644 14680 14676
rect 14640 14516 14680 14644
rect 14640 14484 14644 14516
rect 14676 14484 14680 14516
rect 14640 14356 14680 14484
rect 14640 14324 14644 14356
rect 14676 14324 14680 14356
rect 14640 14276 14680 14324
rect 14640 14244 14644 14276
rect 14676 14244 14680 14276
rect 14640 14196 14680 14244
rect 14640 14164 14644 14196
rect 14676 14164 14680 14196
rect 14640 14116 14680 14164
rect 14640 14084 14644 14116
rect 14676 14084 14680 14116
rect 14640 14036 14680 14084
rect 14640 14004 14644 14036
rect 14676 14004 14680 14036
rect 14640 13956 14680 14004
rect 14640 13924 14644 13956
rect 14676 13924 14680 13956
rect 14640 13876 14680 13924
rect 14640 13844 14644 13876
rect 14676 13844 14680 13876
rect 14640 13796 14680 13844
rect 14640 13764 14644 13796
rect 14676 13764 14680 13796
rect 14640 13716 14680 13764
rect 14640 13684 14644 13716
rect 14676 13684 14680 13716
rect 14640 13636 14680 13684
rect 14640 13604 14644 13636
rect 14676 13604 14680 13636
rect 14640 13556 14680 13604
rect 14640 13524 14644 13556
rect 14676 13524 14680 13556
rect 14640 13476 14680 13524
rect 14640 13444 14644 13476
rect 14676 13444 14680 13476
rect 14640 13396 14680 13444
rect 14640 13364 14644 13396
rect 14676 13364 14680 13396
rect 14640 13316 14680 13364
rect 14640 13284 14644 13316
rect 14676 13284 14680 13316
rect 14640 13236 14680 13284
rect 14640 13204 14644 13236
rect 14676 13204 14680 13236
rect 14640 13156 14680 13204
rect 14640 13124 14644 13156
rect 14676 13124 14680 13156
rect 14640 13076 14680 13124
rect 14640 13044 14644 13076
rect 14676 13044 14680 13076
rect 14640 12996 14680 13044
rect 14640 12964 14644 12996
rect 14676 12964 14680 12996
rect 14640 12916 14680 12964
rect 14640 12884 14644 12916
rect 14676 12884 14680 12916
rect 14640 12836 14680 12884
rect 14640 12804 14644 12836
rect 14676 12804 14680 12836
rect 14640 12756 14680 12804
rect 14640 12724 14644 12756
rect 14676 12724 14680 12756
rect 14640 12676 14680 12724
rect 14640 12644 14644 12676
rect 14676 12644 14680 12676
rect 14640 12596 14680 12644
rect 14640 12564 14644 12596
rect 14676 12564 14680 12596
rect 14640 12516 14680 12564
rect 14640 12484 14644 12516
rect 14676 12484 14680 12516
rect 14640 12436 14680 12484
rect 14640 12404 14644 12436
rect 14676 12404 14680 12436
rect 14640 12356 14680 12404
rect 14640 12324 14644 12356
rect 14676 12324 14680 12356
rect 14640 12276 14680 12324
rect 14640 12244 14644 12276
rect 14676 12244 14680 12276
rect 14640 12196 14680 12244
rect 14640 12164 14644 12196
rect 14676 12164 14680 12196
rect 14640 12116 14680 12164
rect 14640 12084 14644 12116
rect 14676 12084 14680 12116
rect 14640 12036 14680 12084
rect 14640 12004 14644 12036
rect 14676 12004 14680 12036
rect 14640 11956 14680 12004
rect 14640 11924 14644 11956
rect 14676 11924 14680 11956
rect 14640 11796 14680 11924
rect 14640 11764 14644 11796
rect 14676 11764 14680 11796
rect 14640 11636 14680 11764
rect 14640 11604 14644 11636
rect 14676 11604 14680 11636
rect 14640 11556 14680 11604
rect 14640 11524 14644 11556
rect 14676 11524 14680 11556
rect 14640 11476 14680 11524
rect 14640 11444 14644 11476
rect 14676 11444 14680 11476
rect 14640 11396 14680 11444
rect 14640 11364 14644 11396
rect 14676 11364 14680 11396
rect 14640 11316 14680 11364
rect 14640 11284 14644 11316
rect 14676 11284 14680 11316
rect 14640 11236 14680 11284
rect 14640 11204 14644 11236
rect 14676 11204 14680 11236
rect 14640 11156 14680 11204
rect 14640 11124 14644 11156
rect 14676 11124 14680 11156
rect 14640 11076 14680 11124
rect 14640 11044 14644 11076
rect 14676 11044 14680 11076
rect 14640 10996 14680 11044
rect 14640 10964 14644 10996
rect 14676 10964 14680 10996
rect 14640 10916 14680 10964
rect 14640 10884 14644 10916
rect 14676 10884 14680 10916
rect 14640 10836 14680 10884
rect 14640 10804 14644 10836
rect 14676 10804 14680 10836
rect 14640 10756 14680 10804
rect 14640 10724 14644 10756
rect 14676 10724 14680 10756
rect 14640 10676 14680 10724
rect 14640 10644 14644 10676
rect 14676 10644 14680 10676
rect 14640 10596 14680 10644
rect 14640 10564 14644 10596
rect 14676 10564 14680 10596
rect 14640 10516 14680 10564
rect 14640 10484 14644 10516
rect 14676 10484 14680 10516
rect 14640 10436 14680 10484
rect 14640 10404 14644 10436
rect 14676 10404 14680 10436
rect 14640 10356 14680 10404
rect 14640 10324 14644 10356
rect 14676 10324 14680 10356
rect 14640 10276 14680 10324
rect 14640 10244 14644 10276
rect 14676 10244 14680 10276
rect 14640 10196 14680 10244
rect 14640 10164 14644 10196
rect 14676 10164 14680 10196
rect 14640 10116 14680 10164
rect 14640 10084 14644 10116
rect 14676 10084 14680 10116
rect 14640 10036 14680 10084
rect 14640 10004 14644 10036
rect 14676 10004 14680 10036
rect 14640 9956 14680 10004
rect 14640 9924 14644 9956
rect 14676 9924 14680 9956
rect 14640 9876 14680 9924
rect 14640 9844 14644 9876
rect 14676 9844 14680 9876
rect 14640 9796 14680 9844
rect 14640 9764 14644 9796
rect 14676 9764 14680 9796
rect 14640 9716 14680 9764
rect 14640 9684 14644 9716
rect 14676 9684 14680 9716
rect 14640 9636 14680 9684
rect 14640 9604 14644 9636
rect 14676 9604 14680 9636
rect 14640 9556 14680 9604
rect 14640 9524 14644 9556
rect 14676 9524 14680 9556
rect 14640 9476 14680 9524
rect 14640 9444 14644 9476
rect 14676 9444 14680 9476
rect 14640 9396 14680 9444
rect 14640 9364 14644 9396
rect 14676 9364 14680 9396
rect 14640 9316 14680 9364
rect 14640 9284 14644 9316
rect 14676 9284 14680 9316
rect 14640 9236 14680 9284
rect 14640 9204 14644 9236
rect 14676 9204 14680 9236
rect 14640 9156 14680 9204
rect 14640 9124 14644 9156
rect 14676 9124 14680 9156
rect 14640 9076 14680 9124
rect 14640 9044 14644 9076
rect 14676 9044 14680 9076
rect 14640 8996 14680 9044
rect 14640 8964 14644 8996
rect 14676 8964 14680 8996
rect 14640 8916 14680 8964
rect 14640 8884 14644 8916
rect 14676 8884 14680 8916
rect 14640 8836 14680 8884
rect 14640 8804 14644 8836
rect 14676 8804 14680 8836
rect 14640 8756 14680 8804
rect 14640 8724 14644 8756
rect 14676 8724 14680 8756
rect 14640 8676 14680 8724
rect 14640 8644 14644 8676
rect 14676 8644 14680 8676
rect 14640 8596 14680 8644
rect 14640 8564 14644 8596
rect 14676 8564 14680 8596
rect 14640 8516 14680 8564
rect 14640 8484 14644 8516
rect 14676 8484 14680 8516
rect 14640 8436 14680 8484
rect 14640 8404 14644 8436
rect 14676 8404 14680 8436
rect 14640 8356 14680 8404
rect 14640 8324 14644 8356
rect 14676 8324 14680 8356
rect 14640 8276 14680 8324
rect 14640 8244 14644 8276
rect 14676 8244 14680 8276
rect 14640 8196 14680 8244
rect 14640 8164 14644 8196
rect 14676 8164 14680 8196
rect 14640 8116 14680 8164
rect 14640 8084 14644 8116
rect 14676 8084 14680 8116
rect 14640 8036 14680 8084
rect 14640 8004 14644 8036
rect 14676 8004 14680 8036
rect 14640 7956 14680 8004
rect 14640 7924 14644 7956
rect 14676 7924 14680 7956
rect 14640 7876 14680 7924
rect 14640 7844 14644 7876
rect 14676 7844 14680 7876
rect 14640 7796 14680 7844
rect 14640 7764 14644 7796
rect 14676 7764 14680 7796
rect 14640 7716 14680 7764
rect 14640 7684 14644 7716
rect 14676 7684 14680 7716
rect 14640 7636 14680 7684
rect 14640 7604 14644 7636
rect 14676 7604 14680 7636
rect 14640 7556 14680 7604
rect 14640 7524 14644 7556
rect 14676 7524 14680 7556
rect 14640 7476 14680 7524
rect 14640 7444 14644 7476
rect 14676 7444 14680 7476
rect 14640 7396 14680 7444
rect 14640 7364 14644 7396
rect 14676 7364 14680 7396
rect 14640 7316 14680 7364
rect 14640 7284 14644 7316
rect 14676 7284 14680 7316
rect 14640 7236 14680 7284
rect 14640 7204 14644 7236
rect 14676 7204 14680 7236
rect 14640 7156 14680 7204
rect 14640 7124 14644 7156
rect 14676 7124 14680 7156
rect 14640 7076 14680 7124
rect 14640 7044 14644 7076
rect 14676 7044 14680 7076
rect 14640 6996 14680 7044
rect 14640 6964 14644 6996
rect 14676 6964 14680 6996
rect 14640 6916 14680 6964
rect 14640 6884 14644 6916
rect 14676 6884 14680 6916
rect 14640 6836 14680 6884
rect 14640 6804 14644 6836
rect 14676 6804 14680 6836
rect 14640 6756 14680 6804
rect 14640 6724 14644 6756
rect 14676 6724 14680 6756
rect 14640 6676 14680 6724
rect 14640 6644 14644 6676
rect 14676 6644 14680 6676
rect 14640 6596 14680 6644
rect 14640 6564 14644 6596
rect 14676 6564 14680 6596
rect 14640 6516 14680 6564
rect 14640 6484 14644 6516
rect 14676 6484 14680 6516
rect 14640 6436 14680 6484
rect 14640 6404 14644 6436
rect 14676 6404 14680 6436
rect 14640 6356 14680 6404
rect 14640 6324 14644 6356
rect 14676 6324 14680 6356
rect 14640 6276 14680 6324
rect 14640 6244 14644 6276
rect 14676 6244 14680 6276
rect 14640 6196 14680 6244
rect 14640 6164 14644 6196
rect 14676 6164 14680 6196
rect 14640 6116 14680 6164
rect 14640 6084 14644 6116
rect 14676 6084 14680 6116
rect 14640 6036 14680 6084
rect 14640 6004 14644 6036
rect 14676 6004 14680 6036
rect 14640 5956 14680 6004
rect 14640 5924 14644 5956
rect 14676 5924 14680 5956
rect 14640 5876 14680 5924
rect 14640 5844 14644 5876
rect 14676 5844 14680 5876
rect 14640 5796 14680 5844
rect 14640 5764 14644 5796
rect 14676 5764 14680 5796
rect 14640 5716 14680 5764
rect 14640 5684 14644 5716
rect 14676 5684 14680 5716
rect 14640 5636 14680 5684
rect 14640 5604 14644 5636
rect 14676 5604 14680 5636
rect 14640 5556 14680 5604
rect 14640 5524 14644 5556
rect 14676 5524 14680 5556
rect 14640 5476 14680 5524
rect 14640 5444 14644 5476
rect 14676 5444 14680 5476
rect 14640 5396 14680 5444
rect 14640 5364 14644 5396
rect 14676 5364 14680 5396
rect 14640 5316 14680 5364
rect 14640 5284 14644 5316
rect 14676 5284 14680 5316
rect 14640 5236 14680 5284
rect 14640 5204 14644 5236
rect 14676 5204 14680 5236
rect 14640 5156 14680 5204
rect 14640 5124 14644 5156
rect 14676 5124 14680 5156
rect 14640 5076 14680 5124
rect 14640 5044 14644 5076
rect 14676 5044 14680 5076
rect 14640 4996 14680 5044
rect 14640 4964 14644 4996
rect 14676 4964 14680 4996
rect 14640 4916 14680 4964
rect 14640 4884 14644 4916
rect 14676 4884 14680 4916
rect 14640 4836 14680 4884
rect 14640 4804 14644 4836
rect 14676 4804 14680 4836
rect 14640 4676 14680 4804
rect 14640 4644 14644 4676
rect 14676 4644 14680 4676
rect 14640 4516 14680 4644
rect 14640 4484 14644 4516
rect 14676 4484 14680 4516
rect 14640 4436 14680 4484
rect 14640 4404 14644 4436
rect 14676 4404 14680 4436
rect 14640 4356 14680 4404
rect 14640 4324 14644 4356
rect 14676 4324 14680 4356
rect 14640 4276 14680 4324
rect 14640 4244 14644 4276
rect 14676 4244 14680 4276
rect 14640 4196 14680 4244
rect 14640 4164 14644 4196
rect 14676 4164 14680 4196
rect 14640 4116 14680 4164
rect 14640 4084 14644 4116
rect 14676 4084 14680 4116
rect 14640 4036 14680 4084
rect 14640 4004 14644 4036
rect 14676 4004 14680 4036
rect 14640 3956 14680 4004
rect 14640 3924 14644 3956
rect 14676 3924 14680 3956
rect 14640 3876 14680 3924
rect 14640 3844 14644 3876
rect 14676 3844 14680 3876
rect 14640 3796 14680 3844
rect 14640 3764 14644 3796
rect 14676 3764 14680 3796
rect 14640 3716 14680 3764
rect 14640 3684 14644 3716
rect 14676 3684 14680 3716
rect 14640 3636 14680 3684
rect 14640 3604 14644 3636
rect 14676 3604 14680 3636
rect 14640 3556 14680 3604
rect 14640 3524 14644 3556
rect 14676 3524 14680 3556
rect 14640 3476 14680 3524
rect 14640 3444 14644 3476
rect 14676 3444 14680 3476
rect 14640 3396 14680 3444
rect 14640 3364 14644 3396
rect 14676 3364 14680 3396
rect 14640 3316 14680 3364
rect 14640 3284 14644 3316
rect 14676 3284 14680 3316
rect 14640 3236 14680 3284
rect 14640 3204 14644 3236
rect 14676 3204 14680 3236
rect 14640 3156 14680 3204
rect 14640 3124 14644 3156
rect 14676 3124 14680 3156
rect 14640 3076 14680 3124
rect 14640 3044 14644 3076
rect 14676 3044 14680 3076
rect 14640 2996 14680 3044
rect 14640 2964 14644 2996
rect 14676 2964 14680 2996
rect 14640 2916 14680 2964
rect 14640 2884 14644 2916
rect 14676 2884 14680 2916
rect 14640 2836 14680 2884
rect 14640 2804 14644 2836
rect 14676 2804 14680 2836
rect 14640 2756 14680 2804
rect 14640 2724 14644 2756
rect 14676 2724 14680 2756
rect 14640 2676 14680 2724
rect 14640 2644 14644 2676
rect 14676 2644 14680 2676
rect 14640 2596 14680 2644
rect 14640 2564 14644 2596
rect 14676 2564 14680 2596
rect 14640 2516 14680 2564
rect 14640 2484 14644 2516
rect 14676 2484 14680 2516
rect 14640 2436 14680 2484
rect 14640 2404 14644 2436
rect 14676 2404 14680 2436
rect 14640 2356 14680 2404
rect 14640 2324 14644 2356
rect 14676 2324 14680 2356
rect 14640 2276 14680 2324
rect 14640 2244 14644 2276
rect 14676 2244 14680 2276
rect 14640 2196 14680 2244
rect 14640 2164 14644 2196
rect 14676 2164 14680 2196
rect 14640 2116 14680 2164
rect 14640 2084 14644 2116
rect 14676 2084 14680 2116
rect 14640 1956 14680 2084
rect 14640 1924 14644 1956
rect 14676 1924 14680 1956
rect 14640 1796 14680 1924
rect 14640 1764 14644 1796
rect 14676 1764 14680 1796
rect 14640 1716 14680 1764
rect 14640 1684 14644 1716
rect 14676 1684 14680 1716
rect 14640 1636 14680 1684
rect 14640 1604 14644 1636
rect 14676 1604 14680 1636
rect 14640 1556 14680 1604
rect 14640 1524 14644 1556
rect 14676 1524 14680 1556
rect 14640 1476 14680 1524
rect 14640 1444 14644 1476
rect 14676 1444 14680 1476
rect 14640 1396 14680 1444
rect 14640 1364 14644 1396
rect 14676 1364 14680 1396
rect 14640 1316 14680 1364
rect 14640 1284 14644 1316
rect 14676 1284 14680 1316
rect 14640 1236 14680 1284
rect 14640 1204 14644 1236
rect 14676 1204 14680 1236
rect 14640 1156 14680 1204
rect 14640 1124 14644 1156
rect 14676 1124 14680 1156
rect 14640 1076 14680 1124
rect 14640 1044 14644 1076
rect 14676 1044 14680 1076
rect 14640 996 14680 1044
rect 14640 964 14644 996
rect 14676 964 14680 996
rect 14640 916 14680 964
rect 14640 884 14644 916
rect 14676 884 14680 916
rect 14640 836 14680 884
rect 14640 804 14644 836
rect 14676 804 14680 836
rect 14640 756 14680 804
rect 14640 724 14644 756
rect 14676 724 14680 756
rect 14640 676 14680 724
rect 14640 644 14644 676
rect 14676 644 14680 676
rect 14640 596 14680 644
rect 14640 564 14644 596
rect 14676 564 14680 596
rect 14640 516 14680 564
rect 14640 484 14644 516
rect 14676 484 14680 516
rect 14480 244 14484 436
rect 14516 244 14520 436
rect 14480 240 14520 244
rect 14640 436 14680 484
rect 14720 14436 14760 15960
rect 14720 14404 14724 14436
rect 14756 14404 14760 14436
rect 14720 11876 14760 14404
rect 14720 11844 14724 11876
rect 14756 11844 14760 11876
rect 14720 4596 14760 11844
rect 14720 4564 14724 4596
rect 14756 4564 14760 4596
rect 14720 2036 14760 4564
rect 14720 2004 14724 2036
rect 14756 2004 14760 2036
rect 14720 480 14760 2004
rect 14800 15956 14840 15960
rect 14800 15924 14804 15956
rect 14836 15924 14840 15956
rect 14800 15876 14840 15924
rect 14800 15844 14804 15876
rect 14836 15844 14840 15876
rect 14800 15796 14840 15844
rect 14800 15764 14804 15796
rect 14836 15764 14840 15796
rect 14800 15716 14840 15764
rect 14800 15684 14804 15716
rect 14836 15684 14840 15716
rect 14800 15636 14840 15684
rect 14800 15604 14804 15636
rect 14836 15604 14840 15636
rect 14800 15556 14840 15604
rect 14800 15524 14804 15556
rect 14836 15524 14840 15556
rect 14800 15476 14840 15524
rect 14800 15444 14804 15476
rect 14836 15444 14840 15476
rect 14800 15396 14840 15444
rect 14800 15364 14804 15396
rect 14836 15364 14840 15396
rect 14800 15316 14840 15364
rect 14800 15284 14804 15316
rect 14836 15284 14840 15316
rect 14800 15236 14840 15284
rect 14800 15204 14804 15236
rect 14836 15204 14840 15236
rect 14800 15156 14840 15204
rect 14800 15124 14804 15156
rect 14836 15124 14840 15156
rect 14800 15076 14840 15124
rect 14800 15044 14804 15076
rect 14836 15044 14840 15076
rect 14800 14996 14840 15044
rect 14800 14964 14804 14996
rect 14836 14964 14840 14996
rect 14800 14916 14840 14964
rect 14800 14884 14804 14916
rect 14836 14884 14840 14916
rect 14800 14836 14840 14884
rect 14800 14804 14804 14836
rect 14836 14804 14840 14836
rect 14800 14756 14840 14804
rect 14800 14724 14804 14756
rect 14836 14724 14840 14756
rect 14800 14676 14840 14724
rect 14800 14644 14804 14676
rect 14836 14644 14840 14676
rect 14800 14516 14840 14644
rect 14800 14484 14804 14516
rect 14836 14484 14840 14516
rect 14800 14436 14840 14484
rect 14800 14404 14804 14436
rect 14836 14404 14840 14436
rect 14800 14356 14840 14404
rect 14800 14324 14804 14356
rect 14836 14324 14840 14356
rect 14800 14276 14840 14324
rect 14800 14244 14804 14276
rect 14836 14244 14840 14276
rect 14800 14196 14840 14244
rect 14800 14164 14804 14196
rect 14836 14164 14840 14196
rect 14800 14116 14840 14164
rect 14800 14084 14804 14116
rect 14836 14084 14840 14116
rect 14800 14036 14840 14084
rect 14800 14004 14804 14036
rect 14836 14004 14840 14036
rect 14800 13956 14840 14004
rect 14800 13924 14804 13956
rect 14836 13924 14840 13956
rect 14800 13876 14840 13924
rect 14800 13844 14804 13876
rect 14836 13844 14840 13876
rect 14800 13796 14840 13844
rect 14800 13764 14804 13796
rect 14836 13764 14840 13796
rect 14800 13716 14840 13764
rect 14800 13684 14804 13716
rect 14836 13684 14840 13716
rect 14800 13636 14840 13684
rect 14800 13604 14804 13636
rect 14836 13604 14840 13636
rect 14800 13556 14840 13604
rect 14800 13524 14804 13556
rect 14836 13524 14840 13556
rect 14800 13476 14840 13524
rect 14800 13444 14804 13476
rect 14836 13444 14840 13476
rect 14800 13396 14840 13444
rect 14800 13364 14804 13396
rect 14836 13364 14840 13396
rect 14800 13316 14840 13364
rect 14800 13284 14804 13316
rect 14836 13284 14840 13316
rect 14800 13236 14840 13284
rect 14800 13204 14804 13236
rect 14836 13204 14840 13236
rect 14800 13156 14840 13204
rect 14800 13124 14804 13156
rect 14836 13124 14840 13156
rect 14800 13076 14840 13124
rect 14800 13044 14804 13076
rect 14836 13044 14840 13076
rect 14800 12996 14840 13044
rect 14800 12964 14804 12996
rect 14836 12964 14840 12996
rect 14800 12916 14840 12964
rect 14800 12884 14804 12916
rect 14836 12884 14840 12916
rect 14800 12836 14840 12884
rect 14800 12804 14804 12836
rect 14836 12804 14840 12836
rect 14800 12756 14840 12804
rect 14800 12724 14804 12756
rect 14836 12724 14840 12756
rect 14800 12676 14840 12724
rect 14800 12644 14804 12676
rect 14836 12644 14840 12676
rect 14800 12596 14840 12644
rect 14800 12564 14804 12596
rect 14836 12564 14840 12596
rect 14800 12516 14840 12564
rect 14800 12484 14804 12516
rect 14836 12484 14840 12516
rect 14800 12436 14840 12484
rect 14800 12404 14804 12436
rect 14836 12404 14840 12436
rect 14800 12356 14840 12404
rect 14800 12324 14804 12356
rect 14836 12324 14840 12356
rect 14800 12276 14840 12324
rect 14800 12244 14804 12276
rect 14836 12244 14840 12276
rect 14800 12196 14840 12244
rect 14800 12164 14804 12196
rect 14836 12164 14840 12196
rect 14800 12116 14840 12164
rect 14800 12084 14804 12116
rect 14836 12084 14840 12116
rect 14800 12036 14840 12084
rect 14800 12004 14804 12036
rect 14836 12004 14840 12036
rect 14800 11956 14840 12004
rect 14800 11924 14804 11956
rect 14836 11924 14840 11956
rect 14800 11876 14840 11924
rect 14800 11844 14804 11876
rect 14836 11844 14840 11876
rect 14800 11796 14840 11844
rect 14800 11764 14804 11796
rect 14836 11764 14840 11796
rect 14800 11636 14840 11764
rect 14800 11604 14804 11636
rect 14836 11604 14840 11636
rect 14800 11556 14840 11604
rect 14800 11524 14804 11556
rect 14836 11524 14840 11556
rect 14800 11476 14840 11524
rect 14800 11444 14804 11476
rect 14836 11444 14840 11476
rect 14800 11396 14840 11444
rect 14800 11364 14804 11396
rect 14836 11364 14840 11396
rect 14800 11316 14840 11364
rect 14800 11284 14804 11316
rect 14836 11284 14840 11316
rect 14800 11236 14840 11284
rect 14800 11204 14804 11236
rect 14836 11204 14840 11236
rect 14800 11156 14840 11204
rect 14800 11124 14804 11156
rect 14836 11124 14840 11156
rect 14800 11076 14840 11124
rect 14800 11044 14804 11076
rect 14836 11044 14840 11076
rect 14800 10996 14840 11044
rect 14800 10964 14804 10996
rect 14836 10964 14840 10996
rect 14800 10916 14840 10964
rect 14800 10884 14804 10916
rect 14836 10884 14840 10916
rect 14800 10836 14840 10884
rect 14800 10804 14804 10836
rect 14836 10804 14840 10836
rect 14800 10756 14840 10804
rect 14800 10724 14804 10756
rect 14836 10724 14840 10756
rect 14800 10676 14840 10724
rect 14800 10644 14804 10676
rect 14836 10644 14840 10676
rect 14800 10596 14840 10644
rect 14800 10564 14804 10596
rect 14836 10564 14840 10596
rect 14800 10516 14840 10564
rect 14800 10484 14804 10516
rect 14836 10484 14840 10516
rect 14800 10436 14840 10484
rect 14800 10404 14804 10436
rect 14836 10404 14840 10436
rect 14800 10356 14840 10404
rect 14800 10324 14804 10356
rect 14836 10324 14840 10356
rect 14800 10276 14840 10324
rect 14800 10244 14804 10276
rect 14836 10244 14840 10276
rect 14800 10196 14840 10244
rect 14800 10164 14804 10196
rect 14836 10164 14840 10196
rect 14800 10116 14840 10164
rect 14800 10084 14804 10116
rect 14836 10084 14840 10116
rect 14800 10036 14840 10084
rect 14800 10004 14804 10036
rect 14836 10004 14840 10036
rect 14800 9956 14840 10004
rect 14800 9924 14804 9956
rect 14836 9924 14840 9956
rect 14800 9876 14840 9924
rect 14800 9844 14804 9876
rect 14836 9844 14840 9876
rect 14800 9796 14840 9844
rect 14800 9764 14804 9796
rect 14836 9764 14840 9796
rect 14800 9716 14840 9764
rect 14800 9684 14804 9716
rect 14836 9684 14840 9716
rect 14800 9636 14840 9684
rect 14800 9604 14804 9636
rect 14836 9604 14840 9636
rect 14800 9556 14840 9604
rect 14800 9524 14804 9556
rect 14836 9524 14840 9556
rect 14800 9476 14840 9524
rect 14800 9444 14804 9476
rect 14836 9444 14840 9476
rect 14800 9396 14840 9444
rect 14800 9364 14804 9396
rect 14836 9364 14840 9396
rect 14800 9316 14840 9364
rect 14800 9284 14804 9316
rect 14836 9284 14840 9316
rect 14800 9236 14840 9284
rect 14800 9204 14804 9236
rect 14836 9204 14840 9236
rect 14800 9156 14840 9204
rect 14800 9124 14804 9156
rect 14836 9124 14840 9156
rect 14800 9076 14840 9124
rect 14800 9044 14804 9076
rect 14836 9044 14840 9076
rect 14800 8996 14840 9044
rect 14800 8964 14804 8996
rect 14836 8964 14840 8996
rect 14800 8916 14840 8964
rect 14800 8884 14804 8916
rect 14836 8884 14840 8916
rect 14800 8836 14840 8884
rect 14800 8804 14804 8836
rect 14836 8804 14840 8836
rect 14800 8756 14840 8804
rect 14800 8724 14804 8756
rect 14836 8724 14840 8756
rect 14800 8676 14840 8724
rect 14800 8644 14804 8676
rect 14836 8644 14840 8676
rect 14800 8596 14840 8644
rect 14800 8564 14804 8596
rect 14836 8564 14840 8596
rect 14800 8516 14840 8564
rect 14800 8484 14804 8516
rect 14836 8484 14840 8516
rect 14800 8436 14840 8484
rect 14800 8404 14804 8436
rect 14836 8404 14840 8436
rect 14800 8356 14840 8404
rect 14800 8324 14804 8356
rect 14836 8324 14840 8356
rect 14800 8276 14840 8324
rect 14800 8244 14804 8276
rect 14836 8244 14840 8276
rect 14800 8196 14840 8244
rect 14800 8164 14804 8196
rect 14836 8164 14840 8196
rect 14800 8116 14840 8164
rect 14800 8084 14804 8116
rect 14836 8084 14840 8116
rect 14800 8036 14840 8084
rect 14800 8004 14804 8036
rect 14836 8004 14840 8036
rect 14800 7956 14840 8004
rect 14800 7924 14804 7956
rect 14836 7924 14840 7956
rect 14800 7876 14840 7924
rect 14800 7844 14804 7876
rect 14836 7844 14840 7876
rect 14800 7796 14840 7844
rect 14800 7764 14804 7796
rect 14836 7764 14840 7796
rect 14800 7716 14840 7764
rect 14800 7684 14804 7716
rect 14836 7684 14840 7716
rect 14800 7636 14840 7684
rect 14800 7604 14804 7636
rect 14836 7604 14840 7636
rect 14800 7556 14840 7604
rect 14800 7524 14804 7556
rect 14836 7524 14840 7556
rect 14800 7476 14840 7524
rect 14800 7444 14804 7476
rect 14836 7444 14840 7476
rect 14800 7396 14840 7444
rect 14800 7364 14804 7396
rect 14836 7364 14840 7396
rect 14800 7316 14840 7364
rect 14800 7284 14804 7316
rect 14836 7284 14840 7316
rect 14800 7236 14840 7284
rect 14800 7204 14804 7236
rect 14836 7204 14840 7236
rect 14800 7156 14840 7204
rect 14800 7124 14804 7156
rect 14836 7124 14840 7156
rect 14800 7076 14840 7124
rect 14800 7044 14804 7076
rect 14836 7044 14840 7076
rect 14800 6996 14840 7044
rect 14800 6964 14804 6996
rect 14836 6964 14840 6996
rect 14800 6916 14840 6964
rect 14800 6884 14804 6916
rect 14836 6884 14840 6916
rect 14800 6836 14840 6884
rect 14800 6804 14804 6836
rect 14836 6804 14840 6836
rect 14800 6756 14840 6804
rect 14800 6724 14804 6756
rect 14836 6724 14840 6756
rect 14800 6676 14840 6724
rect 14800 6644 14804 6676
rect 14836 6644 14840 6676
rect 14800 6596 14840 6644
rect 14800 6564 14804 6596
rect 14836 6564 14840 6596
rect 14800 6516 14840 6564
rect 14800 6484 14804 6516
rect 14836 6484 14840 6516
rect 14800 6436 14840 6484
rect 14800 6404 14804 6436
rect 14836 6404 14840 6436
rect 14800 6356 14840 6404
rect 14800 6324 14804 6356
rect 14836 6324 14840 6356
rect 14800 6276 14840 6324
rect 14800 6244 14804 6276
rect 14836 6244 14840 6276
rect 14800 6196 14840 6244
rect 14800 6164 14804 6196
rect 14836 6164 14840 6196
rect 14800 6116 14840 6164
rect 14800 6084 14804 6116
rect 14836 6084 14840 6116
rect 14800 6036 14840 6084
rect 14800 6004 14804 6036
rect 14836 6004 14840 6036
rect 14800 5956 14840 6004
rect 14800 5924 14804 5956
rect 14836 5924 14840 5956
rect 14800 5876 14840 5924
rect 14800 5844 14804 5876
rect 14836 5844 14840 5876
rect 14800 5796 14840 5844
rect 14800 5764 14804 5796
rect 14836 5764 14840 5796
rect 14800 5716 14840 5764
rect 14800 5684 14804 5716
rect 14836 5684 14840 5716
rect 14800 5636 14840 5684
rect 14800 5604 14804 5636
rect 14836 5604 14840 5636
rect 14800 5556 14840 5604
rect 14800 5524 14804 5556
rect 14836 5524 14840 5556
rect 14800 5476 14840 5524
rect 14800 5444 14804 5476
rect 14836 5444 14840 5476
rect 14800 5396 14840 5444
rect 14800 5364 14804 5396
rect 14836 5364 14840 5396
rect 14800 5316 14840 5364
rect 14800 5284 14804 5316
rect 14836 5284 14840 5316
rect 14800 5236 14840 5284
rect 14800 5204 14804 5236
rect 14836 5204 14840 5236
rect 14800 5156 14840 5204
rect 14800 5124 14804 5156
rect 14836 5124 14840 5156
rect 14800 5076 14840 5124
rect 14800 5044 14804 5076
rect 14836 5044 14840 5076
rect 14800 4996 14840 5044
rect 14800 4964 14804 4996
rect 14836 4964 14840 4996
rect 14800 4916 14840 4964
rect 14800 4884 14804 4916
rect 14836 4884 14840 4916
rect 14800 4836 14840 4884
rect 14800 4804 14804 4836
rect 14836 4804 14840 4836
rect 14800 4676 14840 4804
rect 14800 4644 14804 4676
rect 14836 4644 14840 4676
rect 14800 4596 14840 4644
rect 14800 4564 14804 4596
rect 14836 4564 14840 4596
rect 14800 4516 14840 4564
rect 14800 4484 14804 4516
rect 14836 4484 14840 4516
rect 14800 4436 14840 4484
rect 14800 4404 14804 4436
rect 14836 4404 14840 4436
rect 14800 4356 14840 4404
rect 14800 4324 14804 4356
rect 14836 4324 14840 4356
rect 14800 4276 14840 4324
rect 14800 4244 14804 4276
rect 14836 4244 14840 4276
rect 14800 4196 14840 4244
rect 14800 4164 14804 4196
rect 14836 4164 14840 4196
rect 14800 4116 14840 4164
rect 14800 4084 14804 4116
rect 14836 4084 14840 4116
rect 14800 4036 14840 4084
rect 14800 4004 14804 4036
rect 14836 4004 14840 4036
rect 14800 3956 14840 4004
rect 14800 3924 14804 3956
rect 14836 3924 14840 3956
rect 14800 3876 14840 3924
rect 14800 3844 14804 3876
rect 14836 3844 14840 3876
rect 14800 3796 14840 3844
rect 14800 3764 14804 3796
rect 14836 3764 14840 3796
rect 14800 3716 14840 3764
rect 14800 3684 14804 3716
rect 14836 3684 14840 3716
rect 14800 3636 14840 3684
rect 14800 3604 14804 3636
rect 14836 3604 14840 3636
rect 14800 3556 14840 3604
rect 14800 3524 14804 3556
rect 14836 3524 14840 3556
rect 14800 3476 14840 3524
rect 14800 3444 14804 3476
rect 14836 3444 14840 3476
rect 14800 3396 14840 3444
rect 14800 3364 14804 3396
rect 14836 3364 14840 3396
rect 14800 3316 14840 3364
rect 14800 3284 14804 3316
rect 14836 3284 14840 3316
rect 14800 3236 14840 3284
rect 14800 3204 14804 3236
rect 14836 3204 14840 3236
rect 14800 3156 14840 3204
rect 14800 3124 14804 3156
rect 14836 3124 14840 3156
rect 14800 3076 14840 3124
rect 14800 3044 14804 3076
rect 14836 3044 14840 3076
rect 14800 2996 14840 3044
rect 14800 2964 14804 2996
rect 14836 2964 14840 2996
rect 14800 2916 14840 2964
rect 14800 2884 14804 2916
rect 14836 2884 14840 2916
rect 14800 2836 14840 2884
rect 14800 2804 14804 2836
rect 14836 2804 14840 2836
rect 14800 2756 14840 2804
rect 14800 2724 14804 2756
rect 14836 2724 14840 2756
rect 14800 2676 14840 2724
rect 14800 2644 14804 2676
rect 14836 2644 14840 2676
rect 14800 2596 14840 2644
rect 14800 2564 14804 2596
rect 14836 2564 14840 2596
rect 14800 2516 14840 2564
rect 14800 2484 14804 2516
rect 14836 2484 14840 2516
rect 14800 2436 14840 2484
rect 14800 2404 14804 2436
rect 14836 2404 14840 2436
rect 14800 2356 14840 2404
rect 14800 2324 14804 2356
rect 14836 2324 14840 2356
rect 14800 2276 14840 2324
rect 14800 2244 14804 2276
rect 14836 2244 14840 2276
rect 14800 2196 14840 2244
rect 14800 2164 14804 2196
rect 14836 2164 14840 2196
rect 14800 2116 14840 2164
rect 14800 2084 14804 2116
rect 14836 2084 14840 2116
rect 14800 2036 14840 2084
rect 14800 2004 14804 2036
rect 14836 2004 14840 2036
rect 14800 1956 14840 2004
rect 14800 1924 14804 1956
rect 14836 1924 14840 1956
rect 14800 1796 14840 1924
rect 14800 1764 14804 1796
rect 14836 1764 14840 1796
rect 14800 1716 14840 1764
rect 14800 1684 14804 1716
rect 14836 1684 14840 1716
rect 14800 1636 14840 1684
rect 14800 1604 14804 1636
rect 14836 1604 14840 1636
rect 14800 1556 14840 1604
rect 14800 1524 14804 1556
rect 14836 1524 14840 1556
rect 14800 1476 14840 1524
rect 14800 1444 14804 1476
rect 14836 1444 14840 1476
rect 14800 1396 14840 1444
rect 14800 1364 14804 1396
rect 14836 1364 14840 1396
rect 14800 1316 14840 1364
rect 14800 1284 14804 1316
rect 14836 1284 14840 1316
rect 14800 1236 14840 1284
rect 14800 1204 14804 1236
rect 14836 1204 14840 1236
rect 14800 1156 14840 1204
rect 14800 1124 14804 1156
rect 14836 1124 14840 1156
rect 14800 1076 14840 1124
rect 14800 1044 14804 1076
rect 14836 1044 14840 1076
rect 14800 996 14840 1044
rect 14800 964 14804 996
rect 14836 964 14840 996
rect 14800 916 14840 964
rect 14800 884 14804 916
rect 14836 884 14840 916
rect 14800 836 14840 884
rect 14800 804 14804 836
rect 14836 804 14840 836
rect 14800 756 14840 804
rect 14800 724 14804 756
rect 14836 724 14840 756
rect 14800 676 14840 724
rect 14800 644 14804 676
rect 14836 644 14840 676
rect 14800 596 14840 644
rect 14800 564 14804 596
rect 14836 564 14840 596
rect 14800 516 14840 564
rect 14800 484 14804 516
rect 14836 484 14840 516
rect 14640 244 14644 436
rect 14676 244 14680 436
rect 14640 240 14680 244
rect 14800 436 14840 484
rect 14880 14596 14920 15960
rect 14880 14564 14884 14596
rect 14916 14564 14920 14596
rect 14880 11716 14920 14564
rect 14880 11684 14884 11716
rect 14916 11684 14920 11716
rect 14880 4756 14920 11684
rect 14880 4724 14884 4756
rect 14916 4724 14920 4756
rect 14880 1876 14920 4724
rect 14880 1844 14884 1876
rect 14916 1844 14920 1876
rect 14880 480 14920 1844
rect 14960 15956 15000 15960
rect 14960 15924 14964 15956
rect 14996 15924 15000 15956
rect 14960 15876 15000 15924
rect 14960 15844 14964 15876
rect 14996 15844 15000 15876
rect 14960 15796 15000 15844
rect 14960 15764 14964 15796
rect 14996 15764 15000 15796
rect 14960 15716 15000 15764
rect 14960 15684 14964 15716
rect 14996 15684 15000 15716
rect 14960 15636 15000 15684
rect 14960 15604 14964 15636
rect 14996 15604 15000 15636
rect 14960 15556 15000 15604
rect 14960 15524 14964 15556
rect 14996 15524 15000 15556
rect 14960 15476 15000 15524
rect 14960 15444 14964 15476
rect 14996 15444 15000 15476
rect 14960 15396 15000 15444
rect 14960 15364 14964 15396
rect 14996 15364 15000 15396
rect 14960 15316 15000 15364
rect 14960 15284 14964 15316
rect 14996 15284 15000 15316
rect 14960 15236 15000 15284
rect 14960 15204 14964 15236
rect 14996 15204 15000 15236
rect 14960 15156 15000 15204
rect 14960 15124 14964 15156
rect 14996 15124 15000 15156
rect 14960 15076 15000 15124
rect 14960 15044 14964 15076
rect 14996 15044 15000 15076
rect 14960 14996 15000 15044
rect 14960 14964 14964 14996
rect 14996 14964 15000 14996
rect 14960 14916 15000 14964
rect 14960 14884 14964 14916
rect 14996 14884 15000 14916
rect 14960 14836 15000 14884
rect 14960 14804 14964 14836
rect 14996 14804 15000 14836
rect 14960 14756 15000 14804
rect 14960 14724 14964 14756
rect 14996 14724 15000 14756
rect 14960 14676 15000 14724
rect 14960 14644 14964 14676
rect 14996 14644 15000 14676
rect 14960 14516 15000 14644
rect 14960 14484 14964 14516
rect 14996 14484 15000 14516
rect 14960 14436 15000 14484
rect 14960 14404 14964 14436
rect 14996 14404 15000 14436
rect 14960 14356 15000 14404
rect 14960 14324 14964 14356
rect 14996 14324 15000 14356
rect 14960 14276 15000 14324
rect 14960 14244 14964 14276
rect 14996 14244 15000 14276
rect 14960 14196 15000 14244
rect 14960 14164 14964 14196
rect 14996 14164 15000 14196
rect 14960 14116 15000 14164
rect 14960 14084 14964 14116
rect 14996 14084 15000 14116
rect 14960 14036 15000 14084
rect 14960 14004 14964 14036
rect 14996 14004 15000 14036
rect 14960 13956 15000 14004
rect 14960 13924 14964 13956
rect 14996 13924 15000 13956
rect 14960 13876 15000 13924
rect 14960 13844 14964 13876
rect 14996 13844 15000 13876
rect 14960 13796 15000 13844
rect 14960 13764 14964 13796
rect 14996 13764 15000 13796
rect 14960 13716 15000 13764
rect 14960 13684 14964 13716
rect 14996 13684 15000 13716
rect 14960 13636 15000 13684
rect 14960 13604 14964 13636
rect 14996 13604 15000 13636
rect 14960 13556 15000 13604
rect 14960 13524 14964 13556
rect 14996 13524 15000 13556
rect 14960 13476 15000 13524
rect 14960 13444 14964 13476
rect 14996 13444 15000 13476
rect 14960 13396 15000 13444
rect 14960 13364 14964 13396
rect 14996 13364 15000 13396
rect 14960 13316 15000 13364
rect 14960 13284 14964 13316
rect 14996 13284 15000 13316
rect 14960 13236 15000 13284
rect 14960 13204 14964 13236
rect 14996 13204 15000 13236
rect 14960 13156 15000 13204
rect 14960 13124 14964 13156
rect 14996 13124 15000 13156
rect 14960 13076 15000 13124
rect 14960 13044 14964 13076
rect 14996 13044 15000 13076
rect 14960 12996 15000 13044
rect 14960 12964 14964 12996
rect 14996 12964 15000 12996
rect 14960 12916 15000 12964
rect 14960 12884 14964 12916
rect 14996 12884 15000 12916
rect 14960 12836 15000 12884
rect 14960 12804 14964 12836
rect 14996 12804 15000 12836
rect 14960 12756 15000 12804
rect 14960 12724 14964 12756
rect 14996 12724 15000 12756
rect 14960 12676 15000 12724
rect 14960 12644 14964 12676
rect 14996 12644 15000 12676
rect 14960 12596 15000 12644
rect 14960 12564 14964 12596
rect 14996 12564 15000 12596
rect 14960 12516 15000 12564
rect 14960 12484 14964 12516
rect 14996 12484 15000 12516
rect 14960 12436 15000 12484
rect 14960 12404 14964 12436
rect 14996 12404 15000 12436
rect 14960 12356 15000 12404
rect 14960 12324 14964 12356
rect 14996 12324 15000 12356
rect 14960 12276 15000 12324
rect 14960 12244 14964 12276
rect 14996 12244 15000 12276
rect 14960 12196 15000 12244
rect 14960 12164 14964 12196
rect 14996 12164 15000 12196
rect 14960 12116 15000 12164
rect 14960 12084 14964 12116
rect 14996 12084 15000 12116
rect 14960 12036 15000 12084
rect 14960 12004 14964 12036
rect 14996 12004 15000 12036
rect 14960 11956 15000 12004
rect 14960 11924 14964 11956
rect 14996 11924 15000 11956
rect 14960 11876 15000 11924
rect 14960 11844 14964 11876
rect 14996 11844 15000 11876
rect 14960 11796 15000 11844
rect 14960 11764 14964 11796
rect 14996 11764 15000 11796
rect 14960 11636 15000 11764
rect 14960 11604 14964 11636
rect 14996 11604 15000 11636
rect 14960 11556 15000 11604
rect 14960 11524 14964 11556
rect 14996 11524 15000 11556
rect 14960 11476 15000 11524
rect 14960 11444 14964 11476
rect 14996 11444 15000 11476
rect 14960 11396 15000 11444
rect 14960 11364 14964 11396
rect 14996 11364 15000 11396
rect 14960 11316 15000 11364
rect 14960 11284 14964 11316
rect 14996 11284 15000 11316
rect 14960 11236 15000 11284
rect 14960 11204 14964 11236
rect 14996 11204 15000 11236
rect 14960 11156 15000 11204
rect 14960 11124 14964 11156
rect 14996 11124 15000 11156
rect 14960 11076 15000 11124
rect 14960 11044 14964 11076
rect 14996 11044 15000 11076
rect 14960 10996 15000 11044
rect 14960 10964 14964 10996
rect 14996 10964 15000 10996
rect 14960 10916 15000 10964
rect 14960 10884 14964 10916
rect 14996 10884 15000 10916
rect 14960 10836 15000 10884
rect 14960 10804 14964 10836
rect 14996 10804 15000 10836
rect 14960 10756 15000 10804
rect 14960 10724 14964 10756
rect 14996 10724 15000 10756
rect 14960 10676 15000 10724
rect 14960 10644 14964 10676
rect 14996 10644 15000 10676
rect 14960 10596 15000 10644
rect 14960 10564 14964 10596
rect 14996 10564 15000 10596
rect 14960 10516 15000 10564
rect 14960 10484 14964 10516
rect 14996 10484 15000 10516
rect 14960 10436 15000 10484
rect 14960 10404 14964 10436
rect 14996 10404 15000 10436
rect 14960 10356 15000 10404
rect 14960 10324 14964 10356
rect 14996 10324 15000 10356
rect 14960 10276 15000 10324
rect 14960 10244 14964 10276
rect 14996 10244 15000 10276
rect 14960 10196 15000 10244
rect 14960 10164 14964 10196
rect 14996 10164 15000 10196
rect 14960 10116 15000 10164
rect 14960 10084 14964 10116
rect 14996 10084 15000 10116
rect 14960 10036 15000 10084
rect 14960 10004 14964 10036
rect 14996 10004 15000 10036
rect 14960 9956 15000 10004
rect 14960 9924 14964 9956
rect 14996 9924 15000 9956
rect 14960 9876 15000 9924
rect 14960 9844 14964 9876
rect 14996 9844 15000 9876
rect 14960 9796 15000 9844
rect 14960 9764 14964 9796
rect 14996 9764 15000 9796
rect 14960 9716 15000 9764
rect 14960 9684 14964 9716
rect 14996 9684 15000 9716
rect 14960 9636 15000 9684
rect 14960 9604 14964 9636
rect 14996 9604 15000 9636
rect 14960 9556 15000 9604
rect 14960 9524 14964 9556
rect 14996 9524 15000 9556
rect 14960 9476 15000 9524
rect 14960 9444 14964 9476
rect 14996 9444 15000 9476
rect 14960 9396 15000 9444
rect 14960 9364 14964 9396
rect 14996 9364 15000 9396
rect 14960 9316 15000 9364
rect 14960 9284 14964 9316
rect 14996 9284 15000 9316
rect 14960 9236 15000 9284
rect 14960 9204 14964 9236
rect 14996 9204 15000 9236
rect 14960 9156 15000 9204
rect 14960 9124 14964 9156
rect 14996 9124 15000 9156
rect 14960 9076 15000 9124
rect 14960 9044 14964 9076
rect 14996 9044 15000 9076
rect 14960 8996 15000 9044
rect 14960 8964 14964 8996
rect 14996 8964 15000 8996
rect 14960 8916 15000 8964
rect 14960 8884 14964 8916
rect 14996 8884 15000 8916
rect 14960 8836 15000 8884
rect 14960 8804 14964 8836
rect 14996 8804 15000 8836
rect 14960 8756 15000 8804
rect 14960 8724 14964 8756
rect 14996 8724 15000 8756
rect 14960 8676 15000 8724
rect 14960 8644 14964 8676
rect 14996 8644 15000 8676
rect 14960 8596 15000 8644
rect 14960 8564 14964 8596
rect 14996 8564 15000 8596
rect 14960 8516 15000 8564
rect 14960 8484 14964 8516
rect 14996 8484 15000 8516
rect 14960 8436 15000 8484
rect 14960 8404 14964 8436
rect 14996 8404 15000 8436
rect 14960 8356 15000 8404
rect 14960 8324 14964 8356
rect 14996 8324 15000 8356
rect 14960 8276 15000 8324
rect 14960 8244 14964 8276
rect 14996 8244 15000 8276
rect 14960 8196 15000 8244
rect 14960 8164 14964 8196
rect 14996 8164 15000 8196
rect 14960 8116 15000 8164
rect 14960 8084 14964 8116
rect 14996 8084 15000 8116
rect 14960 8036 15000 8084
rect 14960 8004 14964 8036
rect 14996 8004 15000 8036
rect 14960 7956 15000 8004
rect 14960 7924 14964 7956
rect 14996 7924 15000 7956
rect 14960 7876 15000 7924
rect 14960 7844 14964 7876
rect 14996 7844 15000 7876
rect 14960 7796 15000 7844
rect 14960 7764 14964 7796
rect 14996 7764 15000 7796
rect 14960 7716 15000 7764
rect 14960 7684 14964 7716
rect 14996 7684 15000 7716
rect 14960 7636 15000 7684
rect 14960 7604 14964 7636
rect 14996 7604 15000 7636
rect 14960 7556 15000 7604
rect 14960 7524 14964 7556
rect 14996 7524 15000 7556
rect 14960 7476 15000 7524
rect 14960 7444 14964 7476
rect 14996 7444 15000 7476
rect 14960 7396 15000 7444
rect 14960 7364 14964 7396
rect 14996 7364 15000 7396
rect 14960 7316 15000 7364
rect 14960 7284 14964 7316
rect 14996 7284 15000 7316
rect 14960 7236 15000 7284
rect 14960 7204 14964 7236
rect 14996 7204 15000 7236
rect 14960 7156 15000 7204
rect 14960 7124 14964 7156
rect 14996 7124 15000 7156
rect 14960 7076 15000 7124
rect 14960 7044 14964 7076
rect 14996 7044 15000 7076
rect 14960 6996 15000 7044
rect 14960 6964 14964 6996
rect 14996 6964 15000 6996
rect 14960 6916 15000 6964
rect 14960 6884 14964 6916
rect 14996 6884 15000 6916
rect 14960 6836 15000 6884
rect 14960 6804 14964 6836
rect 14996 6804 15000 6836
rect 14960 6756 15000 6804
rect 14960 6724 14964 6756
rect 14996 6724 15000 6756
rect 14960 6676 15000 6724
rect 14960 6644 14964 6676
rect 14996 6644 15000 6676
rect 14960 6596 15000 6644
rect 14960 6564 14964 6596
rect 14996 6564 15000 6596
rect 14960 6516 15000 6564
rect 14960 6484 14964 6516
rect 14996 6484 15000 6516
rect 14960 6436 15000 6484
rect 14960 6404 14964 6436
rect 14996 6404 15000 6436
rect 14960 6356 15000 6404
rect 14960 6324 14964 6356
rect 14996 6324 15000 6356
rect 14960 6276 15000 6324
rect 14960 6244 14964 6276
rect 14996 6244 15000 6276
rect 14960 6196 15000 6244
rect 14960 6164 14964 6196
rect 14996 6164 15000 6196
rect 14960 6116 15000 6164
rect 14960 6084 14964 6116
rect 14996 6084 15000 6116
rect 14960 6036 15000 6084
rect 14960 6004 14964 6036
rect 14996 6004 15000 6036
rect 14960 5956 15000 6004
rect 14960 5924 14964 5956
rect 14996 5924 15000 5956
rect 14960 5876 15000 5924
rect 14960 5844 14964 5876
rect 14996 5844 15000 5876
rect 14960 5796 15000 5844
rect 14960 5764 14964 5796
rect 14996 5764 15000 5796
rect 14960 5716 15000 5764
rect 14960 5684 14964 5716
rect 14996 5684 15000 5716
rect 14960 5636 15000 5684
rect 14960 5604 14964 5636
rect 14996 5604 15000 5636
rect 14960 5556 15000 5604
rect 14960 5524 14964 5556
rect 14996 5524 15000 5556
rect 14960 5476 15000 5524
rect 14960 5444 14964 5476
rect 14996 5444 15000 5476
rect 14960 5396 15000 5444
rect 14960 5364 14964 5396
rect 14996 5364 15000 5396
rect 14960 5316 15000 5364
rect 14960 5284 14964 5316
rect 14996 5284 15000 5316
rect 14960 5236 15000 5284
rect 14960 5204 14964 5236
rect 14996 5204 15000 5236
rect 14960 5156 15000 5204
rect 14960 5124 14964 5156
rect 14996 5124 15000 5156
rect 14960 5076 15000 5124
rect 14960 5044 14964 5076
rect 14996 5044 15000 5076
rect 14960 4996 15000 5044
rect 14960 4964 14964 4996
rect 14996 4964 15000 4996
rect 14960 4916 15000 4964
rect 14960 4884 14964 4916
rect 14996 4884 15000 4916
rect 14960 4836 15000 4884
rect 14960 4804 14964 4836
rect 14996 4804 15000 4836
rect 14960 4676 15000 4804
rect 14960 4644 14964 4676
rect 14996 4644 15000 4676
rect 14960 4596 15000 4644
rect 14960 4564 14964 4596
rect 14996 4564 15000 4596
rect 14960 4516 15000 4564
rect 14960 4484 14964 4516
rect 14996 4484 15000 4516
rect 14960 4436 15000 4484
rect 14960 4404 14964 4436
rect 14996 4404 15000 4436
rect 14960 4356 15000 4404
rect 14960 4324 14964 4356
rect 14996 4324 15000 4356
rect 14960 4276 15000 4324
rect 14960 4244 14964 4276
rect 14996 4244 15000 4276
rect 14960 4196 15000 4244
rect 14960 4164 14964 4196
rect 14996 4164 15000 4196
rect 14960 4116 15000 4164
rect 14960 4084 14964 4116
rect 14996 4084 15000 4116
rect 14960 4036 15000 4084
rect 14960 4004 14964 4036
rect 14996 4004 15000 4036
rect 14960 3956 15000 4004
rect 14960 3924 14964 3956
rect 14996 3924 15000 3956
rect 14960 3876 15000 3924
rect 14960 3844 14964 3876
rect 14996 3844 15000 3876
rect 14960 3796 15000 3844
rect 14960 3764 14964 3796
rect 14996 3764 15000 3796
rect 14960 3716 15000 3764
rect 14960 3684 14964 3716
rect 14996 3684 15000 3716
rect 14960 3636 15000 3684
rect 14960 3604 14964 3636
rect 14996 3604 15000 3636
rect 14960 3556 15000 3604
rect 14960 3524 14964 3556
rect 14996 3524 15000 3556
rect 14960 3476 15000 3524
rect 14960 3444 14964 3476
rect 14996 3444 15000 3476
rect 14960 3396 15000 3444
rect 14960 3364 14964 3396
rect 14996 3364 15000 3396
rect 14960 3316 15000 3364
rect 14960 3284 14964 3316
rect 14996 3284 15000 3316
rect 14960 3236 15000 3284
rect 14960 3204 14964 3236
rect 14996 3204 15000 3236
rect 14960 3156 15000 3204
rect 14960 3124 14964 3156
rect 14996 3124 15000 3156
rect 14960 3076 15000 3124
rect 14960 3044 14964 3076
rect 14996 3044 15000 3076
rect 14960 2996 15000 3044
rect 14960 2964 14964 2996
rect 14996 2964 15000 2996
rect 14960 2916 15000 2964
rect 14960 2884 14964 2916
rect 14996 2884 15000 2916
rect 14960 2836 15000 2884
rect 14960 2804 14964 2836
rect 14996 2804 15000 2836
rect 14960 2756 15000 2804
rect 14960 2724 14964 2756
rect 14996 2724 15000 2756
rect 14960 2676 15000 2724
rect 14960 2644 14964 2676
rect 14996 2644 15000 2676
rect 14960 2596 15000 2644
rect 14960 2564 14964 2596
rect 14996 2564 15000 2596
rect 14960 2516 15000 2564
rect 14960 2484 14964 2516
rect 14996 2484 15000 2516
rect 14960 2436 15000 2484
rect 14960 2404 14964 2436
rect 14996 2404 15000 2436
rect 14960 2356 15000 2404
rect 14960 2324 14964 2356
rect 14996 2324 15000 2356
rect 14960 2276 15000 2324
rect 14960 2244 14964 2276
rect 14996 2244 15000 2276
rect 14960 2196 15000 2244
rect 14960 2164 14964 2196
rect 14996 2164 15000 2196
rect 14960 2116 15000 2164
rect 14960 2084 14964 2116
rect 14996 2084 15000 2116
rect 14960 2036 15000 2084
rect 14960 2004 14964 2036
rect 14996 2004 15000 2036
rect 14960 1956 15000 2004
rect 14960 1924 14964 1956
rect 14996 1924 15000 1956
rect 14960 1796 15000 1924
rect 14960 1764 14964 1796
rect 14996 1764 15000 1796
rect 14960 1716 15000 1764
rect 14960 1684 14964 1716
rect 14996 1684 15000 1716
rect 14960 1636 15000 1684
rect 14960 1604 14964 1636
rect 14996 1604 15000 1636
rect 14960 1556 15000 1604
rect 14960 1524 14964 1556
rect 14996 1524 15000 1556
rect 14960 1476 15000 1524
rect 14960 1444 14964 1476
rect 14996 1444 15000 1476
rect 14960 1396 15000 1444
rect 14960 1364 14964 1396
rect 14996 1364 15000 1396
rect 14960 1316 15000 1364
rect 14960 1284 14964 1316
rect 14996 1284 15000 1316
rect 14960 1236 15000 1284
rect 14960 1204 14964 1236
rect 14996 1204 15000 1236
rect 14960 1156 15000 1204
rect 14960 1124 14964 1156
rect 14996 1124 15000 1156
rect 14960 1076 15000 1124
rect 14960 1044 14964 1076
rect 14996 1044 15000 1076
rect 14960 996 15000 1044
rect 14960 964 14964 996
rect 14996 964 15000 996
rect 14960 916 15000 964
rect 14960 884 14964 916
rect 14996 884 15000 916
rect 14960 836 15000 884
rect 14960 804 14964 836
rect 14996 804 15000 836
rect 14960 756 15000 804
rect 14960 724 14964 756
rect 14996 724 15000 756
rect 14960 676 15000 724
rect 14960 644 14964 676
rect 14996 644 15000 676
rect 14960 596 15000 644
rect 14960 564 14964 596
rect 14996 564 15000 596
rect 14960 516 15000 564
rect 14960 484 14964 516
rect 14996 484 15000 516
rect 14800 244 14804 436
rect 14836 244 14840 436
rect 14800 240 14840 244
rect 14960 436 15000 484
rect 14960 244 14964 436
rect 14996 244 15000 436
rect 14960 240 15000 244
rect 14400 4 14404 196
rect 14436 4 14440 196
rect 14400 0 14440 4
<< via3 >>
rect 4 15955 36 15956
rect 4 15925 5 15955
rect 5 15925 35 15955
rect 35 15925 36 15955
rect 4 15924 36 15925
rect 4 15875 36 15876
rect 4 15845 5 15875
rect 5 15845 35 15875
rect 35 15845 36 15875
rect 4 15844 36 15845
rect 4 15795 36 15796
rect 4 15765 5 15795
rect 5 15765 35 15795
rect 35 15765 36 15795
rect 4 15764 36 15765
rect 4 15715 36 15716
rect 4 15685 5 15715
rect 5 15685 35 15715
rect 35 15685 36 15715
rect 4 15684 36 15685
rect 4 15635 36 15636
rect 4 15605 5 15635
rect 5 15605 35 15635
rect 35 15605 36 15635
rect 4 15604 36 15605
rect 4 15555 36 15556
rect 4 15525 5 15555
rect 5 15525 35 15555
rect 35 15525 36 15555
rect 4 15524 36 15525
rect 4 15475 36 15476
rect 4 15445 5 15475
rect 5 15445 35 15475
rect 35 15445 36 15475
rect 4 15444 36 15445
rect 4 15395 36 15396
rect 4 15365 5 15395
rect 5 15365 35 15395
rect 35 15365 36 15395
rect 4 15364 36 15365
rect 4 15315 36 15316
rect 4 15285 5 15315
rect 5 15285 35 15315
rect 35 15285 36 15315
rect 4 15284 36 15285
rect 4 15235 36 15236
rect 4 15205 5 15235
rect 5 15205 35 15235
rect 35 15205 36 15235
rect 4 15204 36 15205
rect 4 15155 36 15156
rect 4 15125 5 15155
rect 5 15125 35 15155
rect 35 15125 36 15155
rect 4 15124 36 15125
rect 4 15075 36 15076
rect 4 15045 5 15075
rect 5 15045 35 15075
rect 35 15045 36 15075
rect 4 15044 36 15045
rect 4 14995 36 14996
rect 4 14965 5 14995
rect 5 14965 35 14995
rect 35 14965 36 14995
rect 4 14964 36 14965
rect 4 14915 36 14916
rect 4 14885 5 14915
rect 5 14885 35 14915
rect 35 14885 36 14915
rect 4 14884 36 14885
rect 4 14835 36 14836
rect 4 14805 5 14835
rect 5 14805 35 14835
rect 35 14805 36 14835
rect 4 14804 36 14805
rect 4 14755 36 14756
rect 4 14725 5 14755
rect 5 14725 35 14755
rect 35 14725 36 14755
rect 4 14724 36 14725
rect 4 14675 36 14676
rect 4 14645 5 14675
rect 5 14645 35 14675
rect 35 14645 36 14675
rect 4 14644 36 14645
rect 4 14595 36 14596
rect 4 14565 5 14595
rect 5 14565 35 14595
rect 35 14565 36 14595
rect 4 14564 36 14565
rect 4 14515 36 14516
rect 4 14485 5 14515
rect 5 14485 35 14515
rect 35 14485 36 14515
rect 4 14484 36 14485
rect 4 14435 36 14436
rect 4 14405 5 14435
rect 5 14405 35 14435
rect 35 14405 36 14435
rect 4 14404 36 14405
rect 4 14355 36 14356
rect 4 14325 5 14355
rect 5 14325 35 14355
rect 35 14325 36 14355
rect 4 14324 36 14325
rect 4 14275 36 14276
rect 4 14245 5 14275
rect 5 14245 35 14275
rect 35 14245 36 14275
rect 4 14244 36 14245
rect 4 14195 36 14196
rect 4 14165 5 14195
rect 5 14165 35 14195
rect 35 14165 36 14195
rect 4 14164 36 14165
rect 4 14115 36 14116
rect 4 14085 5 14115
rect 5 14085 35 14115
rect 35 14085 36 14115
rect 4 14084 36 14085
rect 4 14035 36 14036
rect 4 14005 5 14035
rect 5 14005 35 14035
rect 35 14005 36 14035
rect 4 14004 36 14005
rect 4 13955 36 13956
rect 4 13925 5 13955
rect 5 13925 35 13955
rect 35 13925 36 13955
rect 4 13924 36 13925
rect 4 13875 36 13876
rect 4 13845 5 13875
rect 5 13845 35 13875
rect 35 13845 36 13875
rect 4 13844 36 13845
rect 4 13795 36 13796
rect 4 13765 5 13795
rect 5 13765 35 13795
rect 35 13765 36 13795
rect 4 13764 36 13765
rect 4 13715 36 13716
rect 4 13685 5 13715
rect 5 13685 35 13715
rect 35 13685 36 13715
rect 4 13684 36 13685
rect 4 13635 36 13636
rect 4 13605 5 13635
rect 5 13605 35 13635
rect 35 13605 36 13635
rect 4 13604 36 13605
rect 4 13555 36 13556
rect 4 13525 5 13555
rect 5 13525 35 13555
rect 35 13525 36 13555
rect 4 13524 36 13525
rect 4 13475 36 13476
rect 4 13445 5 13475
rect 5 13445 35 13475
rect 35 13445 36 13475
rect 4 13444 36 13445
rect 4 13395 36 13396
rect 4 13365 5 13395
rect 5 13365 35 13395
rect 35 13365 36 13395
rect 4 13364 36 13365
rect 4 13315 36 13316
rect 4 13285 5 13315
rect 5 13285 35 13315
rect 35 13285 36 13315
rect 4 13284 36 13285
rect 4 13235 36 13236
rect 4 13205 5 13235
rect 5 13205 35 13235
rect 35 13205 36 13235
rect 4 13204 36 13205
rect 4 13155 36 13156
rect 4 13125 5 13155
rect 5 13125 35 13155
rect 35 13125 36 13155
rect 4 13124 36 13125
rect 4 13075 36 13076
rect 4 13045 5 13075
rect 5 13045 35 13075
rect 35 13045 36 13075
rect 4 13044 36 13045
rect 4 12995 36 12996
rect 4 12965 5 12995
rect 5 12965 35 12995
rect 35 12965 36 12995
rect 4 12964 36 12965
rect 4 12915 36 12916
rect 4 12885 5 12915
rect 5 12885 35 12915
rect 35 12885 36 12915
rect 4 12884 36 12885
rect 4 12835 36 12836
rect 4 12805 5 12835
rect 5 12805 35 12835
rect 35 12805 36 12835
rect 4 12804 36 12805
rect 4 12755 36 12756
rect 4 12725 5 12755
rect 5 12725 35 12755
rect 35 12725 36 12755
rect 4 12724 36 12725
rect 4 12675 36 12676
rect 4 12645 5 12675
rect 5 12645 35 12675
rect 35 12645 36 12675
rect 4 12644 36 12645
rect 4 12595 36 12596
rect 4 12565 5 12595
rect 5 12565 35 12595
rect 35 12565 36 12595
rect 4 12564 36 12565
rect 4 12515 36 12516
rect 4 12485 5 12515
rect 5 12485 35 12515
rect 35 12485 36 12515
rect 4 12484 36 12485
rect 4 12435 36 12436
rect 4 12405 5 12435
rect 5 12405 35 12435
rect 35 12405 36 12435
rect 4 12404 36 12405
rect 4 12355 36 12356
rect 4 12325 5 12355
rect 5 12325 35 12355
rect 35 12325 36 12355
rect 4 12324 36 12325
rect 4 12275 36 12276
rect 4 12245 5 12275
rect 5 12245 35 12275
rect 35 12245 36 12275
rect 4 12244 36 12245
rect 4 12195 36 12196
rect 4 12165 5 12195
rect 5 12165 35 12195
rect 35 12165 36 12195
rect 4 12164 36 12165
rect 4 12115 36 12116
rect 4 12085 5 12115
rect 5 12085 35 12115
rect 35 12085 36 12115
rect 4 12084 36 12085
rect 4 12035 36 12036
rect 4 12005 5 12035
rect 5 12005 35 12035
rect 35 12005 36 12035
rect 4 12004 36 12005
rect 4 11955 36 11956
rect 4 11925 5 11955
rect 5 11925 35 11955
rect 35 11925 36 11955
rect 4 11924 36 11925
rect 4 11875 36 11876
rect 4 11845 5 11875
rect 5 11845 35 11875
rect 35 11845 36 11875
rect 4 11844 36 11845
rect 4 11795 36 11796
rect 4 11765 5 11795
rect 5 11765 35 11795
rect 35 11765 36 11795
rect 4 11764 36 11765
rect 4 11715 36 11716
rect 4 11685 5 11715
rect 5 11685 35 11715
rect 35 11685 36 11715
rect 4 11684 36 11685
rect 4 11635 36 11636
rect 4 11605 5 11635
rect 5 11605 35 11635
rect 35 11605 36 11635
rect 4 11604 36 11605
rect 4 11555 36 11556
rect 4 11525 5 11555
rect 5 11525 35 11555
rect 35 11525 36 11555
rect 4 11524 36 11525
rect 4 11475 36 11476
rect 4 11445 5 11475
rect 5 11445 35 11475
rect 35 11445 36 11475
rect 4 11444 36 11445
rect 4 11395 36 11396
rect 4 11365 5 11395
rect 5 11365 35 11395
rect 35 11365 36 11395
rect 4 11364 36 11365
rect 4 11235 36 11236
rect 4 11205 5 11235
rect 5 11205 35 11235
rect 35 11205 36 11235
rect 4 11204 36 11205
rect 4 11155 36 11156
rect 4 11125 5 11155
rect 5 11125 35 11155
rect 35 11125 36 11155
rect 4 11124 36 11125
rect 4 11075 36 11076
rect 4 11045 5 11075
rect 5 11045 35 11075
rect 35 11045 36 11075
rect 4 11044 36 11045
rect 4 10995 36 10996
rect 4 10965 5 10995
rect 5 10965 35 10995
rect 35 10965 36 10995
rect 4 10964 36 10965
rect 4 10915 36 10916
rect 4 10885 5 10915
rect 5 10885 35 10915
rect 35 10885 36 10915
rect 4 10884 36 10885
rect 4 10835 36 10836
rect 4 10805 5 10835
rect 5 10805 35 10835
rect 35 10805 36 10835
rect 4 10804 36 10805
rect 4 10755 36 10756
rect 4 10725 5 10755
rect 5 10725 35 10755
rect 35 10725 36 10755
rect 4 10724 36 10725
rect 4 10675 36 10676
rect 4 10645 5 10675
rect 5 10645 35 10675
rect 35 10645 36 10675
rect 4 10644 36 10645
rect 4 10595 36 10596
rect 4 10565 5 10595
rect 5 10565 35 10595
rect 35 10565 36 10595
rect 4 10564 36 10565
rect 4 10515 36 10516
rect 4 10485 5 10515
rect 5 10485 35 10515
rect 35 10485 36 10515
rect 4 10484 36 10485
rect 4 10435 36 10436
rect 4 10405 5 10435
rect 5 10405 35 10435
rect 35 10405 36 10435
rect 4 10404 36 10405
rect 4 10355 36 10356
rect 4 10325 5 10355
rect 5 10325 35 10355
rect 35 10325 36 10355
rect 4 10324 36 10325
rect 4 10275 36 10276
rect 4 10245 5 10275
rect 5 10245 35 10275
rect 35 10245 36 10275
rect 4 10244 36 10245
rect 4 10195 36 10196
rect 4 10165 5 10195
rect 5 10165 35 10195
rect 35 10165 36 10195
rect 4 10164 36 10165
rect 4 10115 36 10116
rect 4 10085 5 10115
rect 5 10085 35 10115
rect 35 10085 36 10115
rect 4 10084 36 10085
rect 4 10035 36 10036
rect 4 10005 5 10035
rect 5 10005 35 10035
rect 35 10005 36 10035
rect 4 10004 36 10005
rect 4 9955 36 9956
rect 4 9925 5 9955
rect 5 9925 35 9955
rect 35 9925 36 9955
rect 4 9924 36 9925
rect 4 9875 36 9876
rect 4 9845 5 9875
rect 5 9845 35 9875
rect 35 9845 36 9875
rect 4 9844 36 9845
rect 4 9795 36 9796
rect 4 9765 5 9795
rect 5 9765 35 9795
rect 35 9765 36 9795
rect 4 9764 36 9765
rect 4 9715 36 9716
rect 4 9685 5 9715
rect 5 9685 35 9715
rect 35 9685 36 9715
rect 4 9684 36 9685
rect 4 9635 36 9636
rect 4 9605 5 9635
rect 5 9605 35 9635
rect 35 9605 36 9635
rect 4 9604 36 9605
rect 4 9555 36 9556
rect 4 9525 5 9555
rect 5 9525 35 9555
rect 35 9525 36 9555
rect 4 9524 36 9525
rect 4 9475 36 9476
rect 4 9445 5 9475
rect 5 9445 35 9475
rect 35 9445 36 9475
rect 4 9444 36 9445
rect 4 9395 36 9396
rect 4 9365 5 9395
rect 5 9365 35 9395
rect 35 9365 36 9395
rect 4 9364 36 9365
rect 4 9315 36 9316
rect 4 9285 5 9315
rect 5 9285 35 9315
rect 35 9285 36 9315
rect 4 9284 36 9285
rect 4 9235 36 9236
rect 4 9205 5 9235
rect 5 9205 35 9235
rect 35 9205 36 9235
rect 4 9204 36 9205
rect 4 9155 36 9156
rect 4 9125 5 9155
rect 5 9125 35 9155
rect 35 9125 36 9155
rect 4 9124 36 9125
rect 4 9075 36 9076
rect 4 9045 5 9075
rect 5 9045 35 9075
rect 35 9045 36 9075
rect 4 9044 36 9045
rect 4 8995 36 8996
rect 4 8965 5 8995
rect 5 8965 35 8995
rect 35 8965 36 8995
rect 4 8964 36 8965
rect 4 8915 36 8916
rect 4 8885 5 8915
rect 5 8885 35 8915
rect 35 8885 36 8915
rect 4 8884 36 8885
rect 4 8835 36 8836
rect 4 8805 5 8835
rect 5 8805 35 8835
rect 35 8805 36 8835
rect 4 8804 36 8805
rect 4 8755 36 8756
rect 4 8725 5 8755
rect 5 8725 35 8755
rect 35 8725 36 8755
rect 4 8724 36 8725
rect 4 8675 36 8676
rect 4 8645 5 8675
rect 5 8645 35 8675
rect 35 8645 36 8675
rect 4 8644 36 8645
rect 4 8595 36 8596
rect 4 8565 5 8595
rect 5 8565 35 8595
rect 35 8565 36 8595
rect 4 8564 36 8565
rect 4 8515 36 8516
rect 4 8485 5 8515
rect 5 8485 35 8515
rect 35 8485 36 8515
rect 4 8484 36 8485
rect 4 8355 36 8356
rect 4 8325 5 8355
rect 5 8325 35 8355
rect 35 8325 36 8355
rect 4 8324 36 8325
rect 4 8275 36 8276
rect 4 8245 5 8275
rect 5 8245 35 8275
rect 35 8245 36 8275
rect 4 8244 36 8245
rect 4 8195 36 8196
rect 4 8165 5 8195
rect 5 8165 35 8195
rect 35 8165 36 8195
rect 4 8164 36 8165
rect 4 8115 36 8116
rect 4 8085 5 8115
rect 5 8085 35 8115
rect 35 8085 36 8115
rect 4 8084 36 8085
rect 4 7955 36 7956
rect 4 7925 5 7955
rect 5 7925 35 7955
rect 35 7925 36 7955
rect 4 7924 36 7925
rect 4 7875 36 7876
rect 4 7845 5 7875
rect 5 7845 35 7875
rect 35 7845 36 7875
rect 4 7844 36 7845
rect 4 7795 36 7796
rect 4 7765 5 7795
rect 5 7765 35 7795
rect 35 7765 36 7795
rect 4 7764 36 7765
rect 4 7715 36 7716
rect 4 7685 5 7715
rect 5 7685 35 7715
rect 35 7685 36 7715
rect 4 7684 36 7685
rect 4 7635 36 7636
rect 4 7605 5 7635
rect 5 7605 35 7635
rect 35 7605 36 7635
rect 4 7604 36 7605
rect 4 7555 36 7556
rect 4 7525 5 7555
rect 5 7525 35 7555
rect 35 7525 36 7555
rect 4 7524 36 7525
rect 4 7475 36 7476
rect 4 7445 5 7475
rect 5 7445 35 7475
rect 35 7445 36 7475
rect 4 7444 36 7445
rect 4 7395 36 7396
rect 4 7365 5 7395
rect 5 7365 35 7395
rect 35 7365 36 7395
rect 4 7364 36 7365
rect 4 7315 36 7316
rect 4 7285 5 7315
rect 5 7285 35 7315
rect 35 7285 36 7315
rect 4 7284 36 7285
rect 4 7235 36 7236
rect 4 7205 5 7235
rect 5 7205 35 7235
rect 35 7205 36 7235
rect 4 7204 36 7205
rect 4 7155 36 7156
rect 4 7125 5 7155
rect 5 7125 35 7155
rect 35 7125 36 7155
rect 4 7124 36 7125
rect 4 7075 36 7076
rect 4 7045 5 7075
rect 5 7045 35 7075
rect 35 7045 36 7075
rect 4 7044 36 7045
rect 4 6995 36 6996
rect 4 6965 5 6995
rect 5 6965 35 6995
rect 35 6965 36 6995
rect 4 6964 36 6965
rect 4 6915 36 6916
rect 4 6885 5 6915
rect 5 6885 35 6915
rect 35 6885 36 6915
rect 4 6884 36 6885
rect 4 6835 36 6836
rect 4 6805 5 6835
rect 5 6805 35 6835
rect 35 6805 36 6835
rect 4 6804 36 6805
rect 4 6755 36 6756
rect 4 6725 5 6755
rect 5 6725 35 6755
rect 35 6725 36 6755
rect 4 6724 36 6725
rect 4 6675 36 6676
rect 4 6645 5 6675
rect 5 6645 35 6675
rect 35 6645 36 6675
rect 4 6644 36 6645
rect 4 6595 36 6596
rect 4 6565 5 6595
rect 5 6565 35 6595
rect 35 6565 36 6595
rect 4 6564 36 6565
rect 4 6515 36 6516
rect 4 6485 5 6515
rect 5 6485 35 6515
rect 35 6485 36 6515
rect 4 6484 36 6485
rect 4 6435 36 6436
rect 4 6405 5 6435
rect 5 6405 35 6435
rect 35 6405 36 6435
rect 4 6404 36 6405
rect 4 6355 36 6356
rect 4 6325 5 6355
rect 5 6325 35 6355
rect 35 6325 36 6355
rect 4 6324 36 6325
rect 4 6275 36 6276
rect 4 6245 5 6275
rect 5 6245 35 6275
rect 35 6245 36 6275
rect 4 6244 36 6245
rect 4 6195 36 6196
rect 4 6165 5 6195
rect 5 6165 35 6195
rect 35 6165 36 6195
rect 4 6164 36 6165
rect 4 6115 36 6116
rect 4 6085 5 6115
rect 5 6085 35 6115
rect 35 6085 36 6115
rect 4 6084 36 6085
rect 4 6035 36 6036
rect 4 6005 5 6035
rect 5 6005 35 6035
rect 35 6005 36 6035
rect 4 6004 36 6005
rect 4 5955 36 5956
rect 4 5925 5 5955
rect 5 5925 35 5955
rect 35 5925 36 5955
rect 4 5924 36 5925
rect 4 5875 36 5876
rect 4 5845 5 5875
rect 5 5845 35 5875
rect 35 5845 36 5875
rect 4 5844 36 5845
rect 4 5795 36 5796
rect 4 5765 5 5795
rect 5 5765 35 5795
rect 35 5765 36 5795
rect 4 5764 36 5765
rect 4 5715 36 5716
rect 4 5685 5 5715
rect 5 5685 35 5715
rect 35 5685 36 5715
rect 4 5684 36 5685
rect 4 5635 36 5636
rect 4 5605 5 5635
rect 5 5605 35 5635
rect 35 5605 36 5635
rect 4 5604 36 5605
rect 4 5555 36 5556
rect 4 5525 5 5555
rect 5 5525 35 5555
rect 35 5525 36 5555
rect 4 5524 36 5525
rect 4 5475 36 5476
rect 4 5445 5 5475
rect 5 5445 35 5475
rect 35 5445 36 5475
rect 4 5444 36 5445
rect 4 5395 36 5396
rect 4 5365 5 5395
rect 5 5365 35 5395
rect 35 5365 36 5395
rect 4 5364 36 5365
rect 4 5315 36 5316
rect 4 5285 5 5315
rect 5 5285 35 5315
rect 35 5285 36 5315
rect 4 5284 36 5285
rect 4 5235 36 5236
rect 4 5205 5 5235
rect 5 5205 35 5235
rect 35 5205 36 5235
rect 4 5204 36 5205
rect 4 5075 36 5076
rect 4 5045 5 5075
rect 5 5045 35 5075
rect 35 5045 36 5075
rect 4 5044 36 5045
rect 4 4995 36 4996
rect 4 4965 5 4995
rect 5 4965 35 4995
rect 35 4965 36 4995
rect 4 4964 36 4965
rect 4 4915 36 4916
rect 4 4885 5 4915
rect 5 4885 35 4915
rect 35 4885 36 4915
rect 4 4884 36 4885
rect 4 4835 36 4836
rect 4 4805 5 4835
rect 5 4805 35 4835
rect 35 4805 36 4835
rect 4 4804 36 4805
rect 4 4755 36 4756
rect 4 4725 5 4755
rect 5 4725 35 4755
rect 35 4725 36 4755
rect 4 4724 36 4725
rect 4 4675 36 4676
rect 4 4645 5 4675
rect 5 4645 35 4675
rect 35 4645 36 4675
rect 4 4644 36 4645
rect 4 4595 36 4596
rect 4 4565 5 4595
rect 5 4565 35 4595
rect 35 4565 36 4595
rect 4 4564 36 4565
rect 4 4515 36 4516
rect 4 4485 5 4515
rect 5 4485 35 4515
rect 35 4485 36 4515
rect 4 4484 36 4485
rect 4 4435 36 4436
rect 4 4405 5 4435
rect 5 4405 35 4435
rect 35 4405 36 4435
rect 4 4404 36 4405
rect 4 4355 36 4356
rect 4 4325 5 4355
rect 5 4325 35 4355
rect 35 4325 36 4355
rect 4 4324 36 4325
rect 4 4275 36 4276
rect 4 4245 5 4275
rect 5 4245 35 4275
rect 35 4245 36 4275
rect 4 4244 36 4245
rect 4 4195 36 4196
rect 4 4165 5 4195
rect 5 4165 35 4195
rect 35 4165 36 4195
rect 4 4164 36 4165
rect 4 4115 36 4116
rect 4 4085 5 4115
rect 5 4085 35 4115
rect 35 4085 36 4115
rect 4 4084 36 4085
rect 4 4035 36 4036
rect 4 4005 5 4035
rect 5 4005 35 4035
rect 35 4005 36 4035
rect 4 4004 36 4005
rect 4 3955 36 3956
rect 4 3925 5 3955
rect 5 3925 35 3955
rect 35 3925 36 3955
rect 4 3924 36 3925
rect 4 3875 36 3876
rect 4 3845 5 3875
rect 5 3845 35 3875
rect 35 3845 36 3875
rect 4 3844 36 3845
rect 4 3795 36 3796
rect 4 3765 5 3795
rect 5 3765 35 3795
rect 35 3765 36 3795
rect 4 3764 36 3765
rect 4 3715 36 3716
rect 4 3685 5 3715
rect 5 3685 35 3715
rect 35 3685 36 3715
rect 4 3684 36 3685
rect 4 3635 36 3636
rect 4 3605 5 3635
rect 5 3605 35 3635
rect 35 3605 36 3635
rect 4 3604 36 3605
rect 4 3555 36 3556
rect 4 3525 5 3555
rect 5 3525 35 3555
rect 35 3525 36 3555
rect 4 3524 36 3525
rect 4 3475 36 3476
rect 4 3445 5 3475
rect 5 3445 35 3475
rect 35 3445 36 3475
rect 4 3444 36 3445
rect 4 3395 36 3396
rect 4 3365 5 3395
rect 5 3365 35 3395
rect 35 3365 36 3395
rect 4 3364 36 3365
rect 4 3315 36 3316
rect 4 3285 5 3315
rect 5 3285 35 3315
rect 35 3285 36 3315
rect 4 3284 36 3285
rect 4 3235 36 3236
rect 4 3205 5 3235
rect 5 3205 35 3235
rect 35 3205 36 3235
rect 4 3204 36 3205
rect 4 3155 36 3156
rect 4 3125 5 3155
rect 5 3125 35 3155
rect 35 3125 36 3155
rect 4 3124 36 3125
rect 4 3075 36 3076
rect 4 3045 5 3075
rect 5 3045 35 3075
rect 35 3045 36 3075
rect 4 3044 36 3045
rect 4 2995 36 2996
rect 4 2965 5 2995
rect 5 2965 35 2995
rect 35 2965 36 2995
rect 4 2964 36 2965
rect 4 2915 36 2916
rect 4 2885 5 2915
rect 5 2885 35 2915
rect 35 2885 36 2915
rect 4 2884 36 2885
rect 4 2835 36 2836
rect 4 2805 5 2835
rect 5 2805 35 2835
rect 35 2805 36 2835
rect 4 2804 36 2805
rect 4 2755 36 2756
rect 4 2725 5 2755
rect 5 2725 35 2755
rect 35 2725 36 2755
rect 4 2724 36 2725
rect 4 2675 36 2676
rect 4 2645 5 2675
rect 5 2645 35 2675
rect 35 2645 36 2675
rect 4 2644 36 2645
rect 4 2595 36 2596
rect 4 2565 5 2595
rect 5 2565 35 2595
rect 35 2565 36 2595
rect 4 2564 36 2565
rect 4 2515 36 2516
rect 4 2485 5 2515
rect 5 2485 35 2515
rect 35 2485 36 2515
rect 4 2484 36 2485
rect 4 2435 36 2436
rect 4 2405 5 2435
rect 5 2405 35 2435
rect 35 2405 36 2435
rect 4 2404 36 2405
rect 4 2355 36 2356
rect 4 2325 5 2355
rect 5 2325 35 2355
rect 35 2325 36 2355
rect 4 2324 36 2325
rect 4 2275 36 2276
rect 4 2245 5 2275
rect 5 2245 35 2275
rect 35 2245 36 2275
rect 4 2244 36 2245
rect 4 2195 36 2196
rect 4 2165 5 2195
rect 5 2165 35 2195
rect 35 2165 36 2195
rect 4 2164 36 2165
rect 4 2115 36 2116
rect 4 2085 5 2115
rect 5 2085 35 2115
rect 35 2085 36 2115
rect 4 2084 36 2085
rect 4 2035 36 2036
rect 4 2005 5 2035
rect 5 2005 35 2035
rect 35 2005 36 2035
rect 4 2004 36 2005
rect 4 1955 36 1956
rect 4 1925 5 1955
rect 5 1925 35 1955
rect 35 1925 36 1955
rect 4 1924 36 1925
rect 4 1875 36 1876
rect 4 1845 5 1875
rect 5 1845 35 1875
rect 35 1845 36 1875
rect 4 1844 36 1845
rect 4 1795 36 1796
rect 4 1765 5 1795
rect 5 1765 35 1795
rect 35 1765 36 1795
rect 4 1764 36 1765
rect 4 1715 36 1716
rect 4 1685 5 1715
rect 5 1685 35 1715
rect 35 1685 36 1715
rect 4 1684 36 1685
rect 4 1635 36 1636
rect 4 1605 5 1635
rect 5 1605 35 1635
rect 35 1605 36 1635
rect 4 1604 36 1605
rect 4 1555 36 1556
rect 4 1525 5 1555
rect 5 1525 35 1555
rect 35 1525 36 1555
rect 4 1524 36 1525
rect 4 1475 36 1476
rect 4 1445 5 1475
rect 5 1445 35 1475
rect 35 1445 36 1475
rect 4 1444 36 1445
rect 4 1395 36 1396
rect 4 1365 5 1395
rect 5 1365 35 1395
rect 35 1365 36 1395
rect 4 1364 36 1365
rect 4 1315 36 1316
rect 4 1285 5 1315
rect 5 1285 35 1315
rect 35 1285 36 1315
rect 4 1284 36 1285
rect 4 1235 36 1236
rect 4 1205 5 1235
rect 5 1205 35 1235
rect 35 1205 36 1235
rect 4 1204 36 1205
rect 4 1155 36 1156
rect 4 1125 5 1155
rect 5 1125 35 1155
rect 35 1125 36 1155
rect 4 1124 36 1125
rect 4 1075 36 1076
rect 4 1045 5 1075
rect 5 1045 35 1075
rect 35 1045 36 1075
rect 4 1044 36 1045
rect 4 995 36 996
rect 4 965 5 995
rect 5 965 35 995
rect 35 965 36 995
rect 4 964 36 965
rect 4 915 36 916
rect 4 885 5 915
rect 5 885 35 915
rect 35 885 36 915
rect 4 884 36 885
rect 4 835 36 836
rect 4 805 5 835
rect 5 805 35 835
rect 35 805 36 835
rect 4 804 36 805
rect 4 755 36 756
rect 4 725 5 755
rect 5 725 35 755
rect 35 725 36 755
rect 4 724 36 725
rect 4 675 36 676
rect 4 645 5 675
rect 5 645 35 675
rect 35 645 36 675
rect 4 644 36 645
rect 4 595 36 596
rect 4 565 5 595
rect 5 565 35 595
rect 35 565 36 595
rect 4 564 36 565
rect 4 515 36 516
rect 4 485 5 515
rect 5 485 35 515
rect 35 485 36 515
rect 4 484 36 485
rect 84 11284 116 11316
rect 84 8404 116 8436
rect 84 8004 116 8036
rect 84 5124 116 5156
rect 164 15955 196 15956
rect 164 15925 165 15955
rect 165 15925 195 15955
rect 195 15925 196 15955
rect 164 15924 196 15925
rect 164 15875 196 15876
rect 164 15845 165 15875
rect 165 15845 195 15875
rect 195 15845 196 15875
rect 164 15844 196 15845
rect 164 15795 196 15796
rect 164 15765 165 15795
rect 165 15765 195 15795
rect 195 15765 196 15795
rect 164 15764 196 15765
rect 164 15715 196 15716
rect 164 15685 165 15715
rect 165 15685 195 15715
rect 195 15685 196 15715
rect 164 15684 196 15685
rect 164 15635 196 15636
rect 164 15605 165 15635
rect 165 15605 195 15635
rect 195 15605 196 15635
rect 164 15604 196 15605
rect 164 15555 196 15556
rect 164 15525 165 15555
rect 165 15525 195 15555
rect 195 15525 196 15555
rect 164 15524 196 15525
rect 164 15475 196 15476
rect 164 15445 165 15475
rect 165 15445 195 15475
rect 195 15445 196 15475
rect 164 15444 196 15445
rect 164 15395 196 15396
rect 164 15365 165 15395
rect 165 15365 195 15395
rect 195 15365 196 15395
rect 164 15364 196 15365
rect 164 15315 196 15316
rect 164 15285 165 15315
rect 165 15285 195 15315
rect 195 15285 196 15315
rect 164 15284 196 15285
rect 164 15235 196 15236
rect 164 15205 165 15235
rect 165 15205 195 15235
rect 195 15205 196 15235
rect 164 15204 196 15205
rect 164 15155 196 15156
rect 164 15125 165 15155
rect 165 15125 195 15155
rect 195 15125 196 15155
rect 164 15124 196 15125
rect 164 15075 196 15076
rect 164 15045 165 15075
rect 165 15045 195 15075
rect 195 15045 196 15075
rect 164 15044 196 15045
rect 164 14995 196 14996
rect 164 14965 165 14995
rect 165 14965 195 14995
rect 195 14965 196 14995
rect 164 14964 196 14965
rect 164 14915 196 14916
rect 164 14885 165 14915
rect 165 14885 195 14915
rect 195 14885 196 14915
rect 164 14884 196 14885
rect 164 14835 196 14836
rect 164 14805 165 14835
rect 165 14805 195 14835
rect 195 14805 196 14835
rect 164 14804 196 14805
rect 164 14755 196 14756
rect 164 14725 165 14755
rect 165 14725 195 14755
rect 195 14725 196 14755
rect 164 14724 196 14725
rect 164 14675 196 14676
rect 164 14645 165 14675
rect 165 14645 195 14675
rect 195 14645 196 14675
rect 164 14644 196 14645
rect 164 14595 196 14596
rect 164 14565 165 14595
rect 165 14565 195 14595
rect 195 14565 196 14595
rect 164 14564 196 14565
rect 164 14515 196 14516
rect 164 14485 165 14515
rect 165 14485 195 14515
rect 195 14485 196 14515
rect 164 14484 196 14485
rect 164 14435 196 14436
rect 164 14405 165 14435
rect 165 14405 195 14435
rect 195 14405 196 14435
rect 164 14404 196 14405
rect 164 14355 196 14356
rect 164 14325 165 14355
rect 165 14325 195 14355
rect 195 14325 196 14355
rect 164 14324 196 14325
rect 164 14275 196 14276
rect 164 14245 165 14275
rect 165 14245 195 14275
rect 195 14245 196 14275
rect 164 14244 196 14245
rect 164 14195 196 14196
rect 164 14165 165 14195
rect 165 14165 195 14195
rect 195 14165 196 14195
rect 164 14164 196 14165
rect 164 14115 196 14116
rect 164 14085 165 14115
rect 165 14085 195 14115
rect 195 14085 196 14115
rect 164 14084 196 14085
rect 164 14035 196 14036
rect 164 14005 165 14035
rect 165 14005 195 14035
rect 195 14005 196 14035
rect 164 14004 196 14005
rect 164 13955 196 13956
rect 164 13925 165 13955
rect 165 13925 195 13955
rect 195 13925 196 13955
rect 164 13924 196 13925
rect 164 13875 196 13876
rect 164 13845 165 13875
rect 165 13845 195 13875
rect 195 13845 196 13875
rect 164 13844 196 13845
rect 164 13795 196 13796
rect 164 13765 165 13795
rect 165 13765 195 13795
rect 195 13765 196 13795
rect 164 13764 196 13765
rect 164 13715 196 13716
rect 164 13685 165 13715
rect 165 13685 195 13715
rect 195 13685 196 13715
rect 164 13684 196 13685
rect 164 13635 196 13636
rect 164 13605 165 13635
rect 165 13605 195 13635
rect 195 13605 196 13635
rect 164 13604 196 13605
rect 164 13555 196 13556
rect 164 13525 165 13555
rect 165 13525 195 13555
rect 195 13525 196 13555
rect 164 13524 196 13525
rect 164 13475 196 13476
rect 164 13445 165 13475
rect 165 13445 195 13475
rect 195 13445 196 13475
rect 164 13444 196 13445
rect 164 13395 196 13396
rect 164 13365 165 13395
rect 165 13365 195 13395
rect 195 13365 196 13395
rect 164 13364 196 13365
rect 164 13315 196 13316
rect 164 13285 165 13315
rect 165 13285 195 13315
rect 195 13285 196 13315
rect 164 13284 196 13285
rect 164 13235 196 13236
rect 164 13205 165 13235
rect 165 13205 195 13235
rect 195 13205 196 13235
rect 164 13204 196 13205
rect 164 13155 196 13156
rect 164 13125 165 13155
rect 165 13125 195 13155
rect 195 13125 196 13155
rect 164 13124 196 13125
rect 164 13075 196 13076
rect 164 13045 165 13075
rect 165 13045 195 13075
rect 195 13045 196 13075
rect 164 13044 196 13045
rect 164 12995 196 12996
rect 164 12965 165 12995
rect 165 12965 195 12995
rect 195 12965 196 12995
rect 164 12964 196 12965
rect 164 12915 196 12916
rect 164 12885 165 12915
rect 165 12885 195 12915
rect 195 12885 196 12915
rect 164 12884 196 12885
rect 164 12835 196 12836
rect 164 12805 165 12835
rect 165 12805 195 12835
rect 195 12805 196 12835
rect 164 12804 196 12805
rect 164 12755 196 12756
rect 164 12725 165 12755
rect 165 12725 195 12755
rect 195 12725 196 12755
rect 164 12724 196 12725
rect 164 12675 196 12676
rect 164 12645 165 12675
rect 165 12645 195 12675
rect 195 12645 196 12675
rect 164 12644 196 12645
rect 164 12595 196 12596
rect 164 12565 165 12595
rect 165 12565 195 12595
rect 195 12565 196 12595
rect 164 12564 196 12565
rect 164 12515 196 12516
rect 164 12485 165 12515
rect 165 12485 195 12515
rect 195 12485 196 12515
rect 164 12484 196 12485
rect 164 12435 196 12436
rect 164 12405 165 12435
rect 165 12405 195 12435
rect 195 12405 196 12435
rect 164 12404 196 12405
rect 164 12355 196 12356
rect 164 12325 165 12355
rect 165 12325 195 12355
rect 195 12325 196 12355
rect 164 12324 196 12325
rect 164 12275 196 12276
rect 164 12245 165 12275
rect 165 12245 195 12275
rect 195 12245 196 12275
rect 164 12244 196 12245
rect 164 12195 196 12196
rect 164 12165 165 12195
rect 165 12165 195 12195
rect 195 12165 196 12195
rect 164 12164 196 12165
rect 164 12115 196 12116
rect 164 12085 165 12115
rect 165 12085 195 12115
rect 195 12085 196 12115
rect 164 12084 196 12085
rect 164 12035 196 12036
rect 164 12005 165 12035
rect 165 12005 195 12035
rect 195 12005 196 12035
rect 164 12004 196 12005
rect 164 11955 196 11956
rect 164 11925 165 11955
rect 165 11925 195 11955
rect 195 11925 196 11955
rect 164 11924 196 11925
rect 164 11875 196 11876
rect 164 11845 165 11875
rect 165 11845 195 11875
rect 195 11845 196 11875
rect 164 11844 196 11845
rect 164 11795 196 11796
rect 164 11765 165 11795
rect 165 11765 195 11795
rect 195 11765 196 11795
rect 164 11764 196 11765
rect 164 11715 196 11716
rect 164 11685 165 11715
rect 165 11685 195 11715
rect 195 11685 196 11715
rect 164 11684 196 11685
rect 164 11635 196 11636
rect 164 11605 165 11635
rect 165 11605 195 11635
rect 195 11605 196 11635
rect 164 11604 196 11605
rect 164 11555 196 11556
rect 164 11525 165 11555
rect 165 11525 195 11555
rect 195 11525 196 11555
rect 164 11524 196 11525
rect 164 11475 196 11476
rect 164 11445 165 11475
rect 165 11445 195 11475
rect 195 11445 196 11475
rect 164 11444 196 11445
rect 164 11395 196 11396
rect 164 11365 165 11395
rect 165 11365 195 11395
rect 195 11365 196 11395
rect 164 11364 196 11365
rect 164 11235 196 11236
rect 164 11205 165 11235
rect 165 11205 195 11235
rect 195 11205 196 11235
rect 164 11204 196 11205
rect 164 11155 196 11156
rect 164 11125 165 11155
rect 165 11125 195 11155
rect 195 11125 196 11155
rect 164 11124 196 11125
rect 164 11075 196 11076
rect 164 11045 165 11075
rect 165 11045 195 11075
rect 195 11045 196 11075
rect 164 11044 196 11045
rect 164 10995 196 10996
rect 164 10965 165 10995
rect 165 10965 195 10995
rect 195 10965 196 10995
rect 164 10964 196 10965
rect 164 10915 196 10916
rect 164 10885 165 10915
rect 165 10885 195 10915
rect 195 10885 196 10915
rect 164 10884 196 10885
rect 164 10835 196 10836
rect 164 10805 165 10835
rect 165 10805 195 10835
rect 195 10805 196 10835
rect 164 10804 196 10805
rect 164 10755 196 10756
rect 164 10725 165 10755
rect 165 10725 195 10755
rect 195 10725 196 10755
rect 164 10724 196 10725
rect 164 10675 196 10676
rect 164 10645 165 10675
rect 165 10645 195 10675
rect 195 10645 196 10675
rect 164 10644 196 10645
rect 164 10595 196 10596
rect 164 10565 165 10595
rect 165 10565 195 10595
rect 195 10565 196 10595
rect 164 10564 196 10565
rect 164 10515 196 10516
rect 164 10485 165 10515
rect 165 10485 195 10515
rect 195 10485 196 10515
rect 164 10484 196 10485
rect 164 10435 196 10436
rect 164 10405 165 10435
rect 165 10405 195 10435
rect 195 10405 196 10435
rect 164 10404 196 10405
rect 164 10355 196 10356
rect 164 10325 165 10355
rect 165 10325 195 10355
rect 195 10325 196 10355
rect 164 10324 196 10325
rect 164 10275 196 10276
rect 164 10245 165 10275
rect 165 10245 195 10275
rect 195 10245 196 10275
rect 164 10244 196 10245
rect 164 10195 196 10196
rect 164 10165 165 10195
rect 165 10165 195 10195
rect 195 10165 196 10195
rect 164 10164 196 10165
rect 164 10115 196 10116
rect 164 10085 165 10115
rect 165 10085 195 10115
rect 195 10085 196 10115
rect 164 10084 196 10085
rect 164 10035 196 10036
rect 164 10005 165 10035
rect 165 10005 195 10035
rect 195 10005 196 10035
rect 164 10004 196 10005
rect 164 9955 196 9956
rect 164 9925 165 9955
rect 165 9925 195 9955
rect 195 9925 196 9955
rect 164 9924 196 9925
rect 164 9875 196 9876
rect 164 9845 165 9875
rect 165 9845 195 9875
rect 195 9845 196 9875
rect 164 9844 196 9845
rect 164 9795 196 9796
rect 164 9765 165 9795
rect 165 9765 195 9795
rect 195 9765 196 9795
rect 164 9764 196 9765
rect 164 9715 196 9716
rect 164 9685 165 9715
rect 165 9685 195 9715
rect 195 9685 196 9715
rect 164 9684 196 9685
rect 164 9635 196 9636
rect 164 9605 165 9635
rect 165 9605 195 9635
rect 195 9605 196 9635
rect 164 9604 196 9605
rect 164 9555 196 9556
rect 164 9525 165 9555
rect 165 9525 195 9555
rect 195 9525 196 9555
rect 164 9524 196 9525
rect 164 9475 196 9476
rect 164 9445 165 9475
rect 165 9445 195 9475
rect 195 9445 196 9475
rect 164 9444 196 9445
rect 164 9395 196 9396
rect 164 9365 165 9395
rect 165 9365 195 9395
rect 195 9365 196 9395
rect 164 9364 196 9365
rect 164 9315 196 9316
rect 164 9285 165 9315
rect 165 9285 195 9315
rect 195 9285 196 9315
rect 164 9284 196 9285
rect 164 9235 196 9236
rect 164 9205 165 9235
rect 165 9205 195 9235
rect 195 9205 196 9235
rect 164 9204 196 9205
rect 164 9155 196 9156
rect 164 9125 165 9155
rect 165 9125 195 9155
rect 195 9125 196 9155
rect 164 9124 196 9125
rect 164 9075 196 9076
rect 164 9045 165 9075
rect 165 9045 195 9075
rect 195 9045 196 9075
rect 164 9044 196 9045
rect 164 8995 196 8996
rect 164 8965 165 8995
rect 165 8965 195 8995
rect 195 8965 196 8995
rect 164 8964 196 8965
rect 164 8915 196 8916
rect 164 8885 165 8915
rect 165 8885 195 8915
rect 195 8885 196 8915
rect 164 8884 196 8885
rect 164 8835 196 8836
rect 164 8805 165 8835
rect 165 8805 195 8835
rect 195 8805 196 8835
rect 164 8804 196 8805
rect 164 8755 196 8756
rect 164 8725 165 8755
rect 165 8725 195 8755
rect 195 8725 196 8755
rect 164 8724 196 8725
rect 164 8675 196 8676
rect 164 8645 165 8675
rect 165 8645 195 8675
rect 195 8645 196 8675
rect 164 8644 196 8645
rect 164 8595 196 8596
rect 164 8565 165 8595
rect 165 8565 195 8595
rect 195 8565 196 8595
rect 164 8564 196 8565
rect 164 8515 196 8516
rect 164 8485 165 8515
rect 165 8485 195 8515
rect 195 8485 196 8515
rect 164 8484 196 8485
rect 164 8355 196 8356
rect 164 8325 165 8355
rect 165 8325 195 8355
rect 195 8325 196 8355
rect 164 8324 196 8325
rect 164 8275 196 8276
rect 164 8245 165 8275
rect 165 8245 195 8275
rect 195 8245 196 8275
rect 164 8244 196 8245
rect 164 8195 196 8196
rect 164 8165 165 8195
rect 165 8165 195 8195
rect 195 8165 196 8195
rect 164 8164 196 8165
rect 164 8115 196 8116
rect 164 8085 165 8115
rect 165 8085 195 8115
rect 195 8085 196 8115
rect 164 8084 196 8085
rect 164 7955 196 7956
rect 164 7925 165 7955
rect 165 7925 195 7955
rect 195 7925 196 7955
rect 164 7924 196 7925
rect 164 7875 196 7876
rect 164 7845 165 7875
rect 165 7845 195 7875
rect 195 7845 196 7875
rect 164 7844 196 7845
rect 164 7795 196 7796
rect 164 7765 165 7795
rect 165 7765 195 7795
rect 195 7765 196 7795
rect 164 7764 196 7765
rect 164 7715 196 7716
rect 164 7685 165 7715
rect 165 7685 195 7715
rect 195 7685 196 7715
rect 164 7684 196 7685
rect 164 7635 196 7636
rect 164 7605 165 7635
rect 165 7605 195 7635
rect 195 7605 196 7635
rect 164 7604 196 7605
rect 164 7555 196 7556
rect 164 7525 165 7555
rect 165 7525 195 7555
rect 195 7525 196 7555
rect 164 7524 196 7525
rect 164 7475 196 7476
rect 164 7445 165 7475
rect 165 7445 195 7475
rect 195 7445 196 7475
rect 164 7444 196 7445
rect 164 7395 196 7396
rect 164 7365 165 7395
rect 165 7365 195 7395
rect 195 7365 196 7395
rect 164 7364 196 7365
rect 164 7315 196 7316
rect 164 7285 165 7315
rect 165 7285 195 7315
rect 195 7285 196 7315
rect 164 7284 196 7285
rect 164 7235 196 7236
rect 164 7205 165 7235
rect 165 7205 195 7235
rect 195 7205 196 7235
rect 164 7204 196 7205
rect 164 7155 196 7156
rect 164 7125 165 7155
rect 165 7125 195 7155
rect 195 7125 196 7155
rect 164 7124 196 7125
rect 164 7075 196 7076
rect 164 7045 165 7075
rect 165 7045 195 7075
rect 195 7045 196 7075
rect 164 7044 196 7045
rect 164 6995 196 6996
rect 164 6965 165 6995
rect 165 6965 195 6995
rect 195 6965 196 6995
rect 164 6964 196 6965
rect 164 6915 196 6916
rect 164 6885 165 6915
rect 165 6885 195 6915
rect 195 6885 196 6915
rect 164 6884 196 6885
rect 164 6835 196 6836
rect 164 6805 165 6835
rect 165 6805 195 6835
rect 195 6805 196 6835
rect 164 6804 196 6805
rect 164 6755 196 6756
rect 164 6725 165 6755
rect 165 6725 195 6755
rect 195 6725 196 6755
rect 164 6724 196 6725
rect 164 6675 196 6676
rect 164 6645 165 6675
rect 165 6645 195 6675
rect 195 6645 196 6675
rect 164 6644 196 6645
rect 164 6595 196 6596
rect 164 6565 165 6595
rect 165 6565 195 6595
rect 195 6565 196 6595
rect 164 6564 196 6565
rect 164 6515 196 6516
rect 164 6485 165 6515
rect 165 6485 195 6515
rect 195 6485 196 6515
rect 164 6484 196 6485
rect 164 6435 196 6436
rect 164 6405 165 6435
rect 165 6405 195 6435
rect 195 6405 196 6435
rect 164 6404 196 6405
rect 164 6355 196 6356
rect 164 6325 165 6355
rect 165 6325 195 6355
rect 195 6325 196 6355
rect 164 6324 196 6325
rect 164 6275 196 6276
rect 164 6245 165 6275
rect 165 6245 195 6275
rect 195 6245 196 6275
rect 164 6244 196 6245
rect 164 6195 196 6196
rect 164 6165 165 6195
rect 165 6165 195 6195
rect 195 6165 196 6195
rect 164 6164 196 6165
rect 164 6115 196 6116
rect 164 6085 165 6115
rect 165 6085 195 6115
rect 195 6085 196 6115
rect 164 6084 196 6085
rect 164 6035 196 6036
rect 164 6005 165 6035
rect 165 6005 195 6035
rect 195 6005 196 6035
rect 164 6004 196 6005
rect 164 5955 196 5956
rect 164 5925 165 5955
rect 165 5925 195 5955
rect 195 5925 196 5955
rect 164 5924 196 5925
rect 164 5875 196 5876
rect 164 5845 165 5875
rect 165 5845 195 5875
rect 195 5845 196 5875
rect 164 5844 196 5845
rect 164 5795 196 5796
rect 164 5765 165 5795
rect 165 5765 195 5795
rect 195 5765 196 5795
rect 164 5764 196 5765
rect 164 5715 196 5716
rect 164 5685 165 5715
rect 165 5685 195 5715
rect 195 5685 196 5715
rect 164 5684 196 5685
rect 164 5635 196 5636
rect 164 5605 165 5635
rect 165 5605 195 5635
rect 195 5605 196 5635
rect 164 5604 196 5605
rect 164 5555 196 5556
rect 164 5525 165 5555
rect 165 5525 195 5555
rect 195 5525 196 5555
rect 164 5524 196 5525
rect 164 5475 196 5476
rect 164 5445 165 5475
rect 165 5445 195 5475
rect 195 5445 196 5475
rect 164 5444 196 5445
rect 164 5395 196 5396
rect 164 5365 165 5395
rect 165 5365 195 5395
rect 195 5365 196 5395
rect 164 5364 196 5365
rect 164 5315 196 5316
rect 164 5285 165 5315
rect 165 5285 195 5315
rect 195 5285 196 5315
rect 164 5284 196 5285
rect 164 5235 196 5236
rect 164 5205 165 5235
rect 165 5205 195 5235
rect 195 5205 196 5235
rect 164 5204 196 5205
rect 164 5075 196 5076
rect 164 5045 165 5075
rect 165 5045 195 5075
rect 195 5045 196 5075
rect 164 5044 196 5045
rect 164 4995 196 4996
rect 164 4965 165 4995
rect 165 4965 195 4995
rect 195 4965 196 4995
rect 164 4964 196 4965
rect 164 4915 196 4916
rect 164 4885 165 4915
rect 165 4885 195 4915
rect 195 4885 196 4915
rect 164 4884 196 4885
rect 164 4835 196 4836
rect 164 4805 165 4835
rect 165 4805 195 4835
rect 195 4805 196 4835
rect 164 4804 196 4805
rect 164 4755 196 4756
rect 164 4725 165 4755
rect 165 4725 195 4755
rect 195 4725 196 4755
rect 164 4724 196 4725
rect 164 4675 196 4676
rect 164 4645 165 4675
rect 165 4645 195 4675
rect 195 4645 196 4675
rect 164 4644 196 4645
rect 164 4595 196 4596
rect 164 4565 165 4595
rect 165 4565 195 4595
rect 195 4565 196 4595
rect 164 4564 196 4565
rect 164 4515 196 4516
rect 164 4485 165 4515
rect 165 4485 195 4515
rect 195 4485 196 4515
rect 164 4484 196 4485
rect 164 4435 196 4436
rect 164 4405 165 4435
rect 165 4405 195 4435
rect 195 4405 196 4435
rect 164 4404 196 4405
rect 164 4355 196 4356
rect 164 4325 165 4355
rect 165 4325 195 4355
rect 195 4325 196 4355
rect 164 4324 196 4325
rect 164 4275 196 4276
rect 164 4245 165 4275
rect 165 4245 195 4275
rect 195 4245 196 4275
rect 164 4244 196 4245
rect 164 4195 196 4196
rect 164 4165 165 4195
rect 165 4165 195 4195
rect 195 4165 196 4195
rect 164 4164 196 4165
rect 164 4115 196 4116
rect 164 4085 165 4115
rect 165 4085 195 4115
rect 195 4085 196 4115
rect 164 4084 196 4085
rect 164 4035 196 4036
rect 164 4005 165 4035
rect 165 4005 195 4035
rect 195 4005 196 4035
rect 164 4004 196 4005
rect 164 3955 196 3956
rect 164 3925 165 3955
rect 165 3925 195 3955
rect 195 3925 196 3955
rect 164 3924 196 3925
rect 164 3875 196 3876
rect 164 3845 165 3875
rect 165 3845 195 3875
rect 195 3845 196 3875
rect 164 3844 196 3845
rect 164 3795 196 3796
rect 164 3765 165 3795
rect 165 3765 195 3795
rect 195 3765 196 3795
rect 164 3764 196 3765
rect 164 3715 196 3716
rect 164 3685 165 3715
rect 165 3685 195 3715
rect 195 3685 196 3715
rect 164 3684 196 3685
rect 164 3635 196 3636
rect 164 3605 165 3635
rect 165 3605 195 3635
rect 195 3605 196 3635
rect 164 3604 196 3605
rect 164 3555 196 3556
rect 164 3525 165 3555
rect 165 3525 195 3555
rect 195 3525 196 3555
rect 164 3524 196 3525
rect 164 3475 196 3476
rect 164 3445 165 3475
rect 165 3445 195 3475
rect 195 3445 196 3475
rect 164 3444 196 3445
rect 164 3395 196 3396
rect 164 3365 165 3395
rect 165 3365 195 3395
rect 195 3365 196 3395
rect 164 3364 196 3365
rect 164 3315 196 3316
rect 164 3285 165 3315
rect 165 3285 195 3315
rect 195 3285 196 3315
rect 164 3284 196 3285
rect 164 3235 196 3236
rect 164 3205 165 3235
rect 165 3205 195 3235
rect 195 3205 196 3235
rect 164 3204 196 3205
rect 164 3155 196 3156
rect 164 3125 165 3155
rect 165 3125 195 3155
rect 195 3125 196 3155
rect 164 3124 196 3125
rect 164 3075 196 3076
rect 164 3045 165 3075
rect 165 3045 195 3075
rect 195 3045 196 3075
rect 164 3044 196 3045
rect 164 2995 196 2996
rect 164 2965 165 2995
rect 165 2965 195 2995
rect 195 2965 196 2995
rect 164 2964 196 2965
rect 164 2915 196 2916
rect 164 2885 165 2915
rect 165 2885 195 2915
rect 195 2885 196 2915
rect 164 2884 196 2885
rect 164 2835 196 2836
rect 164 2805 165 2835
rect 165 2805 195 2835
rect 195 2805 196 2835
rect 164 2804 196 2805
rect 164 2755 196 2756
rect 164 2725 165 2755
rect 165 2725 195 2755
rect 195 2725 196 2755
rect 164 2724 196 2725
rect 164 2675 196 2676
rect 164 2645 165 2675
rect 165 2645 195 2675
rect 195 2645 196 2675
rect 164 2644 196 2645
rect 164 2595 196 2596
rect 164 2565 165 2595
rect 165 2565 195 2595
rect 195 2565 196 2595
rect 164 2564 196 2565
rect 164 2515 196 2516
rect 164 2485 165 2515
rect 165 2485 195 2515
rect 195 2485 196 2515
rect 164 2484 196 2485
rect 164 2435 196 2436
rect 164 2405 165 2435
rect 165 2405 195 2435
rect 195 2405 196 2435
rect 164 2404 196 2405
rect 164 2355 196 2356
rect 164 2325 165 2355
rect 165 2325 195 2355
rect 195 2325 196 2355
rect 164 2324 196 2325
rect 164 2275 196 2276
rect 164 2245 165 2275
rect 165 2245 195 2275
rect 195 2245 196 2275
rect 164 2244 196 2245
rect 164 2195 196 2196
rect 164 2165 165 2195
rect 165 2165 195 2195
rect 195 2165 196 2195
rect 164 2164 196 2165
rect 164 2115 196 2116
rect 164 2085 165 2115
rect 165 2085 195 2115
rect 195 2085 196 2115
rect 164 2084 196 2085
rect 164 2035 196 2036
rect 164 2005 165 2035
rect 165 2005 195 2035
rect 195 2005 196 2035
rect 164 2004 196 2005
rect 164 1955 196 1956
rect 164 1925 165 1955
rect 165 1925 195 1955
rect 195 1925 196 1955
rect 164 1924 196 1925
rect 164 1875 196 1876
rect 164 1845 165 1875
rect 165 1845 195 1875
rect 195 1845 196 1875
rect 164 1844 196 1845
rect 164 1795 196 1796
rect 164 1765 165 1795
rect 165 1765 195 1795
rect 195 1765 196 1795
rect 164 1764 196 1765
rect 164 1715 196 1716
rect 164 1685 165 1715
rect 165 1685 195 1715
rect 195 1685 196 1715
rect 164 1684 196 1685
rect 164 1635 196 1636
rect 164 1605 165 1635
rect 165 1605 195 1635
rect 195 1605 196 1635
rect 164 1604 196 1605
rect 164 1555 196 1556
rect 164 1525 165 1555
rect 165 1525 195 1555
rect 195 1525 196 1555
rect 164 1524 196 1525
rect 164 1475 196 1476
rect 164 1445 165 1475
rect 165 1445 195 1475
rect 195 1445 196 1475
rect 164 1444 196 1445
rect 164 1395 196 1396
rect 164 1365 165 1395
rect 165 1365 195 1395
rect 195 1365 196 1395
rect 164 1364 196 1365
rect 164 1315 196 1316
rect 164 1285 165 1315
rect 165 1285 195 1315
rect 195 1285 196 1315
rect 164 1284 196 1285
rect 164 1235 196 1236
rect 164 1205 165 1235
rect 165 1205 195 1235
rect 195 1205 196 1235
rect 164 1204 196 1205
rect 164 1155 196 1156
rect 164 1125 165 1155
rect 165 1125 195 1155
rect 195 1125 196 1155
rect 164 1124 196 1125
rect 164 1075 196 1076
rect 164 1045 165 1075
rect 165 1045 195 1075
rect 195 1045 196 1075
rect 164 1044 196 1045
rect 164 995 196 996
rect 164 965 165 995
rect 165 965 195 995
rect 195 965 196 995
rect 164 964 196 965
rect 164 915 196 916
rect 164 885 165 915
rect 165 885 195 915
rect 195 885 196 915
rect 164 884 196 885
rect 164 835 196 836
rect 164 805 165 835
rect 165 805 195 835
rect 195 805 196 835
rect 164 804 196 805
rect 164 755 196 756
rect 164 725 165 755
rect 165 725 195 755
rect 195 725 196 755
rect 164 724 196 725
rect 164 675 196 676
rect 164 645 165 675
rect 165 645 195 675
rect 195 645 196 675
rect 164 644 196 645
rect 164 595 196 596
rect 164 565 165 595
rect 165 565 195 595
rect 195 565 196 595
rect 164 564 196 565
rect 164 515 196 516
rect 164 485 165 515
rect 165 485 195 515
rect 195 485 196 515
rect 164 484 196 485
rect 4 244 36 436
rect 244 11124 276 11156
rect 244 8564 276 8596
rect 244 7844 276 7876
rect 244 5284 276 5316
rect 324 15955 356 15956
rect 324 15925 325 15955
rect 325 15925 355 15955
rect 355 15925 356 15955
rect 324 15924 356 15925
rect 324 15875 356 15876
rect 324 15845 325 15875
rect 325 15845 355 15875
rect 355 15845 356 15875
rect 324 15844 356 15845
rect 324 15795 356 15796
rect 324 15765 325 15795
rect 325 15765 355 15795
rect 355 15765 356 15795
rect 324 15764 356 15765
rect 324 15715 356 15716
rect 324 15685 325 15715
rect 325 15685 355 15715
rect 355 15685 356 15715
rect 324 15684 356 15685
rect 324 15635 356 15636
rect 324 15605 325 15635
rect 325 15605 355 15635
rect 355 15605 356 15635
rect 324 15604 356 15605
rect 324 15555 356 15556
rect 324 15525 325 15555
rect 325 15525 355 15555
rect 355 15525 356 15555
rect 324 15524 356 15525
rect 324 15475 356 15476
rect 324 15445 325 15475
rect 325 15445 355 15475
rect 355 15445 356 15475
rect 324 15444 356 15445
rect 324 15395 356 15396
rect 324 15365 325 15395
rect 325 15365 355 15395
rect 355 15365 356 15395
rect 324 15364 356 15365
rect 324 15315 356 15316
rect 324 15285 325 15315
rect 325 15285 355 15315
rect 355 15285 356 15315
rect 324 15284 356 15285
rect 324 15235 356 15236
rect 324 15205 325 15235
rect 325 15205 355 15235
rect 355 15205 356 15235
rect 324 15204 356 15205
rect 324 15155 356 15156
rect 324 15125 325 15155
rect 325 15125 355 15155
rect 355 15125 356 15155
rect 324 15124 356 15125
rect 324 15075 356 15076
rect 324 15045 325 15075
rect 325 15045 355 15075
rect 355 15045 356 15075
rect 324 15044 356 15045
rect 324 14995 356 14996
rect 324 14965 325 14995
rect 325 14965 355 14995
rect 355 14965 356 14995
rect 324 14964 356 14965
rect 324 14915 356 14916
rect 324 14885 325 14915
rect 325 14885 355 14915
rect 355 14885 356 14915
rect 324 14884 356 14885
rect 324 14835 356 14836
rect 324 14805 325 14835
rect 325 14805 355 14835
rect 355 14805 356 14835
rect 324 14804 356 14805
rect 324 14755 356 14756
rect 324 14725 325 14755
rect 325 14725 355 14755
rect 355 14725 356 14755
rect 324 14724 356 14725
rect 324 14675 356 14676
rect 324 14645 325 14675
rect 325 14645 355 14675
rect 355 14645 356 14675
rect 324 14644 356 14645
rect 324 14595 356 14596
rect 324 14565 325 14595
rect 325 14565 355 14595
rect 355 14565 356 14595
rect 324 14564 356 14565
rect 324 14515 356 14516
rect 324 14485 325 14515
rect 325 14485 355 14515
rect 355 14485 356 14515
rect 324 14484 356 14485
rect 324 14435 356 14436
rect 324 14405 325 14435
rect 325 14405 355 14435
rect 355 14405 356 14435
rect 324 14404 356 14405
rect 324 14355 356 14356
rect 324 14325 325 14355
rect 325 14325 355 14355
rect 355 14325 356 14355
rect 324 14324 356 14325
rect 324 14275 356 14276
rect 324 14245 325 14275
rect 325 14245 355 14275
rect 355 14245 356 14275
rect 324 14244 356 14245
rect 324 14195 356 14196
rect 324 14165 325 14195
rect 325 14165 355 14195
rect 355 14165 356 14195
rect 324 14164 356 14165
rect 324 14115 356 14116
rect 324 14085 325 14115
rect 325 14085 355 14115
rect 355 14085 356 14115
rect 324 14084 356 14085
rect 324 14035 356 14036
rect 324 14005 325 14035
rect 325 14005 355 14035
rect 355 14005 356 14035
rect 324 14004 356 14005
rect 324 13955 356 13956
rect 324 13925 325 13955
rect 325 13925 355 13955
rect 355 13925 356 13955
rect 324 13924 356 13925
rect 324 13875 356 13876
rect 324 13845 325 13875
rect 325 13845 355 13875
rect 355 13845 356 13875
rect 324 13844 356 13845
rect 324 13795 356 13796
rect 324 13765 325 13795
rect 325 13765 355 13795
rect 355 13765 356 13795
rect 324 13764 356 13765
rect 324 13715 356 13716
rect 324 13685 325 13715
rect 325 13685 355 13715
rect 355 13685 356 13715
rect 324 13684 356 13685
rect 324 13635 356 13636
rect 324 13605 325 13635
rect 325 13605 355 13635
rect 355 13605 356 13635
rect 324 13604 356 13605
rect 324 13555 356 13556
rect 324 13525 325 13555
rect 325 13525 355 13555
rect 355 13525 356 13555
rect 324 13524 356 13525
rect 324 13475 356 13476
rect 324 13445 325 13475
rect 325 13445 355 13475
rect 355 13445 356 13475
rect 324 13444 356 13445
rect 324 13395 356 13396
rect 324 13365 325 13395
rect 325 13365 355 13395
rect 355 13365 356 13395
rect 324 13364 356 13365
rect 324 13315 356 13316
rect 324 13285 325 13315
rect 325 13285 355 13315
rect 355 13285 356 13315
rect 324 13284 356 13285
rect 324 13235 356 13236
rect 324 13205 325 13235
rect 325 13205 355 13235
rect 355 13205 356 13235
rect 324 13204 356 13205
rect 324 13155 356 13156
rect 324 13125 325 13155
rect 325 13125 355 13155
rect 355 13125 356 13155
rect 324 13124 356 13125
rect 324 13075 356 13076
rect 324 13045 325 13075
rect 325 13045 355 13075
rect 355 13045 356 13075
rect 324 13044 356 13045
rect 324 12995 356 12996
rect 324 12965 325 12995
rect 325 12965 355 12995
rect 355 12965 356 12995
rect 324 12964 356 12965
rect 324 12915 356 12916
rect 324 12885 325 12915
rect 325 12885 355 12915
rect 355 12885 356 12915
rect 324 12884 356 12885
rect 324 12835 356 12836
rect 324 12805 325 12835
rect 325 12805 355 12835
rect 355 12805 356 12835
rect 324 12804 356 12805
rect 324 12755 356 12756
rect 324 12725 325 12755
rect 325 12725 355 12755
rect 355 12725 356 12755
rect 324 12724 356 12725
rect 324 12675 356 12676
rect 324 12645 325 12675
rect 325 12645 355 12675
rect 355 12645 356 12675
rect 324 12644 356 12645
rect 324 12595 356 12596
rect 324 12565 325 12595
rect 325 12565 355 12595
rect 355 12565 356 12595
rect 324 12564 356 12565
rect 324 12515 356 12516
rect 324 12485 325 12515
rect 325 12485 355 12515
rect 355 12485 356 12515
rect 324 12484 356 12485
rect 324 12435 356 12436
rect 324 12405 325 12435
rect 325 12405 355 12435
rect 355 12405 356 12435
rect 324 12404 356 12405
rect 324 12355 356 12356
rect 324 12325 325 12355
rect 325 12325 355 12355
rect 355 12325 356 12355
rect 324 12324 356 12325
rect 324 12275 356 12276
rect 324 12245 325 12275
rect 325 12245 355 12275
rect 355 12245 356 12275
rect 324 12244 356 12245
rect 324 12195 356 12196
rect 324 12165 325 12195
rect 325 12165 355 12195
rect 355 12165 356 12195
rect 324 12164 356 12165
rect 324 12115 356 12116
rect 324 12085 325 12115
rect 325 12085 355 12115
rect 355 12085 356 12115
rect 324 12084 356 12085
rect 324 12035 356 12036
rect 324 12005 325 12035
rect 325 12005 355 12035
rect 355 12005 356 12035
rect 324 12004 356 12005
rect 324 11955 356 11956
rect 324 11925 325 11955
rect 325 11925 355 11955
rect 355 11925 356 11955
rect 324 11924 356 11925
rect 324 11875 356 11876
rect 324 11845 325 11875
rect 325 11845 355 11875
rect 355 11845 356 11875
rect 324 11844 356 11845
rect 324 11795 356 11796
rect 324 11765 325 11795
rect 325 11765 355 11795
rect 355 11765 356 11795
rect 324 11764 356 11765
rect 324 11715 356 11716
rect 324 11685 325 11715
rect 325 11685 355 11715
rect 355 11685 356 11715
rect 324 11684 356 11685
rect 324 11635 356 11636
rect 324 11605 325 11635
rect 325 11605 355 11635
rect 355 11605 356 11635
rect 324 11604 356 11605
rect 324 11555 356 11556
rect 324 11525 325 11555
rect 325 11525 355 11555
rect 355 11525 356 11555
rect 324 11524 356 11525
rect 324 11475 356 11476
rect 324 11445 325 11475
rect 325 11445 355 11475
rect 355 11445 356 11475
rect 324 11444 356 11445
rect 324 11395 356 11396
rect 324 11365 325 11395
rect 325 11365 355 11395
rect 355 11365 356 11395
rect 324 11364 356 11365
rect 324 11235 356 11236
rect 324 11205 325 11235
rect 325 11205 355 11235
rect 355 11205 356 11235
rect 324 11204 356 11205
rect 324 11075 356 11076
rect 324 11045 325 11075
rect 325 11045 355 11075
rect 355 11045 356 11075
rect 324 11044 356 11045
rect 324 10995 356 10996
rect 324 10965 325 10995
rect 325 10965 355 10995
rect 355 10965 356 10995
rect 324 10964 356 10965
rect 324 10915 356 10916
rect 324 10885 325 10915
rect 325 10885 355 10915
rect 355 10885 356 10915
rect 324 10884 356 10885
rect 324 10835 356 10836
rect 324 10805 325 10835
rect 325 10805 355 10835
rect 355 10805 356 10835
rect 324 10804 356 10805
rect 324 10755 356 10756
rect 324 10725 325 10755
rect 325 10725 355 10755
rect 355 10725 356 10755
rect 324 10724 356 10725
rect 324 10675 356 10676
rect 324 10645 325 10675
rect 325 10645 355 10675
rect 355 10645 356 10675
rect 324 10644 356 10645
rect 324 10595 356 10596
rect 324 10565 325 10595
rect 325 10565 355 10595
rect 355 10565 356 10595
rect 324 10564 356 10565
rect 324 10515 356 10516
rect 324 10485 325 10515
rect 325 10485 355 10515
rect 355 10485 356 10515
rect 324 10484 356 10485
rect 324 10435 356 10436
rect 324 10405 325 10435
rect 325 10405 355 10435
rect 355 10405 356 10435
rect 324 10404 356 10405
rect 324 10355 356 10356
rect 324 10325 325 10355
rect 325 10325 355 10355
rect 355 10325 356 10355
rect 324 10324 356 10325
rect 324 10275 356 10276
rect 324 10245 325 10275
rect 325 10245 355 10275
rect 355 10245 356 10275
rect 324 10244 356 10245
rect 324 10195 356 10196
rect 324 10165 325 10195
rect 325 10165 355 10195
rect 355 10165 356 10195
rect 324 10164 356 10165
rect 324 10115 356 10116
rect 324 10085 325 10115
rect 325 10085 355 10115
rect 355 10085 356 10115
rect 324 10084 356 10085
rect 324 10035 356 10036
rect 324 10005 325 10035
rect 325 10005 355 10035
rect 355 10005 356 10035
rect 324 10004 356 10005
rect 324 9955 356 9956
rect 324 9925 325 9955
rect 325 9925 355 9955
rect 355 9925 356 9955
rect 324 9924 356 9925
rect 324 9875 356 9876
rect 324 9845 325 9875
rect 325 9845 355 9875
rect 355 9845 356 9875
rect 324 9844 356 9845
rect 324 9795 356 9796
rect 324 9765 325 9795
rect 325 9765 355 9795
rect 355 9765 356 9795
rect 324 9764 356 9765
rect 324 9715 356 9716
rect 324 9685 325 9715
rect 325 9685 355 9715
rect 355 9685 356 9715
rect 324 9684 356 9685
rect 324 9635 356 9636
rect 324 9605 325 9635
rect 325 9605 355 9635
rect 355 9605 356 9635
rect 324 9604 356 9605
rect 324 9555 356 9556
rect 324 9525 325 9555
rect 325 9525 355 9555
rect 355 9525 356 9555
rect 324 9524 356 9525
rect 324 9475 356 9476
rect 324 9445 325 9475
rect 325 9445 355 9475
rect 355 9445 356 9475
rect 324 9444 356 9445
rect 324 9395 356 9396
rect 324 9365 325 9395
rect 325 9365 355 9395
rect 355 9365 356 9395
rect 324 9364 356 9365
rect 324 9315 356 9316
rect 324 9285 325 9315
rect 325 9285 355 9315
rect 355 9285 356 9315
rect 324 9284 356 9285
rect 324 9235 356 9236
rect 324 9205 325 9235
rect 325 9205 355 9235
rect 355 9205 356 9235
rect 324 9204 356 9205
rect 324 9155 356 9156
rect 324 9125 325 9155
rect 325 9125 355 9155
rect 355 9125 356 9155
rect 324 9124 356 9125
rect 324 9075 356 9076
rect 324 9045 325 9075
rect 325 9045 355 9075
rect 355 9045 356 9075
rect 324 9044 356 9045
rect 324 8995 356 8996
rect 324 8965 325 8995
rect 325 8965 355 8995
rect 355 8965 356 8995
rect 324 8964 356 8965
rect 324 8915 356 8916
rect 324 8885 325 8915
rect 325 8885 355 8915
rect 355 8885 356 8915
rect 324 8884 356 8885
rect 324 8835 356 8836
rect 324 8805 325 8835
rect 325 8805 355 8835
rect 355 8805 356 8835
rect 324 8804 356 8805
rect 324 8755 356 8756
rect 324 8725 325 8755
rect 325 8725 355 8755
rect 355 8725 356 8755
rect 324 8724 356 8725
rect 324 8675 356 8676
rect 324 8645 325 8675
rect 325 8645 355 8675
rect 355 8645 356 8675
rect 324 8644 356 8645
rect 324 8515 356 8516
rect 324 8485 325 8515
rect 325 8485 355 8515
rect 355 8485 356 8515
rect 324 8484 356 8485
rect 324 8355 356 8356
rect 324 8325 325 8355
rect 325 8325 355 8355
rect 355 8325 356 8355
rect 324 8324 356 8325
rect 324 8275 356 8276
rect 324 8245 325 8275
rect 325 8245 355 8275
rect 355 8245 356 8275
rect 324 8244 356 8245
rect 324 8195 356 8196
rect 324 8165 325 8195
rect 325 8165 355 8195
rect 355 8165 356 8195
rect 324 8164 356 8165
rect 324 8115 356 8116
rect 324 8085 325 8115
rect 325 8085 355 8115
rect 355 8085 356 8115
rect 324 8084 356 8085
rect 324 7955 356 7956
rect 324 7925 325 7955
rect 325 7925 355 7955
rect 355 7925 356 7955
rect 324 7924 356 7925
rect 324 7795 356 7796
rect 324 7765 325 7795
rect 325 7765 355 7795
rect 355 7765 356 7795
rect 324 7764 356 7765
rect 324 7715 356 7716
rect 324 7685 325 7715
rect 325 7685 355 7715
rect 355 7685 356 7715
rect 324 7684 356 7685
rect 324 7635 356 7636
rect 324 7605 325 7635
rect 325 7605 355 7635
rect 355 7605 356 7635
rect 324 7604 356 7605
rect 324 7555 356 7556
rect 324 7525 325 7555
rect 325 7525 355 7555
rect 355 7525 356 7555
rect 324 7524 356 7525
rect 324 7475 356 7476
rect 324 7445 325 7475
rect 325 7445 355 7475
rect 355 7445 356 7475
rect 324 7444 356 7445
rect 324 7395 356 7396
rect 324 7365 325 7395
rect 325 7365 355 7395
rect 355 7365 356 7395
rect 324 7364 356 7365
rect 324 7315 356 7316
rect 324 7285 325 7315
rect 325 7285 355 7315
rect 355 7285 356 7315
rect 324 7284 356 7285
rect 324 7235 356 7236
rect 324 7205 325 7235
rect 325 7205 355 7235
rect 355 7205 356 7235
rect 324 7204 356 7205
rect 324 7155 356 7156
rect 324 7125 325 7155
rect 325 7125 355 7155
rect 355 7125 356 7155
rect 324 7124 356 7125
rect 324 7075 356 7076
rect 324 7045 325 7075
rect 325 7045 355 7075
rect 355 7045 356 7075
rect 324 7044 356 7045
rect 324 6995 356 6996
rect 324 6965 325 6995
rect 325 6965 355 6995
rect 355 6965 356 6995
rect 324 6964 356 6965
rect 324 6915 356 6916
rect 324 6885 325 6915
rect 325 6885 355 6915
rect 355 6885 356 6915
rect 324 6884 356 6885
rect 324 6835 356 6836
rect 324 6805 325 6835
rect 325 6805 355 6835
rect 355 6805 356 6835
rect 324 6804 356 6805
rect 324 6755 356 6756
rect 324 6725 325 6755
rect 325 6725 355 6755
rect 355 6725 356 6755
rect 324 6724 356 6725
rect 324 6675 356 6676
rect 324 6645 325 6675
rect 325 6645 355 6675
rect 355 6645 356 6675
rect 324 6644 356 6645
rect 324 6595 356 6596
rect 324 6565 325 6595
rect 325 6565 355 6595
rect 355 6565 356 6595
rect 324 6564 356 6565
rect 324 6515 356 6516
rect 324 6485 325 6515
rect 325 6485 355 6515
rect 355 6485 356 6515
rect 324 6484 356 6485
rect 324 6435 356 6436
rect 324 6405 325 6435
rect 325 6405 355 6435
rect 355 6405 356 6435
rect 324 6404 356 6405
rect 324 6355 356 6356
rect 324 6325 325 6355
rect 325 6325 355 6355
rect 355 6325 356 6355
rect 324 6324 356 6325
rect 324 6275 356 6276
rect 324 6245 325 6275
rect 325 6245 355 6275
rect 355 6245 356 6275
rect 324 6244 356 6245
rect 324 6195 356 6196
rect 324 6165 325 6195
rect 325 6165 355 6195
rect 355 6165 356 6195
rect 324 6164 356 6165
rect 324 6115 356 6116
rect 324 6085 325 6115
rect 325 6085 355 6115
rect 355 6085 356 6115
rect 324 6084 356 6085
rect 324 6035 356 6036
rect 324 6005 325 6035
rect 325 6005 355 6035
rect 355 6005 356 6035
rect 324 6004 356 6005
rect 324 5955 356 5956
rect 324 5925 325 5955
rect 325 5925 355 5955
rect 355 5925 356 5955
rect 324 5924 356 5925
rect 324 5875 356 5876
rect 324 5845 325 5875
rect 325 5845 355 5875
rect 355 5845 356 5875
rect 324 5844 356 5845
rect 324 5795 356 5796
rect 324 5765 325 5795
rect 325 5765 355 5795
rect 355 5765 356 5795
rect 324 5764 356 5765
rect 324 5715 356 5716
rect 324 5685 325 5715
rect 325 5685 355 5715
rect 355 5685 356 5715
rect 324 5684 356 5685
rect 324 5635 356 5636
rect 324 5605 325 5635
rect 325 5605 355 5635
rect 355 5605 356 5635
rect 324 5604 356 5605
rect 324 5555 356 5556
rect 324 5525 325 5555
rect 325 5525 355 5555
rect 355 5525 356 5555
rect 324 5524 356 5525
rect 324 5475 356 5476
rect 324 5445 325 5475
rect 325 5445 355 5475
rect 355 5445 356 5475
rect 324 5444 356 5445
rect 324 5395 356 5396
rect 324 5365 325 5395
rect 325 5365 355 5395
rect 355 5365 356 5395
rect 324 5364 356 5365
rect 324 5235 356 5236
rect 324 5205 325 5235
rect 325 5205 355 5235
rect 355 5205 356 5235
rect 324 5204 356 5205
rect 324 5075 356 5076
rect 324 5045 325 5075
rect 325 5045 355 5075
rect 355 5045 356 5075
rect 324 5044 356 5045
rect 324 4995 356 4996
rect 324 4965 325 4995
rect 325 4965 355 4995
rect 355 4965 356 4995
rect 324 4964 356 4965
rect 324 4915 356 4916
rect 324 4885 325 4915
rect 325 4885 355 4915
rect 355 4885 356 4915
rect 324 4884 356 4885
rect 324 4835 356 4836
rect 324 4805 325 4835
rect 325 4805 355 4835
rect 355 4805 356 4835
rect 324 4804 356 4805
rect 324 4755 356 4756
rect 324 4725 325 4755
rect 325 4725 355 4755
rect 355 4725 356 4755
rect 324 4724 356 4725
rect 324 4675 356 4676
rect 324 4645 325 4675
rect 325 4645 355 4675
rect 355 4645 356 4675
rect 324 4644 356 4645
rect 324 4595 356 4596
rect 324 4565 325 4595
rect 325 4565 355 4595
rect 355 4565 356 4595
rect 324 4564 356 4565
rect 324 4515 356 4516
rect 324 4485 325 4515
rect 325 4485 355 4515
rect 355 4485 356 4515
rect 324 4484 356 4485
rect 324 4435 356 4436
rect 324 4405 325 4435
rect 325 4405 355 4435
rect 355 4405 356 4435
rect 324 4404 356 4405
rect 324 4355 356 4356
rect 324 4325 325 4355
rect 325 4325 355 4355
rect 355 4325 356 4355
rect 324 4324 356 4325
rect 324 4275 356 4276
rect 324 4245 325 4275
rect 325 4245 355 4275
rect 355 4245 356 4275
rect 324 4244 356 4245
rect 324 4195 356 4196
rect 324 4165 325 4195
rect 325 4165 355 4195
rect 355 4165 356 4195
rect 324 4164 356 4165
rect 324 4115 356 4116
rect 324 4085 325 4115
rect 325 4085 355 4115
rect 355 4085 356 4115
rect 324 4084 356 4085
rect 324 4035 356 4036
rect 324 4005 325 4035
rect 325 4005 355 4035
rect 355 4005 356 4035
rect 324 4004 356 4005
rect 324 3955 356 3956
rect 324 3925 325 3955
rect 325 3925 355 3955
rect 355 3925 356 3955
rect 324 3924 356 3925
rect 324 3875 356 3876
rect 324 3845 325 3875
rect 325 3845 355 3875
rect 355 3845 356 3875
rect 324 3844 356 3845
rect 324 3795 356 3796
rect 324 3765 325 3795
rect 325 3765 355 3795
rect 355 3765 356 3795
rect 324 3764 356 3765
rect 324 3715 356 3716
rect 324 3685 325 3715
rect 325 3685 355 3715
rect 355 3685 356 3715
rect 324 3684 356 3685
rect 324 3635 356 3636
rect 324 3605 325 3635
rect 325 3605 355 3635
rect 355 3605 356 3635
rect 324 3604 356 3605
rect 324 3555 356 3556
rect 324 3525 325 3555
rect 325 3525 355 3555
rect 355 3525 356 3555
rect 324 3524 356 3525
rect 324 3475 356 3476
rect 324 3445 325 3475
rect 325 3445 355 3475
rect 355 3445 356 3475
rect 324 3444 356 3445
rect 324 3395 356 3396
rect 324 3365 325 3395
rect 325 3365 355 3395
rect 355 3365 356 3395
rect 324 3364 356 3365
rect 324 3315 356 3316
rect 324 3285 325 3315
rect 325 3285 355 3315
rect 355 3285 356 3315
rect 324 3284 356 3285
rect 324 3235 356 3236
rect 324 3205 325 3235
rect 325 3205 355 3235
rect 355 3205 356 3235
rect 324 3204 356 3205
rect 324 3155 356 3156
rect 324 3125 325 3155
rect 325 3125 355 3155
rect 355 3125 356 3155
rect 324 3124 356 3125
rect 324 3075 356 3076
rect 324 3045 325 3075
rect 325 3045 355 3075
rect 355 3045 356 3075
rect 324 3044 356 3045
rect 324 2995 356 2996
rect 324 2965 325 2995
rect 325 2965 355 2995
rect 355 2965 356 2995
rect 324 2964 356 2965
rect 324 2915 356 2916
rect 324 2885 325 2915
rect 325 2885 355 2915
rect 355 2885 356 2915
rect 324 2884 356 2885
rect 324 2835 356 2836
rect 324 2805 325 2835
rect 325 2805 355 2835
rect 355 2805 356 2835
rect 324 2804 356 2805
rect 324 2755 356 2756
rect 324 2725 325 2755
rect 325 2725 355 2755
rect 355 2725 356 2755
rect 324 2724 356 2725
rect 324 2675 356 2676
rect 324 2645 325 2675
rect 325 2645 355 2675
rect 355 2645 356 2675
rect 324 2644 356 2645
rect 324 2595 356 2596
rect 324 2565 325 2595
rect 325 2565 355 2595
rect 355 2565 356 2595
rect 324 2564 356 2565
rect 324 2515 356 2516
rect 324 2485 325 2515
rect 325 2485 355 2515
rect 355 2485 356 2515
rect 324 2484 356 2485
rect 324 2435 356 2436
rect 324 2405 325 2435
rect 325 2405 355 2435
rect 355 2405 356 2435
rect 324 2404 356 2405
rect 324 2355 356 2356
rect 324 2325 325 2355
rect 325 2325 355 2355
rect 355 2325 356 2355
rect 324 2324 356 2325
rect 324 2275 356 2276
rect 324 2245 325 2275
rect 325 2245 355 2275
rect 355 2245 356 2275
rect 324 2244 356 2245
rect 324 2195 356 2196
rect 324 2165 325 2195
rect 325 2165 355 2195
rect 355 2165 356 2195
rect 324 2164 356 2165
rect 324 2115 356 2116
rect 324 2085 325 2115
rect 325 2085 355 2115
rect 355 2085 356 2115
rect 324 2084 356 2085
rect 324 2035 356 2036
rect 324 2005 325 2035
rect 325 2005 355 2035
rect 355 2005 356 2035
rect 324 2004 356 2005
rect 324 1955 356 1956
rect 324 1925 325 1955
rect 325 1925 355 1955
rect 355 1925 356 1955
rect 324 1924 356 1925
rect 324 1875 356 1876
rect 324 1845 325 1875
rect 325 1845 355 1875
rect 355 1845 356 1875
rect 324 1844 356 1845
rect 324 1795 356 1796
rect 324 1765 325 1795
rect 325 1765 355 1795
rect 355 1765 356 1795
rect 324 1764 356 1765
rect 324 1715 356 1716
rect 324 1685 325 1715
rect 325 1685 355 1715
rect 355 1685 356 1715
rect 324 1684 356 1685
rect 324 1635 356 1636
rect 324 1605 325 1635
rect 325 1605 355 1635
rect 355 1605 356 1635
rect 324 1604 356 1605
rect 324 1555 356 1556
rect 324 1525 325 1555
rect 325 1525 355 1555
rect 355 1525 356 1555
rect 324 1524 356 1525
rect 324 1475 356 1476
rect 324 1445 325 1475
rect 325 1445 355 1475
rect 355 1445 356 1475
rect 324 1444 356 1445
rect 324 1395 356 1396
rect 324 1365 325 1395
rect 325 1365 355 1395
rect 355 1365 356 1395
rect 324 1364 356 1365
rect 324 1315 356 1316
rect 324 1285 325 1315
rect 325 1285 355 1315
rect 355 1285 356 1315
rect 324 1284 356 1285
rect 324 1235 356 1236
rect 324 1205 325 1235
rect 325 1205 355 1235
rect 355 1205 356 1235
rect 324 1204 356 1205
rect 324 1155 356 1156
rect 324 1125 325 1155
rect 325 1125 355 1155
rect 355 1125 356 1155
rect 324 1124 356 1125
rect 324 1075 356 1076
rect 324 1045 325 1075
rect 325 1045 355 1075
rect 355 1045 356 1075
rect 324 1044 356 1045
rect 324 995 356 996
rect 324 965 325 995
rect 325 965 355 995
rect 355 965 356 995
rect 324 964 356 965
rect 324 915 356 916
rect 324 885 325 915
rect 325 885 355 915
rect 355 885 356 915
rect 324 884 356 885
rect 324 835 356 836
rect 324 805 325 835
rect 325 805 355 835
rect 355 805 356 835
rect 324 804 356 805
rect 324 755 356 756
rect 324 725 325 755
rect 325 725 355 755
rect 355 725 356 755
rect 324 724 356 725
rect 324 675 356 676
rect 324 645 325 675
rect 325 645 355 675
rect 355 645 356 675
rect 324 644 356 645
rect 324 595 356 596
rect 324 565 325 595
rect 325 565 355 595
rect 355 565 356 595
rect 324 564 356 565
rect 324 515 356 516
rect 324 485 325 515
rect 325 485 355 515
rect 355 485 356 515
rect 324 484 356 485
rect 164 244 196 436
rect 404 9844 436 9876
rect 404 6564 436 6596
rect 484 15955 516 15956
rect 484 15925 485 15955
rect 485 15925 515 15955
rect 515 15925 516 15955
rect 484 15924 516 15925
rect 484 15875 516 15876
rect 484 15845 485 15875
rect 485 15845 515 15875
rect 515 15845 516 15875
rect 484 15844 516 15845
rect 484 15795 516 15796
rect 484 15765 485 15795
rect 485 15765 515 15795
rect 515 15765 516 15795
rect 484 15764 516 15765
rect 484 15715 516 15716
rect 484 15685 485 15715
rect 485 15685 515 15715
rect 515 15685 516 15715
rect 484 15684 516 15685
rect 484 15635 516 15636
rect 484 15605 485 15635
rect 485 15605 515 15635
rect 515 15605 516 15635
rect 484 15604 516 15605
rect 484 15555 516 15556
rect 484 15525 485 15555
rect 485 15525 515 15555
rect 515 15525 516 15555
rect 484 15524 516 15525
rect 484 15475 516 15476
rect 484 15445 485 15475
rect 485 15445 515 15475
rect 515 15445 516 15475
rect 484 15444 516 15445
rect 484 15395 516 15396
rect 484 15365 485 15395
rect 485 15365 515 15395
rect 515 15365 516 15395
rect 484 15364 516 15365
rect 484 15315 516 15316
rect 484 15285 485 15315
rect 485 15285 515 15315
rect 515 15285 516 15315
rect 484 15284 516 15285
rect 484 15235 516 15236
rect 484 15205 485 15235
rect 485 15205 515 15235
rect 515 15205 516 15235
rect 484 15204 516 15205
rect 484 15155 516 15156
rect 484 15125 485 15155
rect 485 15125 515 15155
rect 515 15125 516 15155
rect 484 15124 516 15125
rect 484 15075 516 15076
rect 484 15045 485 15075
rect 485 15045 515 15075
rect 515 15045 516 15075
rect 484 15044 516 15045
rect 484 14995 516 14996
rect 484 14965 485 14995
rect 485 14965 515 14995
rect 515 14965 516 14995
rect 484 14964 516 14965
rect 484 14915 516 14916
rect 484 14885 485 14915
rect 485 14885 515 14915
rect 515 14885 516 14915
rect 484 14884 516 14885
rect 484 14835 516 14836
rect 484 14805 485 14835
rect 485 14805 515 14835
rect 515 14805 516 14835
rect 484 14804 516 14805
rect 484 14755 516 14756
rect 484 14725 485 14755
rect 485 14725 515 14755
rect 515 14725 516 14755
rect 484 14724 516 14725
rect 484 14675 516 14676
rect 484 14645 485 14675
rect 485 14645 515 14675
rect 515 14645 516 14675
rect 484 14644 516 14645
rect 484 14595 516 14596
rect 484 14565 485 14595
rect 485 14565 515 14595
rect 515 14565 516 14595
rect 484 14564 516 14565
rect 484 14515 516 14516
rect 484 14485 485 14515
rect 485 14485 515 14515
rect 515 14485 516 14515
rect 484 14484 516 14485
rect 484 14435 516 14436
rect 484 14405 485 14435
rect 485 14405 515 14435
rect 515 14405 516 14435
rect 484 14404 516 14405
rect 484 14355 516 14356
rect 484 14325 485 14355
rect 485 14325 515 14355
rect 515 14325 516 14355
rect 484 14324 516 14325
rect 484 14275 516 14276
rect 484 14245 485 14275
rect 485 14245 515 14275
rect 515 14245 516 14275
rect 484 14244 516 14245
rect 484 14195 516 14196
rect 484 14165 485 14195
rect 485 14165 515 14195
rect 515 14165 516 14195
rect 484 14164 516 14165
rect 484 14115 516 14116
rect 484 14085 485 14115
rect 485 14085 515 14115
rect 515 14085 516 14115
rect 484 14084 516 14085
rect 484 14035 516 14036
rect 484 14005 485 14035
rect 485 14005 515 14035
rect 515 14005 516 14035
rect 484 14004 516 14005
rect 484 13955 516 13956
rect 484 13925 485 13955
rect 485 13925 515 13955
rect 515 13925 516 13955
rect 484 13924 516 13925
rect 484 13875 516 13876
rect 484 13845 485 13875
rect 485 13845 515 13875
rect 515 13845 516 13875
rect 484 13844 516 13845
rect 484 13795 516 13796
rect 484 13765 485 13795
rect 485 13765 515 13795
rect 515 13765 516 13795
rect 484 13764 516 13765
rect 484 13715 516 13716
rect 484 13685 485 13715
rect 485 13685 515 13715
rect 515 13685 516 13715
rect 484 13684 516 13685
rect 484 13635 516 13636
rect 484 13605 485 13635
rect 485 13605 515 13635
rect 515 13605 516 13635
rect 484 13604 516 13605
rect 484 13555 516 13556
rect 484 13525 485 13555
rect 485 13525 515 13555
rect 515 13525 516 13555
rect 484 13524 516 13525
rect 484 13475 516 13476
rect 484 13445 485 13475
rect 485 13445 515 13475
rect 515 13445 516 13475
rect 484 13444 516 13445
rect 484 13395 516 13396
rect 484 13365 485 13395
rect 485 13365 515 13395
rect 515 13365 516 13395
rect 484 13364 516 13365
rect 484 13315 516 13316
rect 484 13285 485 13315
rect 485 13285 515 13315
rect 515 13285 516 13315
rect 484 13284 516 13285
rect 484 13235 516 13236
rect 484 13205 485 13235
rect 485 13205 515 13235
rect 515 13205 516 13235
rect 484 13204 516 13205
rect 484 13155 516 13156
rect 484 13125 485 13155
rect 485 13125 515 13155
rect 515 13125 516 13155
rect 484 13124 516 13125
rect 484 13075 516 13076
rect 484 13045 485 13075
rect 485 13045 515 13075
rect 515 13045 516 13075
rect 484 13044 516 13045
rect 484 12995 516 12996
rect 484 12965 485 12995
rect 485 12965 515 12995
rect 515 12965 516 12995
rect 484 12964 516 12965
rect 484 12915 516 12916
rect 484 12885 485 12915
rect 485 12885 515 12915
rect 515 12885 516 12915
rect 484 12884 516 12885
rect 484 12835 516 12836
rect 484 12805 485 12835
rect 485 12805 515 12835
rect 515 12805 516 12835
rect 484 12804 516 12805
rect 484 12755 516 12756
rect 484 12725 485 12755
rect 485 12725 515 12755
rect 515 12725 516 12755
rect 484 12724 516 12725
rect 484 12675 516 12676
rect 484 12645 485 12675
rect 485 12645 515 12675
rect 515 12645 516 12675
rect 484 12644 516 12645
rect 484 12595 516 12596
rect 484 12565 485 12595
rect 485 12565 515 12595
rect 515 12565 516 12595
rect 484 12564 516 12565
rect 484 12515 516 12516
rect 484 12485 485 12515
rect 485 12485 515 12515
rect 515 12485 516 12515
rect 484 12484 516 12485
rect 484 12435 516 12436
rect 484 12405 485 12435
rect 485 12405 515 12435
rect 515 12405 516 12435
rect 484 12404 516 12405
rect 484 12355 516 12356
rect 484 12325 485 12355
rect 485 12325 515 12355
rect 515 12325 516 12355
rect 484 12324 516 12325
rect 484 12275 516 12276
rect 484 12245 485 12275
rect 485 12245 515 12275
rect 515 12245 516 12275
rect 484 12244 516 12245
rect 484 12195 516 12196
rect 484 12165 485 12195
rect 485 12165 515 12195
rect 515 12165 516 12195
rect 484 12164 516 12165
rect 484 12115 516 12116
rect 484 12085 485 12115
rect 485 12085 515 12115
rect 515 12085 516 12115
rect 484 12084 516 12085
rect 484 12035 516 12036
rect 484 12005 485 12035
rect 485 12005 515 12035
rect 515 12005 516 12035
rect 484 12004 516 12005
rect 484 11955 516 11956
rect 484 11925 485 11955
rect 485 11925 515 11955
rect 515 11925 516 11955
rect 484 11924 516 11925
rect 484 11875 516 11876
rect 484 11845 485 11875
rect 485 11845 515 11875
rect 515 11845 516 11875
rect 484 11844 516 11845
rect 484 11795 516 11796
rect 484 11765 485 11795
rect 485 11765 515 11795
rect 515 11765 516 11795
rect 484 11764 516 11765
rect 484 11715 516 11716
rect 484 11685 485 11715
rect 485 11685 515 11715
rect 515 11685 516 11715
rect 484 11684 516 11685
rect 484 11635 516 11636
rect 484 11605 485 11635
rect 485 11605 515 11635
rect 515 11605 516 11635
rect 484 11604 516 11605
rect 484 11555 516 11556
rect 484 11525 485 11555
rect 485 11525 515 11555
rect 515 11525 516 11555
rect 484 11524 516 11525
rect 484 11475 516 11476
rect 484 11445 485 11475
rect 485 11445 515 11475
rect 515 11445 516 11475
rect 484 11444 516 11445
rect 484 11395 516 11396
rect 484 11365 485 11395
rect 485 11365 515 11395
rect 515 11365 516 11395
rect 484 11364 516 11365
rect 484 11235 516 11236
rect 484 11205 485 11235
rect 485 11205 515 11235
rect 515 11205 516 11235
rect 484 11204 516 11205
rect 484 11075 516 11076
rect 484 11045 485 11075
rect 485 11045 515 11075
rect 515 11045 516 11075
rect 484 11044 516 11045
rect 484 10995 516 10996
rect 484 10965 485 10995
rect 485 10965 515 10995
rect 515 10965 516 10995
rect 484 10964 516 10965
rect 484 10915 516 10916
rect 484 10885 485 10915
rect 485 10885 515 10915
rect 515 10885 516 10915
rect 484 10884 516 10885
rect 484 10835 516 10836
rect 484 10805 485 10835
rect 485 10805 515 10835
rect 515 10805 516 10835
rect 484 10804 516 10805
rect 484 10755 516 10756
rect 484 10725 485 10755
rect 485 10725 515 10755
rect 515 10725 516 10755
rect 484 10724 516 10725
rect 484 10675 516 10676
rect 484 10645 485 10675
rect 485 10645 515 10675
rect 515 10645 516 10675
rect 484 10644 516 10645
rect 484 10595 516 10596
rect 484 10565 485 10595
rect 485 10565 515 10595
rect 515 10565 516 10595
rect 484 10564 516 10565
rect 484 10515 516 10516
rect 484 10485 485 10515
rect 485 10485 515 10515
rect 515 10485 516 10515
rect 484 10484 516 10485
rect 484 10435 516 10436
rect 484 10405 485 10435
rect 485 10405 515 10435
rect 515 10405 516 10435
rect 484 10404 516 10405
rect 484 10355 516 10356
rect 484 10325 485 10355
rect 485 10325 515 10355
rect 515 10325 516 10355
rect 484 10324 516 10325
rect 484 10275 516 10276
rect 484 10245 485 10275
rect 485 10245 515 10275
rect 515 10245 516 10275
rect 484 10244 516 10245
rect 484 10195 516 10196
rect 484 10165 485 10195
rect 485 10165 515 10195
rect 515 10165 516 10195
rect 484 10164 516 10165
rect 484 10115 516 10116
rect 484 10085 485 10115
rect 485 10085 515 10115
rect 515 10085 516 10115
rect 484 10084 516 10085
rect 484 10035 516 10036
rect 484 10005 485 10035
rect 485 10005 515 10035
rect 515 10005 516 10035
rect 484 10004 516 10005
rect 484 9955 516 9956
rect 484 9925 485 9955
rect 485 9925 515 9955
rect 515 9925 516 9955
rect 484 9924 516 9925
rect 484 9795 516 9796
rect 484 9765 485 9795
rect 485 9765 515 9795
rect 515 9765 516 9795
rect 484 9764 516 9765
rect 484 9715 516 9716
rect 484 9685 485 9715
rect 485 9685 515 9715
rect 515 9685 516 9715
rect 484 9684 516 9685
rect 484 9635 516 9636
rect 484 9605 485 9635
rect 485 9605 515 9635
rect 515 9605 516 9635
rect 484 9604 516 9605
rect 484 9555 516 9556
rect 484 9525 485 9555
rect 485 9525 515 9555
rect 515 9525 516 9555
rect 484 9524 516 9525
rect 484 9475 516 9476
rect 484 9445 485 9475
rect 485 9445 515 9475
rect 515 9445 516 9475
rect 484 9444 516 9445
rect 484 9395 516 9396
rect 484 9365 485 9395
rect 485 9365 515 9395
rect 515 9365 516 9395
rect 484 9364 516 9365
rect 484 9315 516 9316
rect 484 9285 485 9315
rect 485 9285 515 9315
rect 515 9285 516 9315
rect 484 9284 516 9285
rect 484 9235 516 9236
rect 484 9205 485 9235
rect 485 9205 515 9235
rect 515 9205 516 9235
rect 484 9204 516 9205
rect 484 9155 516 9156
rect 484 9125 485 9155
rect 485 9125 515 9155
rect 515 9125 516 9155
rect 484 9124 516 9125
rect 484 9075 516 9076
rect 484 9045 485 9075
rect 485 9045 515 9075
rect 515 9045 516 9075
rect 484 9044 516 9045
rect 484 8995 516 8996
rect 484 8965 485 8995
rect 485 8965 515 8995
rect 515 8965 516 8995
rect 484 8964 516 8965
rect 484 8915 516 8916
rect 484 8885 485 8915
rect 485 8885 515 8915
rect 515 8885 516 8915
rect 484 8884 516 8885
rect 484 8835 516 8836
rect 484 8805 485 8835
rect 485 8805 515 8835
rect 515 8805 516 8835
rect 484 8804 516 8805
rect 484 8755 516 8756
rect 484 8725 485 8755
rect 485 8725 515 8755
rect 515 8725 516 8755
rect 484 8724 516 8725
rect 484 8675 516 8676
rect 484 8645 485 8675
rect 485 8645 515 8675
rect 515 8645 516 8675
rect 484 8644 516 8645
rect 484 8515 516 8516
rect 484 8485 485 8515
rect 485 8485 515 8515
rect 515 8485 516 8515
rect 484 8484 516 8485
rect 484 8355 516 8356
rect 484 8325 485 8355
rect 485 8325 515 8355
rect 515 8325 516 8355
rect 484 8324 516 8325
rect 484 8275 516 8276
rect 484 8245 485 8275
rect 485 8245 515 8275
rect 515 8245 516 8275
rect 484 8244 516 8245
rect 484 8195 516 8196
rect 484 8165 485 8195
rect 485 8165 515 8195
rect 515 8165 516 8195
rect 484 8164 516 8165
rect 484 8115 516 8116
rect 484 8085 485 8115
rect 485 8085 515 8115
rect 515 8085 516 8115
rect 484 8084 516 8085
rect 484 7955 516 7956
rect 484 7925 485 7955
rect 485 7925 515 7955
rect 515 7925 516 7955
rect 484 7924 516 7925
rect 484 7795 516 7796
rect 484 7765 485 7795
rect 485 7765 515 7795
rect 515 7765 516 7795
rect 484 7764 516 7765
rect 484 7715 516 7716
rect 484 7685 485 7715
rect 485 7685 515 7715
rect 515 7685 516 7715
rect 484 7684 516 7685
rect 484 7635 516 7636
rect 484 7605 485 7635
rect 485 7605 515 7635
rect 515 7605 516 7635
rect 484 7604 516 7605
rect 484 7555 516 7556
rect 484 7525 485 7555
rect 485 7525 515 7555
rect 515 7525 516 7555
rect 484 7524 516 7525
rect 484 7475 516 7476
rect 484 7445 485 7475
rect 485 7445 515 7475
rect 515 7445 516 7475
rect 484 7444 516 7445
rect 484 7395 516 7396
rect 484 7365 485 7395
rect 485 7365 515 7395
rect 515 7365 516 7395
rect 484 7364 516 7365
rect 484 7315 516 7316
rect 484 7285 485 7315
rect 485 7285 515 7315
rect 515 7285 516 7315
rect 484 7284 516 7285
rect 484 7235 516 7236
rect 484 7205 485 7235
rect 485 7205 515 7235
rect 515 7205 516 7235
rect 484 7204 516 7205
rect 484 7155 516 7156
rect 484 7125 485 7155
rect 485 7125 515 7155
rect 515 7125 516 7155
rect 484 7124 516 7125
rect 484 7075 516 7076
rect 484 7045 485 7075
rect 485 7045 515 7075
rect 515 7045 516 7075
rect 484 7044 516 7045
rect 484 6995 516 6996
rect 484 6965 485 6995
rect 485 6965 515 6995
rect 515 6965 516 6995
rect 484 6964 516 6965
rect 484 6915 516 6916
rect 484 6885 485 6915
rect 485 6885 515 6915
rect 515 6885 516 6915
rect 484 6884 516 6885
rect 484 6835 516 6836
rect 484 6805 485 6835
rect 485 6805 515 6835
rect 515 6805 516 6835
rect 484 6804 516 6805
rect 484 6755 516 6756
rect 484 6725 485 6755
rect 485 6725 515 6755
rect 515 6725 516 6755
rect 484 6724 516 6725
rect 484 6675 516 6676
rect 484 6645 485 6675
rect 485 6645 515 6675
rect 515 6645 516 6675
rect 484 6644 516 6645
rect 484 6515 516 6516
rect 484 6485 485 6515
rect 485 6485 515 6515
rect 515 6485 516 6515
rect 484 6484 516 6485
rect 484 6435 516 6436
rect 484 6405 485 6435
rect 485 6405 515 6435
rect 515 6405 516 6435
rect 484 6404 516 6405
rect 484 6355 516 6356
rect 484 6325 485 6355
rect 485 6325 515 6355
rect 515 6325 516 6355
rect 484 6324 516 6325
rect 484 6275 516 6276
rect 484 6245 485 6275
rect 485 6245 515 6275
rect 515 6245 516 6275
rect 484 6244 516 6245
rect 484 6195 516 6196
rect 484 6165 485 6195
rect 485 6165 515 6195
rect 515 6165 516 6195
rect 484 6164 516 6165
rect 484 6115 516 6116
rect 484 6085 485 6115
rect 485 6085 515 6115
rect 515 6085 516 6115
rect 484 6084 516 6085
rect 484 6035 516 6036
rect 484 6005 485 6035
rect 485 6005 515 6035
rect 515 6005 516 6035
rect 484 6004 516 6005
rect 484 5955 516 5956
rect 484 5925 485 5955
rect 485 5925 515 5955
rect 515 5925 516 5955
rect 484 5924 516 5925
rect 484 5875 516 5876
rect 484 5845 485 5875
rect 485 5845 515 5875
rect 515 5845 516 5875
rect 484 5844 516 5845
rect 484 5795 516 5796
rect 484 5765 485 5795
rect 485 5765 515 5795
rect 515 5765 516 5795
rect 484 5764 516 5765
rect 484 5715 516 5716
rect 484 5685 485 5715
rect 485 5685 515 5715
rect 515 5685 516 5715
rect 484 5684 516 5685
rect 484 5635 516 5636
rect 484 5605 485 5635
rect 485 5605 515 5635
rect 515 5605 516 5635
rect 484 5604 516 5605
rect 484 5555 516 5556
rect 484 5525 485 5555
rect 485 5525 515 5555
rect 515 5525 516 5555
rect 484 5524 516 5525
rect 484 5475 516 5476
rect 484 5445 485 5475
rect 485 5445 515 5475
rect 515 5445 516 5475
rect 484 5444 516 5445
rect 484 5395 516 5396
rect 484 5365 485 5395
rect 485 5365 515 5395
rect 515 5365 516 5395
rect 484 5364 516 5365
rect 484 5235 516 5236
rect 484 5205 485 5235
rect 485 5205 515 5235
rect 515 5205 516 5235
rect 484 5204 516 5205
rect 484 5075 516 5076
rect 484 5045 485 5075
rect 485 5045 515 5075
rect 515 5045 516 5075
rect 484 5044 516 5045
rect 484 4995 516 4996
rect 484 4965 485 4995
rect 485 4965 515 4995
rect 515 4965 516 4995
rect 484 4964 516 4965
rect 484 4915 516 4916
rect 484 4885 485 4915
rect 485 4885 515 4915
rect 515 4885 516 4915
rect 484 4884 516 4885
rect 484 4835 516 4836
rect 484 4805 485 4835
rect 485 4805 515 4835
rect 515 4805 516 4835
rect 484 4804 516 4805
rect 484 4755 516 4756
rect 484 4725 485 4755
rect 485 4725 515 4755
rect 515 4725 516 4755
rect 484 4724 516 4725
rect 484 4675 516 4676
rect 484 4645 485 4675
rect 485 4645 515 4675
rect 515 4645 516 4675
rect 484 4644 516 4645
rect 484 4595 516 4596
rect 484 4565 485 4595
rect 485 4565 515 4595
rect 515 4565 516 4595
rect 484 4564 516 4565
rect 484 4515 516 4516
rect 484 4485 485 4515
rect 485 4485 515 4515
rect 515 4485 516 4515
rect 484 4484 516 4485
rect 484 4435 516 4436
rect 484 4405 485 4435
rect 485 4405 515 4435
rect 515 4405 516 4435
rect 484 4404 516 4405
rect 484 4355 516 4356
rect 484 4325 485 4355
rect 485 4325 515 4355
rect 515 4325 516 4355
rect 484 4324 516 4325
rect 484 4275 516 4276
rect 484 4245 485 4275
rect 485 4245 515 4275
rect 515 4245 516 4275
rect 484 4244 516 4245
rect 484 4195 516 4196
rect 484 4165 485 4195
rect 485 4165 515 4195
rect 515 4165 516 4195
rect 484 4164 516 4165
rect 484 4115 516 4116
rect 484 4085 485 4115
rect 485 4085 515 4115
rect 515 4085 516 4115
rect 484 4084 516 4085
rect 484 4035 516 4036
rect 484 4005 485 4035
rect 485 4005 515 4035
rect 515 4005 516 4035
rect 484 4004 516 4005
rect 484 3955 516 3956
rect 484 3925 485 3955
rect 485 3925 515 3955
rect 515 3925 516 3955
rect 484 3924 516 3925
rect 484 3875 516 3876
rect 484 3845 485 3875
rect 485 3845 515 3875
rect 515 3845 516 3875
rect 484 3844 516 3845
rect 484 3795 516 3796
rect 484 3765 485 3795
rect 485 3765 515 3795
rect 515 3765 516 3795
rect 484 3764 516 3765
rect 484 3715 516 3716
rect 484 3685 485 3715
rect 485 3685 515 3715
rect 515 3685 516 3715
rect 484 3684 516 3685
rect 484 3635 516 3636
rect 484 3605 485 3635
rect 485 3605 515 3635
rect 515 3605 516 3635
rect 484 3604 516 3605
rect 484 3555 516 3556
rect 484 3525 485 3555
rect 485 3525 515 3555
rect 515 3525 516 3555
rect 484 3524 516 3525
rect 484 3475 516 3476
rect 484 3445 485 3475
rect 485 3445 515 3475
rect 515 3445 516 3475
rect 484 3444 516 3445
rect 484 3395 516 3396
rect 484 3365 485 3395
rect 485 3365 515 3395
rect 515 3365 516 3395
rect 484 3364 516 3365
rect 484 3315 516 3316
rect 484 3285 485 3315
rect 485 3285 515 3315
rect 515 3285 516 3315
rect 484 3284 516 3285
rect 484 3235 516 3236
rect 484 3205 485 3235
rect 485 3205 515 3235
rect 515 3205 516 3235
rect 484 3204 516 3205
rect 484 3155 516 3156
rect 484 3125 485 3155
rect 485 3125 515 3155
rect 515 3125 516 3155
rect 484 3124 516 3125
rect 484 3075 516 3076
rect 484 3045 485 3075
rect 485 3045 515 3075
rect 515 3045 516 3075
rect 484 3044 516 3045
rect 484 2995 516 2996
rect 484 2965 485 2995
rect 485 2965 515 2995
rect 515 2965 516 2995
rect 484 2964 516 2965
rect 484 2915 516 2916
rect 484 2885 485 2915
rect 485 2885 515 2915
rect 515 2885 516 2915
rect 484 2884 516 2885
rect 484 2835 516 2836
rect 484 2805 485 2835
rect 485 2805 515 2835
rect 515 2805 516 2835
rect 484 2804 516 2805
rect 484 2755 516 2756
rect 484 2725 485 2755
rect 485 2725 515 2755
rect 515 2725 516 2755
rect 484 2724 516 2725
rect 484 2675 516 2676
rect 484 2645 485 2675
rect 485 2645 515 2675
rect 515 2645 516 2675
rect 484 2644 516 2645
rect 484 2595 516 2596
rect 484 2565 485 2595
rect 485 2565 515 2595
rect 515 2565 516 2595
rect 484 2564 516 2565
rect 484 2515 516 2516
rect 484 2485 485 2515
rect 485 2485 515 2515
rect 515 2485 516 2515
rect 484 2484 516 2485
rect 484 2435 516 2436
rect 484 2405 485 2435
rect 485 2405 515 2435
rect 515 2405 516 2435
rect 484 2404 516 2405
rect 484 2355 516 2356
rect 484 2325 485 2355
rect 485 2325 515 2355
rect 515 2325 516 2355
rect 484 2324 516 2325
rect 484 2275 516 2276
rect 484 2245 485 2275
rect 485 2245 515 2275
rect 515 2245 516 2275
rect 484 2244 516 2245
rect 484 2195 516 2196
rect 484 2165 485 2195
rect 485 2165 515 2195
rect 515 2165 516 2195
rect 484 2164 516 2165
rect 484 2115 516 2116
rect 484 2085 485 2115
rect 485 2085 515 2115
rect 515 2085 516 2115
rect 484 2084 516 2085
rect 484 2035 516 2036
rect 484 2005 485 2035
rect 485 2005 515 2035
rect 515 2005 516 2035
rect 484 2004 516 2005
rect 484 1955 516 1956
rect 484 1925 485 1955
rect 485 1925 515 1955
rect 515 1925 516 1955
rect 484 1924 516 1925
rect 484 1875 516 1876
rect 484 1845 485 1875
rect 485 1845 515 1875
rect 515 1845 516 1875
rect 484 1844 516 1845
rect 484 1795 516 1796
rect 484 1765 485 1795
rect 485 1765 515 1795
rect 515 1765 516 1795
rect 484 1764 516 1765
rect 484 1715 516 1716
rect 484 1685 485 1715
rect 485 1685 515 1715
rect 515 1685 516 1715
rect 484 1684 516 1685
rect 484 1635 516 1636
rect 484 1605 485 1635
rect 485 1605 515 1635
rect 515 1605 516 1635
rect 484 1604 516 1605
rect 484 1555 516 1556
rect 484 1525 485 1555
rect 485 1525 515 1555
rect 515 1525 516 1555
rect 484 1524 516 1525
rect 484 1475 516 1476
rect 484 1445 485 1475
rect 485 1445 515 1475
rect 515 1445 516 1475
rect 484 1444 516 1445
rect 484 1395 516 1396
rect 484 1365 485 1395
rect 485 1365 515 1395
rect 515 1365 516 1395
rect 484 1364 516 1365
rect 484 1315 516 1316
rect 484 1285 485 1315
rect 485 1285 515 1315
rect 515 1285 516 1315
rect 484 1284 516 1285
rect 484 1235 516 1236
rect 484 1205 485 1235
rect 485 1205 515 1235
rect 515 1205 516 1235
rect 484 1204 516 1205
rect 484 1155 516 1156
rect 484 1125 485 1155
rect 485 1125 515 1155
rect 515 1125 516 1155
rect 484 1124 516 1125
rect 484 1075 516 1076
rect 484 1045 485 1075
rect 485 1045 515 1075
rect 515 1045 516 1075
rect 484 1044 516 1045
rect 484 995 516 996
rect 484 965 485 995
rect 485 965 515 995
rect 515 965 516 995
rect 484 964 516 965
rect 484 915 516 916
rect 484 885 485 915
rect 485 885 515 915
rect 515 885 516 915
rect 484 884 516 885
rect 484 835 516 836
rect 484 805 485 835
rect 485 805 515 835
rect 515 805 516 835
rect 484 804 516 805
rect 484 755 516 756
rect 484 725 485 755
rect 485 725 515 755
rect 515 725 516 755
rect 484 724 516 725
rect 484 675 516 676
rect 484 645 485 675
rect 485 645 515 675
rect 515 645 516 675
rect 484 644 516 645
rect 484 595 516 596
rect 484 565 485 595
rect 485 565 515 595
rect 515 565 516 595
rect 484 564 516 565
rect 14484 15955 14516 15956
rect 14484 15925 14485 15955
rect 14485 15925 14515 15955
rect 14515 15925 14516 15955
rect 14484 15924 14516 15925
rect 14484 15875 14516 15876
rect 14484 15845 14485 15875
rect 14485 15845 14515 15875
rect 14515 15845 14516 15875
rect 14484 15844 14516 15845
rect 14484 15795 14516 15796
rect 14484 15765 14485 15795
rect 14485 15765 14515 15795
rect 14515 15765 14516 15795
rect 14484 15764 14516 15765
rect 14484 15715 14516 15716
rect 14484 15685 14485 15715
rect 14485 15685 14515 15715
rect 14515 15685 14516 15715
rect 14484 15684 14516 15685
rect 14484 15635 14516 15636
rect 14484 15605 14485 15635
rect 14485 15605 14515 15635
rect 14515 15605 14516 15635
rect 14484 15604 14516 15605
rect 14484 15555 14516 15556
rect 14484 15525 14485 15555
rect 14485 15525 14515 15555
rect 14515 15525 14516 15555
rect 14484 15524 14516 15525
rect 14484 15475 14516 15476
rect 14484 15445 14485 15475
rect 14485 15445 14515 15475
rect 14515 15445 14516 15475
rect 14484 15444 14516 15445
rect 14484 15395 14516 15396
rect 14484 15365 14485 15395
rect 14485 15365 14515 15395
rect 14515 15365 14516 15395
rect 14484 15364 14516 15365
rect 14484 15315 14516 15316
rect 14484 15285 14485 15315
rect 14485 15285 14515 15315
rect 14515 15285 14516 15315
rect 14484 15284 14516 15285
rect 14484 15235 14516 15236
rect 14484 15205 14485 15235
rect 14485 15205 14515 15235
rect 14515 15205 14516 15235
rect 14484 15204 14516 15205
rect 14484 15155 14516 15156
rect 14484 15125 14485 15155
rect 14485 15125 14515 15155
rect 14515 15125 14516 15155
rect 14484 15124 14516 15125
rect 14484 15075 14516 15076
rect 14484 15045 14485 15075
rect 14485 15045 14515 15075
rect 14515 15045 14516 15075
rect 14484 15044 14516 15045
rect 14484 14995 14516 14996
rect 14484 14965 14485 14995
rect 14485 14965 14515 14995
rect 14515 14965 14516 14995
rect 14484 14964 14516 14965
rect 14484 14915 14516 14916
rect 14484 14885 14485 14915
rect 14485 14885 14515 14915
rect 14515 14885 14516 14915
rect 14484 14884 14516 14885
rect 14484 14835 14516 14836
rect 14484 14805 14485 14835
rect 14485 14805 14515 14835
rect 14515 14805 14516 14835
rect 14484 14804 14516 14805
rect 14484 14755 14516 14756
rect 14484 14725 14485 14755
rect 14485 14725 14515 14755
rect 14515 14725 14516 14755
rect 14484 14724 14516 14725
rect 14484 14675 14516 14676
rect 14484 14645 14485 14675
rect 14485 14645 14515 14675
rect 14515 14645 14516 14675
rect 14484 14644 14516 14645
rect 14484 14515 14516 14516
rect 14484 14485 14485 14515
rect 14485 14485 14515 14515
rect 14515 14485 14516 14515
rect 14484 14484 14516 14485
rect 14484 14355 14516 14356
rect 14484 14325 14485 14355
rect 14485 14325 14515 14355
rect 14515 14325 14516 14355
rect 14484 14324 14516 14325
rect 14484 14275 14516 14276
rect 14484 14245 14485 14275
rect 14485 14245 14515 14275
rect 14515 14245 14516 14275
rect 14484 14244 14516 14245
rect 14484 14195 14516 14196
rect 14484 14165 14485 14195
rect 14485 14165 14515 14195
rect 14515 14165 14516 14195
rect 14484 14164 14516 14165
rect 14484 14115 14516 14116
rect 14484 14085 14485 14115
rect 14485 14085 14515 14115
rect 14515 14085 14516 14115
rect 14484 14084 14516 14085
rect 14484 14035 14516 14036
rect 14484 14005 14485 14035
rect 14485 14005 14515 14035
rect 14515 14005 14516 14035
rect 14484 14004 14516 14005
rect 14484 13955 14516 13956
rect 14484 13925 14485 13955
rect 14485 13925 14515 13955
rect 14515 13925 14516 13955
rect 14484 13924 14516 13925
rect 14484 13875 14516 13876
rect 14484 13845 14485 13875
rect 14485 13845 14515 13875
rect 14515 13845 14516 13875
rect 14484 13844 14516 13845
rect 14484 13795 14516 13796
rect 14484 13765 14485 13795
rect 14485 13765 14515 13795
rect 14515 13765 14516 13795
rect 14484 13764 14516 13765
rect 14484 13715 14516 13716
rect 14484 13685 14485 13715
rect 14485 13685 14515 13715
rect 14515 13685 14516 13715
rect 14484 13684 14516 13685
rect 14484 13635 14516 13636
rect 14484 13605 14485 13635
rect 14485 13605 14515 13635
rect 14515 13605 14516 13635
rect 14484 13604 14516 13605
rect 14484 13555 14516 13556
rect 14484 13525 14485 13555
rect 14485 13525 14515 13555
rect 14515 13525 14516 13555
rect 14484 13524 14516 13525
rect 14484 13475 14516 13476
rect 14484 13445 14485 13475
rect 14485 13445 14515 13475
rect 14515 13445 14516 13475
rect 14484 13444 14516 13445
rect 14484 13395 14516 13396
rect 14484 13365 14485 13395
rect 14485 13365 14515 13395
rect 14515 13365 14516 13395
rect 14484 13364 14516 13365
rect 14484 13315 14516 13316
rect 14484 13285 14485 13315
rect 14485 13285 14515 13315
rect 14515 13285 14516 13315
rect 14484 13284 14516 13285
rect 14484 13235 14516 13236
rect 14484 13205 14485 13235
rect 14485 13205 14515 13235
rect 14515 13205 14516 13235
rect 14484 13204 14516 13205
rect 14484 13075 14516 13076
rect 14484 13045 14485 13075
rect 14485 13045 14515 13075
rect 14515 13045 14516 13075
rect 14484 13044 14516 13045
rect 14484 12995 14516 12996
rect 14484 12965 14485 12995
rect 14485 12965 14515 12995
rect 14515 12965 14516 12995
rect 14484 12964 14516 12965
rect 14484 12915 14516 12916
rect 14484 12885 14485 12915
rect 14485 12885 14515 12915
rect 14515 12885 14516 12915
rect 14484 12884 14516 12885
rect 14484 12835 14516 12836
rect 14484 12805 14485 12835
rect 14485 12805 14515 12835
rect 14515 12805 14516 12835
rect 14484 12804 14516 12805
rect 14484 12755 14516 12756
rect 14484 12725 14485 12755
rect 14485 12725 14515 12755
rect 14515 12725 14516 12755
rect 14484 12724 14516 12725
rect 14484 12675 14516 12676
rect 14484 12645 14485 12675
rect 14485 12645 14515 12675
rect 14515 12645 14516 12675
rect 14484 12644 14516 12645
rect 14484 12595 14516 12596
rect 14484 12565 14485 12595
rect 14485 12565 14515 12595
rect 14515 12565 14516 12595
rect 14484 12564 14516 12565
rect 14484 12515 14516 12516
rect 14484 12485 14485 12515
rect 14485 12485 14515 12515
rect 14515 12485 14516 12515
rect 14484 12484 14516 12485
rect 14484 12435 14516 12436
rect 14484 12405 14485 12435
rect 14485 12405 14515 12435
rect 14515 12405 14516 12435
rect 14484 12404 14516 12405
rect 14484 12355 14516 12356
rect 14484 12325 14485 12355
rect 14485 12325 14515 12355
rect 14515 12325 14516 12355
rect 14484 12324 14516 12325
rect 14484 12275 14516 12276
rect 14484 12245 14485 12275
rect 14485 12245 14515 12275
rect 14515 12245 14516 12275
rect 14484 12244 14516 12245
rect 14484 12195 14516 12196
rect 14484 12165 14485 12195
rect 14485 12165 14515 12195
rect 14515 12165 14516 12195
rect 14484 12164 14516 12165
rect 14484 12115 14516 12116
rect 14484 12085 14485 12115
rect 14485 12085 14515 12115
rect 14515 12085 14516 12115
rect 14484 12084 14516 12085
rect 14484 12035 14516 12036
rect 14484 12005 14485 12035
rect 14485 12005 14515 12035
rect 14515 12005 14516 12035
rect 14484 12004 14516 12005
rect 14484 11955 14516 11956
rect 14484 11925 14485 11955
rect 14485 11925 14515 11955
rect 14515 11925 14516 11955
rect 14484 11924 14516 11925
rect 14484 11795 14516 11796
rect 14484 11765 14485 11795
rect 14485 11765 14515 11795
rect 14515 11765 14516 11795
rect 14484 11764 14516 11765
rect 14484 11635 14516 11636
rect 14484 11605 14485 11635
rect 14485 11605 14515 11635
rect 14515 11605 14516 11635
rect 14484 11604 14516 11605
rect 14484 11555 14516 11556
rect 14484 11525 14485 11555
rect 14485 11525 14515 11555
rect 14515 11525 14516 11555
rect 14484 11524 14516 11525
rect 14484 11475 14516 11476
rect 14484 11445 14485 11475
rect 14485 11445 14515 11475
rect 14515 11445 14516 11475
rect 14484 11444 14516 11445
rect 14484 11395 14516 11396
rect 14484 11365 14485 11395
rect 14485 11365 14515 11395
rect 14515 11365 14516 11395
rect 14484 11364 14516 11365
rect 14484 11315 14516 11316
rect 14484 11285 14485 11315
rect 14485 11285 14515 11315
rect 14515 11285 14516 11315
rect 14484 11284 14516 11285
rect 14484 11235 14516 11236
rect 14484 11205 14485 11235
rect 14485 11205 14515 11235
rect 14515 11205 14516 11235
rect 14484 11204 14516 11205
rect 14484 11155 14516 11156
rect 14484 11125 14485 11155
rect 14485 11125 14515 11155
rect 14515 11125 14516 11155
rect 14484 11124 14516 11125
rect 14484 11075 14516 11076
rect 14484 11045 14485 11075
rect 14485 11045 14515 11075
rect 14515 11045 14516 11075
rect 14484 11044 14516 11045
rect 14484 10995 14516 10996
rect 14484 10965 14485 10995
rect 14485 10965 14515 10995
rect 14515 10965 14516 10995
rect 14484 10964 14516 10965
rect 14484 10915 14516 10916
rect 14484 10885 14485 10915
rect 14485 10885 14515 10915
rect 14515 10885 14516 10915
rect 14484 10884 14516 10885
rect 14484 10835 14516 10836
rect 14484 10805 14485 10835
rect 14485 10805 14515 10835
rect 14515 10805 14516 10835
rect 14484 10804 14516 10805
rect 14484 10755 14516 10756
rect 14484 10725 14485 10755
rect 14485 10725 14515 10755
rect 14515 10725 14516 10755
rect 14484 10724 14516 10725
rect 14484 10675 14516 10676
rect 14484 10645 14485 10675
rect 14485 10645 14515 10675
rect 14515 10645 14516 10675
rect 14484 10644 14516 10645
rect 14484 10595 14516 10596
rect 14484 10565 14485 10595
rect 14485 10565 14515 10595
rect 14515 10565 14516 10595
rect 14484 10564 14516 10565
rect 14484 10515 14516 10516
rect 14484 10485 14485 10515
rect 14485 10485 14515 10515
rect 14515 10485 14516 10515
rect 14484 10484 14516 10485
rect 14484 10435 14516 10436
rect 14484 10405 14485 10435
rect 14485 10405 14515 10435
rect 14515 10405 14516 10435
rect 14484 10404 14516 10405
rect 14484 10355 14516 10356
rect 14484 10325 14485 10355
rect 14485 10325 14515 10355
rect 14515 10325 14516 10355
rect 14484 10324 14516 10325
rect 14484 10275 14516 10276
rect 14484 10245 14485 10275
rect 14485 10245 14515 10275
rect 14515 10245 14516 10275
rect 14484 10244 14516 10245
rect 14484 10195 14516 10196
rect 14484 10165 14485 10195
rect 14485 10165 14515 10195
rect 14515 10165 14516 10195
rect 14484 10164 14516 10165
rect 14484 10115 14516 10116
rect 14484 10085 14485 10115
rect 14485 10085 14515 10115
rect 14515 10085 14516 10115
rect 14484 10084 14516 10085
rect 14484 10035 14516 10036
rect 14484 10005 14485 10035
rect 14485 10005 14515 10035
rect 14515 10005 14516 10035
rect 14484 10004 14516 10005
rect 14484 9955 14516 9956
rect 14484 9925 14485 9955
rect 14485 9925 14515 9955
rect 14515 9925 14516 9955
rect 14484 9924 14516 9925
rect 14484 9875 14516 9876
rect 14484 9845 14485 9875
rect 14485 9845 14515 9875
rect 14515 9845 14516 9875
rect 14484 9844 14516 9845
rect 14484 9795 14516 9796
rect 14484 9765 14485 9795
rect 14485 9765 14515 9795
rect 14515 9765 14516 9795
rect 14484 9764 14516 9765
rect 14484 9715 14516 9716
rect 14484 9685 14485 9715
rect 14485 9685 14515 9715
rect 14515 9685 14516 9715
rect 14484 9684 14516 9685
rect 14484 9635 14516 9636
rect 14484 9605 14485 9635
rect 14485 9605 14515 9635
rect 14515 9605 14516 9635
rect 14484 9604 14516 9605
rect 14484 9555 14516 9556
rect 14484 9525 14485 9555
rect 14485 9525 14515 9555
rect 14515 9525 14516 9555
rect 14484 9524 14516 9525
rect 14484 9475 14516 9476
rect 14484 9445 14485 9475
rect 14485 9445 14515 9475
rect 14515 9445 14516 9475
rect 14484 9444 14516 9445
rect 14484 9395 14516 9396
rect 14484 9365 14485 9395
rect 14485 9365 14515 9395
rect 14515 9365 14516 9395
rect 14484 9364 14516 9365
rect 14484 9315 14516 9316
rect 14484 9285 14485 9315
rect 14485 9285 14515 9315
rect 14515 9285 14516 9315
rect 14484 9284 14516 9285
rect 14484 9235 14516 9236
rect 14484 9205 14485 9235
rect 14485 9205 14515 9235
rect 14515 9205 14516 9235
rect 14484 9204 14516 9205
rect 14484 9155 14516 9156
rect 14484 9125 14485 9155
rect 14485 9125 14515 9155
rect 14515 9125 14516 9155
rect 14484 9124 14516 9125
rect 14484 9075 14516 9076
rect 14484 9045 14485 9075
rect 14485 9045 14515 9075
rect 14515 9045 14516 9075
rect 14484 9044 14516 9045
rect 14484 8995 14516 8996
rect 14484 8965 14485 8995
rect 14485 8965 14515 8995
rect 14515 8965 14516 8995
rect 14484 8964 14516 8965
rect 14484 8915 14516 8916
rect 14484 8885 14485 8915
rect 14485 8885 14515 8915
rect 14515 8885 14516 8915
rect 14484 8884 14516 8885
rect 14484 8835 14516 8836
rect 14484 8805 14485 8835
rect 14485 8805 14515 8835
rect 14515 8805 14516 8835
rect 14484 8804 14516 8805
rect 14484 8755 14516 8756
rect 14484 8725 14485 8755
rect 14485 8725 14515 8755
rect 14515 8725 14516 8755
rect 14484 8724 14516 8725
rect 14484 8675 14516 8676
rect 14484 8645 14485 8675
rect 14485 8645 14515 8675
rect 14515 8645 14516 8675
rect 14484 8644 14516 8645
rect 14484 8595 14516 8596
rect 14484 8565 14485 8595
rect 14485 8565 14515 8595
rect 14515 8565 14516 8595
rect 14484 8564 14516 8565
rect 14484 8515 14516 8516
rect 14484 8485 14485 8515
rect 14485 8485 14515 8515
rect 14515 8485 14516 8515
rect 14484 8484 14516 8485
rect 14484 8435 14516 8436
rect 14484 8405 14485 8435
rect 14485 8405 14515 8435
rect 14515 8405 14516 8435
rect 14484 8404 14516 8405
rect 14484 8355 14516 8356
rect 14484 8325 14485 8355
rect 14485 8325 14515 8355
rect 14515 8325 14516 8355
rect 14484 8324 14516 8325
rect 14484 8275 14516 8276
rect 14484 8245 14485 8275
rect 14485 8245 14515 8275
rect 14515 8245 14516 8275
rect 14484 8244 14516 8245
rect 14484 8195 14516 8196
rect 14484 8165 14485 8195
rect 14485 8165 14515 8195
rect 14515 8165 14516 8195
rect 14484 8164 14516 8165
rect 14484 8115 14516 8116
rect 14484 8085 14485 8115
rect 14485 8085 14515 8115
rect 14515 8085 14516 8115
rect 14484 8084 14516 8085
rect 14484 8035 14516 8036
rect 14484 8005 14485 8035
rect 14485 8005 14515 8035
rect 14515 8005 14516 8035
rect 14484 8004 14516 8005
rect 14484 7955 14516 7956
rect 14484 7925 14485 7955
rect 14485 7925 14515 7955
rect 14515 7925 14516 7955
rect 14484 7924 14516 7925
rect 14484 7875 14516 7876
rect 14484 7845 14485 7875
rect 14485 7845 14515 7875
rect 14515 7845 14516 7875
rect 14484 7844 14516 7845
rect 14484 7795 14516 7796
rect 14484 7765 14485 7795
rect 14485 7765 14515 7795
rect 14515 7765 14516 7795
rect 14484 7764 14516 7765
rect 14484 7715 14516 7716
rect 14484 7685 14485 7715
rect 14485 7685 14515 7715
rect 14515 7685 14516 7715
rect 14484 7684 14516 7685
rect 14484 7635 14516 7636
rect 14484 7605 14485 7635
rect 14485 7605 14515 7635
rect 14515 7605 14516 7635
rect 14484 7604 14516 7605
rect 14484 7555 14516 7556
rect 14484 7525 14485 7555
rect 14485 7525 14515 7555
rect 14515 7525 14516 7555
rect 14484 7524 14516 7525
rect 14484 7475 14516 7476
rect 14484 7445 14485 7475
rect 14485 7445 14515 7475
rect 14515 7445 14516 7475
rect 14484 7444 14516 7445
rect 14484 7395 14516 7396
rect 14484 7365 14485 7395
rect 14485 7365 14515 7395
rect 14515 7365 14516 7395
rect 14484 7364 14516 7365
rect 14484 7315 14516 7316
rect 14484 7285 14485 7315
rect 14485 7285 14515 7315
rect 14515 7285 14516 7315
rect 14484 7284 14516 7285
rect 14484 7235 14516 7236
rect 14484 7205 14485 7235
rect 14485 7205 14515 7235
rect 14515 7205 14516 7235
rect 14484 7204 14516 7205
rect 14484 7155 14516 7156
rect 14484 7125 14485 7155
rect 14485 7125 14515 7155
rect 14515 7125 14516 7155
rect 14484 7124 14516 7125
rect 14484 7075 14516 7076
rect 14484 7045 14485 7075
rect 14485 7045 14515 7075
rect 14515 7045 14516 7075
rect 14484 7044 14516 7045
rect 14484 6995 14516 6996
rect 14484 6965 14485 6995
rect 14485 6965 14515 6995
rect 14515 6965 14516 6995
rect 14484 6964 14516 6965
rect 14484 6915 14516 6916
rect 14484 6885 14485 6915
rect 14485 6885 14515 6915
rect 14515 6885 14516 6915
rect 14484 6884 14516 6885
rect 14484 6835 14516 6836
rect 14484 6805 14485 6835
rect 14485 6805 14515 6835
rect 14515 6805 14516 6835
rect 14484 6804 14516 6805
rect 14484 6755 14516 6756
rect 14484 6725 14485 6755
rect 14485 6725 14515 6755
rect 14515 6725 14516 6755
rect 14484 6724 14516 6725
rect 14484 6675 14516 6676
rect 14484 6645 14485 6675
rect 14485 6645 14515 6675
rect 14515 6645 14516 6675
rect 14484 6644 14516 6645
rect 14484 6595 14516 6596
rect 14484 6565 14485 6595
rect 14485 6565 14515 6595
rect 14515 6565 14516 6595
rect 14484 6564 14516 6565
rect 14484 6515 14516 6516
rect 14484 6485 14485 6515
rect 14485 6485 14515 6515
rect 14515 6485 14516 6515
rect 14484 6484 14516 6485
rect 14484 6435 14516 6436
rect 14484 6405 14485 6435
rect 14485 6405 14515 6435
rect 14515 6405 14516 6435
rect 14484 6404 14516 6405
rect 14484 6355 14516 6356
rect 14484 6325 14485 6355
rect 14485 6325 14515 6355
rect 14515 6325 14516 6355
rect 14484 6324 14516 6325
rect 14484 6275 14516 6276
rect 14484 6245 14485 6275
rect 14485 6245 14515 6275
rect 14515 6245 14516 6275
rect 14484 6244 14516 6245
rect 14484 6195 14516 6196
rect 14484 6165 14485 6195
rect 14485 6165 14515 6195
rect 14515 6165 14516 6195
rect 14484 6164 14516 6165
rect 14484 6115 14516 6116
rect 14484 6085 14485 6115
rect 14485 6085 14515 6115
rect 14515 6085 14516 6115
rect 14484 6084 14516 6085
rect 14484 6035 14516 6036
rect 14484 6005 14485 6035
rect 14485 6005 14515 6035
rect 14515 6005 14516 6035
rect 14484 6004 14516 6005
rect 14484 5955 14516 5956
rect 14484 5925 14485 5955
rect 14485 5925 14515 5955
rect 14515 5925 14516 5955
rect 14484 5924 14516 5925
rect 14484 5875 14516 5876
rect 14484 5845 14485 5875
rect 14485 5845 14515 5875
rect 14515 5845 14516 5875
rect 14484 5844 14516 5845
rect 14484 5795 14516 5796
rect 14484 5765 14485 5795
rect 14485 5765 14515 5795
rect 14515 5765 14516 5795
rect 14484 5764 14516 5765
rect 14484 5715 14516 5716
rect 14484 5685 14485 5715
rect 14485 5685 14515 5715
rect 14515 5685 14516 5715
rect 14484 5684 14516 5685
rect 14484 5635 14516 5636
rect 14484 5605 14485 5635
rect 14485 5605 14515 5635
rect 14515 5605 14516 5635
rect 14484 5604 14516 5605
rect 14484 5555 14516 5556
rect 14484 5525 14485 5555
rect 14485 5525 14515 5555
rect 14515 5525 14516 5555
rect 14484 5524 14516 5525
rect 14484 5475 14516 5476
rect 14484 5445 14485 5475
rect 14485 5445 14515 5475
rect 14515 5445 14516 5475
rect 14484 5444 14516 5445
rect 14484 5395 14516 5396
rect 14484 5365 14485 5395
rect 14485 5365 14515 5395
rect 14515 5365 14516 5395
rect 14484 5364 14516 5365
rect 14484 5315 14516 5316
rect 14484 5285 14485 5315
rect 14485 5285 14515 5315
rect 14515 5285 14516 5315
rect 14484 5284 14516 5285
rect 14484 5235 14516 5236
rect 14484 5205 14485 5235
rect 14485 5205 14515 5235
rect 14515 5205 14516 5235
rect 14484 5204 14516 5205
rect 14484 5155 14516 5156
rect 14484 5125 14485 5155
rect 14485 5125 14515 5155
rect 14515 5125 14516 5155
rect 14484 5124 14516 5125
rect 14484 5075 14516 5076
rect 14484 5045 14485 5075
rect 14485 5045 14515 5075
rect 14515 5045 14516 5075
rect 14484 5044 14516 5045
rect 14484 4995 14516 4996
rect 14484 4965 14485 4995
rect 14485 4965 14515 4995
rect 14515 4965 14516 4995
rect 14484 4964 14516 4965
rect 14484 4915 14516 4916
rect 14484 4885 14485 4915
rect 14485 4885 14515 4915
rect 14515 4885 14516 4915
rect 14484 4884 14516 4885
rect 14484 4835 14516 4836
rect 14484 4805 14485 4835
rect 14485 4805 14515 4835
rect 14515 4805 14516 4835
rect 14484 4804 14516 4805
rect 14484 4675 14516 4676
rect 14484 4645 14485 4675
rect 14485 4645 14515 4675
rect 14515 4645 14516 4675
rect 14484 4644 14516 4645
rect 14484 4515 14516 4516
rect 14484 4485 14485 4515
rect 14485 4485 14515 4515
rect 14515 4485 14516 4515
rect 14484 4484 14516 4485
rect 14484 4435 14516 4436
rect 14484 4405 14485 4435
rect 14485 4405 14515 4435
rect 14515 4405 14516 4435
rect 14484 4404 14516 4405
rect 14484 4355 14516 4356
rect 14484 4325 14485 4355
rect 14485 4325 14515 4355
rect 14515 4325 14516 4355
rect 14484 4324 14516 4325
rect 14484 4275 14516 4276
rect 14484 4245 14485 4275
rect 14485 4245 14515 4275
rect 14515 4245 14516 4275
rect 14484 4244 14516 4245
rect 14484 4195 14516 4196
rect 14484 4165 14485 4195
rect 14485 4165 14515 4195
rect 14515 4165 14516 4195
rect 14484 4164 14516 4165
rect 14484 4115 14516 4116
rect 14484 4085 14485 4115
rect 14485 4085 14515 4115
rect 14515 4085 14516 4115
rect 14484 4084 14516 4085
rect 14484 4035 14516 4036
rect 14484 4005 14485 4035
rect 14485 4005 14515 4035
rect 14515 4005 14516 4035
rect 14484 4004 14516 4005
rect 14484 3955 14516 3956
rect 14484 3925 14485 3955
rect 14485 3925 14515 3955
rect 14515 3925 14516 3955
rect 14484 3924 14516 3925
rect 14484 3875 14516 3876
rect 14484 3845 14485 3875
rect 14485 3845 14515 3875
rect 14515 3845 14516 3875
rect 14484 3844 14516 3845
rect 14484 3795 14516 3796
rect 14484 3765 14485 3795
rect 14485 3765 14515 3795
rect 14515 3765 14516 3795
rect 14484 3764 14516 3765
rect 14484 3715 14516 3716
rect 14484 3685 14485 3715
rect 14485 3685 14515 3715
rect 14515 3685 14516 3715
rect 14484 3684 14516 3685
rect 14484 3635 14516 3636
rect 14484 3605 14485 3635
rect 14485 3605 14515 3635
rect 14515 3605 14516 3635
rect 14484 3604 14516 3605
rect 14484 3555 14516 3556
rect 14484 3525 14485 3555
rect 14485 3525 14515 3555
rect 14515 3525 14516 3555
rect 14484 3524 14516 3525
rect 14484 3475 14516 3476
rect 14484 3445 14485 3475
rect 14485 3445 14515 3475
rect 14515 3445 14516 3475
rect 14484 3444 14516 3445
rect 14484 3395 14516 3396
rect 14484 3365 14485 3395
rect 14485 3365 14515 3395
rect 14515 3365 14516 3395
rect 14484 3364 14516 3365
rect 14484 3235 14516 3236
rect 14484 3205 14485 3235
rect 14485 3205 14515 3235
rect 14515 3205 14516 3235
rect 14484 3204 14516 3205
rect 14484 3155 14516 3156
rect 14484 3125 14485 3155
rect 14485 3125 14515 3155
rect 14515 3125 14516 3155
rect 14484 3124 14516 3125
rect 14484 3075 14516 3076
rect 14484 3045 14485 3075
rect 14485 3045 14515 3075
rect 14515 3045 14516 3075
rect 14484 3044 14516 3045
rect 14484 2995 14516 2996
rect 14484 2965 14485 2995
rect 14485 2965 14515 2995
rect 14515 2965 14516 2995
rect 14484 2964 14516 2965
rect 14484 2915 14516 2916
rect 14484 2885 14485 2915
rect 14485 2885 14515 2915
rect 14515 2885 14516 2915
rect 14484 2884 14516 2885
rect 14484 2835 14516 2836
rect 14484 2805 14485 2835
rect 14485 2805 14515 2835
rect 14515 2805 14516 2835
rect 14484 2804 14516 2805
rect 14484 2755 14516 2756
rect 14484 2725 14485 2755
rect 14485 2725 14515 2755
rect 14515 2725 14516 2755
rect 14484 2724 14516 2725
rect 14484 2675 14516 2676
rect 14484 2645 14485 2675
rect 14485 2645 14515 2675
rect 14515 2645 14516 2675
rect 14484 2644 14516 2645
rect 14484 2595 14516 2596
rect 14484 2565 14485 2595
rect 14485 2565 14515 2595
rect 14515 2565 14516 2595
rect 14484 2564 14516 2565
rect 14484 2515 14516 2516
rect 14484 2485 14485 2515
rect 14485 2485 14515 2515
rect 14515 2485 14516 2515
rect 14484 2484 14516 2485
rect 14484 2435 14516 2436
rect 14484 2405 14485 2435
rect 14485 2405 14515 2435
rect 14515 2405 14516 2435
rect 14484 2404 14516 2405
rect 14484 2355 14516 2356
rect 14484 2325 14485 2355
rect 14485 2325 14515 2355
rect 14515 2325 14516 2355
rect 14484 2324 14516 2325
rect 14484 2275 14516 2276
rect 14484 2245 14485 2275
rect 14485 2245 14515 2275
rect 14515 2245 14516 2275
rect 14484 2244 14516 2245
rect 14484 2195 14516 2196
rect 14484 2165 14485 2195
rect 14485 2165 14515 2195
rect 14515 2165 14516 2195
rect 14484 2164 14516 2165
rect 14484 2115 14516 2116
rect 14484 2085 14485 2115
rect 14485 2085 14515 2115
rect 14515 2085 14516 2115
rect 14484 2084 14516 2085
rect 14484 1955 14516 1956
rect 14484 1925 14485 1955
rect 14485 1925 14515 1955
rect 14515 1925 14516 1955
rect 14484 1924 14516 1925
rect 14484 1795 14516 1796
rect 14484 1765 14485 1795
rect 14485 1765 14515 1795
rect 14515 1765 14516 1795
rect 14484 1764 14516 1765
rect 14484 1715 14516 1716
rect 14484 1685 14485 1715
rect 14485 1685 14515 1715
rect 14515 1685 14516 1715
rect 14484 1684 14516 1685
rect 14484 1635 14516 1636
rect 14484 1605 14485 1635
rect 14485 1605 14515 1635
rect 14515 1605 14516 1635
rect 14484 1604 14516 1605
rect 14484 1555 14516 1556
rect 14484 1525 14485 1555
rect 14485 1525 14515 1555
rect 14515 1525 14516 1555
rect 14484 1524 14516 1525
rect 14484 1475 14516 1476
rect 14484 1445 14485 1475
rect 14485 1445 14515 1475
rect 14515 1445 14516 1475
rect 14484 1444 14516 1445
rect 14484 1395 14516 1396
rect 14484 1365 14485 1395
rect 14485 1365 14515 1395
rect 14515 1365 14516 1395
rect 14484 1364 14516 1365
rect 14484 1315 14516 1316
rect 14484 1285 14485 1315
rect 14485 1285 14515 1315
rect 14515 1285 14516 1315
rect 14484 1284 14516 1285
rect 14484 1235 14516 1236
rect 14484 1205 14485 1235
rect 14485 1205 14515 1235
rect 14515 1205 14516 1235
rect 14484 1204 14516 1205
rect 14484 1155 14516 1156
rect 14484 1125 14485 1155
rect 14485 1125 14515 1155
rect 14515 1125 14516 1155
rect 14484 1124 14516 1125
rect 14484 1075 14516 1076
rect 14484 1045 14485 1075
rect 14485 1045 14515 1075
rect 14515 1045 14516 1075
rect 14484 1044 14516 1045
rect 14484 995 14516 996
rect 14484 965 14485 995
rect 14485 965 14515 995
rect 14515 965 14516 995
rect 14484 964 14516 965
rect 14484 915 14516 916
rect 14484 885 14485 915
rect 14485 885 14515 915
rect 14515 885 14516 915
rect 14484 884 14516 885
rect 14484 835 14516 836
rect 14484 805 14485 835
rect 14485 805 14515 835
rect 14515 805 14516 835
rect 14484 804 14516 805
rect 14484 755 14516 756
rect 14484 725 14485 755
rect 14485 725 14515 755
rect 14515 725 14516 755
rect 14484 724 14516 725
rect 14484 675 14516 676
rect 14484 645 14485 675
rect 14485 645 14515 675
rect 14515 645 14516 675
rect 14484 644 14516 645
rect 14484 595 14516 596
rect 14484 565 14485 595
rect 14485 565 14515 595
rect 14515 565 14516 595
rect 14484 564 14516 565
rect 484 515 516 516
rect 484 485 485 515
rect 485 485 515 515
rect 515 485 516 515
rect 484 484 516 485
rect 324 244 356 436
rect 484 244 516 436
rect 564 4 596 196
rect 14484 515 14516 516
rect 14484 485 14485 515
rect 14485 485 14515 515
rect 14515 485 14516 515
rect 14484 484 14516 485
rect 14564 13124 14596 13156
rect 14564 3284 14596 3316
rect 14644 15955 14676 15956
rect 14644 15925 14645 15955
rect 14645 15925 14675 15955
rect 14675 15925 14676 15955
rect 14644 15924 14676 15925
rect 14644 15875 14676 15876
rect 14644 15845 14645 15875
rect 14645 15845 14675 15875
rect 14675 15845 14676 15875
rect 14644 15844 14676 15845
rect 14644 15795 14676 15796
rect 14644 15765 14645 15795
rect 14645 15765 14675 15795
rect 14675 15765 14676 15795
rect 14644 15764 14676 15765
rect 14644 15715 14676 15716
rect 14644 15685 14645 15715
rect 14645 15685 14675 15715
rect 14675 15685 14676 15715
rect 14644 15684 14676 15685
rect 14644 15635 14676 15636
rect 14644 15605 14645 15635
rect 14645 15605 14675 15635
rect 14675 15605 14676 15635
rect 14644 15604 14676 15605
rect 14644 15555 14676 15556
rect 14644 15525 14645 15555
rect 14645 15525 14675 15555
rect 14675 15525 14676 15555
rect 14644 15524 14676 15525
rect 14644 15475 14676 15476
rect 14644 15445 14645 15475
rect 14645 15445 14675 15475
rect 14675 15445 14676 15475
rect 14644 15444 14676 15445
rect 14644 15395 14676 15396
rect 14644 15365 14645 15395
rect 14645 15365 14675 15395
rect 14675 15365 14676 15395
rect 14644 15364 14676 15365
rect 14644 15315 14676 15316
rect 14644 15285 14645 15315
rect 14645 15285 14675 15315
rect 14675 15285 14676 15315
rect 14644 15284 14676 15285
rect 14644 15235 14676 15236
rect 14644 15205 14645 15235
rect 14645 15205 14675 15235
rect 14675 15205 14676 15235
rect 14644 15204 14676 15205
rect 14644 15155 14676 15156
rect 14644 15125 14645 15155
rect 14645 15125 14675 15155
rect 14675 15125 14676 15155
rect 14644 15124 14676 15125
rect 14644 15075 14676 15076
rect 14644 15045 14645 15075
rect 14645 15045 14675 15075
rect 14675 15045 14676 15075
rect 14644 15044 14676 15045
rect 14644 14995 14676 14996
rect 14644 14965 14645 14995
rect 14645 14965 14675 14995
rect 14675 14965 14676 14995
rect 14644 14964 14676 14965
rect 14644 14915 14676 14916
rect 14644 14885 14645 14915
rect 14645 14885 14675 14915
rect 14675 14885 14676 14915
rect 14644 14884 14676 14885
rect 14644 14835 14676 14836
rect 14644 14805 14645 14835
rect 14645 14805 14675 14835
rect 14675 14805 14676 14835
rect 14644 14804 14676 14805
rect 14644 14755 14676 14756
rect 14644 14725 14645 14755
rect 14645 14725 14675 14755
rect 14675 14725 14676 14755
rect 14644 14724 14676 14725
rect 14644 14675 14676 14676
rect 14644 14645 14645 14675
rect 14645 14645 14675 14675
rect 14675 14645 14676 14675
rect 14644 14644 14676 14645
rect 14644 14515 14676 14516
rect 14644 14485 14645 14515
rect 14645 14485 14675 14515
rect 14675 14485 14676 14515
rect 14644 14484 14676 14485
rect 14644 14355 14676 14356
rect 14644 14325 14645 14355
rect 14645 14325 14675 14355
rect 14675 14325 14676 14355
rect 14644 14324 14676 14325
rect 14644 14275 14676 14276
rect 14644 14245 14645 14275
rect 14645 14245 14675 14275
rect 14675 14245 14676 14275
rect 14644 14244 14676 14245
rect 14644 14195 14676 14196
rect 14644 14165 14645 14195
rect 14645 14165 14675 14195
rect 14675 14165 14676 14195
rect 14644 14164 14676 14165
rect 14644 14115 14676 14116
rect 14644 14085 14645 14115
rect 14645 14085 14675 14115
rect 14675 14085 14676 14115
rect 14644 14084 14676 14085
rect 14644 14035 14676 14036
rect 14644 14005 14645 14035
rect 14645 14005 14675 14035
rect 14675 14005 14676 14035
rect 14644 14004 14676 14005
rect 14644 13955 14676 13956
rect 14644 13925 14645 13955
rect 14645 13925 14675 13955
rect 14675 13925 14676 13955
rect 14644 13924 14676 13925
rect 14644 13875 14676 13876
rect 14644 13845 14645 13875
rect 14645 13845 14675 13875
rect 14675 13845 14676 13875
rect 14644 13844 14676 13845
rect 14644 13795 14676 13796
rect 14644 13765 14645 13795
rect 14645 13765 14675 13795
rect 14675 13765 14676 13795
rect 14644 13764 14676 13765
rect 14644 13715 14676 13716
rect 14644 13685 14645 13715
rect 14645 13685 14675 13715
rect 14675 13685 14676 13715
rect 14644 13684 14676 13685
rect 14644 13635 14676 13636
rect 14644 13605 14645 13635
rect 14645 13605 14675 13635
rect 14675 13605 14676 13635
rect 14644 13604 14676 13605
rect 14644 13555 14676 13556
rect 14644 13525 14645 13555
rect 14645 13525 14675 13555
rect 14675 13525 14676 13555
rect 14644 13524 14676 13525
rect 14644 13475 14676 13476
rect 14644 13445 14645 13475
rect 14645 13445 14675 13475
rect 14675 13445 14676 13475
rect 14644 13444 14676 13445
rect 14644 13395 14676 13396
rect 14644 13365 14645 13395
rect 14645 13365 14675 13395
rect 14675 13365 14676 13395
rect 14644 13364 14676 13365
rect 14644 13315 14676 13316
rect 14644 13285 14645 13315
rect 14645 13285 14675 13315
rect 14675 13285 14676 13315
rect 14644 13284 14676 13285
rect 14644 13235 14676 13236
rect 14644 13205 14645 13235
rect 14645 13205 14675 13235
rect 14675 13205 14676 13235
rect 14644 13204 14676 13205
rect 14644 13155 14676 13156
rect 14644 13125 14645 13155
rect 14645 13125 14675 13155
rect 14675 13125 14676 13155
rect 14644 13124 14676 13125
rect 14644 13075 14676 13076
rect 14644 13045 14645 13075
rect 14645 13045 14675 13075
rect 14675 13045 14676 13075
rect 14644 13044 14676 13045
rect 14644 12995 14676 12996
rect 14644 12965 14645 12995
rect 14645 12965 14675 12995
rect 14675 12965 14676 12995
rect 14644 12964 14676 12965
rect 14644 12915 14676 12916
rect 14644 12885 14645 12915
rect 14645 12885 14675 12915
rect 14675 12885 14676 12915
rect 14644 12884 14676 12885
rect 14644 12835 14676 12836
rect 14644 12805 14645 12835
rect 14645 12805 14675 12835
rect 14675 12805 14676 12835
rect 14644 12804 14676 12805
rect 14644 12755 14676 12756
rect 14644 12725 14645 12755
rect 14645 12725 14675 12755
rect 14675 12725 14676 12755
rect 14644 12724 14676 12725
rect 14644 12675 14676 12676
rect 14644 12645 14645 12675
rect 14645 12645 14675 12675
rect 14675 12645 14676 12675
rect 14644 12644 14676 12645
rect 14644 12595 14676 12596
rect 14644 12565 14645 12595
rect 14645 12565 14675 12595
rect 14675 12565 14676 12595
rect 14644 12564 14676 12565
rect 14644 12515 14676 12516
rect 14644 12485 14645 12515
rect 14645 12485 14675 12515
rect 14675 12485 14676 12515
rect 14644 12484 14676 12485
rect 14644 12435 14676 12436
rect 14644 12405 14645 12435
rect 14645 12405 14675 12435
rect 14675 12405 14676 12435
rect 14644 12404 14676 12405
rect 14644 12355 14676 12356
rect 14644 12325 14645 12355
rect 14645 12325 14675 12355
rect 14675 12325 14676 12355
rect 14644 12324 14676 12325
rect 14644 12275 14676 12276
rect 14644 12245 14645 12275
rect 14645 12245 14675 12275
rect 14675 12245 14676 12275
rect 14644 12244 14676 12245
rect 14644 12195 14676 12196
rect 14644 12165 14645 12195
rect 14645 12165 14675 12195
rect 14675 12165 14676 12195
rect 14644 12164 14676 12165
rect 14644 12115 14676 12116
rect 14644 12085 14645 12115
rect 14645 12085 14675 12115
rect 14675 12085 14676 12115
rect 14644 12084 14676 12085
rect 14644 12035 14676 12036
rect 14644 12005 14645 12035
rect 14645 12005 14675 12035
rect 14675 12005 14676 12035
rect 14644 12004 14676 12005
rect 14644 11955 14676 11956
rect 14644 11925 14645 11955
rect 14645 11925 14675 11955
rect 14675 11925 14676 11955
rect 14644 11924 14676 11925
rect 14644 11795 14676 11796
rect 14644 11765 14645 11795
rect 14645 11765 14675 11795
rect 14675 11765 14676 11795
rect 14644 11764 14676 11765
rect 14644 11635 14676 11636
rect 14644 11605 14645 11635
rect 14645 11605 14675 11635
rect 14675 11605 14676 11635
rect 14644 11604 14676 11605
rect 14644 11555 14676 11556
rect 14644 11525 14645 11555
rect 14645 11525 14675 11555
rect 14675 11525 14676 11555
rect 14644 11524 14676 11525
rect 14644 11475 14676 11476
rect 14644 11445 14645 11475
rect 14645 11445 14675 11475
rect 14675 11445 14676 11475
rect 14644 11444 14676 11445
rect 14644 11395 14676 11396
rect 14644 11365 14645 11395
rect 14645 11365 14675 11395
rect 14675 11365 14676 11395
rect 14644 11364 14676 11365
rect 14644 11315 14676 11316
rect 14644 11285 14645 11315
rect 14645 11285 14675 11315
rect 14675 11285 14676 11315
rect 14644 11284 14676 11285
rect 14644 11235 14676 11236
rect 14644 11205 14645 11235
rect 14645 11205 14675 11235
rect 14675 11205 14676 11235
rect 14644 11204 14676 11205
rect 14644 11155 14676 11156
rect 14644 11125 14645 11155
rect 14645 11125 14675 11155
rect 14675 11125 14676 11155
rect 14644 11124 14676 11125
rect 14644 11075 14676 11076
rect 14644 11045 14645 11075
rect 14645 11045 14675 11075
rect 14675 11045 14676 11075
rect 14644 11044 14676 11045
rect 14644 10995 14676 10996
rect 14644 10965 14645 10995
rect 14645 10965 14675 10995
rect 14675 10965 14676 10995
rect 14644 10964 14676 10965
rect 14644 10915 14676 10916
rect 14644 10885 14645 10915
rect 14645 10885 14675 10915
rect 14675 10885 14676 10915
rect 14644 10884 14676 10885
rect 14644 10835 14676 10836
rect 14644 10805 14645 10835
rect 14645 10805 14675 10835
rect 14675 10805 14676 10835
rect 14644 10804 14676 10805
rect 14644 10755 14676 10756
rect 14644 10725 14645 10755
rect 14645 10725 14675 10755
rect 14675 10725 14676 10755
rect 14644 10724 14676 10725
rect 14644 10675 14676 10676
rect 14644 10645 14645 10675
rect 14645 10645 14675 10675
rect 14675 10645 14676 10675
rect 14644 10644 14676 10645
rect 14644 10595 14676 10596
rect 14644 10565 14645 10595
rect 14645 10565 14675 10595
rect 14675 10565 14676 10595
rect 14644 10564 14676 10565
rect 14644 10515 14676 10516
rect 14644 10485 14645 10515
rect 14645 10485 14675 10515
rect 14675 10485 14676 10515
rect 14644 10484 14676 10485
rect 14644 10435 14676 10436
rect 14644 10405 14645 10435
rect 14645 10405 14675 10435
rect 14675 10405 14676 10435
rect 14644 10404 14676 10405
rect 14644 10355 14676 10356
rect 14644 10325 14645 10355
rect 14645 10325 14675 10355
rect 14675 10325 14676 10355
rect 14644 10324 14676 10325
rect 14644 10275 14676 10276
rect 14644 10245 14645 10275
rect 14645 10245 14675 10275
rect 14675 10245 14676 10275
rect 14644 10244 14676 10245
rect 14644 10195 14676 10196
rect 14644 10165 14645 10195
rect 14645 10165 14675 10195
rect 14675 10165 14676 10195
rect 14644 10164 14676 10165
rect 14644 10115 14676 10116
rect 14644 10085 14645 10115
rect 14645 10085 14675 10115
rect 14675 10085 14676 10115
rect 14644 10084 14676 10085
rect 14644 10035 14676 10036
rect 14644 10005 14645 10035
rect 14645 10005 14675 10035
rect 14675 10005 14676 10035
rect 14644 10004 14676 10005
rect 14644 9955 14676 9956
rect 14644 9925 14645 9955
rect 14645 9925 14675 9955
rect 14675 9925 14676 9955
rect 14644 9924 14676 9925
rect 14644 9875 14676 9876
rect 14644 9845 14645 9875
rect 14645 9845 14675 9875
rect 14675 9845 14676 9875
rect 14644 9844 14676 9845
rect 14644 9795 14676 9796
rect 14644 9765 14645 9795
rect 14645 9765 14675 9795
rect 14675 9765 14676 9795
rect 14644 9764 14676 9765
rect 14644 9715 14676 9716
rect 14644 9685 14645 9715
rect 14645 9685 14675 9715
rect 14675 9685 14676 9715
rect 14644 9684 14676 9685
rect 14644 9635 14676 9636
rect 14644 9605 14645 9635
rect 14645 9605 14675 9635
rect 14675 9605 14676 9635
rect 14644 9604 14676 9605
rect 14644 9555 14676 9556
rect 14644 9525 14645 9555
rect 14645 9525 14675 9555
rect 14675 9525 14676 9555
rect 14644 9524 14676 9525
rect 14644 9475 14676 9476
rect 14644 9445 14645 9475
rect 14645 9445 14675 9475
rect 14675 9445 14676 9475
rect 14644 9444 14676 9445
rect 14644 9395 14676 9396
rect 14644 9365 14645 9395
rect 14645 9365 14675 9395
rect 14675 9365 14676 9395
rect 14644 9364 14676 9365
rect 14644 9315 14676 9316
rect 14644 9285 14645 9315
rect 14645 9285 14675 9315
rect 14675 9285 14676 9315
rect 14644 9284 14676 9285
rect 14644 9235 14676 9236
rect 14644 9205 14645 9235
rect 14645 9205 14675 9235
rect 14675 9205 14676 9235
rect 14644 9204 14676 9205
rect 14644 9155 14676 9156
rect 14644 9125 14645 9155
rect 14645 9125 14675 9155
rect 14675 9125 14676 9155
rect 14644 9124 14676 9125
rect 14644 9075 14676 9076
rect 14644 9045 14645 9075
rect 14645 9045 14675 9075
rect 14675 9045 14676 9075
rect 14644 9044 14676 9045
rect 14644 8995 14676 8996
rect 14644 8965 14645 8995
rect 14645 8965 14675 8995
rect 14675 8965 14676 8995
rect 14644 8964 14676 8965
rect 14644 8915 14676 8916
rect 14644 8885 14645 8915
rect 14645 8885 14675 8915
rect 14675 8885 14676 8915
rect 14644 8884 14676 8885
rect 14644 8835 14676 8836
rect 14644 8805 14645 8835
rect 14645 8805 14675 8835
rect 14675 8805 14676 8835
rect 14644 8804 14676 8805
rect 14644 8755 14676 8756
rect 14644 8725 14645 8755
rect 14645 8725 14675 8755
rect 14675 8725 14676 8755
rect 14644 8724 14676 8725
rect 14644 8675 14676 8676
rect 14644 8645 14645 8675
rect 14645 8645 14675 8675
rect 14675 8645 14676 8675
rect 14644 8644 14676 8645
rect 14644 8595 14676 8596
rect 14644 8565 14645 8595
rect 14645 8565 14675 8595
rect 14675 8565 14676 8595
rect 14644 8564 14676 8565
rect 14644 8515 14676 8516
rect 14644 8485 14645 8515
rect 14645 8485 14675 8515
rect 14675 8485 14676 8515
rect 14644 8484 14676 8485
rect 14644 8435 14676 8436
rect 14644 8405 14645 8435
rect 14645 8405 14675 8435
rect 14675 8405 14676 8435
rect 14644 8404 14676 8405
rect 14644 8355 14676 8356
rect 14644 8325 14645 8355
rect 14645 8325 14675 8355
rect 14675 8325 14676 8355
rect 14644 8324 14676 8325
rect 14644 8275 14676 8276
rect 14644 8245 14645 8275
rect 14645 8245 14675 8275
rect 14675 8245 14676 8275
rect 14644 8244 14676 8245
rect 14644 8195 14676 8196
rect 14644 8165 14645 8195
rect 14645 8165 14675 8195
rect 14675 8165 14676 8195
rect 14644 8164 14676 8165
rect 14644 8115 14676 8116
rect 14644 8085 14645 8115
rect 14645 8085 14675 8115
rect 14675 8085 14676 8115
rect 14644 8084 14676 8085
rect 14644 8035 14676 8036
rect 14644 8005 14645 8035
rect 14645 8005 14675 8035
rect 14675 8005 14676 8035
rect 14644 8004 14676 8005
rect 14644 7955 14676 7956
rect 14644 7925 14645 7955
rect 14645 7925 14675 7955
rect 14675 7925 14676 7955
rect 14644 7924 14676 7925
rect 14644 7875 14676 7876
rect 14644 7845 14645 7875
rect 14645 7845 14675 7875
rect 14675 7845 14676 7875
rect 14644 7844 14676 7845
rect 14644 7795 14676 7796
rect 14644 7765 14645 7795
rect 14645 7765 14675 7795
rect 14675 7765 14676 7795
rect 14644 7764 14676 7765
rect 14644 7715 14676 7716
rect 14644 7685 14645 7715
rect 14645 7685 14675 7715
rect 14675 7685 14676 7715
rect 14644 7684 14676 7685
rect 14644 7635 14676 7636
rect 14644 7605 14645 7635
rect 14645 7605 14675 7635
rect 14675 7605 14676 7635
rect 14644 7604 14676 7605
rect 14644 7555 14676 7556
rect 14644 7525 14645 7555
rect 14645 7525 14675 7555
rect 14675 7525 14676 7555
rect 14644 7524 14676 7525
rect 14644 7475 14676 7476
rect 14644 7445 14645 7475
rect 14645 7445 14675 7475
rect 14675 7445 14676 7475
rect 14644 7444 14676 7445
rect 14644 7395 14676 7396
rect 14644 7365 14645 7395
rect 14645 7365 14675 7395
rect 14675 7365 14676 7395
rect 14644 7364 14676 7365
rect 14644 7315 14676 7316
rect 14644 7285 14645 7315
rect 14645 7285 14675 7315
rect 14675 7285 14676 7315
rect 14644 7284 14676 7285
rect 14644 7235 14676 7236
rect 14644 7205 14645 7235
rect 14645 7205 14675 7235
rect 14675 7205 14676 7235
rect 14644 7204 14676 7205
rect 14644 7155 14676 7156
rect 14644 7125 14645 7155
rect 14645 7125 14675 7155
rect 14675 7125 14676 7155
rect 14644 7124 14676 7125
rect 14644 7075 14676 7076
rect 14644 7045 14645 7075
rect 14645 7045 14675 7075
rect 14675 7045 14676 7075
rect 14644 7044 14676 7045
rect 14644 6995 14676 6996
rect 14644 6965 14645 6995
rect 14645 6965 14675 6995
rect 14675 6965 14676 6995
rect 14644 6964 14676 6965
rect 14644 6915 14676 6916
rect 14644 6885 14645 6915
rect 14645 6885 14675 6915
rect 14675 6885 14676 6915
rect 14644 6884 14676 6885
rect 14644 6835 14676 6836
rect 14644 6805 14645 6835
rect 14645 6805 14675 6835
rect 14675 6805 14676 6835
rect 14644 6804 14676 6805
rect 14644 6755 14676 6756
rect 14644 6725 14645 6755
rect 14645 6725 14675 6755
rect 14675 6725 14676 6755
rect 14644 6724 14676 6725
rect 14644 6675 14676 6676
rect 14644 6645 14645 6675
rect 14645 6645 14675 6675
rect 14675 6645 14676 6675
rect 14644 6644 14676 6645
rect 14644 6595 14676 6596
rect 14644 6565 14645 6595
rect 14645 6565 14675 6595
rect 14675 6565 14676 6595
rect 14644 6564 14676 6565
rect 14644 6515 14676 6516
rect 14644 6485 14645 6515
rect 14645 6485 14675 6515
rect 14675 6485 14676 6515
rect 14644 6484 14676 6485
rect 14644 6435 14676 6436
rect 14644 6405 14645 6435
rect 14645 6405 14675 6435
rect 14675 6405 14676 6435
rect 14644 6404 14676 6405
rect 14644 6355 14676 6356
rect 14644 6325 14645 6355
rect 14645 6325 14675 6355
rect 14675 6325 14676 6355
rect 14644 6324 14676 6325
rect 14644 6275 14676 6276
rect 14644 6245 14645 6275
rect 14645 6245 14675 6275
rect 14675 6245 14676 6275
rect 14644 6244 14676 6245
rect 14644 6195 14676 6196
rect 14644 6165 14645 6195
rect 14645 6165 14675 6195
rect 14675 6165 14676 6195
rect 14644 6164 14676 6165
rect 14644 6115 14676 6116
rect 14644 6085 14645 6115
rect 14645 6085 14675 6115
rect 14675 6085 14676 6115
rect 14644 6084 14676 6085
rect 14644 6035 14676 6036
rect 14644 6005 14645 6035
rect 14645 6005 14675 6035
rect 14675 6005 14676 6035
rect 14644 6004 14676 6005
rect 14644 5955 14676 5956
rect 14644 5925 14645 5955
rect 14645 5925 14675 5955
rect 14675 5925 14676 5955
rect 14644 5924 14676 5925
rect 14644 5875 14676 5876
rect 14644 5845 14645 5875
rect 14645 5845 14675 5875
rect 14675 5845 14676 5875
rect 14644 5844 14676 5845
rect 14644 5795 14676 5796
rect 14644 5765 14645 5795
rect 14645 5765 14675 5795
rect 14675 5765 14676 5795
rect 14644 5764 14676 5765
rect 14644 5715 14676 5716
rect 14644 5685 14645 5715
rect 14645 5685 14675 5715
rect 14675 5685 14676 5715
rect 14644 5684 14676 5685
rect 14644 5635 14676 5636
rect 14644 5605 14645 5635
rect 14645 5605 14675 5635
rect 14675 5605 14676 5635
rect 14644 5604 14676 5605
rect 14644 5555 14676 5556
rect 14644 5525 14645 5555
rect 14645 5525 14675 5555
rect 14675 5525 14676 5555
rect 14644 5524 14676 5525
rect 14644 5475 14676 5476
rect 14644 5445 14645 5475
rect 14645 5445 14675 5475
rect 14675 5445 14676 5475
rect 14644 5444 14676 5445
rect 14644 5395 14676 5396
rect 14644 5365 14645 5395
rect 14645 5365 14675 5395
rect 14675 5365 14676 5395
rect 14644 5364 14676 5365
rect 14644 5315 14676 5316
rect 14644 5285 14645 5315
rect 14645 5285 14675 5315
rect 14675 5285 14676 5315
rect 14644 5284 14676 5285
rect 14644 5235 14676 5236
rect 14644 5205 14645 5235
rect 14645 5205 14675 5235
rect 14675 5205 14676 5235
rect 14644 5204 14676 5205
rect 14644 5155 14676 5156
rect 14644 5125 14645 5155
rect 14645 5125 14675 5155
rect 14675 5125 14676 5155
rect 14644 5124 14676 5125
rect 14644 5075 14676 5076
rect 14644 5045 14645 5075
rect 14645 5045 14675 5075
rect 14675 5045 14676 5075
rect 14644 5044 14676 5045
rect 14644 4995 14676 4996
rect 14644 4965 14645 4995
rect 14645 4965 14675 4995
rect 14675 4965 14676 4995
rect 14644 4964 14676 4965
rect 14644 4915 14676 4916
rect 14644 4885 14645 4915
rect 14645 4885 14675 4915
rect 14675 4885 14676 4915
rect 14644 4884 14676 4885
rect 14644 4835 14676 4836
rect 14644 4805 14645 4835
rect 14645 4805 14675 4835
rect 14675 4805 14676 4835
rect 14644 4804 14676 4805
rect 14644 4675 14676 4676
rect 14644 4645 14645 4675
rect 14645 4645 14675 4675
rect 14675 4645 14676 4675
rect 14644 4644 14676 4645
rect 14644 4515 14676 4516
rect 14644 4485 14645 4515
rect 14645 4485 14675 4515
rect 14675 4485 14676 4515
rect 14644 4484 14676 4485
rect 14644 4435 14676 4436
rect 14644 4405 14645 4435
rect 14645 4405 14675 4435
rect 14675 4405 14676 4435
rect 14644 4404 14676 4405
rect 14644 4355 14676 4356
rect 14644 4325 14645 4355
rect 14645 4325 14675 4355
rect 14675 4325 14676 4355
rect 14644 4324 14676 4325
rect 14644 4275 14676 4276
rect 14644 4245 14645 4275
rect 14645 4245 14675 4275
rect 14675 4245 14676 4275
rect 14644 4244 14676 4245
rect 14644 4195 14676 4196
rect 14644 4165 14645 4195
rect 14645 4165 14675 4195
rect 14675 4165 14676 4195
rect 14644 4164 14676 4165
rect 14644 4115 14676 4116
rect 14644 4085 14645 4115
rect 14645 4085 14675 4115
rect 14675 4085 14676 4115
rect 14644 4084 14676 4085
rect 14644 4035 14676 4036
rect 14644 4005 14645 4035
rect 14645 4005 14675 4035
rect 14675 4005 14676 4035
rect 14644 4004 14676 4005
rect 14644 3955 14676 3956
rect 14644 3925 14645 3955
rect 14645 3925 14675 3955
rect 14675 3925 14676 3955
rect 14644 3924 14676 3925
rect 14644 3875 14676 3876
rect 14644 3845 14645 3875
rect 14645 3845 14675 3875
rect 14675 3845 14676 3875
rect 14644 3844 14676 3845
rect 14644 3795 14676 3796
rect 14644 3765 14645 3795
rect 14645 3765 14675 3795
rect 14675 3765 14676 3795
rect 14644 3764 14676 3765
rect 14644 3715 14676 3716
rect 14644 3685 14645 3715
rect 14645 3685 14675 3715
rect 14675 3685 14676 3715
rect 14644 3684 14676 3685
rect 14644 3635 14676 3636
rect 14644 3605 14645 3635
rect 14645 3605 14675 3635
rect 14675 3605 14676 3635
rect 14644 3604 14676 3605
rect 14644 3555 14676 3556
rect 14644 3525 14645 3555
rect 14645 3525 14675 3555
rect 14675 3525 14676 3555
rect 14644 3524 14676 3525
rect 14644 3475 14676 3476
rect 14644 3445 14645 3475
rect 14645 3445 14675 3475
rect 14675 3445 14676 3475
rect 14644 3444 14676 3445
rect 14644 3395 14676 3396
rect 14644 3365 14645 3395
rect 14645 3365 14675 3395
rect 14675 3365 14676 3395
rect 14644 3364 14676 3365
rect 14644 3315 14676 3316
rect 14644 3285 14645 3315
rect 14645 3285 14675 3315
rect 14675 3285 14676 3315
rect 14644 3284 14676 3285
rect 14644 3235 14676 3236
rect 14644 3205 14645 3235
rect 14645 3205 14675 3235
rect 14675 3205 14676 3235
rect 14644 3204 14676 3205
rect 14644 3155 14676 3156
rect 14644 3125 14645 3155
rect 14645 3125 14675 3155
rect 14675 3125 14676 3155
rect 14644 3124 14676 3125
rect 14644 3075 14676 3076
rect 14644 3045 14645 3075
rect 14645 3045 14675 3075
rect 14675 3045 14676 3075
rect 14644 3044 14676 3045
rect 14644 2995 14676 2996
rect 14644 2965 14645 2995
rect 14645 2965 14675 2995
rect 14675 2965 14676 2995
rect 14644 2964 14676 2965
rect 14644 2915 14676 2916
rect 14644 2885 14645 2915
rect 14645 2885 14675 2915
rect 14675 2885 14676 2915
rect 14644 2884 14676 2885
rect 14644 2835 14676 2836
rect 14644 2805 14645 2835
rect 14645 2805 14675 2835
rect 14675 2805 14676 2835
rect 14644 2804 14676 2805
rect 14644 2755 14676 2756
rect 14644 2725 14645 2755
rect 14645 2725 14675 2755
rect 14675 2725 14676 2755
rect 14644 2724 14676 2725
rect 14644 2675 14676 2676
rect 14644 2645 14645 2675
rect 14645 2645 14675 2675
rect 14675 2645 14676 2675
rect 14644 2644 14676 2645
rect 14644 2595 14676 2596
rect 14644 2565 14645 2595
rect 14645 2565 14675 2595
rect 14675 2565 14676 2595
rect 14644 2564 14676 2565
rect 14644 2515 14676 2516
rect 14644 2485 14645 2515
rect 14645 2485 14675 2515
rect 14675 2485 14676 2515
rect 14644 2484 14676 2485
rect 14644 2435 14676 2436
rect 14644 2405 14645 2435
rect 14645 2405 14675 2435
rect 14675 2405 14676 2435
rect 14644 2404 14676 2405
rect 14644 2355 14676 2356
rect 14644 2325 14645 2355
rect 14645 2325 14675 2355
rect 14675 2325 14676 2355
rect 14644 2324 14676 2325
rect 14644 2275 14676 2276
rect 14644 2245 14645 2275
rect 14645 2245 14675 2275
rect 14675 2245 14676 2275
rect 14644 2244 14676 2245
rect 14644 2195 14676 2196
rect 14644 2165 14645 2195
rect 14645 2165 14675 2195
rect 14675 2165 14676 2195
rect 14644 2164 14676 2165
rect 14644 2115 14676 2116
rect 14644 2085 14645 2115
rect 14645 2085 14675 2115
rect 14675 2085 14676 2115
rect 14644 2084 14676 2085
rect 14644 1955 14676 1956
rect 14644 1925 14645 1955
rect 14645 1925 14675 1955
rect 14675 1925 14676 1955
rect 14644 1924 14676 1925
rect 14644 1795 14676 1796
rect 14644 1765 14645 1795
rect 14645 1765 14675 1795
rect 14675 1765 14676 1795
rect 14644 1764 14676 1765
rect 14644 1715 14676 1716
rect 14644 1685 14645 1715
rect 14645 1685 14675 1715
rect 14675 1685 14676 1715
rect 14644 1684 14676 1685
rect 14644 1635 14676 1636
rect 14644 1605 14645 1635
rect 14645 1605 14675 1635
rect 14675 1605 14676 1635
rect 14644 1604 14676 1605
rect 14644 1555 14676 1556
rect 14644 1525 14645 1555
rect 14645 1525 14675 1555
rect 14675 1525 14676 1555
rect 14644 1524 14676 1525
rect 14644 1475 14676 1476
rect 14644 1445 14645 1475
rect 14645 1445 14675 1475
rect 14675 1445 14676 1475
rect 14644 1444 14676 1445
rect 14644 1395 14676 1396
rect 14644 1365 14645 1395
rect 14645 1365 14675 1395
rect 14675 1365 14676 1395
rect 14644 1364 14676 1365
rect 14644 1315 14676 1316
rect 14644 1285 14645 1315
rect 14645 1285 14675 1315
rect 14675 1285 14676 1315
rect 14644 1284 14676 1285
rect 14644 1235 14676 1236
rect 14644 1205 14645 1235
rect 14645 1205 14675 1235
rect 14675 1205 14676 1235
rect 14644 1204 14676 1205
rect 14644 1155 14676 1156
rect 14644 1125 14645 1155
rect 14645 1125 14675 1155
rect 14675 1125 14676 1155
rect 14644 1124 14676 1125
rect 14644 1075 14676 1076
rect 14644 1045 14645 1075
rect 14645 1045 14675 1075
rect 14675 1045 14676 1075
rect 14644 1044 14676 1045
rect 14644 995 14676 996
rect 14644 965 14645 995
rect 14645 965 14675 995
rect 14675 965 14676 995
rect 14644 964 14676 965
rect 14644 915 14676 916
rect 14644 885 14645 915
rect 14645 885 14675 915
rect 14675 885 14676 915
rect 14644 884 14676 885
rect 14644 835 14676 836
rect 14644 805 14645 835
rect 14645 805 14675 835
rect 14675 805 14676 835
rect 14644 804 14676 805
rect 14644 755 14676 756
rect 14644 725 14645 755
rect 14645 725 14675 755
rect 14675 725 14676 755
rect 14644 724 14676 725
rect 14644 675 14676 676
rect 14644 645 14645 675
rect 14645 645 14675 675
rect 14675 645 14676 675
rect 14644 644 14676 645
rect 14644 595 14676 596
rect 14644 565 14645 595
rect 14645 565 14675 595
rect 14675 565 14676 595
rect 14644 564 14676 565
rect 14644 515 14676 516
rect 14644 485 14645 515
rect 14645 485 14675 515
rect 14675 485 14676 515
rect 14644 484 14676 485
rect 14484 244 14516 436
rect 14724 14404 14756 14436
rect 14724 11844 14756 11876
rect 14724 4564 14756 4596
rect 14724 2004 14756 2036
rect 14804 15955 14836 15956
rect 14804 15925 14805 15955
rect 14805 15925 14835 15955
rect 14835 15925 14836 15955
rect 14804 15924 14836 15925
rect 14804 15875 14836 15876
rect 14804 15845 14805 15875
rect 14805 15845 14835 15875
rect 14835 15845 14836 15875
rect 14804 15844 14836 15845
rect 14804 15795 14836 15796
rect 14804 15765 14805 15795
rect 14805 15765 14835 15795
rect 14835 15765 14836 15795
rect 14804 15764 14836 15765
rect 14804 15715 14836 15716
rect 14804 15685 14805 15715
rect 14805 15685 14835 15715
rect 14835 15685 14836 15715
rect 14804 15684 14836 15685
rect 14804 15635 14836 15636
rect 14804 15605 14805 15635
rect 14805 15605 14835 15635
rect 14835 15605 14836 15635
rect 14804 15604 14836 15605
rect 14804 15555 14836 15556
rect 14804 15525 14805 15555
rect 14805 15525 14835 15555
rect 14835 15525 14836 15555
rect 14804 15524 14836 15525
rect 14804 15475 14836 15476
rect 14804 15445 14805 15475
rect 14805 15445 14835 15475
rect 14835 15445 14836 15475
rect 14804 15444 14836 15445
rect 14804 15395 14836 15396
rect 14804 15365 14805 15395
rect 14805 15365 14835 15395
rect 14835 15365 14836 15395
rect 14804 15364 14836 15365
rect 14804 15315 14836 15316
rect 14804 15285 14805 15315
rect 14805 15285 14835 15315
rect 14835 15285 14836 15315
rect 14804 15284 14836 15285
rect 14804 15235 14836 15236
rect 14804 15205 14805 15235
rect 14805 15205 14835 15235
rect 14835 15205 14836 15235
rect 14804 15204 14836 15205
rect 14804 15155 14836 15156
rect 14804 15125 14805 15155
rect 14805 15125 14835 15155
rect 14835 15125 14836 15155
rect 14804 15124 14836 15125
rect 14804 15075 14836 15076
rect 14804 15045 14805 15075
rect 14805 15045 14835 15075
rect 14835 15045 14836 15075
rect 14804 15044 14836 15045
rect 14804 14995 14836 14996
rect 14804 14965 14805 14995
rect 14805 14965 14835 14995
rect 14835 14965 14836 14995
rect 14804 14964 14836 14965
rect 14804 14915 14836 14916
rect 14804 14885 14805 14915
rect 14805 14885 14835 14915
rect 14835 14885 14836 14915
rect 14804 14884 14836 14885
rect 14804 14835 14836 14836
rect 14804 14805 14805 14835
rect 14805 14805 14835 14835
rect 14835 14805 14836 14835
rect 14804 14804 14836 14805
rect 14804 14755 14836 14756
rect 14804 14725 14805 14755
rect 14805 14725 14835 14755
rect 14835 14725 14836 14755
rect 14804 14724 14836 14725
rect 14804 14675 14836 14676
rect 14804 14645 14805 14675
rect 14805 14645 14835 14675
rect 14835 14645 14836 14675
rect 14804 14644 14836 14645
rect 14804 14515 14836 14516
rect 14804 14485 14805 14515
rect 14805 14485 14835 14515
rect 14835 14485 14836 14515
rect 14804 14484 14836 14485
rect 14804 14435 14836 14436
rect 14804 14405 14805 14435
rect 14805 14405 14835 14435
rect 14835 14405 14836 14435
rect 14804 14404 14836 14405
rect 14804 14355 14836 14356
rect 14804 14325 14805 14355
rect 14805 14325 14835 14355
rect 14835 14325 14836 14355
rect 14804 14324 14836 14325
rect 14804 14275 14836 14276
rect 14804 14245 14805 14275
rect 14805 14245 14835 14275
rect 14835 14245 14836 14275
rect 14804 14244 14836 14245
rect 14804 14195 14836 14196
rect 14804 14165 14805 14195
rect 14805 14165 14835 14195
rect 14835 14165 14836 14195
rect 14804 14164 14836 14165
rect 14804 14115 14836 14116
rect 14804 14085 14805 14115
rect 14805 14085 14835 14115
rect 14835 14085 14836 14115
rect 14804 14084 14836 14085
rect 14804 14035 14836 14036
rect 14804 14005 14805 14035
rect 14805 14005 14835 14035
rect 14835 14005 14836 14035
rect 14804 14004 14836 14005
rect 14804 13955 14836 13956
rect 14804 13925 14805 13955
rect 14805 13925 14835 13955
rect 14835 13925 14836 13955
rect 14804 13924 14836 13925
rect 14804 13875 14836 13876
rect 14804 13845 14805 13875
rect 14805 13845 14835 13875
rect 14835 13845 14836 13875
rect 14804 13844 14836 13845
rect 14804 13795 14836 13796
rect 14804 13765 14805 13795
rect 14805 13765 14835 13795
rect 14835 13765 14836 13795
rect 14804 13764 14836 13765
rect 14804 13715 14836 13716
rect 14804 13685 14805 13715
rect 14805 13685 14835 13715
rect 14835 13685 14836 13715
rect 14804 13684 14836 13685
rect 14804 13635 14836 13636
rect 14804 13605 14805 13635
rect 14805 13605 14835 13635
rect 14835 13605 14836 13635
rect 14804 13604 14836 13605
rect 14804 13555 14836 13556
rect 14804 13525 14805 13555
rect 14805 13525 14835 13555
rect 14835 13525 14836 13555
rect 14804 13524 14836 13525
rect 14804 13475 14836 13476
rect 14804 13445 14805 13475
rect 14805 13445 14835 13475
rect 14835 13445 14836 13475
rect 14804 13444 14836 13445
rect 14804 13395 14836 13396
rect 14804 13365 14805 13395
rect 14805 13365 14835 13395
rect 14835 13365 14836 13395
rect 14804 13364 14836 13365
rect 14804 13315 14836 13316
rect 14804 13285 14805 13315
rect 14805 13285 14835 13315
rect 14835 13285 14836 13315
rect 14804 13284 14836 13285
rect 14804 13235 14836 13236
rect 14804 13205 14805 13235
rect 14805 13205 14835 13235
rect 14835 13205 14836 13235
rect 14804 13204 14836 13205
rect 14804 13155 14836 13156
rect 14804 13125 14805 13155
rect 14805 13125 14835 13155
rect 14835 13125 14836 13155
rect 14804 13124 14836 13125
rect 14804 13075 14836 13076
rect 14804 13045 14805 13075
rect 14805 13045 14835 13075
rect 14835 13045 14836 13075
rect 14804 13044 14836 13045
rect 14804 12995 14836 12996
rect 14804 12965 14805 12995
rect 14805 12965 14835 12995
rect 14835 12965 14836 12995
rect 14804 12964 14836 12965
rect 14804 12915 14836 12916
rect 14804 12885 14805 12915
rect 14805 12885 14835 12915
rect 14835 12885 14836 12915
rect 14804 12884 14836 12885
rect 14804 12835 14836 12836
rect 14804 12805 14805 12835
rect 14805 12805 14835 12835
rect 14835 12805 14836 12835
rect 14804 12804 14836 12805
rect 14804 12755 14836 12756
rect 14804 12725 14805 12755
rect 14805 12725 14835 12755
rect 14835 12725 14836 12755
rect 14804 12724 14836 12725
rect 14804 12675 14836 12676
rect 14804 12645 14805 12675
rect 14805 12645 14835 12675
rect 14835 12645 14836 12675
rect 14804 12644 14836 12645
rect 14804 12595 14836 12596
rect 14804 12565 14805 12595
rect 14805 12565 14835 12595
rect 14835 12565 14836 12595
rect 14804 12564 14836 12565
rect 14804 12515 14836 12516
rect 14804 12485 14805 12515
rect 14805 12485 14835 12515
rect 14835 12485 14836 12515
rect 14804 12484 14836 12485
rect 14804 12435 14836 12436
rect 14804 12405 14805 12435
rect 14805 12405 14835 12435
rect 14835 12405 14836 12435
rect 14804 12404 14836 12405
rect 14804 12355 14836 12356
rect 14804 12325 14805 12355
rect 14805 12325 14835 12355
rect 14835 12325 14836 12355
rect 14804 12324 14836 12325
rect 14804 12275 14836 12276
rect 14804 12245 14805 12275
rect 14805 12245 14835 12275
rect 14835 12245 14836 12275
rect 14804 12244 14836 12245
rect 14804 12195 14836 12196
rect 14804 12165 14805 12195
rect 14805 12165 14835 12195
rect 14835 12165 14836 12195
rect 14804 12164 14836 12165
rect 14804 12115 14836 12116
rect 14804 12085 14805 12115
rect 14805 12085 14835 12115
rect 14835 12085 14836 12115
rect 14804 12084 14836 12085
rect 14804 12035 14836 12036
rect 14804 12005 14805 12035
rect 14805 12005 14835 12035
rect 14835 12005 14836 12035
rect 14804 12004 14836 12005
rect 14804 11955 14836 11956
rect 14804 11925 14805 11955
rect 14805 11925 14835 11955
rect 14835 11925 14836 11955
rect 14804 11924 14836 11925
rect 14804 11875 14836 11876
rect 14804 11845 14805 11875
rect 14805 11845 14835 11875
rect 14835 11845 14836 11875
rect 14804 11844 14836 11845
rect 14804 11795 14836 11796
rect 14804 11765 14805 11795
rect 14805 11765 14835 11795
rect 14835 11765 14836 11795
rect 14804 11764 14836 11765
rect 14804 11635 14836 11636
rect 14804 11605 14805 11635
rect 14805 11605 14835 11635
rect 14835 11605 14836 11635
rect 14804 11604 14836 11605
rect 14804 11555 14836 11556
rect 14804 11525 14805 11555
rect 14805 11525 14835 11555
rect 14835 11525 14836 11555
rect 14804 11524 14836 11525
rect 14804 11475 14836 11476
rect 14804 11445 14805 11475
rect 14805 11445 14835 11475
rect 14835 11445 14836 11475
rect 14804 11444 14836 11445
rect 14804 11395 14836 11396
rect 14804 11365 14805 11395
rect 14805 11365 14835 11395
rect 14835 11365 14836 11395
rect 14804 11364 14836 11365
rect 14804 11315 14836 11316
rect 14804 11285 14805 11315
rect 14805 11285 14835 11315
rect 14835 11285 14836 11315
rect 14804 11284 14836 11285
rect 14804 11235 14836 11236
rect 14804 11205 14805 11235
rect 14805 11205 14835 11235
rect 14835 11205 14836 11235
rect 14804 11204 14836 11205
rect 14804 11155 14836 11156
rect 14804 11125 14805 11155
rect 14805 11125 14835 11155
rect 14835 11125 14836 11155
rect 14804 11124 14836 11125
rect 14804 11075 14836 11076
rect 14804 11045 14805 11075
rect 14805 11045 14835 11075
rect 14835 11045 14836 11075
rect 14804 11044 14836 11045
rect 14804 10995 14836 10996
rect 14804 10965 14805 10995
rect 14805 10965 14835 10995
rect 14835 10965 14836 10995
rect 14804 10964 14836 10965
rect 14804 10915 14836 10916
rect 14804 10885 14805 10915
rect 14805 10885 14835 10915
rect 14835 10885 14836 10915
rect 14804 10884 14836 10885
rect 14804 10835 14836 10836
rect 14804 10805 14805 10835
rect 14805 10805 14835 10835
rect 14835 10805 14836 10835
rect 14804 10804 14836 10805
rect 14804 10755 14836 10756
rect 14804 10725 14805 10755
rect 14805 10725 14835 10755
rect 14835 10725 14836 10755
rect 14804 10724 14836 10725
rect 14804 10675 14836 10676
rect 14804 10645 14805 10675
rect 14805 10645 14835 10675
rect 14835 10645 14836 10675
rect 14804 10644 14836 10645
rect 14804 10595 14836 10596
rect 14804 10565 14805 10595
rect 14805 10565 14835 10595
rect 14835 10565 14836 10595
rect 14804 10564 14836 10565
rect 14804 10515 14836 10516
rect 14804 10485 14805 10515
rect 14805 10485 14835 10515
rect 14835 10485 14836 10515
rect 14804 10484 14836 10485
rect 14804 10435 14836 10436
rect 14804 10405 14805 10435
rect 14805 10405 14835 10435
rect 14835 10405 14836 10435
rect 14804 10404 14836 10405
rect 14804 10355 14836 10356
rect 14804 10325 14805 10355
rect 14805 10325 14835 10355
rect 14835 10325 14836 10355
rect 14804 10324 14836 10325
rect 14804 10275 14836 10276
rect 14804 10245 14805 10275
rect 14805 10245 14835 10275
rect 14835 10245 14836 10275
rect 14804 10244 14836 10245
rect 14804 10195 14836 10196
rect 14804 10165 14805 10195
rect 14805 10165 14835 10195
rect 14835 10165 14836 10195
rect 14804 10164 14836 10165
rect 14804 10115 14836 10116
rect 14804 10085 14805 10115
rect 14805 10085 14835 10115
rect 14835 10085 14836 10115
rect 14804 10084 14836 10085
rect 14804 10035 14836 10036
rect 14804 10005 14805 10035
rect 14805 10005 14835 10035
rect 14835 10005 14836 10035
rect 14804 10004 14836 10005
rect 14804 9955 14836 9956
rect 14804 9925 14805 9955
rect 14805 9925 14835 9955
rect 14835 9925 14836 9955
rect 14804 9924 14836 9925
rect 14804 9875 14836 9876
rect 14804 9845 14805 9875
rect 14805 9845 14835 9875
rect 14835 9845 14836 9875
rect 14804 9844 14836 9845
rect 14804 9795 14836 9796
rect 14804 9765 14805 9795
rect 14805 9765 14835 9795
rect 14835 9765 14836 9795
rect 14804 9764 14836 9765
rect 14804 9715 14836 9716
rect 14804 9685 14805 9715
rect 14805 9685 14835 9715
rect 14835 9685 14836 9715
rect 14804 9684 14836 9685
rect 14804 9635 14836 9636
rect 14804 9605 14805 9635
rect 14805 9605 14835 9635
rect 14835 9605 14836 9635
rect 14804 9604 14836 9605
rect 14804 9555 14836 9556
rect 14804 9525 14805 9555
rect 14805 9525 14835 9555
rect 14835 9525 14836 9555
rect 14804 9524 14836 9525
rect 14804 9475 14836 9476
rect 14804 9445 14805 9475
rect 14805 9445 14835 9475
rect 14835 9445 14836 9475
rect 14804 9444 14836 9445
rect 14804 9395 14836 9396
rect 14804 9365 14805 9395
rect 14805 9365 14835 9395
rect 14835 9365 14836 9395
rect 14804 9364 14836 9365
rect 14804 9315 14836 9316
rect 14804 9285 14805 9315
rect 14805 9285 14835 9315
rect 14835 9285 14836 9315
rect 14804 9284 14836 9285
rect 14804 9235 14836 9236
rect 14804 9205 14805 9235
rect 14805 9205 14835 9235
rect 14835 9205 14836 9235
rect 14804 9204 14836 9205
rect 14804 9155 14836 9156
rect 14804 9125 14805 9155
rect 14805 9125 14835 9155
rect 14835 9125 14836 9155
rect 14804 9124 14836 9125
rect 14804 9075 14836 9076
rect 14804 9045 14805 9075
rect 14805 9045 14835 9075
rect 14835 9045 14836 9075
rect 14804 9044 14836 9045
rect 14804 8995 14836 8996
rect 14804 8965 14805 8995
rect 14805 8965 14835 8995
rect 14835 8965 14836 8995
rect 14804 8964 14836 8965
rect 14804 8915 14836 8916
rect 14804 8885 14805 8915
rect 14805 8885 14835 8915
rect 14835 8885 14836 8915
rect 14804 8884 14836 8885
rect 14804 8835 14836 8836
rect 14804 8805 14805 8835
rect 14805 8805 14835 8835
rect 14835 8805 14836 8835
rect 14804 8804 14836 8805
rect 14804 8755 14836 8756
rect 14804 8725 14805 8755
rect 14805 8725 14835 8755
rect 14835 8725 14836 8755
rect 14804 8724 14836 8725
rect 14804 8675 14836 8676
rect 14804 8645 14805 8675
rect 14805 8645 14835 8675
rect 14835 8645 14836 8675
rect 14804 8644 14836 8645
rect 14804 8595 14836 8596
rect 14804 8565 14805 8595
rect 14805 8565 14835 8595
rect 14835 8565 14836 8595
rect 14804 8564 14836 8565
rect 14804 8515 14836 8516
rect 14804 8485 14805 8515
rect 14805 8485 14835 8515
rect 14835 8485 14836 8515
rect 14804 8484 14836 8485
rect 14804 8435 14836 8436
rect 14804 8405 14805 8435
rect 14805 8405 14835 8435
rect 14835 8405 14836 8435
rect 14804 8404 14836 8405
rect 14804 8355 14836 8356
rect 14804 8325 14805 8355
rect 14805 8325 14835 8355
rect 14835 8325 14836 8355
rect 14804 8324 14836 8325
rect 14804 8275 14836 8276
rect 14804 8245 14805 8275
rect 14805 8245 14835 8275
rect 14835 8245 14836 8275
rect 14804 8244 14836 8245
rect 14804 8195 14836 8196
rect 14804 8165 14805 8195
rect 14805 8165 14835 8195
rect 14835 8165 14836 8195
rect 14804 8164 14836 8165
rect 14804 8115 14836 8116
rect 14804 8085 14805 8115
rect 14805 8085 14835 8115
rect 14835 8085 14836 8115
rect 14804 8084 14836 8085
rect 14804 8035 14836 8036
rect 14804 8005 14805 8035
rect 14805 8005 14835 8035
rect 14835 8005 14836 8035
rect 14804 8004 14836 8005
rect 14804 7955 14836 7956
rect 14804 7925 14805 7955
rect 14805 7925 14835 7955
rect 14835 7925 14836 7955
rect 14804 7924 14836 7925
rect 14804 7875 14836 7876
rect 14804 7845 14805 7875
rect 14805 7845 14835 7875
rect 14835 7845 14836 7875
rect 14804 7844 14836 7845
rect 14804 7795 14836 7796
rect 14804 7765 14805 7795
rect 14805 7765 14835 7795
rect 14835 7765 14836 7795
rect 14804 7764 14836 7765
rect 14804 7715 14836 7716
rect 14804 7685 14805 7715
rect 14805 7685 14835 7715
rect 14835 7685 14836 7715
rect 14804 7684 14836 7685
rect 14804 7635 14836 7636
rect 14804 7605 14805 7635
rect 14805 7605 14835 7635
rect 14835 7605 14836 7635
rect 14804 7604 14836 7605
rect 14804 7555 14836 7556
rect 14804 7525 14805 7555
rect 14805 7525 14835 7555
rect 14835 7525 14836 7555
rect 14804 7524 14836 7525
rect 14804 7475 14836 7476
rect 14804 7445 14805 7475
rect 14805 7445 14835 7475
rect 14835 7445 14836 7475
rect 14804 7444 14836 7445
rect 14804 7395 14836 7396
rect 14804 7365 14805 7395
rect 14805 7365 14835 7395
rect 14835 7365 14836 7395
rect 14804 7364 14836 7365
rect 14804 7315 14836 7316
rect 14804 7285 14805 7315
rect 14805 7285 14835 7315
rect 14835 7285 14836 7315
rect 14804 7284 14836 7285
rect 14804 7235 14836 7236
rect 14804 7205 14805 7235
rect 14805 7205 14835 7235
rect 14835 7205 14836 7235
rect 14804 7204 14836 7205
rect 14804 7155 14836 7156
rect 14804 7125 14805 7155
rect 14805 7125 14835 7155
rect 14835 7125 14836 7155
rect 14804 7124 14836 7125
rect 14804 7075 14836 7076
rect 14804 7045 14805 7075
rect 14805 7045 14835 7075
rect 14835 7045 14836 7075
rect 14804 7044 14836 7045
rect 14804 6995 14836 6996
rect 14804 6965 14805 6995
rect 14805 6965 14835 6995
rect 14835 6965 14836 6995
rect 14804 6964 14836 6965
rect 14804 6915 14836 6916
rect 14804 6885 14805 6915
rect 14805 6885 14835 6915
rect 14835 6885 14836 6915
rect 14804 6884 14836 6885
rect 14804 6835 14836 6836
rect 14804 6805 14805 6835
rect 14805 6805 14835 6835
rect 14835 6805 14836 6835
rect 14804 6804 14836 6805
rect 14804 6755 14836 6756
rect 14804 6725 14805 6755
rect 14805 6725 14835 6755
rect 14835 6725 14836 6755
rect 14804 6724 14836 6725
rect 14804 6675 14836 6676
rect 14804 6645 14805 6675
rect 14805 6645 14835 6675
rect 14835 6645 14836 6675
rect 14804 6644 14836 6645
rect 14804 6595 14836 6596
rect 14804 6565 14805 6595
rect 14805 6565 14835 6595
rect 14835 6565 14836 6595
rect 14804 6564 14836 6565
rect 14804 6515 14836 6516
rect 14804 6485 14805 6515
rect 14805 6485 14835 6515
rect 14835 6485 14836 6515
rect 14804 6484 14836 6485
rect 14804 6435 14836 6436
rect 14804 6405 14805 6435
rect 14805 6405 14835 6435
rect 14835 6405 14836 6435
rect 14804 6404 14836 6405
rect 14804 6355 14836 6356
rect 14804 6325 14805 6355
rect 14805 6325 14835 6355
rect 14835 6325 14836 6355
rect 14804 6324 14836 6325
rect 14804 6275 14836 6276
rect 14804 6245 14805 6275
rect 14805 6245 14835 6275
rect 14835 6245 14836 6275
rect 14804 6244 14836 6245
rect 14804 6195 14836 6196
rect 14804 6165 14805 6195
rect 14805 6165 14835 6195
rect 14835 6165 14836 6195
rect 14804 6164 14836 6165
rect 14804 6115 14836 6116
rect 14804 6085 14805 6115
rect 14805 6085 14835 6115
rect 14835 6085 14836 6115
rect 14804 6084 14836 6085
rect 14804 6035 14836 6036
rect 14804 6005 14805 6035
rect 14805 6005 14835 6035
rect 14835 6005 14836 6035
rect 14804 6004 14836 6005
rect 14804 5955 14836 5956
rect 14804 5925 14805 5955
rect 14805 5925 14835 5955
rect 14835 5925 14836 5955
rect 14804 5924 14836 5925
rect 14804 5875 14836 5876
rect 14804 5845 14805 5875
rect 14805 5845 14835 5875
rect 14835 5845 14836 5875
rect 14804 5844 14836 5845
rect 14804 5795 14836 5796
rect 14804 5765 14805 5795
rect 14805 5765 14835 5795
rect 14835 5765 14836 5795
rect 14804 5764 14836 5765
rect 14804 5715 14836 5716
rect 14804 5685 14805 5715
rect 14805 5685 14835 5715
rect 14835 5685 14836 5715
rect 14804 5684 14836 5685
rect 14804 5635 14836 5636
rect 14804 5605 14805 5635
rect 14805 5605 14835 5635
rect 14835 5605 14836 5635
rect 14804 5604 14836 5605
rect 14804 5555 14836 5556
rect 14804 5525 14805 5555
rect 14805 5525 14835 5555
rect 14835 5525 14836 5555
rect 14804 5524 14836 5525
rect 14804 5475 14836 5476
rect 14804 5445 14805 5475
rect 14805 5445 14835 5475
rect 14835 5445 14836 5475
rect 14804 5444 14836 5445
rect 14804 5395 14836 5396
rect 14804 5365 14805 5395
rect 14805 5365 14835 5395
rect 14835 5365 14836 5395
rect 14804 5364 14836 5365
rect 14804 5315 14836 5316
rect 14804 5285 14805 5315
rect 14805 5285 14835 5315
rect 14835 5285 14836 5315
rect 14804 5284 14836 5285
rect 14804 5235 14836 5236
rect 14804 5205 14805 5235
rect 14805 5205 14835 5235
rect 14835 5205 14836 5235
rect 14804 5204 14836 5205
rect 14804 5155 14836 5156
rect 14804 5125 14805 5155
rect 14805 5125 14835 5155
rect 14835 5125 14836 5155
rect 14804 5124 14836 5125
rect 14804 5075 14836 5076
rect 14804 5045 14805 5075
rect 14805 5045 14835 5075
rect 14835 5045 14836 5075
rect 14804 5044 14836 5045
rect 14804 4995 14836 4996
rect 14804 4965 14805 4995
rect 14805 4965 14835 4995
rect 14835 4965 14836 4995
rect 14804 4964 14836 4965
rect 14804 4915 14836 4916
rect 14804 4885 14805 4915
rect 14805 4885 14835 4915
rect 14835 4885 14836 4915
rect 14804 4884 14836 4885
rect 14804 4835 14836 4836
rect 14804 4805 14805 4835
rect 14805 4805 14835 4835
rect 14835 4805 14836 4835
rect 14804 4804 14836 4805
rect 14804 4675 14836 4676
rect 14804 4645 14805 4675
rect 14805 4645 14835 4675
rect 14835 4645 14836 4675
rect 14804 4644 14836 4645
rect 14804 4595 14836 4596
rect 14804 4565 14805 4595
rect 14805 4565 14835 4595
rect 14835 4565 14836 4595
rect 14804 4564 14836 4565
rect 14804 4515 14836 4516
rect 14804 4485 14805 4515
rect 14805 4485 14835 4515
rect 14835 4485 14836 4515
rect 14804 4484 14836 4485
rect 14804 4435 14836 4436
rect 14804 4405 14805 4435
rect 14805 4405 14835 4435
rect 14835 4405 14836 4435
rect 14804 4404 14836 4405
rect 14804 4355 14836 4356
rect 14804 4325 14805 4355
rect 14805 4325 14835 4355
rect 14835 4325 14836 4355
rect 14804 4324 14836 4325
rect 14804 4275 14836 4276
rect 14804 4245 14805 4275
rect 14805 4245 14835 4275
rect 14835 4245 14836 4275
rect 14804 4244 14836 4245
rect 14804 4195 14836 4196
rect 14804 4165 14805 4195
rect 14805 4165 14835 4195
rect 14835 4165 14836 4195
rect 14804 4164 14836 4165
rect 14804 4115 14836 4116
rect 14804 4085 14805 4115
rect 14805 4085 14835 4115
rect 14835 4085 14836 4115
rect 14804 4084 14836 4085
rect 14804 4035 14836 4036
rect 14804 4005 14805 4035
rect 14805 4005 14835 4035
rect 14835 4005 14836 4035
rect 14804 4004 14836 4005
rect 14804 3955 14836 3956
rect 14804 3925 14805 3955
rect 14805 3925 14835 3955
rect 14835 3925 14836 3955
rect 14804 3924 14836 3925
rect 14804 3875 14836 3876
rect 14804 3845 14805 3875
rect 14805 3845 14835 3875
rect 14835 3845 14836 3875
rect 14804 3844 14836 3845
rect 14804 3795 14836 3796
rect 14804 3765 14805 3795
rect 14805 3765 14835 3795
rect 14835 3765 14836 3795
rect 14804 3764 14836 3765
rect 14804 3715 14836 3716
rect 14804 3685 14805 3715
rect 14805 3685 14835 3715
rect 14835 3685 14836 3715
rect 14804 3684 14836 3685
rect 14804 3635 14836 3636
rect 14804 3605 14805 3635
rect 14805 3605 14835 3635
rect 14835 3605 14836 3635
rect 14804 3604 14836 3605
rect 14804 3555 14836 3556
rect 14804 3525 14805 3555
rect 14805 3525 14835 3555
rect 14835 3525 14836 3555
rect 14804 3524 14836 3525
rect 14804 3475 14836 3476
rect 14804 3445 14805 3475
rect 14805 3445 14835 3475
rect 14835 3445 14836 3475
rect 14804 3444 14836 3445
rect 14804 3395 14836 3396
rect 14804 3365 14805 3395
rect 14805 3365 14835 3395
rect 14835 3365 14836 3395
rect 14804 3364 14836 3365
rect 14804 3315 14836 3316
rect 14804 3285 14805 3315
rect 14805 3285 14835 3315
rect 14835 3285 14836 3315
rect 14804 3284 14836 3285
rect 14804 3235 14836 3236
rect 14804 3205 14805 3235
rect 14805 3205 14835 3235
rect 14835 3205 14836 3235
rect 14804 3204 14836 3205
rect 14804 3155 14836 3156
rect 14804 3125 14805 3155
rect 14805 3125 14835 3155
rect 14835 3125 14836 3155
rect 14804 3124 14836 3125
rect 14804 3075 14836 3076
rect 14804 3045 14805 3075
rect 14805 3045 14835 3075
rect 14835 3045 14836 3075
rect 14804 3044 14836 3045
rect 14804 2995 14836 2996
rect 14804 2965 14805 2995
rect 14805 2965 14835 2995
rect 14835 2965 14836 2995
rect 14804 2964 14836 2965
rect 14804 2915 14836 2916
rect 14804 2885 14805 2915
rect 14805 2885 14835 2915
rect 14835 2885 14836 2915
rect 14804 2884 14836 2885
rect 14804 2835 14836 2836
rect 14804 2805 14805 2835
rect 14805 2805 14835 2835
rect 14835 2805 14836 2835
rect 14804 2804 14836 2805
rect 14804 2755 14836 2756
rect 14804 2725 14805 2755
rect 14805 2725 14835 2755
rect 14835 2725 14836 2755
rect 14804 2724 14836 2725
rect 14804 2675 14836 2676
rect 14804 2645 14805 2675
rect 14805 2645 14835 2675
rect 14835 2645 14836 2675
rect 14804 2644 14836 2645
rect 14804 2595 14836 2596
rect 14804 2565 14805 2595
rect 14805 2565 14835 2595
rect 14835 2565 14836 2595
rect 14804 2564 14836 2565
rect 14804 2515 14836 2516
rect 14804 2485 14805 2515
rect 14805 2485 14835 2515
rect 14835 2485 14836 2515
rect 14804 2484 14836 2485
rect 14804 2435 14836 2436
rect 14804 2405 14805 2435
rect 14805 2405 14835 2435
rect 14835 2405 14836 2435
rect 14804 2404 14836 2405
rect 14804 2355 14836 2356
rect 14804 2325 14805 2355
rect 14805 2325 14835 2355
rect 14835 2325 14836 2355
rect 14804 2324 14836 2325
rect 14804 2275 14836 2276
rect 14804 2245 14805 2275
rect 14805 2245 14835 2275
rect 14835 2245 14836 2275
rect 14804 2244 14836 2245
rect 14804 2195 14836 2196
rect 14804 2165 14805 2195
rect 14805 2165 14835 2195
rect 14835 2165 14836 2195
rect 14804 2164 14836 2165
rect 14804 2115 14836 2116
rect 14804 2085 14805 2115
rect 14805 2085 14835 2115
rect 14835 2085 14836 2115
rect 14804 2084 14836 2085
rect 14804 2035 14836 2036
rect 14804 2005 14805 2035
rect 14805 2005 14835 2035
rect 14835 2005 14836 2035
rect 14804 2004 14836 2005
rect 14804 1955 14836 1956
rect 14804 1925 14805 1955
rect 14805 1925 14835 1955
rect 14835 1925 14836 1955
rect 14804 1924 14836 1925
rect 14804 1795 14836 1796
rect 14804 1765 14805 1795
rect 14805 1765 14835 1795
rect 14835 1765 14836 1795
rect 14804 1764 14836 1765
rect 14804 1715 14836 1716
rect 14804 1685 14805 1715
rect 14805 1685 14835 1715
rect 14835 1685 14836 1715
rect 14804 1684 14836 1685
rect 14804 1635 14836 1636
rect 14804 1605 14805 1635
rect 14805 1605 14835 1635
rect 14835 1605 14836 1635
rect 14804 1604 14836 1605
rect 14804 1555 14836 1556
rect 14804 1525 14805 1555
rect 14805 1525 14835 1555
rect 14835 1525 14836 1555
rect 14804 1524 14836 1525
rect 14804 1475 14836 1476
rect 14804 1445 14805 1475
rect 14805 1445 14835 1475
rect 14835 1445 14836 1475
rect 14804 1444 14836 1445
rect 14804 1395 14836 1396
rect 14804 1365 14805 1395
rect 14805 1365 14835 1395
rect 14835 1365 14836 1395
rect 14804 1364 14836 1365
rect 14804 1315 14836 1316
rect 14804 1285 14805 1315
rect 14805 1285 14835 1315
rect 14835 1285 14836 1315
rect 14804 1284 14836 1285
rect 14804 1235 14836 1236
rect 14804 1205 14805 1235
rect 14805 1205 14835 1235
rect 14835 1205 14836 1235
rect 14804 1204 14836 1205
rect 14804 1155 14836 1156
rect 14804 1125 14805 1155
rect 14805 1125 14835 1155
rect 14835 1125 14836 1155
rect 14804 1124 14836 1125
rect 14804 1075 14836 1076
rect 14804 1045 14805 1075
rect 14805 1045 14835 1075
rect 14835 1045 14836 1075
rect 14804 1044 14836 1045
rect 14804 995 14836 996
rect 14804 965 14805 995
rect 14805 965 14835 995
rect 14835 965 14836 995
rect 14804 964 14836 965
rect 14804 915 14836 916
rect 14804 885 14805 915
rect 14805 885 14835 915
rect 14835 885 14836 915
rect 14804 884 14836 885
rect 14804 835 14836 836
rect 14804 805 14805 835
rect 14805 805 14835 835
rect 14835 805 14836 835
rect 14804 804 14836 805
rect 14804 755 14836 756
rect 14804 725 14805 755
rect 14805 725 14835 755
rect 14835 725 14836 755
rect 14804 724 14836 725
rect 14804 675 14836 676
rect 14804 645 14805 675
rect 14805 645 14835 675
rect 14835 645 14836 675
rect 14804 644 14836 645
rect 14804 595 14836 596
rect 14804 565 14805 595
rect 14805 565 14835 595
rect 14835 565 14836 595
rect 14804 564 14836 565
rect 14804 515 14836 516
rect 14804 485 14805 515
rect 14805 485 14835 515
rect 14835 485 14836 515
rect 14804 484 14836 485
rect 14644 244 14676 436
rect 14884 14564 14916 14596
rect 14884 11684 14916 11716
rect 14884 4724 14916 4756
rect 14884 1844 14916 1876
rect 14964 15955 14996 15956
rect 14964 15925 14965 15955
rect 14965 15925 14995 15955
rect 14995 15925 14996 15955
rect 14964 15924 14996 15925
rect 14964 15875 14996 15876
rect 14964 15845 14965 15875
rect 14965 15845 14995 15875
rect 14995 15845 14996 15875
rect 14964 15844 14996 15845
rect 14964 15795 14996 15796
rect 14964 15765 14965 15795
rect 14965 15765 14995 15795
rect 14995 15765 14996 15795
rect 14964 15764 14996 15765
rect 14964 15715 14996 15716
rect 14964 15685 14965 15715
rect 14965 15685 14995 15715
rect 14995 15685 14996 15715
rect 14964 15684 14996 15685
rect 14964 15635 14996 15636
rect 14964 15605 14965 15635
rect 14965 15605 14995 15635
rect 14995 15605 14996 15635
rect 14964 15604 14996 15605
rect 14964 15555 14996 15556
rect 14964 15525 14965 15555
rect 14965 15525 14995 15555
rect 14995 15525 14996 15555
rect 14964 15524 14996 15525
rect 14964 15475 14996 15476
rect 14964 15445 14965 15475
rect 14965 15445 14995 15475
rect 14995 15445 14996 15475
rect 14964 15444 14996 15445
rect 14964 15395 14996 15396
rect 14964 15365 14965 15395
rect 14965 15365 14995 15395
rect 14995 15365 14996 15395
rect 14964 15364 14996 15365
rect 14964 15315 14996 15316
rect 14964 15285 14965 15315
rect 14965 15285 14995 15315
rect 14995 15285 14996 15315
rect 14964 15284 14996 15285
rect 14964 15235 14996 15236
rect 14964 15205 14965 15235
rect 14965 15205 14995 15235
rect 14995 15205 14996 15235
rect 14964 15204 14996 15205
rect 14964 15155 14996 15156
rect 14964 15125 14965 15155
rect 14965 15125 14995 15155
rect 14995 15125 14996 15155
rect 14964 15124 14996 15125
rect 14964 15075 14996 15076
rect 14964 15045 14965 15075
rect 14965 15045 14995 15075
rect 14995 15045 14996 15075
rect 14964 15044 14996 15045
rect 14964 14995 14996 14996
rect 14964 14965 14965 14995
rect 14965 14965 14995 14995
rect 14995 14965 14996 14995
rect 14964 14964 14996 14965
rect 14964 14915 14996 14916
rect 14964 14885 14965 14915
rect 14965 14885 14995 14915
rect 14995 14885 14996 14915
rect 14964 14884 14996 14885
rect 14964 14835 14996 14836
rect 14964 14805 14965 14835
rect 14965 14805 14995 14835
rect 14995 14805 14996 14835
rect 14964 14804 14996 14805
rect 14964 14755 14996 14756
rect 14964 14725 14965 14755
rect 14965 14725 14995 14755
rect 14995 14725 14996 14755
rect 14964 14724 14996 14725
rect 14964 14675 14996 14676
rect 14964 14645 14965 14675
rect 14965 14645 14995 14675
rect 14995 14645 14996 14675
rect 14964 14644 14996 14645
rect 14964 14515 14996 14516
rect 14964 14485 14965 14515
rect 14965 14485 14995 14515
rect 14995 14485 14996 14515
rect 14964 14484 14996 14485
rect 14964 14435 14996 14436
rect 14964 14405 14965 14435
rect 14965 14405 14995 14435
rect 14995 14405 14996 14435
rect 14964 14404 14996 14405
rect 14964 14355 14996 14356
rect 14964 14325 14965 14355
rect 14965 14325 14995 14355
rect 14995 14325 14996 14355
rect 14964 14324 14996 14325
rect 14964 14275 14996 14276
rect 14964 14245 14965 14275
rect 14965 14245 14995 14275
rect 14995 14245 14996 14275
rect 14964 14244 14996 14245
rect 14964 14195 14996 14196
rect 14964 14165 14965 14195
rect 14965 14165 14995 14195
rect 14995 14165 14996 14195
rect 14964 14164 14996 14165
rect 14964 14115 14996 14116
rect 14964 14085 14965 14115
rect 14965 14085 14995 14115
rect 14995 14085 14996 14115
rect 14964 14084 14996 14085
rect 14964 14035 14996 14036
rect 14964 14005 14965 14035
rect 14965 14005 14995 14035
rect 14995 14005 14996 14035
rect 14964 14004 14996 14005
rect 14964 13955 14996 13956
rect 14964 13925 14965 13955
rect 14965 13925 14995 13955
rect 14995 13925 14996 13955
rect 14964 13924 14996 13925
rect 14964 13875 14996 13876
rect 14964 13845 14965 13875
rect 14965 13845 14995 13875
rect 14995 13845 14996 13875
rect 14964 13844 14996 13845
rect 14964 13795 14996 13796
rect 14964 13765 14965 13795
rect 14965 13765 14995 13795
rect 14995 13765 14996 13795
rect 14964 13764 14996 13765
rect 14964 13715 14996 13716
rect 14964 13685 14965 13715
rect 14965 13685 14995 13715
rect 14995 13685 14996 13715
rect 14964 13684 14996 13685
rect 14964 13635 14996 13636
rect 14964 13605 14965 13635
rect 14965 13605 14995 13635
rect 14995 13605 14996 13635
rect 14964 13604 14996 13605
rect 14964 13555 14996 13556
rect 14964 13525 14965 13555
rect 14965 13525 14995 13555
rect 14995 13525 14996 13555
rect 14964 13524 14996 13525
rect 14964 13475 14996 13476
rect 14964 13445 14965 13475
rect 14965 13445 14995 13475
rect 14995 13445 14996 13475
rect 14964 13444 14996 13445
rect 14964 13395 14996 13396
rect 14964 13365 14965 13395
rect 14965 13365 14995 13395
rect 14995 13365 14996 13395
rect 14964 13364 14996 13365
rect 14964 13315 14996 13316
rect 14964 13285 14965 13315
rect 14965 13285 14995 13315
rect 14995 13285 14996 13315
rect 14964 13284 14996 13285
rect 14964 13235 14996 13236
rect 14964 13205 14965 13235
rect 14965 13205 14995 13235
rect 14995 13205 14996 13235
rect 14964 13204 14996 13205
rect 14964 13155 14996 13156
rect 14964 13125 14965 13155
rect 14965 13125 14995 13155
rect 14995 13125 14996 13155
rect 14964 13124 14996 13125
rect 14964 13075 14996 13076
rect 14964 13045 14965 13075
rect 14965 13045 14995 13075
rect 14995 13045 14996 13075
rect 14964 13044 14996 13045
rect 14964 12995 14996 12996
rect 14964 12965 14965 12995
rect 14965 12965 14995 12995
rect 14995 12965 14996 12995
rect 14964 12964 14996 12965
rect 14964 12915 14996 12916
rect 14964 12885 14965 12915
rect 14965 12885 14995 12915
rect 14995 12885 14996 12915
rect 14964 12884 14996 12885
rect 14964 12835 14996 12836
rect 14964 12805 14965 12835
rect 14965 12805 14995 12835
rect 14995 12805 14996 12835
rect 14964 12804 14996 12805
rect 14964 12755 14996 12756
rect 14964 12725 14965 12755
rect 14965 12725 14995 12755
rect 14995 12725 14996 12755
rect 14964 12724 14996 12725
rect 14964 12675 14996 12676
rect 14964 12645 14965 12675
rect 14965 12645 14995 12675
rect 14995 12645 14996 12675
rect 14964 12644 14996 12645
rect 14964 12595 14996 12596
rect 14964 12565 14965 12595
rect 14965 12565 14995 12595
rect 14995 12565 14996 12595
rect 14964 12564 14996 12565
rect 14964 12515 14996 12516
rect 14964 12485 14965 12515
rect 14965 12485 14995 12515
rect 14995 12485 14996 12515
rect 14964 12484 14996 12485
rect 14964 12435 14996 12436
rect 14964 12405 14965 12435
rect 14965 12405 14995 12435
rect 14995 12405 14996 12435
rect 14964 12404 14996 12405
rect 14964 12355 14996 12356
rect 14964 12325 14965 12355
rect 14965 12325 14995 12355
rect 14995 12325 14996 12355
rect 14964 12324 14996 12325
rect 14964 12275 14996 12276
rect 14964 12245 14965 12275
rect 14965 12245 14995 12275
rect 14995 12245 14996 12275
rect 14964 12244 14996 12245
rect 14964 12195 14996 12196
rect 14964 12165 14965 12195
rect 14965 12165 14995 12195
rect 14995 12165 14996 12195
rect 14964 12164 14996 12165
rect 14964 12115 14996 12116
rect 14964 12085 14965 12115
rect 14965 12085 14995 12115
rect 14995 12085 14996 12115
rect 14964 12084 14996 12085
rect 14964 12035 14996 12036
rect 14964 12005 14965 12035
rect 14965 12005 14995 12035
rect 14995 12005 14996 12035
rect 14964 12004 14996 12005
rect 14964 11955 14996 11956
rect 14964 11925 14965 11955
rect 14965 11925 14995 11955
rect 14995 11925 14996 11955
rect 14964 11924 14996 11925
rect 14964 11875 14996 11876
rect 14964 11845 14965 11875
rect 14965 11845 14995 11875
rect 14995 11845 14996 11875
rect 14964 11844 14996 11845
rect 14964 11795 14996 11796
rect 14964 11765 14965 11795
rect 14965 11765 14995 11795
rect 14995 11765 14996 11795
rect 14964 11764 14996 11765
rect 14964 11635 14996 11636
rect 14964 11605 14965 11635
rect 14965 11605 14995 11635
rect 14995 11605 14996 11635
rect 14964 11604 14996 11605
rect 14964 11555 14996 11556
rect 14964 11525 14965 11555
rect 14965 11525 14995 11555
rect 14995 11525 14996 11555
rect 14964 11524 14996 11525
rect 14964 11475 14996 11476
rect 14964 11445 14965 11475
rect 14965 11445 14995 11475
rect 14995 11445 14996 11475
rect 14964 11444 14996 11445
rect 14964 11395 14996 11396
rect 14964 11365 14965 11395
rect 14965 11365 14995 11395
rect 14995 11365 14996 11395
rect 14964 11364 14996 11365
rect 14964 11315 14996 11316
rect 14964 11285 14965 11315
rect 14965 11285 14995 11315
rect 14995 11285 14996 11315
rect 14964 11284 14996 11285
rect 14964 11235 14996 11236
rect 14964 11205 14965 11235
rect 14965 11205 14995 11235
rect 14995 11205 14996 11235
rect 14964 11204 14996 11205
rect 14964 11155 14996 11156
rect 14964 11125 14965 11155
rect 14965 11125 14995 11155
rect 14995 11125 14996 11155
rect 14964 11124 14996 11125
rect 14964 11075 14996 11076
rect 14964 11045 14965 11075
rect 14965 11045 14995 11075
rect 14995 11045 14996 11075
rect 14964 11044 14996 11045
rect 14964 10995 14996 10996
rect 14964 10965 14965 10995
rect 14965 10965 14995 10995
rect 14995 10965 14996 10995
rect 14964 10964 14996 10965
rect 14964 10915 14996 10916
rect 14964 10885 14965 10915
rect 14965 10885 14995 10915
rect 14995 10885 14996 10915
rect 14964 10884 14996 10885
rect 14964 10835 14996 10836
rect 14964 10805 14965 10835
rect 14965 10805 14995 10835
rect 14995 10805 14996 10835
rect 14964 10804 14996 10805
rect 14964 10755 14996 10756
rect 14964 10725 14965 10755
rect 14965 10725 14995 10755
rect 14995 10725 14996 10755
rect 14964 10724 14996 10725
rect 14964 10675 14996 10676
rect 14964 10645 14965 10675
rect 14965 10645 14995 10675
rect 14995 10645 14996 10675
rect 14964 10644 14996 10645
rect 14964 10595 14996 10596
rect 14964 10565 14965 10595
rect 14965 10565 14995 10595
rect 14995 10565 14996 10595
rect 14964 10564 14996 10565
rect 14964 10515 14996 10516
rect 14964 10485 14965 10515
rect 14965 10485 14995 10515
rect 14995 10485 14996 10515
rect 14964 10484 14996 10485
rect 14964 10435 14996 10436
rect 14964 10405 14965 10435
rect 14965 10405 14995 10435
rect 14995 10405 14996 10435
rect 14964 10404 14996 10405
rect 14964 10355 14996 10356
rect 14964 10325 14965 10355
rect 14965 10325 14995 10355
rect 14995 10325 14996 10355
rect 14964 10324 14996 10325
rect 14964 10275 14996 10276
rect 14964 10245 14965 10275
rect 14965 10245 14995 10275
rect 14995 10245 14996 10275
rect 14964 10244 14996 10245
rect 14964 10195 14996 10196
rect 14964 10165 14965 10195
rect 14965 10165 14995 10195
rect 14995 10165 14996 10195
rect 14964 10164 14996 10165
rect 14964 10115 14996 10116
rect 14964 10085 14965 10115
rect 14965 10085 14995 10115
rect 14995 10085 14996 10115
rect 14964 10084 14996 10085
rect 14964 10035 14996 10036
rect 14964 10005 14965 10035
rect 14965 10005 14995 10035
rect 14995 10005 14996 10035
rect 14964 10004 14996 10005
rect 14964 9955 14996 9956
rect 14964 9925 14965 9955
rect 14965 9925 14995 9955
rect 14995 9925 14996 9955
rect 14964 9924 14996 9925
rect 14964 9875 14996 9876
rect 14964 9845 14965 9875
rect 14965 9845 14995 9875
rect 14995 9845 14996 9875
rect 14964 9844 14996 9845
rect 14964 9795 14996 9796
rect 14964 9765 14965 9795
rect 14965 9765 14995 9795
rect 14995 9765 14996 9795
rect 14964 9764 14996 9765
rect 14964 9715 14996 9716
rect 14964 9685 14965 9715
rect 14965 9685 14995 9715
rect 14995 9685 14996 9715
rect 14964 9684 14996 9685
rect 14964 9635 14996 9636
rect 14964 9605 14965 9635
rect 14965 9605 14995 9635
rect 14995 9605 14996 9635
rect 14964 9604 14996 9605
rect 14964 9555 14996 9556
rect 14964 9525 14965 9555
rect 14965 9525 14995 9555
rect 14995 9525 14996 9555
rect 14964 9524 14996 9525
rect 14964 9475 14996 9476
rect 14964 9445 14965 9475
rect 14965 9445 14995 9475
rect 14995 9445 14996 9475
rect 14964 9444 14996 9445
rect 14964 9395 14996 9396
rect 14964 9365 14965 9395
rect 14965 9365 14995 9395
rect 14995 9365 14996 9395
rect 14964 9364 14996 9365
rect 14964 9315 14996 9316
rect 14964 9285 14965 9315
rect 14965 9285 14995 9315
rect 14995 9285 14996 9315
rect 14964 9284 14996 9285
rect 14964 9235 14996 9236
rect 14964 9205 14965 9235
rect 14965 9205 14995 9235
rect 14995 9205 14996 9235
rect 14964 9204 14996 9205
rect 14964 9155 14996 9156
rect 14964 9125 14965 9155
rect 14965 9125 14995 9155
rect 14995 9125 14996 9155
rect 14964 9124 14996 9125
rect 14964 9075 14996 9076
rect 14964 9045 14965 9075
rect 14965 9045 14995 9075
rect 14995 9045 14996 9075
rect 14964 9044 14996 9045
rect 14964 8995 14996 8996
rect 14964 8965 14965 8995
rect 14965 8965 14995 8995
rect 14995 8965 14996 8995
rect 14964 8964 14996 8965
rect 14964 8915 14996 8916
rect 14964 8885 14965 8915
rect 14965 8885 14995 8915
rect 14995 8885 14996 8915
rect 14964 8884 14996 8885
rect 14964 8835 14996 8836
rect 14964 8805 14965 8835
rect 14965 8805 14995 8835
rect 14995 8805 14996 8835
rect 14964 8804 14996 8805
rect 14964 8755 14996 8756
rect 14964 8725 14965 8755
rect 14965 8725 14995 8755
rect 14995 8725 14996 8755
rect 14964 8724 14996 8725
rect 14964 8675 14996 8676
rect 14964 8645 14965 8675
rect 14965 8645 14995 8675
rect 14995 8645 14996 8675
rect 14964 8644 14996 8645
rect 14964 8595 14996 8596
rect 14964 8565 14965 8595
rect 14965 8565 14995 8595
rect 14995 8565 14996 8595
rect 14964 8564 14996 8565
rect 14964 8515 14996 8516
rect 14964 8485 14965 8515
rect 14965 8485 14995 8515
rect 14995 8485 14996 8515
rect 14964 8484 14996 8485
rect 14964 8435 14996 8436
rect 14964 8405 14965 8435
rect 14965 8405 14995 8435
rect 14995 8405 14996 8435
rect 14964 8404 14996 8405
rect 14964 8355 14996 8356
rect 14964 8325 14965 8355
rect 14965 8325 14995 8355
rect 14995 8325 14996 8355
rect 14964 8324 14996 8325
rect 14964 8275 14996 8276
rect 14964 8245 14965 8275
rect 14965 8245 14995 8275
rect 14995 8245 14996 8275
rect 14964 8244 14996 8245
rect 14964 8195 14996 8196
rect 14964 8165 14965 8195
rect 14965 8165 14995 8195
rect 14995 8165 14996 8195
rect 14964 8164 14996 8165
rect 14964 8115 14996 8116
rect 14964 8085 14965 8115
rect 14965 8085 14995 8115
rect 14995 8085 14996 8115
rect 14964 8084 14996 8085
rect 14964 8035 14996 8036
rect 14964 8005 14965 8035
rect 14965 8005 14995 8035
rect 14995 8005 14996 8035
rect 14964 8004 14996 8005
rect 14964 7955 14996 7956
rect 14964 7925 14965 7955
rect 14965 7925 14995 7955
rect 14995 7925 14996 7955
rect 14964 7924 14996 7925
rect 14964 7875 14996 7876
rect 14964 7845 14965 7875
rect 14965 7845 14995 7875
rect 14995 7845 14996 7875
rect 14964 7844 14996 7845
rect 14964 7795 14996 7796
rect 14964 7765 14965 7795
rect 14965 7765 14995 7795
rect 14995 7765 14996 7795
rect 14964 7764 14996 7765
rect 14964 7715 14996 7716
rect 14964 7685 14965 7715
rect 14965 7685 14995 7715
rect 14995 7685 14996 7715
rect 14964 7684 14996 7685
rect 14964 7635 14996 7636
rect 14964 7605 14965 7635
rect 14965 7605 14995 7635
rect 14995 7605 14996 7635
rect 14964 7604 14996 7605
rect 14964 7555 14996 7556
rect 14964 7525 14965 7555
rect 14965 7525 14995 7555
rect 14995 7525 14996 7555
rect 14964 7524 14996 7525
rect 14964 7475 14996 7476
rect 14964 7445 14965 7475
rect 14965 7445 14995 7475
rect 14995 7445 14996 7475
rect 14964 7444 14996 7445
rect 14964 7395 14996 7396
rect 14964 7365 14965 7395
rect 14965 7365 14995 7395
rect 14995 7365 14996 7395
rect 14964 7364 14996 7365
rect 14964 7315 14996 7316
rect 14964 7285 14965 7315
rect 14965 7285 14995 7315
rect 14995 7285 14996 7315
rect 14964 7284 14996 7285
rect 14964 7235 14996 7236
rect 14964 7205 14965 7235
rect 14965 7205 14995 7235
rect 14995 7205 14996 7235
rect 14964 7204 14996 7205
rect 14964 7155 14996 7156
rect 14964 7125 14965 7155
rect 14965 7125 14995 7155
rect 14995 7125 14996 7155
rect 14964 7124 14996 7125
rect 14964 7075 14996 7076
rect 14964 7045 14965 7075
rect 14965 7045 14995 7075
rect 14995 7045 14996 7075
rect 14964 7044 14996 7045
rect 14964 6995 14996 6996
rect 14964 6965 14965 6995
rect 14965 6965 14995 6995
rect 14995 6965 14996 6995
rect 14964 6964 14996 6965
rect 14964 6915 14996 6916
rect 14964 6885 14965 6915
rect 14965 6885 14995 6915
rect 14995 6885 14996 6915
rect 14964 6884 14996 6885
rect 14964 6835 14996 6836
rect 14964 6805 14965 6835
rect 14965 6805 14995 6835
rect 14995 6805 14996 6835
rect 14964 6804 14996 6805
rect 14964 6755 14996 6756
rect 14964 6725 14965 6755
rect 14965 6725 14995 6755
rect 14995 6725 14996 6755
rect 14964 6724 14996 6725
rect 14964 6675 14996 6676
rect 14964 6645 14965 6675
rect 14965 6645 14995 6675
rect 14995 6645 14996 6675
rect 14964 6644 14996 6645
rect 14964 6595 14996 6596
rect 14964 6565 14965 6595
rect 14965 6565 14995 6595
rect 14995 6565 14996 6595
rect 14964 6564 14996 6565
rect 14964 6515 14996 6516
rect 14964 6485 14965 6515
rect 14965 6485 14995 6515
rect 14995 6485 14996 6515
rect 14964 6484 14996 6485
rect 14964 6435 14996 6436
rect 14964 6405 14965 6435
rect 14965 6405 14995 6435
rect 14995 6405 14996 6435
rect 14964 6404 14996 6405
rect 14964 6355 14996 6356
rect 14964 6325 14965 6355
rect 14965 6325 14995 6355
rect 14995 6325 14996 6355
rect 14964 6324 14996 6325
rect 14964 6275 14996 6276
rect 14964 6245 14965 6275
rect 14965 6245 14995 6275
rect 14995 6245 14996 6275
rect 14964 6244 14996 6245
rect 14964 6195 14996 6196
rect 14964 6165 14965 6195
rect 14965 6165 14995 6195
rect 14995 6165 14996 6195
rect 14964 6164 14996 6165
rect 14964 6115 14996 6116
rect 14964 6085 14965 6115
rect 14965 6085 14995 6115
rect 14995 6085 14996 6115
rect 14964 6084 14996 6085
rect 14964 6035 14996 6036
rect 14964 6005 14965 6035
rect 14965 6005 14995 6035
rect 14995 6005 14996 6035
rect 14964 6004 14996 6005
rect 14964 5955 14996 5956
rect 14964 5925 14965 5955
rect 14965 5925 14995 5955
rect 14995 5925 14996 5955
rect 14964 5924 14996 5925
rect 14964 5875 14996 5876
rect 14964 5845 14965 5875
rect 14965 5845 14995 5875
rect 14995 5845 14996 5875
rect 14964 5844 14996 5845
rect 14964 5795 14996 5796
rect 14964 5765 14965 5795
rect 14965 5765 14995 5795
rect 14995 5765 14996 5795
rect 14964 5764 14996 5765
rect 14964 5715 14996 5716
rect 14964 5685 14965 5715
rect 14965 5685 14995 5715
rect 14995 5685 14996 5715
rect 14964 5684 14996 5685
rect 14964 5635 14996 5636
rect 14964 5605 14965 5635
rect 14965 5605 14995 5635
rect 14995 5605 14996 5635
rect 14964 5604 14996 5605
rect 14964 5555 14996 5556
rect 14964 5525 14965 5555
rect 14965 5525 14995 5555
rect 14995 5525 14996 5555
rect 14964 5524 14996 5525
rect 14964 5475 14996 5476
rect 14964 5445 14965 5475
rect 14965 5445 14995 5475
rect 14995 5445 14996 5475
rect 14964 5444 14996 5445
rect 14964 5395 14996 5396
rect 14964 5365 14965 5395
rect 14965 5365 14995 5395
rect 14995 5365 14996 5395
rect 14964 5364 14996 5365
rect 14964 5315 14996 5316
rect 14964 5285 14965 5315
rect 14965 5285 14995 5315
rect 14995 5285 14996 5315
rect 14964 5284 14996 5285
rect 14964 5235 14996 5236
rect 14964 5205 14965 5235
rect 14965 5205 14995 5235
rect 14995 5205 14996 5235
rect 14964 5204 14996 5205
rect 14964 5155 14996 5156
rect 14964 5125 14965 5155
rect 14965 5125 14995 5155
rect 14995 5125 14996 5155
rect 14964 5124 14996 5125
rect 14964 5075 14996 5076
rect 14964 5045 14965 5075
rect 14965 5045 14995 5075
rect 14995 5045 14996 5075
rect 14964 5044 14996 5045
rect 14964 4995 14996 4996
rect 14964 4965 14965 4995
rect 14965 4965 14995 4995
rect 14995 4965 14996 4995
rect 14964 4964 14996 4965
rect 14964 4915 14996 4916
rect 14964 4885 14965 4915
rect 14965 4885 14995 4915
rect 14995 4885 14996 4915
rect 14964 4884 14996 4885
rect 14964 4835 14996 4836
rect 14964 4805 14965 4835
rect 14965 4805 14995 4835
rect 14995 4805 14996 4835
rect 14964 4804 14996 4805
rect 14964 4675 14996 4676
rect 14964 4645 14965 4675
rect 14965 4645 14995 4675
rect 14995 4645 14996 4675
rect 14964 4644 14996 4645
rect 14964 4595 14996 4596
rect 14964 4565 14965 4595
rect 14965 4565 14995 4595
rect 14995 4565 14996 4595
rect 14964 4564 14996 4565
rect 14964 4515 14996 4516
rect 14964 4485 14965 4515
rect 14965 4485 14995 4515
rect 14995 4485 14996 4515
rect 14964 4484 14996 4485
rect 14964 4435 14996 4436
rect 14964 4405 14965 4435
rect 14965 4405 14995 4435
rect 14995 4405 14996 4435
rect 14964 4404 14996 4405
rect 14964 4355 14996 4356
rect 14964 4325 14965 4355
rect 14965 4325 14995 4355
rect 14995 4325 14996 4355
rect 14964 4324 14996 4325
rect 14964 4275 14996 4276
rect 14964 4245 14965 4275
rect 14965 4245 14995 4275
rect 14995 4245 14996 4275
rect 14964 4244 14996 4245
rect 14964 4195 14996 4196
rect 14964 4165 14965 4195
rect 14965 4165 14995 4195
rect 14995 4165 14996 4195
rect 14964 4164 14996 4165
rect 14964 4115 14996 4116
rect 14964 4085 14965 4115
rect 14965 4085 14995 4115
rect 14995 4085 14996 4115
rect 14964 4084 14996 4085
rect 14964 4035 14996 4036
rect 14964 4005 14965 4035
rect 14965 4005 14995 4035
rect 14995 4005 14996 4035
rect 14964 4004 14996 4005
rect 14964 3955 14996 3956
rect 14964 3925 14965 3955
rect 14965 3925 14995 3955
rect 14995 3925 14996 3955
rect 14964 3924 14996 3925
rect 14964 3875 14996 3876
rect 14964 3845 14965 3875
rect 14965 3845 14995 3875
rect 14995 3845 14996 3875
rect 14964 3844 14996 3845
rect 14964 3795 14996 3796
rect 14964 3765 14965 3795
rect 14965 3765 14995 3795
rect 14995 3765 14996 3795
rect 14964 3764 14996 3765
rect 14964 3715 14996 3716
rect 14964 3685 14965 3715
rect 14965 3685 14995 3715
rect 14995 3685 14996 3715
rect 14964 3684 14996 3685
rect 14964 3635 14996 3636
rect 14964 3605 14965 3635
rect 14965 3605 14995 3635
rect 14995 3605 14996 3635
rect 14964 3604 14996 3605
rect 14964 3555 14996 3556
rect 14964 3525 14965 3555
rect 14965 3525 14995 3555
rect 14995 3525 14996 3555
rect 14964 3524 14996 3525
rect 14964 3475 14996 3476
rect 14964 3445 14965 3475
rect 14965 3445 14995 3475
rect 14995 3445 14996 3475
rect 14964 3444 14996 3445
rect 14964 3395 14996 3396
rect 14964 3365 14965 3395
rect 14965 3365 14995 3395
rect 14995 3365 14996 3395
rect 14964 3364 14996 3365
rect 14964 3315 14996 3316
rect 14964 3285 14965 3315
rect 14965 3285 14995 3315
rect 14995 3285 14996 3315
rect 14964 3284 14996 3285
rect 14964 3235 14996 3236
rect 14964 3205 14965 3235
rect 14965 3205 14995 3235
rect 14995 3205 14996 3235
rect 14964 3204 14996 3205
rect 14964 3155 14996 3156
rect 14964 3125 14965 3155
rect 14965 3125 14995 3155
rect 14995 3125 14996 3155
rect 14964 3124 14996 3125
rect 14964 3075 14996 3076
rect 14964 3045 14965 3075
rect 14965 3045 14995 3075
rect 14995 3045 14996 3075
rect 14964 3044 14996 3045
rect 14964 2995 14996 2996
rect 14964 2965 14965 2995
rect 14965 2965 14995 2995
rect 14995 2965 14996 2995
rect 14964 2964 14996 2965
rect 14964 2915 14996 2916
rect 14964 2885 14965 2915
rect 14965 2885 14995 2915
rect 14995 2885 14996 2915
rect 14964 2884 14996 2885
rect 14964 2835 14996 2836
rect 14964 2805 14965 2835
rect 14965 2805 14995 2835
rect 14995 2805 14996 2835
rect 14964 2804 14996 2805
rect 14964 2755 14996 2756
rect 14964 2725 14965 2755
rect 14965 2725 14995 2755
rect 14995 2725 14996 2755
rect 14964 2724 14996 2725
rect 14964 2675 14996 2676
rect 14964 2645 14965 2675
rect 14965 2645 14995 2675
rect 14995 2645 14996 2675
rect 14964 2644 14996 2645
rect 14964 2595 14996 2596
rect 14964 2565 14965 2595
rect 14965 2565 14995 2595
rect 14995 2565 14996 2595
rect 14964 2564 14996 2565
rect 14964 2515 14996 2516
rect 14964 2485 14965 2515
rect 14965 2485 14995 2515
rect 14995 2485 14996 2515
rect 14964 2484 14996 2485
rect 14964 2435 14996 2436
rect 14964 2405 14965 2435
rect 14965 2405 14995 2435
rect 14995 2405 14996 2435
rect 14964 2404 14996 2405
rect 14964 2355 14996 2356
rect 14964 2325 14965 2355
rect 14965 2325 14995 2355
rect 14995 2325 14996 2355
rect 14964 2324 14996 2325
rect 14964 2275 14996 2276
rect 14964 2245 14965 2275
rect 14965 2245 14995 2275
rect 14995 2245 14996 2275
rect 14964 2244 14996 2245
rect 14964 2195 14996 2196
rect 14964 2165 14965 2195
rect 14965 2165 14995 2195
rect 14995 2165 14996 2195
rect 14964 2164 14996 2165
rect 14964 2115 14996 2116
rect 14964 2085 14965 2115
rect 14965 2085 14995 2115
rect 14995 2085 14996 2115
rect 14964 2084 14996 2085
rect 14964 2035 14996 2036
rect 14964 2005 14965 2035
rect 14965 2005 14995 2035
rect 14995 2005 14996 2035
rect 14964 2004 14996 2005
rect 14964 1955 14996 1956
rect 14964 1925 14965 1955
rect 14965 1925 14995 1955
rect 14995 1925 14996 1955
rect 14964 1924 14996 1925
rect 14964 1795 14996 1796
rect 14964 1765 14965 1795
rect 14965 1765 14995 1795
rect 14995 1765 14996 1795
rect 14964 1764 14996 1765
rect 14964 1715 14996 1716
rect 14964 1685 14965 1715
rect 14965 1685 14995 1715
rect 14995 1685 14996 1715
rect 14964 1684 14996 1685
rect 14964 1635 14996 1636
rect 14964 1605 14965 1635
rect 14965 1605 14995 1635
rect 14995 1605 14996 1635
rect 14964 1604 14996 1605
rect 14964 1555 14996 1556
rect 14964 1525 14965 1555
rect 14965 1525 14995 1555
rect 14995 1525 14996 1555
rect 14964 1524 14996 1525
rect 14964 1475 14996 1476
rect 14964 1445 14965 1475
rect 14965 1445 14995 1475
rect 14995 1445 14996 1475
rect 14964 1444 14996 1445
rect 14964 1395 14996 1396
rect 14964 1365 14965 1395
rect 14965 1365 14995 1395
rect 14995 1365 14996 1395
rect 14964 1364 14996 1365
rect 14964 1315 14996 1316
rect 14964 1285 14965 1315
rect 14965 1285 14995 1315
rect 14995 1285 14996 1315
rect 14964 1284 14996 1285
rect 14964 1235 14996 1236
rect 14964 1205 14965 1235
rect 14965 1205 14995 1235
rect 14995 1205 14996 1235
rect 14964 1204 14996 1205
rect 14964 1155 14996 1156
rect 14964 1125 14965 1155
rect 14965 1125 14995 1155
rect 14995 1125 14996 1155
rect 14964 1124 14996 1125
rect 14964 1075 14996 1076
rect 14964 1045 14965 1075
rect 14965 1045 14995 1075
rect 14995 1045 14996 1075
rect 14964 1044 14996 1045
rect 14964 995 14996 996
rect 14964 965 14965 995
rect 14965 965 14995 995
rect 14995 965 14996 995
rect 14964 964 14996 965
rect 14964 915 14996 916
rect 14964 885 14965 915
rect 14965 885 14995 915
rect 14995 885 14996 915
rect 14964 884 14996 885
rect 14964 835 14996 836
rect 14964 805 14965 835
rect 14965 805 14995 835
rect 14995 805 14996 835
rect 14964 804 14996 805
rect 14964 755 14996 756
rect 14964 725 14965 755
rect 14965 725 14995 755
rect 14995 725 14996 755
rect 14964 724 14996 725
rect 14964 675 14996 676
rect 14964 645 14965 675
rect 14965 645 14995 675
rect 14995 645 14996 675
rect 14964 644 14996 645
rect 14964 595 14996 596
rect 14964 565 14965 595
rect 14965 565 14995 595
rect 14995 565 14996 595
rect 14964 564 14996 565
rect 14964 515 14996 516
rect 14964 485 14965 515
rect 14965 485 14995 515
rect 14995 485 14996 515
rect 14964 484 14996 485
rect 14804 244 14836 436
rect 14964 244 14996 436
rect 14404 4 14436 196
<< metal4 >>
rect 0 15956 520 15960
rect 0 15924 4 15956
rect 36 15924 164 15956
rect 196 15924 324 15956
rect 356 15924 484 15956
rect 516 15924 520 15956
rect 0 15920 520 15924
rect 14480 15956 15000 15960
rect 14480 15924 14484 15956
rect 14516 15924 14644 15956
rect 14676 15924 14804 15956
rect 14836 15924 14964 15956
rect 14996 15924 15000 15956
rect 14480 15920 15000 15924
rect 0 15876 680 15880
rect 0 15844 4 15876
rect 36 15844 164 15876
rect 196 15844 324 15876
rect 356 15844 484 15876
rect 516 15844 680 15876
rect 0 15840 680 15844
rect 14320 15876 15000 15880
rect 14320 15844 14484 15876
rect 14516 15844 14644 15876
rect 14676 15844 14804 15876
rect 14836 15844 14964 15876
rect 14996 15844 15000 15876
rect 14320 15840 15000 15844
rect 0 15796 680 15800
rect 0 15764 4 15796
rect 36 15764 164 15796
rect 196 15764 324 15796
rect 356 15764 484 15796
rect 516 15764 680 15796
rect 0 15760 680 15764
rect 14320 15796 15000 15800
rect 14320 15764 14484 15796
rect 14516 15764 14644 15796
rect 14676 15764 14804 15796
rect 14836 15764 14964 15796
rect 14996 15764 15000 15796
rect 14320 15760 15000 15764
rect 0 15716 680 15720
rect 0 15684 4 15716
rect 36 15684 164 15716
rect 196 15684 324 15716
rect 356 15684 484 15716
rect 516 15684 680 15716
rect 0 15680 680 15684
rect 14320 15716 15000 15720
rect 14320 15684 14484 15716
rect 14516 15684 14644 15716
rect 14676 15684 14804 15716
rect 14836 15684 14964 15716
rect 14996 15684 15000 15716
rect 14320 15680 15000 15684
rect 0 15636 680 15640
rect 0 15604 4 15636
rect 36 15604 164 15636
rect 196 15604 324 15636
rect 356 15604 484 15636
rect 516 15604 680 15636
rect 0 15600 680 15604
rect 14320 15636 15000 15640
rect 14320 15604 14484 15636
rect 14516 15604 14644 15636
rect 14676 15604 14804 15636
rect 14836 15604 14964 15636
rect 14996 15604 15000 15636
rect 14320 15600 15000 15604
rect 0 15556 680 15560
rect 0 15524 4 15556
rect 36 15524 164 15556
rect 196 15524 324 15556
rect 356 15524 484 15556
rect 516 15524 680 15556
rect 0 15520 680 15524
rect 14320 15556 15000 15560
rect 14320 15524 14484 15556
rect 14516 15524 14644 15556
rect 14676 15524 14804 15556
rect 14836 15524 14964 15556
rect 14996 15524 15000 15556
rect 14320 15520 15000 15524
rect 0 15476 520 15480
rect 0 15444 4 15476
rect 36 15444 164 15476
rect 196 15444 324 15476
rect 356 15444 484 15476
rect 516 15444 520 15476
rect 0 15440 520 15444
rect 14480 15476 15000 15480
rect 14480 15444 14484 15476
rect 14516 15444 14644 15476
rect 14676 15444 14804 15476
rect 14836 15444 14964 15476
rect 14996 15444 15000 15476
rect 14480 15440 15000 15444
rect 0 15396 520 15400
rect 0 15364 4 15396
rect 36 15364 164 15396
rect 196 15364 324 15396
rect 356 15364 484 15396
rect 516 15364 520 15396
rect 0 15360 520 15364
rect 14480 15396 15000 15400
rect 14480 15364 14484 15396
rect 14516 15364 14644 15396
rect 14676 15364 14804 15396
rect 14836 15364 14964 15396
rect 14996 15364 15000 15396
rect 14480 15360 15000 15364
rect 0 15316 520 15320
rect 0 15284 4 15316
rect 36 15284 164 15316
rect 196 15284 324 15316
rect 356 15284 484 15316
rect 516 15284 520 15316
rect 0 15280 520 15284
rect 14480 15316 15000 15320
rect 14480 15284 14484 15316
rect 14516 15284 14644 15316
rect 14676 15284 14804 15316
rect 14836 15284 14964 15316
rect 14996 15284 15000 15316
rect 14480 15280 15000 15284
rect 0 15236 680 15240
rect 0 15204 4 15236
rect 36 15204 164 15236
rect 196 15204 324 15236
rect 356 15204 484 15236
rect 516 15204 680 15236
rect 0 15200 680 15204
rect 14320 15236 15000 15240
rect 14320 15204 14484 15236
rect 14516 15204 14644 15236
rect 14676 15204 14804 15236
rect 14836 15204 14964 15236
rect 14996 15204 15000 15236
rect 14320 15200 15000 15204
rect 0 15156 680 15160
rect 0 15124 4 15156
rect 36 15124 164 15156
rect 196 15124 324 15156
rect 356 15124 484 15156
rect 516 15124 680 15156
rect 0 15120 680 15124
rect 14320 15156 15000 15160
rect 14320 15124 14484 15156
rect 14516 15124 14644 15156
rect 14676 15124 14804 15156
rect 14836 15124 14964 15156
rect 14996 15124 15000 15156
rect 14320 15120 15000 15124
rect 0 15076 680 15080
rect 0 15044 4 15076
rect 36 15044 164 15076
rect 196 15044 324 15076
rect 356 15044 484 15076
rect 516 15044 680 15076
rect 0 15040 680 15044
rect 14320 15076 15000 15080
rect 14320 15044 14484 15076
rect 14516 15044 14644 15076
rect 14676 15044 14804 15076
rect 14836 15044 14964 15076
rect 14996 15044 15000 15076
rect 14320 15040 15000 15044
rect 0 14996 680 15000
rect 0 14964 4 14996
rect 36 14964 164 14996
rect 196 14964 324 14996
rect 356 14964 484 14996
rect 516 14964 680 14996
rect 0 14960 680 14964
rect 14320 14996 15000 15000
rect 14320 14964 14484 14996
rect 14516 14964 14644 14996
rect 14676 14964 14804 14996
rect 14836 14964 14964 14996
rect 14996 14964 15000 14996
rect 14320 14960 15000 14964
rect 0 14916 680 14920
rect 0 14884 4 14916
rect 36 14884 164 14916
rect 196 14884 324 14916
rect 356 14884 484 14916
rect 516 14884 680 14916
rect 0 14880 680 14884
rect 14320 14916 15000 14920
rect 14320 14884 14484 14916
rect 14516 14884 14644 14916
rect 14676 14884 14804 14916
rect 14836 14884 14964 14916
rect 14996 14884 15000 14916
rect 14320 14880 15000 14884
rect 0 14836 520 14840
rect 0 14804 4 14836
rect 36 14804 164 14836
rect 196 14804 324 14836
rect 356 14804 484 14836
rect 516 14804 520 14836
rect 0 14800 520 14804
rect 14480 14836 15000 14840
rect 14480 14804 14484 14836
rect 14516 14804 14644 14836
rect 14676 14804 14804 14836
rect 14836 14804 14964 14836
rect 14996 14804 15000 14836
rect 14480 14800 15000 14804
rect 0 14756 520 14760
rect 0 14724 4 14756
rect 36 14724 164 14756
rect 196 14724 324 14756
rect 356 14724 484 14756
rect 516 14724 520 14756
rect 0 14720 520 14724
rect 14480 14756 15000 14760
rect 14480 14724 14484 14756
rect 14516 14724 14644 14756
rect 14676 14724 14804 14756
rect 14836 14724 14964 14756
rect 14996 14724 15000 14756
rect 14480 14720 15000 14724
rect 0 14676 680 14680
rect 0 14644 4 14676
rect 36 14644 164 14676
rect 196 14644 324 14676
rect 356 14644 484 14676
rect 516 14644 680 14676
rect 0 14640 680 14644
rect 14360 14676 15000 14680
rect 14360 14644 14484 14676
rect 14516 14644 14644 14676
rect 14676 14644 14804 14676
rect 14836 14644 14964 14676
rect 14996 14644 15000 14676
rect 14360 14640 15000 14644
rect 0 14596 520 14600
rect 0 14564 4 14596
rect 36 14564 164 14596
rect 196 14564 324 14596
rect 356 14564 484 14596
rect 516 14564 520 14596
rect 0 14560 520 14564
rect 14320 14596 14920 14600
rect 14320 14564 14884 14596
rect 14916 14564 14920 14596
rect 14320 14560 14920 14564
rect 0 14516 680 14520
rect 0 14484 4 14516
rect 36 14484 164 14516
rect 196 14484 324 14516
rect 356 14484 484 14516
rect 516 14484 680 14516
rect 0 14480 680 14484
rect 14320 14516 15000 14520
rect 14320 14484 14484 14516
rect 14516 14484 14644 14516
rect 14676 14484 14804 14516
rect 14836 14484 14964 14516
rect 14996 14484 15000 14516
rect 14320 14480 15000 14484
rect 0 14436 520 14440
rect 0 14404 4 14436
rect 36 14404 164 14436
rect 196 14404 324 14436
rect 356 14404 484 14436
rect 516 14404 520 14436
rect 0 14400 520 14404
rect 14320 14436 14760 14440
rect 14320 14404 14724 14436
rect 14756 14404 14760 14436
rect 14320 14400 14760 14404
rect 14800 14436 15000 14440
rect 14800 14404 14804 14436
rect 14836 14404 14964 14436
rect 14996 14404 15000 14436
rect 14800 14400 15000 14404
rect 0 14356 680 14360
rect 0 14324 4 14356
rect 36 14324 164 14356
rect 196 14324 324 14356
rect 356 14324 484 14356
rect 516 14324 680 14356
rect 0 14320 680 14324
rect 14320 14356 15000 14360
rect 14320 14324 14484 14356
rect 14516 14324 14644 14356
rect 14676 14324 14804 14356
rect 14836 14324 14964 14356
rect 14996 14324 15000 14356
rect 14320 14320 15000 14324
rect 0 14276 520 14280
rect 0 14244 4 14276
rect 36 14244 164 14276
rect 196 14244 324 14276
rect 356 14244 484 14276
rect 516 14244 520 14276
rect 0 14240 520 14244
rect 14480 14276 15000 14280
rect 14480 14244 14484 14276
rect 14516 14244 14644 14276
rect 14676 14244 14804 14276
rect 14836 14244 14964 14276
rect 14996 14244 15000 14276
rect 14480 14240 15000 14244
rect 0 14196 520 14200
rect 0 14164 4 14196
rect 36 14164 164 14196
rect 196 14164 324 14196
rect 356 14164 484 14196
rect 516 14164 520 14196
rect 0 14160 520 14164
rect 14480 14196 15000 14200
rect 14480 14164 14484 14196
rect 14516 14164 14644 14196
rect 14676 14164 14804 14196
rect 14836 14164 14964 14196
rect 14996 14164 15000 14196
rect 14480 14160 15000 14164
rect 0 14116 520 14120
rect 0 14084 4 14116
rect 36 14084 164 14116
rect 196 14084 324 14116
rect 356 14084 484 14116
rect 516 14084 520 14116
rect 0 14080 520 14084
rect 14480 14116 15000 14120
rect 14480 14084 14484 14116
rect 14516 14084 14644 14116
rect 14676 14084 14804 14116
rect 14836 14084 14964 14116
rect 14996 14084 15000 14116
rect 14480 14080 15000 14084
rect 0 14036 520 14040
rect 0 14004 4 14036
rect 36 14004 164 14036
rect 196 14004 324 14036
rect 356 14004 484 14036
rect 516 14004 520 14036
rect 0 14000 520 14004
rect 14480 14036 15000 14040
rect 14480 14004 14484 14036
rect 14516 14004 14644 14036
rect 14676 14004 14804 14036
rect 14836 14004 14964 14036
rect 14996 14004 15000 14036
rect 14480 14000 15000 14004
rect 0 13956 520 13960
rect 0 13924 4 13956
rect 36 13924 164 13956
rect 196 13924 324 13956
rect 356 13924 484 13956
rect 516 13924 520 13956
rect 0 13920 520 13924
rect 14480 13956 15000 13960
rect 14480 13924 14484 13956
rect 14516 13924 14644 13956
rect 14676 13924 14804 13956
rect 14836 13924 14964 13956
rect 14996 13924 15000 13956
rect 14480 13920 15000 13924
rect 0 13876 520 13880
rect 0 13844 4 13876
rect 36 13844 164 13876
rect 196 13844 324 13876
rect 356 13844 484 13876
rect 516 13844 520 13876
rect 0 13840 520 13844
rect 14480 13876 15000 13880
rect 14480 13844 14484 13876
rect 14516 13844 14644 13876
rect 14676 13844 14804 13876
rect 14836 13844 14964 13876
rect 14996 13844 15000 13876
rect 14480 13840 15000 13844
rect 0 13796 520 13800
rect 0 13764 4 13796
rect 36 13764 164 13796
rect 196 13764 324 13796
rect 356 13764 484 13796
rect 516 13764 520 13796
rect 0 13760 520 13764
rect 14480 13796 15000 13800
rect 14480 13764 14484 13796
rect 14516 13764 14644 13796
rect 14676 13764 14804 13796
rect 14836 13764 14964 13796
rect 14996 13764 15000 13796
rect 14480 13760 15000 13764
rect 0 13716 520 13720
rect 0 13684 4 13716
rect 36 13684 164 13716
rect 196 13684 324 13716
rect 356 13684 484 13716
rect 516 13684 520 13716
rect 0 13680 520 13684
rect 14480 13716 15000 13720
rect 14480 13684 14484 13716
rect 14516 13684 14644 13716
rect 14676 13684 14804 13716
rect 14836 13684 14964 13716
rect 14996 13684 15000 13716
rect 14480 13680 15000 13684
rect 0 13636 520 13640
rect 0 13604 4 13636
rect 36 13604 164 13636
rect 196 13604 324 13636
rect 356 13604 484 13636
rect 516 13604 520 13636
rect 0 13600 520 13604
rect 14480 13636 15000 13640
rect 14480 13604 14484 13636
rect 14516 13604 14644 13636
rect 14676 13604 14804 13636
rect 14836 13604 14964 13636
rect 14996 13604 15000 13636
rect 14480 13600 15000 13604
rect 0 13556 520 13560
rect 0 13524 4 13556
rect 36 13524 164 13556
rect 196 13524 324 13556
rect 356 13524 484 13556
rect 516 13524 520 13556
rect 0 13520 520 13524
rect 14480 13556 15000 13560
rect 14480 13524 14484 13556
rect 14516 13524 14644 13556
rect 14676 13524 14804 13556
rect 14836 13524 14964 13556
rect 14996 13524 15000 13556
rect 14480 13520 15000 13524
rect 0 13476 520 13480
rect 0 13444 4 13476
rect 36 13444 164 13476
rect 196 13444 324 13476
rect 356 13444 484 13476
rect 516 13444 520 13476
rect 0 13440 520 13444
rect 14480 13476 15000 13480
rect 14480 13444 14484 13476
rect 14516 13444 14644 13476
rect 14676 13444 14804 13476
rect 14836 13444 14964 13476
rect 14996 13444 15000 13476
rect 14480 13440 15000 13444
rect 0 13396 520 13400
rect 0 13364 4 13396
rect 36 13364 164 13396
rect 196 13364 324 13396
rect 356 13364 484 13396
rect 516 13364 520 13396
rect 0 13360 520 13364
rect 14480 13396 15000 13400
rect 14480 13364 14484 13396
rect 14516 13364 14644 13396
rect 14676 13364 14804 13396
rect 14836 13364 14964 13396
rect 14996 13364 15000 13396
rect 14480 13360 15000 13364
rect 0 13316 520 13320
rect 0 13284 4 13316
rect 36 13284 164 13316
rect 196 13284 324 13316
rect 356 13284 484 13316
rect 516 13284 520 13316
rect 0 13280 520 13284
rect 14480 13316 15000 13320
rect 14480 13284 14484 13316
rect 14516 13284 14644 13316
rect 14676 13284 14804 13316
rect 14836 13284 14964 13316
rect 14996 13284 15000 13316
rect 14480 13280 15000 13284
rect 0 13236 520 13240
rect 0 13204 4 13236
rect 36 13204 164 13236
rect 196 13204 324 13236
rect 356 13204 484 13236
rect 516 13204 520 13236
rect 0 13200 520 13204
rect 14480 13236 15000 13240
rect 14480 13204 14484 13236
rect 14516 13204 14644 13236
rect 14676 13204 14804 13236
rect 14836 13204 14964 13236
rect 14996 13204 15000 13236
rect 14480 13200 15000 13204
rect 0 13156 520 13160
rect 0 13124 4 13156
rect 36 13124 164 13156
rect 196 13124 324 13156
rect 356 13124 484 13156
rect 516 13124 520 13156
rect 0 13120 520 13124
rect 14360 13156 14600 13160
rect 14360 13124 14564 13156
rect 14596 13124 14600 13156
rect 14360 13120 14600 13124
rect 14640 13156 15000 13160
rect 14640 13124 14644 13156
rect 14676 13124 14804 13156
rect 14836 13124 14964 13156
rect 14996 13124 15000 13156
rect 14640 13120 15000 13124
rect 0 13076 520 13080
rect 0 13044 4 13076
rect 36 13044 164 13076
rect 196 13044 324 13076
rect 356 13044 484 13076
rect 516 13044 520 13076
rect 0 13040 520 13044
rect 14480 13076 15000 13080
rect 14480 13044 14484 13076
rect 14516 13044 14644 13076
rect 14676 13044 14804 13076
rect 14836 13044 14964 13076
rect 14996 13044 15000 13076
rect 14480 13040 15000 13044
rect 0 12996 520 13000
rect 0 12964 4 12996
rect 36 12964 164 12996
rect 196 12964 324 12996
rect 356 12964 484 12996
rect 516 12964 520 12996
rect 0 12960 520 12964
rect 14480 12996 15000 13000
rect 14480 12964 14484 12996
rect 14516 12964 14644 12996
rect 14676 12964 14804 12996
rect 14836 12964 14964 12996
rect 14996 12964 15000 12996
rect 14480 12960 15000 12964
rect 0 12916 520 12920
rect 0 12884 4 12916
rect 36 12884 164 12916
rect 196 12884 324 12916
rect 356 12884 484 12916
rect 516 12884 520 12916
rect 0 12880 520 12884
rect 14480 12916 15000 12920
rect 14480 12884 14484 12916
rect 14516 12884 14644 12916
rect 14676 12884 14804 12916
rect 14836 12884 14964 12916
rect 14996 12884 15000 12916
rect 14480 12880 15000 12884
rect 0 12836 520 12840
rect 0 12804 4 12836
rect 36 12804 164 12836
rect 196 12804 324 12836
rect 356 12804 484 12836
rect 516 12804 520 12836
rect 0 12800 520 12804
rect 14480 12836 15000 12840
rect 14480 12804 14484 12836
rect 14516 12804 14644 12836
rect 14676 12804 14804 12836
rect 14836 12804 14964 12836
rect 14996 12804 15000 12836
rect 14480 12800 15000 12804
rect 0 12756 520 12760
rect 0 12724 4 12756
rect 36 12724 164 12756
rect 196 12724 324 12756
rect 356 12724 484 12756
rect 516 12724 520 12756
rect 0 12720 520 12724
rect 14480 12756 15000 12760
rect 14480 12724 14484 12756
rect 14516 12724 14644 12756
rect 14676 12724 14804 12756
rect 14836 12724 14964 12756
rect 14996 12724 15000 12756
rect 14480 12720 15000 12724
rect 0 12676 520 12680
rect 0 12644 4 12676
rect 36 12644 164 12676
rect 196 12644 324 12676
rect 356 12644 484 12676
rect 516 12644 520 12676
rect 0 12640 520 12644
rect 14480 12676 15000 12680
rect 14480 12644 14484 12676
rect 14516 12644 14644 12676
rect 14676 12644 14804 12676
rect 14836 12644 14964 12676
rect 14996 12644 15000 12676
rect 14480 12640 15000 12644
rect 0 12596 520 12600
rect 0 12564 4 12596
rect 36 12564 164 12596
rect 196 12564 324 12596
rect 356 12564 484 12596
rect 516 12564 520 12596
rect 0 12560 520 12564
rect 14480 12596 15000 12600
rect 14480 12564 14484 12596
rect 14516 12564 14644 12596
rect 14676 12564 14804 12596
rect 14836 12564 14964 12596
rect 14996 12564 15000 12596
rect 14480 12560 15000 12564
rect 0 12516 520 12520
rect 0 12484 4 12516
rect 36 12484 164 12516
rect 196 12484 324 12516
rect 356 12484 484 12516
rect 516 12484 520 12516
rect 0 12480 520 12484
rect 14480 12516 15000 12520
rect 14480 12484 14484 12516
rect 14516 12484 14644 12516
rect 14676 12484 14804 12516
rect 14836 12484 14964 12516
rect 14996 12484 15000 12516
rect 14480 12480 15000 12484
rect 0 12436 520 12440
rect 0 12404 4 12436
rect 36 12404 164 12436
rect 196 12404 324 12436
rect 356 12404 484 12436
rect 516 12404 520 12436
rect 0 12400 520 12404
rect 14480 12436 15000 12440
rect 14480 12404 14484 12436
rect 14516 12404 14644 12436
rect 14676 12404 14804 12436
rect 14836 12404 14964 12436
rect 14996 12404 15000 12436
rect 14480 12400 15000 12404
rect 0 12356 520 12360
rect 0 12324 4 12356
rect 36 12324 164 12356
rect 196 12324 324 12356
rect 356 12324 484 12356
rect 516 12324 520 12356
rect 0 12320 520 12324
rect 14480 12356 15000 12360
rect 14480 12324 14484 12356
rect 14516 12324 14644 12356
rect 14676 12324 14804 12356
rect 14836 12324 14964 12356
rect 14996 12324 15000 12356
rect 14480 12320 15000 12324
rect 0 12276 520 12280
rect 0 12244 4 12276
rect 36 12244 164 12276
rect 196 12244 324 12276
rect 356 12244 484 12276
rect 516 12244 520 12276
rect 0 12240 520 12244
rect 14480 12276 15000 12280
rect 14480 12244 14484 12276
rect 14516 12244 14644 12276
rect 14676 12244 14804 12276
rect 14836 12244 14964 12276
rect 14996 12244 15000 12276
rect 14480 12240 15000 12244
rect 0 12196 520 12200
rect 0 12164 4 12196
rect 36 12164 164 12196
rect 196 12164 324 12196
rect 356 12164 484 12196
rect 516 12164 520 12196
rect 0 12160 520 12164
rect 14480 12196 15000 12200
rect 14480 12164 14484 12196
rect 14516 12164 14644 12196
rect 14676 12164 14804 12196
rect 14836 12164 14964 12196
rect 14996 12164 15000 12196
rect 14480 12160 15000 12164
rect 0 12116 520 12120
rect 0 12084 4 12116
rect 36 12084 164 12116
rect 196 12084 324 12116
rect 356 12084 484 12116
rect 516 12084 520 12116
rect 0 12080 520 12084
rect 14480 12116 15000 12120
rect 14480 12084 14484 12116
rect 14516 12084 14644 12116
rect 14676 12084 14804 12116
rect 14836 12084 14964 12116
rect 14996 12084 15000 12116
rect 14480 12080 15000 12084
rect 0 12036 520 12040
rect 0 12004 4 12036
rect 36 12004 164 12036
rect 196 12004 324 12036
rect 356 12004 484 12036
rect 516 12004 520 12036
rect 0 12000 520 12004
rect 14480 12036 15000 12040
rect 14480 12004 14484 12036
rect 14516 12004 14644 12036
rect 14676 12004 14804 12036
rect 14836 12004 14964 12036
rect 14996 12004 15000 12036
rect 14480 12000 15000 12004
rect 0 11956 680 11960
rect 0 11924 4 11956
rect 36 11924 164 11956
rect 196 11924 324 11956
rect 356 11924 484 11956
rect 516 11924 680 11956
rect 0 11920 680 11924
rect 14360 11956 15000 11960
rect 14360 11924 14484 11956
rect 14516 11924 14644 11956
rect 14676 11924 14804 11956
rect 14836 11924 14964 11956
rect 14996 11924 15000 11956
rect 14360 11920 15000 11924
rect 0 11876 520 11880
rect 0 11844 4 11876
rect 36 11844 164 11876
rect 196 11844 324 11876
rect 356 11844 484 11876
rect 516 11844 520 11876
rect 0 11840 520 11844
rect 14320 11876 14760 11880
rect 14320 11844 14724 11876
rect 14756 11844 14760 11876
rect 14320 11840 14760 11844
rect 14800 11876 15000 11880
rect 14800 11844 14804 11876
rect 14836 11844 14964 11876
rect 14996 11844 15000 11876
rect 14800 11840 15000 11844
rect 0 11796 680 11800
rect 0 11764 4 11796
rect 36 11764 164 11796
rect 196 11764 324 11796
rect 356 11764 484 11796
rect 516 11764 680 11796
rect 0 11760 680 11764
rect 14360 11796 15000 11800
rect 14360 11764 14484 11796
rect 14516 11764 14644 11796
rect 14676 11764 14804 11796
rect 14836 11764 14964 11796
rect 14996 11764 15000 11796
rect 14360 11760 15000 11764
rect 0 11716 520 11720
rect 0 11684 4 11716
rect 36 11684 164 11716
rect 196 11684 324 11716
rect 356 11684 484 11716
rect 516 11684 520 11716
rect 0 11680 520 11684
rect 14320 11716 14920 11720
rect 14320 11684 14884 11716
rect 14916 11684 14920 11716
rect 14320 11680 14920 11684
rect 0 11636 680 11640
rect 0 11604 4 11636
rect 36 11604 164 11636
rect 196 11604 324 11636
rect 356 11604 484 11636
rect 516 11604 680 11636
rect 0 11600 680 11604
rect 14360 11636 15000 11640
rect 14360 11604 14484 11636
rect 14516 11604 14644 11636
rect 14676 11604 14804 11636
rect 14836 11604 14964 11636
rect 14996 11604 15000 11636
rect 14360 11600 15000 11604
rect 0 11556 520 11560
rect 0 11524 4 11556
rect 36 11524 164 11556
rect 196 11524 324 11556
rect 356 11524 484 11556
rect 516 11524 520 11556
rect 0 11520 520 11524
rect 14480 11556 15000 11560
rect 14480 11524 14484 11556
rect 14516 11524 14644 11556
rect 14676 11524 14804 11556
rect 14836 11524 14964 11556
rect 14996 11524 15000 11556
rect 14480 11520 15000 11524
rect 0 11476 520 11480
rect 0 11444 4 11476
rect 36 11444 164 11476
rect 196 11444 324 11476
rect 356 11444 484 11476
rect 516 11444 520 11476
rect 0 11440 520 11444
rect 14480 11476 15000 11480
rect 14480 11444 14484 11476
rect 14516 11444 14644 11476
rect 14676 11444 14804 11476
rect 14836 11444 14964 11476
rect 14996 11444 15000 11476
rect 14480 11440 15000 11444
rect 0 11396 680 11400
rect 0 11364 4 11396
rect 36 11364 164 11396
rect 196 11364 324 11396
rect 356 11364 484 11396
rect 516 11364 680 11396
rect 0 11360 680 11364
rect 14320 11396 15000 11400
rect 14320 11364 14484 11396
rect 14516 11364 14644 11396
rect 14676 11364 14804 11396
rect 14836 11364 14964 11396
rect 14996 11364 15000 11396
rect 14320 11360 15000 11364
rect 80 11316 680 11320
rect 80 11284 84 11316
rect 116 11284 680 11316
rect 80 11280 680 11284
rect 14480 11316 15000 11320
rect 14480 11284 14484 11316
rect 14516 11284 14644 11316
rect 14676 11284 14804 11316
rect 14836 11284 14964 11316
rect 14996 11284 15000 11316
rect 14480 11280 15000 11284
rect 0 11236 680 11240
rect 0 11204 4 11236
rect 36 11204 164 11236
rect 196 11204 324 11236
rect 356 11204 484 11236
rect 516 11204 680 11236
rect 0 11200 680 11204
rect 14320 11236 15000 11240
rect 14320 11204 14484 11236
rect 14516 11204 14644 11236
rect 14676 11204 14804 11236
rect 14836 11204 14964 11236
rect 14996 11204 15000 11236
rect 14320 11200 15000 11204
rect 0 11156 200 11160
rect 0 11124 4 11156
rect 36 11124 164 11156
rect 196 11124 200 11156
rect 0 11120 200 11124
rect 240 11156 680 11160
rect 240 11124 244 11156
rect 276 11124 680 11156
rect 240 11120 680 11124
rect 14480 11156 15000 11160
rect 14480 11124 14484 11156
rect 14516 11124 14644 11156
rect 14676 11124 14804 11156
rect 14836 11124 14964 11156
rect 14996 11124 15000 11156
rect 14480 11120 15000 11124
rect 0 11076 520 11080
rect 0 11044 4 11076
rect 36 11044 164 11076
rect 196 11044 324 11076
rect 356 11044 484 11076
rect 516 11044 520 11076
rect 0 11040 520 11044
rect 14320 11076 15000 11080
rect 14320 11044 14484 11076
rect 14516 11044 14644 11076
rect 14676 11044 14804 11076
rect 14836 11044 14964 11076
rect 14996 11044 15000 11076
rect 14320 11040 15000 11044
rect 0 10996 520 11000
rect 0 10964 4 10996
rect 36 10964 164 10996
rect 196 10964 324 10996
rect 356 10964 484 10996
rect 516 10964 520 10996
rect 0 10960 520 10964
rect 14480 10996 15000 11000
rect 14480 10964 14484 10996
rect 14516 10964 14644 10996
rect 14676 10964 14804 10996
rect 14836 10964 14964 10996
rect 14996 10964 15000 10996
rect 14480 10960 15000 10964
rect 0 10916 520 10920
rect 0 10884 4 10916
rect 36 10884 164 10916
rect 196 10884 324 10916
rect 356 10884 484 10916
rect 516 10884 520 10916
rect 0 10880 520 10884
rect 14480 10916 15000 10920
rect 14480 10884 14484 10916
rect 14516 10884 14644 10916
rect 14676 10884 14804 10916
rect 14836 10884 14964 10916
rect 14996 10884 15000 10916
rect 14480 10880 15000 10884
rect 0 10836 520 10840
rect 0 10804 4 10836
rect 36 10804 164 10836
rect 196 10804 324 10836
rect 356 10804 484 10836
rect 516 10804 520 10836
rect 0 10800 520 10804
rect 14480 10836 15000 10840
rect 14480 10804 14484 10836
rect 14516 10804 14644 10836
rect 14676 10804 14804 10836
rect 14836 10804 14964 10836
rect 14996 10804 15000 10836
rect 14480 10800 15000 10804
rect 0 10756 520 10760
rect 0 10724 4 10756
rect 36 10724 164 10756
rect 196 10724 324 10756
rect 356 10724 484 10756
rect 516 10724 520 10756
rect 0 10720 520 10724
rect 14480 10756 15000 10760
rect 14480 10724 14484 10756
rect 14516 10724 14644 10756
rect 14676 10724 14804 10756
rect 14836 10724 14964 10756
rect 14996 10724 15000 10756
rect 14480 10720 15000 10724
rect 0 10676 520 10680
rect 0 10644 4 10676
rect 36 10644 164 10676
rect 196 10644 324 10676
rect 356 10644 484 10676
rect 516 10644 520 10676
rect 0 10640 520 10644
rect 14480 10676 15000 10680
rect 14480 10644 14484 10676
rect 14516 10644 14644 10676
rect 14676 10644 14804 10676
rect 14836 10644 14964 10676
rect 14996 10644 15000 10676
rect 14480 10640 15000 10644
rect 0 10596 520 10600
rect 0 10564 4 10596
rect 36 10564 164 10596
rect 196 10564 324 10596
rect 356 10564 484 10596
rect 516 10564 520 10596
rect 0 10560 520 10564
rect 14480 10596 15000 10600
rect 14480 10564 14484 10596
rect 14516 10564 14644 10596
rect 14676 10564 14804 10596
rect 14836 10564 14964 10596
rect 14996 10564 15000 10596
rect 14480 10560 15000 10564
rect 0 10516 520 10520
rect 0 10484 4 10516
rect 36 10484 164 10516
rect 196 10484 324 10516
rect 356 10484 484 10516
rect 516 10484 520 10516
rect 0 10480 520 10484
rect 14480 10516 15000 10520
rect 14480 10484 14484 10516
rect 14516 10484 14644 10516
rect 14676 10484 14804 10516
rect 14836 10484 14964 10516
rect 14996 10484 15000 10516
rect 14480 10480 15000 10484
rect 0 10436 520 10440
rect 0 10404 4 10436
rect 36 10404 164 10436
rect 196 10404 324 10436
rect 356 10404 484 10436
rect 516 10404 520 10436
rect 0 10400 520 10404
rect 14480 10436 15000 10440
rect 14480 10404 14484 10436
rect 14516 10404 14644 10436
rect 14676 10404 14804 10436
rect 14836 10404 14964 10436
rect 14996 10404 15000 10436
rect 14480 10400 15000 10404
rect 0 10356 520 10360
rect 0 10324 4 10356
rect 36 10324 164 10356
rect 196 10324 324 10356
rect 356 10324 484 10356
rect 516 10324 520 10356
rect 0 10320 520 10324
rect 14480 10356 15000 10360
rect 14480 10324 14484 10356
rect 14516 10324 14644 10356
rect 14676 10324 14804 10356
rect 14836 10324 14964 10356
rect 14996 10324 15000 10356
rect 14480 10320 15000 10324
rect 0 10276 520 10280
rect 0 10244 4 10276
rect 36 10244 164 10276
rect 196 10244 324 10276
rect 356 10244 484 10276
rect 516 10244 520 10276
rect 0 10240 520 10244
rect 14480 10276 15000 10280
rect 14480 10244 14484 10276
rect 14516 10244 14644 10276
rect 14676 10244 14804 10276
rect 14836 10244 14964 10276
rect 14996 10244 15000 10276
rect 14480 10240 15000 10244
rect 0 10196 520 10200
rect 0 10164 4 10196
rect 36 10164 164 10196
rect 196 10164 324 10196
rect 356 10164 484 10196
rect 516 10164 520 10196
rect 0 10160 520 10164
rect 14480 10196 15000 10200
rect 14480 10164 14484 10196
rect 14516 10164 14644 10196
rect 14676 10164 14804 10196
rect 14836 10164 14964 10196
rect 14996 10164 15000 10196
rect 14480 10160 15000 10164
rect 0 10116 520 10120
rect 0 10084 4 10116
rect 36 10084 164 10116
rect 196 10084 324 10116
rect 356 10084 484 10116
rect 516 10084 520 10116
rect 0 10080 520 10084
rect 14480 10116 15000 10120
rect 14480 10084 14484 10116
rect 14516 10084 14644 10116
rect 14676 10084 14804 10116
rect 14836 10084 14964 10116
rect 14996 10084 15000 10116
rect 14480 10080 15000 10084
rect 0 10036 520 10040
rect 0 10004 4 10036
rect 36 10004 164 10036
rect 196 10004 324 10036
rect 356 10004 484 10036
rect 516 10004 520 10036
rect 0 10000 520 10004
rect 14480 10036 15000 10040
rect 14480 10004 14484 10036
rect 14516 10004 14644 10036
rect 14676 10004 14804 10036
rect 14836 10004 14964 10036
rect 14996 10004 15000 10036
rect 14480 10000 15000 10004
rect 0 9956 520 9960
rect 0 9924 4 9956
rect 36 9924 164 9956
rect 196 9924 324 9956
rect 356 9924 484 9956
rect 516 9924 520 9956
rect 0 9920 520 9924
rect 14480 9956 15000 9960
rect 14480 9924 14484 9956
rect 14516 9924 14644 9956
rect 14676 9924 14804 9956
rect 14836 9924 14964 9956
rect 14996 9924 15000 9956
rect 14480 9920 15000 9924
rect 0 9876 360 9880
rect 0 9844 4 9876
rect 36 9844 164 9876
rect 196 9844 324 9876
rect 356 9844 360 9876
rect 0 9840 360 9844
rect 400 9876 680 9880
rect 400 9844 404 9876
rect 436 9844 680 9876
rect 400 9840 680 9844
rect 14480 9876 15000 9880
rect 14480 9844 14484 9876
rect 14516 9844 14644 9876
rect 14676 9844 14804 9876
rect 14836 9844 14964 9876
rect 14996 9844 15000 9876
rect 14480 9840 15000 9844
rect 0 9796 520 9800
rect 0 9764 4 9796
rect 36 9764 164 9796
rect 196 9764 324 9796
rect 356 9764 484 9796
rect 516 9764 520 9796
rect 0 9760 520 9764
rect 14480 9796 15000 9800
rect 14480 9764 14484 9796
rect 14516 9764 14644 9796
rect 14676 9764 14804 9796
rect 14836 9764 14964 9796
rect 14996 9764 15000 9796
rect 14480 9760 15000 9764
rect 0 9716 520 9720
rect 0 9684 4 9716
rect 36 9684 164 9716
rect 196 9684 324 9716
rect 356 9684 484 9716
rect 516 9684 520 9716
rect 0 9680 520 9684
rect 14480 9716 15000 9720
rect 14480 9684 14484 9716
rect 14516 9684 14644 9716
rect 14676 9684 14804 9716
rect 14836 9684 14964 9716
rect 14996 9684 15000 9716
rect 14480 9680 15000 9684
rect 0 9636 520 9640
rect 0 9604 4 9636
rect 36 9604 164 9636
rect 196 9604 324 9636
rect 356 9604 484 9636
rect 516 9604 520 9636
rect 0 9600 520 9604
rect 14480 9636 15000 9640
rect 14480 9604 14484 9636
rect 14516 9604 14644 9636
rect 14676 9604 14804 9636
rect 14836 9604 14964 9636
rect 14996 9604 15000 9636
rect 14480 9600 15000 9604
rect 0 9556 520 9560
rect 0 9524 4 9556
rect 36 9524 164 9556
rect 196 9524 324 9556
rect 356 9524 484 9556
rect 516 9524 520 9556
rect 0 9520 520 9524
rect 14480 9556 15000 9560
rect 14480 9524 14484 9556
rect 14516 9524 14644 9556
rect 14676 9524 14804 9556
rect 14836 9524 14964 9556
rect 14996 9524 15000 9556
rect 14480 9520 15000 9524
rect 0 9476 520 9480
rect 0 9444 4 9476
rect 36 9444 164 9476
rect 196 9444 324 9476
rect 356 9444 484 9476
rect 516 9444 520 9476
rect 0 9440 520 9444
rect 14480 9476 15000 9480
rect 14480 9444 14484 9476
rect 14516 9444 14644 9476
rect 14676 9444 14804 9476
rect 14836 9444 14964 9476
rect 14996 9444 15000 9476
rect 14480 9440 15000 9444
rect 0 9396 520 9400
rect 0 9364 4 9396
rect 36 9364 164 9396
rect 196 9364 324 9396
rect 356 9364 484 9396
rect 516 9364 520 9396
rect 0 9360 520 9364
rect 14480 9396 15000 9400
rect 14480 9364 14484 9396
rect 14516 9364 14644 9396
rect 14676 9364 14804 9396
rect 14836 9364 14964 9396
rect 14996 9364 15000 9396
rect 14480 9360 15000 9364
rect 0 9316 520 9320
rect 0 9284 4 9316
rect 36 9284 164 9316
rect 196 9284 324 9316
rect 356 9284 484 9316
rect 516 9284 520 9316
rect 0 9280 520 9284
rect 14480 9316 15000 9320
rect 14480 9284 14484 9316
rect 14516 9284 14644 9316
rect 14676 9284 14804 9316
rect 14836 9284 14964 9316
rect 14996 9284 15000 9316
rect 14480 9280 15000 9284
rect 0 9236 520 9240
rect 0 9204 4 9236
rect 36 9204 164 9236
rect 196 9204 324 9236
rect 356 9204 484 9236
rect 516 9204 520 9236
rect 0 9200 520 9204
rect 14480 9236 15000 9240
rect 14480 9204 14484 9236
rect 14516 9204 14644 9236
rect 14676 9204 14804 9236
rect 14836 9204 14964 9236
rect 14996 9204 15000 9236
rect 14480 9200 15000 9204
rect 0 9156 520 9160
rect 0 9124 4 9156
rect 36 9124 164 9156
rect 196 9124 324 9156
rect 356 9124 484 9156
rect 516 9124 520 9156
rect 0 9120 520 9124
rect 14480 9156 15000 9160
rect 14480 9124 14484 9156
rect 14516 9124 14644 9156
rect 14676 9124 14804 9156
rect 14836 9124 14964 9156
rect 14996 9124 15000 9156
rect 14480 9120 15000 9124
rect 0 9076 520 9080
rect 0 9044 4 9076
rect 36 9044 164 9076
rect 196 9044 324 9076
rect 356 9044 484 9076
rect 516 9044 520 9076
rect 0 9040 520 9044
rect 14480 9076 15000 9080
rect 14480 9044 14484 9076
rect 14516 9044 14644 9076
rect 14676 9044 14804 9076
rect 14836 9044 14964 9076
rect 14996 9044 15000 9076
rect 14480 9040 15000 9044
rect 0 8996 520 9000
rect 0 8964 4 8996
rect 36 8964 164 8996
rect 196 8964 324 8996
rect 356 8964 484 8996
rect 516 8964 520 8996
rect 0 8960 520 8964
rect 14480 8996 15000 9000
rect 14480 8964 14484 8996
rect 14516 8964 14644 8996
rect 14676 8964 14804 8996
rect 14836 8964 14964 8996
rect 14996 8964 15000 8996
rect 14480 8960 15000 8964
rect 0 8916 520 8920
rect 0 8884 4 8916
rect 36 8884 164 8916
rect 196 8884 324 8916
rect 356 8884 484 8916
rect 516 8884 520 8916
rect 0 8880 520 8884
rect 14480 8916 15000 8920
rect 14480 8884 14484 8916
rect 14516 8884 14644 8916
rect 14676 8884 14804 8916
rect 14836 8884 14964 8916
rect 14996 8884 15000 8916
rect 14480 8880 15000 8884
rect 0 8836 520 8840
rect 0 8804 4 8836
rect 36 8804 164 8836
rect 196 8804 324 8836
rect 356 8804 484 8836
rect 516 8804 520 8836
rect 0 8800 520 8804
rect 14480 8836 15000 8840
rect 14480 8804 14484 8836
rect 14516 8804 14644 8836
rect 14676 8804 14804 8836
rect 14836 8804 14964 8836
rect 14996 8804 15000 8836
rect 14480 8800 15000 8804
rect 0 8756 520 8760
rect 0 8724 4 8756
rect 36 8724 164 8756
rect 196 8724 324 8756
rect 356 8724 484 8756
rect 516 8724 520 8756
rect 0 8720 520 8724
rect 14480 8756 15000 8760
rect 14480 8724 14484 8756
rect 14516 8724 14644 8756
rect 14676 8724 14804 8756
rect 14836 8724 14964 8756
rect 14996 8724 15000 8756
rect 14480 8720 15000 8724
rect 0 8676 680 8680
rect 0 8644 4 8676
rect 36 8644 164 8676
rect 196 8644 324 8676
rect 356 8644 484 8676
rect 516 8644 680 8676
rect 0 8640 680 8644
rect 14320 8676 15000 8680
rect 14320 8644 14484 8676
rect 14516 8644 14644 8676
rect 14676 8644 14804 8676
rect 14836 8644 14964 8676
rect 14996 8644 15000 8676
rect 14320 8640 15000 8644
rect 0 8596 200 8600
rect 0 8564 4 8596
rect 36 8564 164 8596
rect 196 8564 200 8596
rect 0 8560 200 8564
rect 240 8596 680 8600
rect 240 8564 244 8596
rect 276 8564 680 8596
rect 240 8560 680 8564
rect 14480 8596 15000 8600
rect 14480 8564 14484 8596
rect 14516 8564 14644 8596
rect 14676 8564 14804 8596
rect 14836 8564 14964 8596
rect 14996 8564 15000 8596
rect 14480 8560 15000 8564
rect 0 8516 680 8520
rect 0 8484 4 8516
rect 36 8484 164 8516
rect 196 8484 324 8516
rect 356 8484 484 8516
rect 516 8484 680 8516
rect 0 8480 680 8484
rect 14320 8516 15000 8520
rect 14320 8484 14484 8516
rect 14516 8484 14644 8516
rect 14676 8484 14804 8516
rect 14836 8484 14964 8516
rect 14996 8484 15000 8516
rect 14320 8480 15000 8484
rect 80 8436 680 8440
rect 80 8404 84 8436
rect 116 8404 680 8436
rect 80 8400 680 8404
rect 14480 8436 15000 8440
rect 14480 8404 14484 8436
rect 14516 8404 14644 8436
rect 14676 8404 14804 8436
rect 14836 8404 14964 8436
rect 14996 8404 15000 8436
rect 14480 8400 15000 8404
rect 0 8356 680 8360
rect 0 8324 4 8356
rect 36 8324 164 8356
rect 196 8324 324 8356
rect 356 8324 484 8356
rect 516 8324 680 8356
rect 0 8320 680 8324
rect 14320 8356 15000 8360
rect 14320 8324 14484 8356
rect 14516 8324 14644 8356
rect 14676 8324 14804 8356
rect 14836 8324 14964 8356
rect 14996 8324 15000 8356
rect 14320 8320 15000 8324
rect 0 8276 520 8280
rect 0 8244 4 8276
rect 36 8244 164 8276
rect 196 8244 324 8276
rect 356 8244 484 8276
rect 516 8244 520 8276
rect 0 8240 520 8244
rect 14480 8276 15000 8280
rect 14480 8244 14484 8276
rect 14516 8244 14644 8276
rect 14676 8244 14804 8276
rect 14836 8244 14964 8276
rect 14996 8244 15000 8276
rect 14480 8240 15000 8244
rect 0 8196 520 8200
rect 0 8164 4 8196
rect 36 8164 164 8196
rect 196 8164 324 8196
rect 356 8164 484 8196
rect 516 8164 520 8196
rect 0 8160 520 8164
rect 14480 8196 15000 8200
rect 14480 8164 14484 8196
rect 14516 8164 14644 8196
rect 14676 8164 14804 8196
rect 14836 8164 14964 8196
rect 14996 8164 15000 8196
rect 14480 8160 15000 8164
rect 0 8116 680 8120
rect 0 8084 4 8116
rect 36 8084 164 8116
rect 196 8084 324 8116
rect 356 8084 484 8116
rect 516 8084 680 8116
rect 0 8080 680 8084
rect 14320 8116 15000 8120
rect 14320 8084 14484 8116
rect 14516 8084 14644 8116
rect 14676 8084 14804 8116
rect 14836 8084 14964 8116
rect 14996 8084 15000 8116
rect 14320 8080 15000 8084
rect 80 8036 680 8040
rect 80 8004 84 8036
rect 116 8004 680 8036
rect 80 8000 680 8004
rect 14480 8036 15000 8040
rect 14480 8004 14484 8036
rect 14516 8004 14644 8036
rect 14676 8004 14804 8036
rect 14836 8004 14964 8036
rect 14996 8004 15000 8036
rect 14480 8000 15000 8004
rect 0 7956 680 7960
rect 0 7924 4 7956
rect 36 7924 164 7956
rect 196 7924 324 7956
rect 356 7924 484 7956
rect 516 7924 680 7956
rect 0 7920 680 7924
rect 14320 7956 15000 7960
rect 14320 7924 14484 7956
rect 14516 7924 14644 7956
rect 14676 7924 14804 7956
rect 14836 7924 14964 7956
rect 14996 7924 15000 7956
rect 14320 7920 15000 7924
rect 0 7876 200 7880
rect 0 7844 4 7876
rect 36 7844 164 7876
rect 196 7844 200 7876
rect 0 7840 200 7844
rect 240 7876 680 7880
rect 240 7844 244 7876
rect 276 7844 680 7876
rect 240 7840 680 7844
rect 14480 7876 15000 7880
rect 14480 7844 14484 7876
rect 14516 7844 14644 7876
rect 14676 7844 14804 7876
rect 14836 7844 14964 7876
rect 14996 7844 15000 7876
rect 14480 7840 15000 7844
rect 0 7796 680 7800
rect 0 7764 4 7796
rect 36 7764 164 7796
rect 196 7764 324 7796
rect 356 7764 484 7796
rect 516 7764 680 7796
rect 0 7760 680 7764
rect 14320 7796 15000 7800
rect 14320 7764 14484 7796
rect 14516 7764 14644 7796
rect 14676 7764 14804 7796
rect 14836 7764 14964 7796
rect 14996 7764 15000 7796
rect 14320 7760 15000 7764
rect 0 7716 520 7720
rect 0 7684 4 7716
rect 36 7684 164 7716
rect 196 7684 324 7716
rect 356 7684 484 7716
rect 516 7684 520 7716
rect 0 7680 520 7684
rect 14480 7716 15000 7720
rect 14480 7684 14484 7716
rect 14516 7684 14644 7716
rect 14676 7684 14804 7716
rect 14836 7684 14964 7716
rect 14996 7684 15000 7716
rect 14480 7680 15000 7684
rect 0 7636 520 7640
rect 0 7604 4 7636
rect 36 7604 164 7636
rect 196 7604 324 7636
rect 356 7604 484 7636
rect 516 7604 520 7636
rect 0 7600 520 7604
rect 14480 7636 15000 7640
rect 14480 7604 14484 7636
rect 14516 7604 14644 7636
rect 14676 7604 14804 7636
rect 14836 7604 14964 7636
rect 14996 7604 15000 7636
rect 14480 7600 15000 7604
rect 0 7556 520 7560
rect 0 7524 4 7556
rect 36 7524 164 7556
rect 196 7524 324 7556
rect 356 7524 484 7556
rect 516 7524 520 7556
rect 0 7520 520 7524
rect 14480 7556 15000 7560
rect 14480 7524 14484 7556
rect 14516 7524 14644 7556
rect 14676 7524 14804 7556
rect 14836 7524 14964 7556
rect 14996 7524 15000 7556
rect 14480 7520 15000 7524
rect 0 7476 520 7480
rect 0 7444 4 7476
rect 36 7444 164 7476
rect 196 7444 324 7476
rect 356 7444 484 7476
rect 516 7444 520 7476
rect 0 7440 520 7444
rect 14480 7476 15000 7480
rect 14480 7444 14484 7476
rect 14516 7444 14644 7476
rect 14676 7444 14804 7476
rect 14836 7444 14964 7476
rect 14996 7444 15000 7476
rect 14480 7440 15000 7444
rect 0 7396 520 7400
rect 0 7364 4 7396
rect 36 7364 164 7396
rect 196 7364 324 7396
rect 356 7364 484 7396
rect 516 7364 520 7396
rect 0 7360 520 7364
rect 14480 7396 15000 7400
rect 14480 7364 14484 7396
rect 14516 7364 14644 7396
rect 14676 7364 14804 7396
rect 14836 7364 14964 7396
rect 14996 7364 15000 7396
rect 14480 7360 15000 7364
rect 0 7316 520 7320
rect 0 7284 4 7316
rect 36 7284 164 7316
rect 196 7284 324 7316
rect 356 7284 484 7316
rect 516 7284 520 7316
rect 0 7280 520 7284
rect 14480 7316 15000 7320
rect 14480 7284 14484 7316
rect 14516 7284 14644 7316
rect 14676 7284 14804 7316
rect 14836 7284 14964 7316
rect 14996 7284 15000 7316
rect 14480 7280 15000 7284
rect 0 7236 520 7240
rect 0 7204 4 7236
rect 36 7204 164 7236
rect 196 7204 324 7236
rect 356 7204 484 7236
rect 516 7204 520 7236
rect 0 7200 520 7204
rect 14480 7236 15000 7240
rect 14480 7204 14484 7236
rect 14516 7204 14644 7236
rect 14676 7204 14804 7236
rect 14836 7204 14964 7236
rect 14996 7204 15000 7236
rect 14480 7200 15000 7204
rect 0 7156 520 7160
rect 0 7124 4 7156
rect 36 7124 164 7156
rect 196 7124 324 7156
rect 356 7124 484 7156
rect 516 7124 520 7156
rect 0 7120 520 7124
rect 14480 7156 15000 7160
rect 14480 7124 14484 7156
rect 14516 7124 14644 7156
rect 14676 7124 14804 7156
rect 14836 7124 14964 7156
rect 14996 7124 15000 7156
rect 14480 7120 15000 7124
rect 0 7076 520 7080
rect 0 7044 4 7076
rect 36 7044 164 7076
rect 196 7044 324 7076
rect 356 7044 484 7076
rect 516 7044 520 7076
rect 0 7040 520 7044
rect 14480 7076 15000 7080
rect 14480 7044 14484 7076
rect 14516 7044 14644 7076
rect 14676 7044 14804 7076
rect 14836 7044 14964 7076
rect 14996 7044 15000 7076
rect 14480 7040 15000 7044
rect 0 6996 520 7000
rect 0 6964 4 6996
rect 36 6964 164 6996
rect 196 6964 324 6996
rect 356 6964 484 6996
rect 516 6964 520 6996
rect 0 6960 520 6964
rect 14480 6996 15000 7000
rect 14480 6964 14484 6996
rect 14516 6964 14644 6996
rect 14676 6964 14804 6996
rect 14836 6964 14964 6996
rect 14996 6964 15000 6996
rect 14480 6960 15000 6964
rect 0 6916 520 6920
rect 0 6884 4 6916
rect 36 6884 164 6916
rect 196 6884 324 6916
rect 356 6884 484 6916
rect 516 6884 520 6916
rect 0 6880 520 6884
rect 14480 6916 15000 6920
rect 14480 6884 14484 6916
rect 14516 6884 14644 6916
rect 14676 6884 14804 6916
rect 14836 6884 14964 6916
rect 14996 6884 15000 6916
rect 14480 6880 15000 6884
rect 0 6836 520 6840
rect 0 6804 4 6836
rect 36 6804 164 6836
rect 196 6804 324 6836
rect 356 6804 484 6836
rect 516 6804 520 6836
rect 0 6800 520 6804
rect 14480 6836 15000 6840
rect 14480 6804 14484 6836
rect 14516 6804 14644 6836
rect 14676 6804 14804 6836
rect 14836 6804 14964 6836
rect 14996 6804 15000 6836
rect 14480 6800 15000 6804
rect 0 6756 520 6760
rect 0 6724 4 6756
rect 36 6724 164 6756
rect 196 6724 324 6756
rect 356 6724 484 6756
rect 516 6724 520 6756
rect 0 6720 520 6724
rect 14480 6756 15000 6760
rect 14480 6724 14484 6756
rect 14516 6724 14644 6756
rect 14676 6724 14804 6756
rect 14836 6724 14964 6756
rect 14996 6724 15000 6756
rect 14480 6720 15000 6724
rect 0 6676 520 6680
rect 0 6644 4 6676
rect 36 6644 164 6676
rect 196 6644 324 6676
rect 356 6644 484 6676
rect 516 6644 520 6676
rect 0 6640 520 6644
rect 14480 6676 15000 6680
rect 14480 6644 14484 6676
rect 14516 6644 14644 6676
rect 14676 6644 14804 6676
rect 14836 6644 14964 6676
rect 14996 6644 15000 6676
rect 14480 6640 15000 6644
rect 0 6596 360 6600
rect 0 6564 4 6596
rect 36 6564 164 6596
rect 196 6564 324 6596
rect 356 6564 360 6596
rect 0 6560 360 6564
rect 400 6596 680 6600
rect 400 6564 404 6596
rect 436 6564 680 6596
rect 400 6560 680 6564
rect 14480 6596 15000 6600
rect 14480 6564 14484 6596
rect 14516 6564 14644 6596
rect 14676 6564 14804 6596
rect 14836 6564 14964 6596
rect 14996 6564 15000 6596
rect 14480 6560 15000 6564
rect 0 6516 520 6520
rect 0 6484 4 6516
rect 36 6484 164 6516
rect 196 6484 324 6516
rect 356 6484 484 6516
rect 516 6484 520 6516
rect 0 6480 520 6484
rect 14480 6516 15000 6520
rect 14480 6484 14484 6516
rect 14516 6484 14644 6516
rect 14676 6484 14804 6516
rect 14836 6484 14964 6516
rect 14996 6484 15000 6516
rect 14480 6480 15000 6484
rect 0 6436 520 6440
rect 0 6404 4 6436
rect 36 6404 164 6436
rect 196 6404 324 6436
rect 356 6404 484 6436
rect 516 6404 520 6436
rect 0 6400 520 6404
rect 14480 6436 15000 6440
rect 14480 6404 14484 6436
rect 14516 6404 14644 6436
rect 14676 6404 14804 6436
rect 14836 6404 14964 6436
rect 14996 6404 15000 6436
rect 14480 6400 15000 6404
rect 0 6356 520 6360
rect 0 6324 4 6356
rect 36 6324 164 6356
rect 196 6324 324 6356
rect 356 6324 484 6356
rect 516 6324 520 6356
rect 0 6320 520 6324
rect 14480 6356 15000 6360
rect 14480 6324 14484 6356
rect 14516 6324 14644 6356
rect 14676 6324 14804 6356
rect 14836 6324 14964 6356
rect 14996 6324 15000 6356
rect 14480 6320 15000 6324
rect 0 6276 520 6280
rect 0 6244 4 6276
rect 36 6244 164 6276
rect 196 6244 324 6276
rect 356 6244 484 6276
rect 516 6244 520 6276
rect 0 6240 520 6244
rect 14480 6276 15000 6280
rect 14480 6244 14484 6276
rect 14516 6244 14644 6276
rect 14676 6244 14804 6276
rect 14836 6244 14964 6276
rect 14996 6244 15000 6276
rect 14480 6240 15000 6244
rect 0 6196 520 6200
rect 0 6164 4 6196
rect 36 6164 164 6196
rect 196 6164 324 6196
rect 356 6164 484 6196
rect 516 6164 520 6196
rect 0 6160 520 6164
rect 14480 6196 15000 6200
rect 14480 6164 14484 6196
rect 14516 6164 14644 6196
rect 14676 6164 14804 6196
rect 14836 6164 14964 6196
rect 14996 6164 15000 6196
rect 14480 6160 15000 6164
rect 0 6116 520 6120
rect 0 6084 4 6116
rect 36 6084 164 6116
rect 196 6084 324 6116
rect 356 6084 484 6116
rect 516 6084 520 6116
rect 0 6080 520 6084
rect 14480 6116 15000 6120
rect 14480 6084 14484 6116
rect 14516 6084 14644 6116
rect 14676 6084 14804 6116
rect 14836 6084 14964 6116
rect 14996 6084 15000 6116
rect 14480 6080 15000 6084
rect 0 6036 520 6040
rect 0 6004 4 6036
rect 36 6004 164 6036
rect 196 6004 324 6036
rect 356 6004 484 6036
rect 516 6004 520 6036
rect 0 6000 520 6004
rect 14480 6036 15000 6040
rect 14480 6004 14484 6036
rect 14516 6004 14644 6036
rect 14676 6004 14804 6036
rect 14836 6004 14964 6036
rect 14996 6004 15000 6036
rect 14480 6000 15000 6004
rect 0 5956 520 5960
rect 0 5924 4 5956
rect 36 5924 164 5956
rect 196 5924 324 5956
rect 356 5924 484 5956
rect 516 5924 520 5956
rect 0 5920 520 5924
rect 14480 5956 15000 5960
rect 14480 5924 14484 5956
rect 14516 5924 14644 5956
rect 14676 5924 14804 5956
rect 14836 5924 14964 5956
rect 14996 5924 15000 5956
rect 14480 5920 15000 5924
rect 0 5876 520 5880
rect 0 5844 4 5876
rect 36 5844 164 5876
rect 196 5844 324 5876
rect 356 5844 484 5876
rect 516 5844 520 5876
rect 0 5840 520 5844
rect 14480 5876 15000 5880
rect 14480 5844 14484 5876
rect 14516 5844 14644 5876
rect 14676 5844 14804 5876
rect 14836 5844 14964 5876
rect 14996 5844 15000 5876
rect 14480 5840 15000 5844
rect 0 5796 520 5800
rect 0 5764 4 5796
rect 36 5764 164 5796
rect 196 5764 324 5796
rect 356 5764 484 5796
rect 516 5764 520 5796
rect 0 5760 520 5764
rect 14480 5796 15000 5800
rect 14480 5764 14484 5796
rect 14516 5764 14644 5796
rect 14676 5764 14804 5796
rect 14836 5764 14964 5796
rect 14996 5764 15000 5796
rect 14480 5760 15000 5764
rect 0 5716 520 5720
rect 0 5684 4 5716
rect 36 5684 164 5716
rect 196 5684 324 5716
rect 356 5684 484 5716
rect 516 5684 520 5716
rect 0 5680 520 5684
rect 14480 5716 15000 5720
rect 14480 5684 14484 5716
rect 14516 5684 14644 5716
rect 14676 5684 14804 5716
rect 14836 5684 14964 5716
rect 14996 5684 15000 5716
rect 14480 5680 15000 5684
rect 0 5636 520 5640
rect 0 5604 4 5636
rect 36 5604 164 5636
rect 196 5604 324 5636
rect 356 5604 484 5636
rect 516 5604 520 5636
rect 0 5600 520 5604
rect 14480 5636 15000 5640
rect 14480 5604 14484 5636
rect 14516 5604 14644 5636
rect 14676 5604 14804 5636
rect 14836 5604 14964 5636
rect 14996 5604 15000 5636
rect 14480 5600 15000 5604
rect 0 5556 520 5560
rect 0 5524 4 5556
rect 36 5524 164 5556
rect 196 5524 324 5556
rect 356 5524 484 5556
rect 516 5524 520 5556
rect 0 5520 520 5524
rect 14480 5556 15000 5560
rect 14480 5524 14484 5556
rect 14516 5524 14644 5556
rect 14676 5524 14804 5556
rect 14836 5524 14964 5556
rect 14996 5524 15000 5556
rect 14480 5520 15000 5524
rect 0 5476 520 5480
rect 0 5444 4 5476
rect 36 5444 164 5476
rect 196 5444 324 5476
rect 356 5444 484 5476
rect 516 5444 520 5476
rect 0 5440 520 5444
rect 14480 5476 15000 5480
rect 14480 5444 14484 5476
rect 14516 5444 14644 5476
rect 14676 5444 14804 5476
rect 14836 5444 14964 5476
rect 14996 5444 15000 5476
rect 14480 5440 15000 5444
rect 0 5396 680 5400
rect 0 5364 4 5396
rect 36 5364 164 5396
rect 196 5364 324 5396
rect 356 5364 484 5396
rect 516 5364 680 5396
rect 0 5360 680 5364
rect 14320 5396 15000 5400
rect 14320 5364 14484 5396
rect 14516 5364 14644 5396
rect 14676 5364 14804 5396
rect 14836 5364 14964 5396
rect 14996 5364 15000 5396
rect 14320 5360 15000 5364
rect 0 5316 200 5320
rect 0 5284 4 5316
rect 36 5284 164 5316
rect 196 5284 200 5316
rect 0 5280 200 5284
rect 240 5316 680 5320
rect 240 5284 244 5316
rect 276 5284 680 5316
rect 240 5280 680 5284
rect 14480 5316 15000 5320
rect 14480 5284 14484 5316
rect 14516 5284 14644 5316
rect 14676 5284 14804 5316
rect 14836 5284 14964 5316
rect 14996 5284 15000 5316
rect 14480 5280 15000 5284
rect 0 5236 680 5240
rect 0 5204 4 5236
rect 36 5204 164 5236
rect 196 5204 324 5236
rect 356 5204 484 5236
rect 516 5204 680 5236
rect 0 5200 680 5204
rect 14320 5236 15000 5240
rect 14320 5204 14484 5236
rect 14516 5204 14644 5236
rect 14676 5204 14804 5236
rect 14836 5204 14964 5236
rect 14996 5204 15000 5236
rect 14320 5200 15000 5204
rect 80 5156 680 5160
rect 80 5124 84 5156
rect 116 5124 680 5156
rect 80 5120 680 5124
rect 14480 5156 15000 5160
rect 14480 5124 14484 5156
rect 14516 5124 14644 5156
rect 14676 5124 14804 5156
rect 14836 5124 14964 5156
rect 14996 5124 15000 5156
rect 14480 5120 15000 5124
rect 0 5076 680 5080
rect 0 5044 4 5076
rect 36 5044 164 5076
rect 196 5044 324 5076
rect 356 5044 484 5076
rect 516 5044 680 5076
rect 0 5040 680 5044
rect 14320 5076 15000 5080
rect 14320 5044 14484 5076
rect 14516 5044 14644 5076
rect 14676 5044 14804 5076
rect 14836 5044 14964 5076
rect 14996 5044 15000 5076
rect 14320 5040 15000 5044
rect 0 4996 520 5000
rect 0 4964 4 4996
rect 36 4964 164 4996
rect 196 4964 324 4996
rect 356 4964 484 4996
rect 516 4964 520 4996
rect 0 4960 520 4964
rect 14480 4996 15000 5000
rect 14480 4964 14484 4996
rect 14516 4964 14644 4996
rect 14676 4964 14804 4996
rect 14836 4964 14964 4996
rect 14996 4964 15000 4996
rect 14480 4960 15000 4964
rect 0 4916 520 4920
rect 0 4884 4 4916
rect 36 4884 164 4916
rect 196 4884 324 4916
rect 356 4884 484 4916
rect 516 4884 520 4916
rect 0 4880 520 4884
rect 14480 4916 15000 4920
rect 14480 4884 14484 4916
rect 14516 4884 14644 4916
rect 14676 4884 14804 4916
rect 14836 4884 14964 4916
rect 14996 4884 15000 4916
rect 14480 4880 15000 4884
rect 0 4836 680 4840
rect 0 4804 4 4836
rect 36 4804 164 4836
rect 196 4804 324 4836
rect 356 4804 484 4836
rect 516 4804 680 4836
rect 0 4800 680 4804
rect 14320 4836 15000 4840
rect 14320 4804 14484 4836
rect 14516 4804 14644 4836
rect 14676 4804 14804 4836
rect 14836 4804 14964 4836
rect 14996 4804 15000 4836
rect 14320 4800 15000 4804
rect 0 4756 520 4760
rect 0 4724 4 4756
rect 36 4724 164 4756
rect 196 4724 324 4756
rect 356 4724 484 4756
rect 516 4724 520 4756
rect 0 4720 520 4724
rect 14320 4756 15000 4760
rect 14320 4724 14884 4756
rect 14916 4724 15000 4756
rect 14320 4720 15000 4724
rect 0 4676 680 4680
rect 0 4644 4 4676
rect 36 4644 164 4676
rect 196 4644 324 4676
rect 356 4644 484 4676
rect 516 4644 680 4676
rect 0 4640 680 4644
rect 14320 4676 15000 4680
rect 14320 4644 14484 4676
rect 14516 4644 14644 4676
rect 14676 4644 14804 4676
rect 14836 4644 14964 4676
rect 14996 4644 15000 4676
rect 14320 4640 15000 4644
rect 0 4596 520 4600
rect 0 4564 4 4596
rect 36 4564 164 4596
rect 196 4564 324 4596
rect 356 4564 484 4596
rect 516 4564 520 4596
rect 0 4560 520 4564
rect 14320 4596 14760 4600
rect 14320 4564 14724 4596
rect 14756 4564 14760 4596
rect 14320 4560 14760 4564
rect 14800 4596 15000 4600
rect 14800 4564 14804 4596
rect 14836 4564 14964 4596
rect 14996 4564 15000 4596
rect 14800 4560 15000 4564
rect 0 4516 680 4520
rect 0 4484 4 4516
rect 36 4484 164 4516
rect 196 4484 324 4516
rect 356 4484 484 4516
rect 516 4484 680 4516
rect 0 4480 680 4484
rect 14320 4516 15000 4520
rect 14320 4484 14484 4516
rect 14516 4484 14644 4516
rect 14676 4484 14804 4516
rect 14836 4484 14964 4516
rect 14996 4484 15000 4516
rect 14320 4480 15000 4484
rect 0 4436 520 4440
rect 0 4404 4 4436
rect 36 4404 164 4436
rect 196 4404 324 4436
rect 356 4404 484 4436
rect 516 4404 520 4436
rect 0 4400 520 4404
rect 14480 4436 15000 4440
rect 14480 4404 14484 4436
rect 14516 4404 14644 4436
rect 14676 4404 14804 4436
rect 14836 4404 14964 4436
rect 14996 4404 15000 4436
rect 14480 4400 15000 4404
rect 0 4356 520 4360
rect 0 4324 4 4356
rect 36 4324 164 4356
rect 196 4324 324 4356
rect 356 4324 484 4356
rect 516 4324 520 4356
rect 0 4320 520 4324
rect 14480 4356 15000 4360
rect 14480 4324 14484 4356
rect 14516 4324 14644 4356
rect 14676 4324 14804 4356
rect 14836 4324 14964 4356
rect 14996 4324 15000 4356
rect 14480 4320 15000 4324
rect 0 4276 520 4280
rect 0 4244 4 4276
rect 36 4244 164 4276
rect 196 4244 324 4276
rect 356 4244 484 4276
rect 516 4244 520 4276
rect 0 4240 520 4244
rect 14480 4276 15000 4280
rect 14480 4244 14484 4276
rect 14516 4244 14644 4276
rect 14676 4244 14804 4276
rect 14836 4244 14964 4276
rect 14996 4244 15000 4276
rect 14480 4240 15000 4244
rect 0 4196 520 4200
rect 0 4164 4 4196
rect 36 4164 164 4196
rect 196 4164 324 4196
rect 356 4164 484 4196
rect 516 4164 520 4196
rect 0 4160 520 4164
rect 14480 4196 15000 4200
rect 14480 4164 14484 4196
rect 14516 4164 14644 4196
rect 14676 4164 14804 4196
rect 14836 4164 14964 4196
rect 14996 4164 15000 4196
rect 14480 4160 15000 4164
rect 0 4116 520 4120
rect 0 4084 4 4116
rect 36 4084 164 4116
rect 196 4084 324 4116
rect 356 4084 484 4116
rect 516 4084 520 4116
rect 0 4080 520 4084
rect 14480 4116 15000 4120
rect 14480 4084 14484 4116
rect 14516 4084 14644 4116
rect 14676 4084 14804 4116
rect 14836 4084 14964 4116
rect 14996 4084 15000 4116
rect 14480 4080 15000 4084
rect 0 4036 520 4040
rect 0 4004 4 4036
rect 36 4004 164 4036
rect 196 4004 324 4036
rect 356 4004 484 4036
rect 516 4004 520 4036
rect 0 4000 520 4004
rect 14480 4036 15000 4040
rect 14480 4004 14484 4036
rect 14516 4004 14644 4036
rect 14676 4004 14804 4036
rect 14836 4004 14964 4036
rect 14996 4004 15000 4036
rect 14480 4000 15000 4004
rect 0 3956 520 3960
rect 0 3924 4 3956
rect 36 3924 164 3956
rect 196 3924 324 3956
rect 356 3924 484 3956
rect 516 3924 520 3956
rect 0 3920 520 3924
rect 14480 3956 15000 3960
rect 14480 3924 14484 3956
rect 14516 3924 14644 3956
rect 14676 3924 14804 3956
rect 14836 3924 14964 3956
rect 14996 3924 15000 3956
rect 14480 3920 15000 3924
rect 0 3876 520 3880
rect 0 3844 4 3876
rect 36 3844 164 3876
rect 196 3844 324 3876
rect 356 3844 484 3876
rect 516 3844 520 3876
rect 0 3840 520 3844
rect 14480 3876 15000 3880
rect 14480 3844 14484 3876
rect 14516 3844 14644 3876
rect 14676 3844 14804 3876
rect 14836 3844 14964 3876
rect 14996 3844 15000 3876
rect 14480 3840 15000 3844
rect 0 3796 520 3800
rect 0 3764 4 3796
rect 36 3764 164 3796
rect 196 3764 324 3796
rect 356 3764 484 3796
rect 516 3764 520 3796
rect 0 3760 520 3764
rect 14480 3796 15000 3800
rect 14480 3764 14484 3796
rect 14516 3764 14644 3796
rect 14676 3764 14804 3796
rect 14836 3764 14964 3796
rect 14996 3764 15000 3796
rect 14480 3760 15000 3764
rect 0 3716 520 3720
rect 0 3684 4 3716
rect 36 3684 164 3716
rect 196 3684 324 3716
rect 356 3684 484 3716
rect 516 3684 520 3716
rect 0 3680 520 3684
rect 14480 3716 15000 3720
rect 14480 3684 14484 3716
rect 14516 3684 14644 3716
rect 14676 3684 14804 3716
rect 14836 3684 14964 3716
rect 14996 3684 15000 3716
rect 14480 3680 15000 3684
rect 0 3636 520 3640
rect 0 3604 4 3636
rect 36 3604 164 3636
rect 196 3604 324 3636
rect 356 3604 484 3636
rect 516 3604 520 3636
rect 0 3600 520 3604
rect 14480 3636 15000 3640
rect 14480 3604 14484 3636
rect 14516 3604 14644 3636
rect 14676 3604 14804 3636
rect 14836 3604 14964 3636
rect 14996 3604 15000 3636
rect 14480 3600 15000 3604
rect 0 3556 520 3560
rect 0 3524 4 3556
rect 36 3524 164 3556
rect 196 3524 324 3556
rect 356 3524 484 3556
rect 516 3524 520 3556
rect 0 3520 520 3524
rect 14480 3556 15000 3560
rect 14480 3524 14484 3556
rect 14516 3524 14644 3556
rect 14676 3524 14804 3556
rect 14836 3524 14964 3556
rect 14996 3524 15000 3556
rect 14480 3520 15000 3524
rect 0 3476 520 3480
rect 0 3444 4 3476
rect 36 3444 164 3476
rect 196 3444 324 3476
rect 356 3444 484 3476
rect 516 3444 520 3476
rect 0 3440 520 3444
rect 14480 3476 15000 3480
rect 14480 3444 14484 3476
rect 14516 3444 14644 3476
rect 14676 3444 14804 3476
rect 14836 3444 14964 3476
rect 14996 3444 15000 3476
rect 14480 3440 15000 3444
rect 0 3396 520 3400
rect 0 3364 4 3396
rect 36 3364 164 3396
rect 196 3364 324 3396
rect 356 3364 484 3396
rect 516 3364 520 3396
rect 0 3360 520 3364
rect 14480 3396 15000 3400
rect 14480 3364 14484 3396
rect 14516 3364 14644 3396
rect 14676 3364 14804 3396
rect 14836 3364 14964 3396
rect 14996 3364 15000 3396
rect 14480 3360 15000 3364
rect 0 3316 520 3320
rect 0 3284 4 3316
rect 36 3284 164 3316
rect 196 3284 324 3316
rect 356 3284 484 3316
rect 516 3284 520 3316
rect 0 3280 520 3284
rect 14320 3316 14600 3320
rect 14320 3284 14564 3316
rect 14596 3284 14600 3316
rect 14320 3280 14600 3284
rect 14640 3316 15000 3320
rect 14640 3284 14644 3316
rect 14676 3284 14804 3316
rect 14836 3284 14964 3316
rect 14996 3284 15000 3316
rect 14640 3280 15000 3284
rect 0 3236 520 3240
rect 0 3204 4 3236
rect 36 3204 164 3236
rect 196 3204 324 3236
rect 356 3204 484 3236
rect 516 3204 520 3236
rect 0 3200 520 3204
rect 14480 3236 15000 3240
rect 14480 3204 14484 3236
rect 14516 3204 14644 3236
rect 14676 3204 14804 3236
rect 14836 3204 14964 3236
rect 14996 3204 15000 3236
rect 14480 3200 15000 3204
rect 0 3156 520 3160
rect 0 3124 4 3156
rect 36 3124 164 3156
rect 196 3124 324 3156
rect 356 3124 484 3156
rect 516 3124 520 3156
rect 0 3120 520 3124
rect 14480 3156 15000 3160
rect 14480 3124 14484 3156
rect 14516 3124 14644 3156
rect 14676 3124 14804 3156
rect 14836 3124 14964 3156
rect 14996 3124 15000 3156
rect 14480 3120 15000 3124
rect 0 3076 520 3080
rect 0 3044 4 3076
rect 36 3044 164 3076
rect 196 3044 324 3076
rect 356 3044 484 3076
rect 516 3044 520 3076
rect 0 3040 520 3044
rect 14480 3076 15000 3080
rect 14480 3044 14484 3076
rect 14516 3044 14644 3076
rect 14676 3044 14804 3076
rect 14836 3044 14964 3076
rect 14996 3044 15000 3076
rect 14480 3040 15000 3044
rect 0 2996 520 3000
rect 0 2964 4 2996
rect 36 2964 164 2996
rect 196 2964 324 2996
rect 356 2964 484 2996
rect 516 2964 520 2996
rect 0 2960 520 2964
rect 14480 2996 15000 3000
rect 14480 2964 14484 2996
rect 14516 2964 14644 2996
rect 14676 2964 14804 2996
rect 14836 2964 14964 2996
rect 14996 2964 15000 2996
rect 14480 2960 15000 2964
rect 0 2916 520 2920
rect 0 2884 4 2916
rect 36 2884 164 2916
rect 196 2884 324 2916
rect 356 2884 484 2916
rect 516 2884 520 2916
rect 0 2880 520 2884
rect 14480 2916 15000 2920
rect 14480 2884 14484 2916
rect 14516 2884 14644 2916
rect 14676 2884 14804 2916
rect 14836 2884 14964 2916
rect 14996 2884 15000 2916
rect 14480 2880 15000 2884
rect 0 2836 520 2840
rect 0 2804 4 2836
rect 36 2804 164 2836
rect 196 2804 324 2836
rect 356 2804 484 2836
rect 516 2804 520 2836
rect 0 2800 520 2804
rect 14480 2836 15000 2840
rect 14480 2804 14484 2836
rect 14516 2804 14644 2836
rect 14676 2804 14804 2836
rect 14836 2804 14964 2836
rect 14996 2804 15000 2836
rect 14480 2800 15000 2804
rect 0 2756 520 2760
rect 0 2724 4 2756
rect 36 2724 164 2756
rect 196 2724 324 2756
rect 356 2724 484 2756
rect 516 2724 520 2756
rect 0 2720 520 2724
rect 14480 2756 15000 2760
rect 14480 2724 14484 2756
rect 14516 2724 14644 2756
rect 14676 2724 14804 2756
rect 14836 2724 14964 2756
rect 14996 2724 15000 2756
rect 14480 2720 15000 2724
rect 0 2676 520 2680
rect 0 2644 4 2676
rect 36 2644 164 2676
rect 196 2644 324 2676
rect 356 2644 484 2676
rect 516 2644 520 2676
rect 0 2640 520 2644
rect 14480 2676 15000 2680
rect 14480 2644 14484 2676
rect 14516 2644 14644 2676
rect 14676 2644 14804 2676
rect 14836 2644 14964 2676
rect 14996 2644 15000 2676
rect 14480 2640 15000 2644
rect 0 2596 520 2600
rect 0 2564 4 2596
rect 36 2564 164 2596
rect 196 2564 324 2596
rect 356 2564 484 2596
rect 516 2564 520 2596
rect 0 2560 520 2564
rect 14480 2596 15000 2600
rect 14480 2564 14484 2596
rect 14516 2564 14644 2596
rect 14676 2564 14804 2596
rect 14836 2564 14964 2596
rect 14996 2564 15000 2596
rect 14480 2560 15000 2564
rect 0 2516 520 2520
rect 0 2484 4 2516
rect 36 2484 164 2516
rect 196 2484 324 2516
rect 356 2484 484 2516
rect 516 2484 520 2516
rect 0 2480 520 2484
rect 14480 2516 15000 2520
rect 14480 2484 14484 2516
rect 14516 2484 14644 2516
rect 14676 2484 14804 2516
rect 14836 2484 14964 2516
rect 14996 2484 15000 2516
rect 14480 2480 15000 2484
rect 0 2436 520 2440
rect 0 2404 4 2436
rect 36 2404 164 2436
rect 196 2404 324 2436
rect 356 2404 484 2436
rect 516 2404 520 2436
rect 0 2400 520 2404
rect 14480 2436 15000 2440
rect 14480 2404 14484 2436
rect 14516 2404 14644 2436
rect 14676 2404 14804 2436
rect 14836 2404 14964 2436
rect 14996 2404 15000 2436
rect 14480 2400 15000 2404
rect 0 2356 520 2360
rect 0 2324 4 2356
rect 36 2324 164 2356
rect 196 2324 324 2356
rect 356 2324 484 2356
rect 516 2324 520 2356
rect 0 2320 520 2324
rect 14480 2356 15000 2360
rect 14480 2324 14484 2356
rect 14516 2324 14644 2356
rect 14676 2324 14804 2356
rect 14836 2324 14964 2356
rect 14996 2324 15000 2356
rect 14480 2320 15000 2324
rect 0 2276 520 2280
rect 0 2244 4 2276
rect 36 2244 164 2276
rect 196 2244 324 2276
rect 356 2244 484 2276
rect 516 2244 520 2276
rect 0 2240 520 2244
rect 14480 2276 15000 2280
rect 14480 2244 14484 2276
rect 14516 2244 14644 2276
rect 14676 2244 14804 2276
rect 14836 2244 14964 2276
rect 14996 2244 15000 2276
rect 14480 2240 15000 2244
rect 0 2196 520 2200
rect 0 2164 4 2196
rect 36 2164 164 2196
rect 196 2164 324 2196
rect 356 2164 484 2196
rect 516 2164 520 2196
rect 0 2160 520 2164
rect 14480 2196 15000 2200
rect 14480 2164 14484 2196
rect 14516 2164 14644 2196
rect 14676 2164 14804 2196
rect 14836 2164 14964 2196
rect 14996 2164 15000 2196
rect 14480 2160 15000 2164
rect 0 2116 680 2120
rect 0 2084 4 2116
rect 36 2084 164 2116
rect 196 2084 324 2116
rect 356 2084 484 2116
rect 516 2084 680 2116
rect 0 2080 680 2084
rect 14360 2116 15000 2120
rect 14360 2084 14484 2116
rect 14516 2084 14644 2116
rect 14676 2084 14804 2116
rect 14836 2084 14964 2116
rect 14996 2084 15000 2116
rect 14360 2080 15000 2084
rect 0 2036 520 2040
rect 0 2004 4 2036
rect 36 2004 164 2036
rect 196 2004 324 2036
rect 356 2004 484 2036
rect 516 2004 520 2036
rect 0 2000 520 2004
rect 14320 2036 14760 2040
rect 14320 2004 14724 2036
rect 14756 2004 14760 2036
rect 14320 2000 14760 2004
rect 14800 2036 15000 2040
rect 14800 2004 14804 2036
rect 14836 2004 14964 2036
rect 14996 2004 15000 2036
rect 14800 2000 15000 2004
rect 0 1956 680 1960
rect 0 1924 4 1956
rect 36 1924 164 1956
rect 196 1924 324 1956
rect 356 1924 484 1956
rect 516 1924 680 1956
rect 0 1920 680 1924
rect 14320 1956 15000 1960
rect 14320 1924 14484 1956
rect 14516 1924 14644 1956
rect 14676 1924 14804 1956
rect 14836 1924 14964 1956
rect 14996 1924 15000 1956
rect 14320 1920 15000 1924
rect 0 1876 520 1880
rect 0 1844 4 1876
rect 36 1844 164 1876
rect 196 1844 324 1876
rect 356 1844 484 1876
rect 516 1844 520 1876
rect 0 1840 520 1844
rect 14320 1876 15000 1880
rect 14320 1844 14884 1876
rect 14916 1844 15000 1876
rect 14320 1840 15000 1844
rect 0 1796 680 1800
rect 0 1764 4 1796
rect 36 1764 164 1796
rect 196 1764 324 1796
rect 356 1764 484 1796
rect 516 1764 680 1796
rect 0 1760 680 1764
rect 14320 1796 15000 1800
rect 14320 1764 14484 1796
rect 14516 1764 14644 1796
rect 14676 1764 14804 1796
rect 14836 1764 14964 1796
rect 14996 1764 15000 1796
rect 14320 1760 15000 1764
rect 0 1716 520 1720
rect 0 1684 4 1716
rect 36 1684 164 1716
rect 196 1684 324 1716
rect 356 1684 484 1716
rect 516 1684 520 1716
rect 0 1680 520 1684
rect 14480 1716 15000 1720
rect 14480 1684 14484 1716
rect 14516 1684 14644 1716
rect 14676 1684 14804 1716
rect 14836 1684 14964 1716
rect 14996 1684 15000 1716
rect 14480 1680 15000 1684
rect 0 1636 520 1640
rect 0 1604 4 1636
rect 36 1604 164 1636
rect 196 1604 324 1636
rect 356 1604 484 1636
rect 516 1604 520 1636
rect 0 1600 520 1604
rect 14480 1636 15000 1640
rect 14480 1604 14484 1636
rect 14516 1604 14644 1636
rect 14676 1604 14804 1636
rect 14836 1604 14964 1636
rect 14996 1604 15000 1636
rect 14480 1600 15000 1604
rect 0 1556 680 1560
rect 0 1524 4 1556
rect 36 1524 164 1556
rect 196 1524 324 1556
rect 356 1524 484 1556
rect 516 1524 680 1556
rect 0 1520 680 1524
rect 14320 1556 15000 1560
rect 14320 1524 14484 1556
rect 14516 1524 14644 1556
rect 14676 1524 14804 1556
rect 14836 1524 14964 1556
rect 14996 1524 15000 1556
rect 14320 1520 15000 1524
rect 0 1476 680 1480
rect 0 1444 4 1476
rect 36 1444 164 1476
rect 196 1444 324 1476
rect 356 1444 484 1476
rect 516 1444 680 1476
rect 0 1440 680 1444
rect 14320 1476 15000 1480
rect 14320 1444 14484 1476
rect 14516 1444 14644 1476
rect 14676 1444 14804 1476
rect 14836 1444 14964 1476
rect 14996 1444 15000 1476
rect 14320 1440 15000 1444
rect 0 1396 680 1400
rect 0 1364 4 1396
rect 36 1364 164 1396
rect 196 1364 324 1396
rect 356 1364 484 1396
rect 516 1364 680 1396
rect 0 1360 680 1364
rect 14320 1396 15000 1400
rect 14320 1364 14484 1396
rect 14516 1364 14644 1396
rect 14676 1364 14804 1396
rect 14836 1364 14964 1396
rect 14996 1364 15000 1396
rect 14320 1360 15000 1364
rect 0 1316 680 1320
rect 0 1284 4 1316
rect 36 1284 164 1316
rect 196 1284 324 1316
rect 356 1284 484 1316
rect 516 1284 680 1316
rect 0 1280 680 1284
rect 14320 1316 15000 1320
rect 14320 1284 14484 1316
rect 14516 1284 14644 1316
rect 14676 1284 14804 1316
rect 14836 1284 14964 1316
rect 14996 1284 15000 1316
rect 14320 1280 15000 1284
rect 0 1236 680 1240
rect 0 1204 4 1236
rect 36 1204 164 1236
rect 196 1204 324 1236
rect 356 1204 484 1236
rect 516 1204 680 1236
rect 0 1200 680 1204
rect 14320 1236 15000 1240
rect 14320 1204 14484 1236
rect 14516 1204 14644 1236
rect 14676 1204 14804 1236
rect 14836 1204 14964 1236
rect 14996 1204 15000 1236
rect 14320 1200 15000 1204
rect 0 1156 520 1160
rect 0 1124 4 1156
rect 36 1124 164 1156
rect 196 1124 324 1156
rect 356 1124 484 1156
rect 516 1124 520 1156
rect 0 1120 520 1124
rect 14480 1156 15000 1160
rect 14480 1124 14484 1156
rect 14516 1124 14644 1156
rect 14676 1124 14804 1156
rect 14836 1124 14964 1156
rect 14996 1124 15000 1156
rect 14480 1120 15000 1124
rect 0 1076 520 1080
rect 0 1044 4 1076
rect 36 1044 164 1076
rect 196 1044 324 1076
rect 356 1044 484 1076
rect 516 1044 520 1076
rect 0 1040 520 1044
rect 14480 1076 15000 1080
rect 14480 1044 14484 1076
rect 14516 1044 14644 1076
rect 14676 1044 14804 1076
rect 14836 1044 14964 1076
rect 14996 1044 15000 1076
rect 14480 1040 15000 1044
rect 0 996 520 1000
rect 0 964 4 996
rect 36 964 164 996
rect 196 964 324 996
rect 356 964 484 996
rect 516 964 520 996
rect 0 960 520 964
rect 14480 996 15000 1000
rect 14480 964 14484 996
rect 14516 964 14644 996
rect 14676 964 14804 996
rect 14836 964 14964 996
rect 14996 964 15000 996
rect 14480 960 15000 964
rect 0 916 680 920
rect 0 884 4 916
rect 36 884 164 916
rect 196 884 324 916
rect 356 884 484 916
rect 516 884 680 916
rect 0 880 680 884
rect 14320 916 15000 920
rect 14320 884 14484 916
rect 14516 884 14644 916
rect 14676 884 14804 916
rect 14836 884 14964 916
rect 14996 884 15000 916
rect 14320 880 15000 884
rect 0 836 680 840
rect 0 804 4 836
rect 36 804 164 836
rect 196 804 324 836
rect 356 804 484 836
rect 516 804 680 836
rect 0 800 680 804
rect 14320 836 15000 840
rect 14320 804 14484 836
rect 14516 804 14644 836
rect 14676 804 14804 836
rect 14836 804 14964 836
rect 14996 804 15000 836
rect 14320 800 15000 804
rect 0 756 680 760
rect 0 724 4 756
rect 36 724 164 756
rect 196 724 324 756
rect 356 724 484 756
rect 516 724 680 756
rect 0 720 680 724
rect 14320 756 15000 760
rect 14320 724 14484 756
rect 14516 724 14644 756
rect 14676 724 14804 756
rect 14836 724 14964 756
rect 14996 724 15000 756
rect 14320 720 15000 724
rect 0 676 680 680
rect 0 644 4 676
rect 36 644 164 676
rect 196 644 324 676
rect 356 644 484 676
rect 516 644 680 676
rect 0 640 680 644
rect 14320 676 15000 680
rect 14320 644 14484 676
rect 14516 644 14644 676
rect 14676 644 14804 676
rect 14836 644 14964 676
rect 14996 644 15000 676
rect 14320 640 15000 644
rect 0 596 680 600
rect 0 564 4 596
rect 36 564 164 596
rect 196 564 324 596
rect 356 564 484 596
rect 516 564 680 596
rect 0 560 680 564
rect 14320 596 15000 600
rect 14320 564 14484 596
rect 14516 564 14644 596
rect 14676 564 14804 596
rect 14836 564 14964 596
rect 14996 564 15000 596
rect 14320 560 15000 564
rect 0 516 520 520
rect 0 484 4 516
rect 36 484 164 516
rect 196 484 324 516
rect 356 484 484 516
rect 516 484 520 516
rect 0 480 520 484
rect 14480 516 15000 520
rect 14480 484 14484 516
rect 14516 484 14644 516
rect 14676 484 14804 516
rect 14836 484 14964 516
rect 14996 484 15000 516
rect 14480 480 15000 484
rect 0 436 15000 440
rect 0 244 4 436
rect 36 244 164 436
rect 196 244 324 436
rect 356 244 484 436
rect 516 244 14484 436
rect 14516 244 14644 436
rect 14676 244 14804 436
rect 14836 244 14964 436
rect 14996 244 15000 436
rect 0 240 15000 244
rect 0 196 15000 200
rect 0 4 564 196
rect 596 4 14404 196
rect 14436 4 15000 196
rect 0 0 15000 4
use cap1_10_core  p2
timestamp 1638207275
transform 1 0 7000 0 1 1000
box -6440 680 7440 3920
use cap1_10_core  m2
timestamp 1638207275
transform 1 0 7000 0 1 4280
box -6440 680 7440 3920
use cap1_10_core  m1
timestamp 1638207275
transform 1 0 7000 0 1 7560
box -6440 680 7440 3920
use cap1_10_core  p1
timestamp 1638207275
transform 1 0 7000 0 1 10840
box -6440 680 7440 3920
use cap1_10_dummy  dummy2
timestamp 1637451829
transform 1 0 7000 0 1 -200
box -6440 680 7440 1840
use cap1_10_dummy  dummy1
timestamp 1637451829
transform 1 0 7000 0 1 14120
box -6440 680 7440 1840
<< labels >>
rlabel metal3 14880 15920 14920 15960 0 ip
port 0 nsew
rlabel metal3 14560 15920 14600 15960 0 xp
port 1 nsew
rlabel metal3 14720 15920 14760 15960 0 om
port 2 nsew
rlabel metal3 80 15920 120 15960 0 im
port 3 nsew
rlabel metal3 400 15920 440 15960 0 xm
port 4 nsew
rlabel metal3 240 15920 280 15960 0 op
port 5 nsew
rlabel metal4 0 240 40 440 0 gnda
port 6 nsew
rlabel metal4 0 0 40 200 0 vssa
port 7 nsew
<< end >>
