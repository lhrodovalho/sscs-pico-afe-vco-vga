* OpAmp open-loop dc testbench

* Include SkyWater sky130 device models
.lib "/usr/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice" tt
.param mc_mm_switch=0
.include "../mag/opamp_core.spice"

* supply voltages
vdda  vdda 0 1.0
vssa  vssa 0 0.0

* input signals
vin in gnda 0
eip ip gnda in gnda  0.5
eim im gnda in gnda -0.5
egnda gnda vssa ib vssa 1

* DUT
x0 im ip out ib q vdda bp vddx gnda vssa xn xp x y z opamp_core
ib vdda ib 2n

.option gmin=1e-14
.control

	op
	print gpa gpb gnb gna i(vdda)

	dc vin -1m 1m 10u
	plot in out
	plot abs(deriv(out)) ylog

.endc

.end
