magic
tech sky130A
timestamp 1638390070
<< nwell >>
rect 60 1980 4140 2940
rect 60 860 4140 1820
<< nmos >>
rect 260 280 1060 380
rect 1220 280 2020 380
rect 2180 280 2980 380
rect 3140 280 3940 380
rect 260 80 1060 180
rect 1220 80 2020 180
rect 2180 80 2980 180
rect 3140 80 3940 180
<< pmoslvt >>
rect 260 2540 1060 2840
rect 1220 2540 2020 2840
rect 2180 2540 2980 2840
rect 3140 2540 3940 2840
rect 260 2160 1060 2460
rect 1220 2160 2020 2460
rect 2180 2160 2980 2460
rect 3140 2160 3940 2460
rect 260 1420 1060 1720
rect 1220 1420 2020 1720
rect 2180 1420 2980 1720
rect 3140 1420 3940 1720
rect 260 1040 1060 1340
rect 1220 1040 2020 1340
rect 2180 1040 2980 1340
rect 3140 1040 3940 1340
<< ndiff >>
rect 160 370 260 380
rect 160 290 165 370
rect 195 290 260 370
rect 160 280 260 290
rect 1060 370 1220 380
rect 1060 290 1125 370
rect 1155 290 1220 370
rect 1060 280 1220 290
rect 2020 370 2180 380
rect 2020 290 2085 370
rect 2115 290 2180 370
rect 2020 280 2180 290
rect 2980 370 3140 380
rect 2980 290 3045 370
rect 3075 290 3140 370
rect 2980 280 3140 290
rect 3940 370 4040 380
rect 3940 290 4005 370
rect 4035 290 4040 370
rect 3940 280 4040 290
rect 160 170 260 180
rect 160 90 165 170
rect 195 90 260 170
rect 160 80 260 90
rect 1060 170 1220 180
rect 1060 90 1125 170
rect 1155 90 1220 170
rect 1060 80 1220 90
rect 2020 170 2180 180
rect 2020 90 2085 170
rect 2115 90 2180 170
rect 2020 80 2180 90
rect 2980 170 3140 180
rect 2980 90 3045 170
rect 3075 90 3140 170
rect 2980 80 3140 90
rect 3940 170 4040 180
rect 3940 90 4005 170
rect 4035 90 4040 170
rect 3940 80 4040 90
<< pdiff >>
rect 160 2830 260 2840
rect 160 2550 165 2830
rect 195 2550 260 2830
rect 160 2540 260 2550
rect 1060 2830 1220 2840
rect 1060 2550 1125 2830
rect 1155 2550 1220 2830
rect 1060 2540 1220 2550
rect 2020 2830 2180 2840
rect 2020 2550 2085 2830
rect 2115 2550 2180 2830
rect 2020 2540 2180 2550
rect 2980 2830 3140 2840
rect 2980 2550 3045 2830
rect 3075 2550 3140 2830
rect 2980 2540 3140 2550
rect 3940 2830 4040 2840
rect 3940 2550 4005 2830
rect 4035 2550 4040 2830
rect 3940 2540 4040 2550
rect 160 2450 260 2460
rect 160 2170 165 2450
rect 195 2170 260 2450
rect 160 2160 260 2170
rect 1060 2450 1220 2460
rect 1060 2170 1125 2450
rect 1155 2170 1220 2450
rect 1060 2160 1220 2170
rect 2020 2450 2180 2460
rect 2020 2170 2085 2450
rect 2115 2170 2180 2450
rect 2020 2160 2180 2170
rect 2980 2450 3140 2460
rect 2980 2170 3045 2450
rect 3075 2170 3140 2450
rect 2980 2160 3140 2170
rect 3940 2450 4040 2460
rect 3940 2170 4005 2450
rect 4035 2170 4040 2450
rect 3940 2160 4040 2170
rect 160 1710 260 1720
rect 160 1430 165 1710
rect 195 1430 260 1710
rect 160 1420 260 1430
rect 1060 1710 1220 1720
rect 1060 1430 1125 1710
rect 1155 1430 1220 1710
rect 1060 1420 1220 1430
rect 2020 1710 2180 1720
rect 2020 1430 2085 1710
rect 2115 1430 2180 1710
rect 2020 1420 2180 1430
rect 2980 1710 3140 1720
rect 2980 1430 3045 1710
rect 3075 1430 3140 1710
rect 2980 1420 3140 1430
rect 3940 1710 4040 1720
rect 3940 1430 4005 1710
rect 4035 1430 4040 1710
rect 3940 1420 4040 1430
rect 160 1330 260 1340
rect 160 1050 165 1330
rect 195 1050 260 1330
rect 160 1040 260 1050
rect 1060 1330 1220 1340
rect 1060 1050 1125 1330
rect 1155 1050 1220 1330
rect 1060 1040 1220 1050
rect 2020 1330 2180 1340
rect 2020 1050 2085 1330
rect 2115 1050 2180 1330
rect 2020 1040 2180 1050
rect 2980 1330 3140 1340
rect 2980 1050 3045 1330
rect 3075 1050 3140 1330
rect 2980 1040 3140 1050
rect 3940 1330 4040 1340
rect 3940 1050 4005 1330
rect 4035 1050 4040 1330
rect 3940 1040 4040 1050
<< ndiffc >>
rect 165 290 195 370
rect 1125 290 1155 370
rect 2085 290 2115 370
rect 3045 290 3075 370
rect 4005 290 4035 370
rect 165 90 195 170
rect 1125 90 1155 170
rect 2085 90 2115 170
rect 3045 90 3075 170
rect 4005 90 4035 170
<< pdiffc >>
rect 165 2550 195 2830
rect 1125 2550 1155 2830
rect 2085 2550 2115 2830
rect 3045 2550 3075 2830
rect 4005 2550 4035 2830
rect 165 2170 195 2450
rect 1125 2170 1155 2450
rect 2085 2170 2115 2450
rect 3045 2170 3075 2450
rect 4005 2170 4035 2450
rect 165 1430 195 1710
rect 1125 1430 1155 1710
rect 2085 1430 2115 1710
rect 3045 1430 3075 1710
rect 4005 1430 4035 1710
rect 165 1050 195 1330
rect 1125 1050 1155 1330
rect 2085 1050 2115 1330
rect 3045 1050 3075 1330
rect 4005 1050 4035 1330
<< psubdiff >>
rect 0 2960 60 3000
rect 4140 2960 4200 3000
rect 0 2940 40 2960
rect 4160 2940 4200 2960
rect 0 1960 40 1980
rect 4160 1960 4200 1980
rect 0 1920 60 1960
rect 4120 1920 4200 1960
rect 0 1840 60 1880
rect 4120 1840 4200 1880
rect 0 1820 40 1840
rect 4160 1820 4200 1840
rect 0 840 40 860
rect 4160 840 4200 860
rect 0 800 60 840
rect 4140 800 4200 840
rect 0 480 60 520
rect 4140 480 4200 520
rect 0 460 40 480
rect 4160 460 4200 480
rect 0 40 40 60
rect 4160 40 4200 60
rect 0 0 60 40
rect 4140 0 4200 40
<< nsubdiff >>
rect 80 2880 140 2920
rect 4060 2880 4120 2920
rect 80 2860 120 2880
rect 4080 2860 4120 2880
rect 80 2040 120 2060
rect 4080 2040 4120 2060
rect 80 2000 140 2040
rect 4060 2000 4120 2040
rect 80 1760 140 1800
rect 4060 1760 4120 1800
rect 80 1740 120 1760
rect 4080 1740 4120 1760
rect 80 920 120 960
rect 4080 920 4120 960
rect 80 880 140 920
rect 4060 880 4120 920
<< psubdiffcont >>
rect 60 2960 4140 3000
rect 0 1980 40 2940
rect 4160 1980 4200 2940
rect 60 1920 4120 1960
rect 60 1840 4120 1880
rect 0 860 40 1820
rect 4160 860 4200 1820
rect 60 800 4140 840
rect 60 480 4140 520
rect 0 60 40 460
rect 4160 60 4200 460
rect 60 0 4140 40
<< nsubdiffcont >>
rect 140 2880 4060 2920
rect 80 2060 120 2860
rect 4080 2060 4120 2860
rect 140 2000 4060 2040
rect 140 1760 4060 1800
rect 80 960 120 1740
rect 4080 960 4120 1740
rect 140 880 4060 920
<< poly >>
rect 260 2840 1060 2860
rect 1220 2840 2020 2860
rect 2180 2840 2980 2860
rect 3140 2840 3940 2860
rect 260 2460 1060 2540
rect 1220 2460 2020 2540
rect 2180 2460 2980 2540
rect 3140 2460 3940 2540
rect 260 2115 1060 2160
rect 260 2085 270 2115
rect 1050 2085 1060 2115
rect 260 2080 1060 2085
rect 1220 2115 2020 2160
rect 1220 2085 1230 2115
rect 2010 2085 2020 2115
rect 1220 2080 2020 2085
rect 2180 2115 2980 2160
rect 2180 2085 2190 2115
rect 2970 2085 2980 2115
rect 2180 2080 2980 2085
rect 3140 2115 3940 2160
rect 3140 2085 3150 2115
rect 3930 2085 3940 2115
rect 3140 2080 3940 2085
rect 260 1720 1060 1740
rect 1220 1720 2020 1740
rect 2180 1720 2980 1740
rect 3140 1720 3940 1740
rect 260 1340 1060 1420
rect 1220 1340 2020 1420
rect 2180 1340 2980 1420
rect 3140 1340 3940 1420
rect 260 995 1060 1040
rect 260 965 270 995
rect 1050 965 1060 995
rect 260 960 1060 965
rect 1220 995 2020 1040
rect 1220 965 1230 995
rect 2010 965 2020 995
rect 1220 960 2020 965
rect 2180 995 2980 1040
rect 2180 965 2190 995
rect 2970 965 2980 995
rect 2180 960 2980 965
rect 3140 995 3940 1040
rect 3140 965 3150 995
rect 3930 965 3940 995
rect 3140 960 3940 965
rect 260 435 1060 440
rect 260 405 270 435
rect 1050 405 1060 435
rect 260 380 1060 405
rect 1220 435 2020 440
rect 1220 405 1230 435
rect 2010 405 2020 435
rect 1220 380 2020 405
rect 2180 435 2980 440
rect 2180 405 2190 435
rect 2970 405 2980 435
rect 2180 380 2980 405
rect 3140 435 3940 440
rect 3140 405 3150 435
rect 3930 405 3940 435
rect 3140 380 3940 405
rect 260 180 1060 280
rect 1220 180 2020 280
rect 2180 180 2980 280
rect 3140 180 3940 280
rect 260 60 1060 80
rect 1220 60 2020 80
rect 2180 60 2980 80
rect 3140 60 3940 80
<< polycont >>
rect 270 2085 1050 2115
rect 1230 2085 2010 2115
rect 2190 2085 2970 2115
rect 3150 2085 3930 2115
rect 270 965 1050 995
rect 1230 965 2010 995
rect 2190 965 2970 995
rect 3150 965 3930 995
rect 270 405 1050 435
rect 1230 405 2010 435
rect 2190 405 2970 435
rect 3150 405 3930 435
<< locali >>
rect 0 2960 60 3000
rect 4140 2960 4200 3000
rect 0 2940 40 2960
rect 4160 2940 4200 2960
rect 80 2880 140 2920
rect 4060 2880 4120 2920
rect 80 2860 120 2880
rect 160 2830 200 2840
rect 160 2550 165 2830
rect 195 2550 200 2830
rect 160 2540 200 2550
rect 1120 2830 1160 2840
rect 1120 2550 1125 2830
rect 1155 2550 1160 2830
rect 1120 2540 1160 2550
rect 2080 2830 2120 2880
rect 4080 2860 4120 2880
rect 2080 2550 2085 2830
rect 2115 2550 2120 2830
rect 2080 2520 2120 2550
rect 3040 2830 3080 2840
rect 3040 2550 3045 2830
rect 3075 2550 3080 2830
rect 3040 2540 3080 2550
rect 4000 2830 4040 2840
rect 4000 2550 4005 2830
rect 4035 2550 4040 2830
rect 4000 2540 4040 2550
rect 1120 2480 3080 2520
rect 160 2450 200 2460
rect 160 2170 165 2450
rect 195 2170 200 2450
rect 160 2160 200 2170
rect 1120 2450 1160 2480
rect 1120 2170 1125 2450
rect 1155 2170 1160 2450
rect 1120 2160 1160 2170
rect 2080 2450 2120 2460
rect 2080 2170 2085 2450
rect 2115 2170 2120 2450
rect 2080 2160 2120 2170
rect 3040 2450 3080 2480
rect 3040 2170 3045 2450
rect 3075 2170 3080 2450
rect 3040 2160 3080 2170
rect 4000 2450 4040 2460
rect 4000 2170 4005 2450
rect 4035 2170 4040 2450
rect 4000 2160 4040 2170
rect 260 2115 1060 2120
rect 260 2085 270 2115
rect 1050 2085 1060 2115
rect 260 2080 1060 2085
rect 1220 2115 2020 2120
rect 1220 2085 1230 2115
rect 2010 2085 2020 2115
rect 1220 2080 2020 2085
rect 2180 2115 2980 2120
rect 2180 2085 2190 2115
rect 2970 2085 2980 2115
rect 2180 2080 2980 2085
rect 3140 2115 3940 2120
rect 3140 2085 3150 2115
rect 3930 2085 3940 2115
rect 3140 2080 3940 2085
rect 80 2040 120 2060
rect 4080 2040 4120 2060
rect 80 2000 140 2040
rect 4060 2000 4120 2040
rect 0 1960 40 1980
rect 4160 1960 4200 1980
rect 0 1920 60 1960
rect 4120 1920 4200 1960
rect 0 1880 40 1920
rect 4160 1880 4200 1920
rect 0 1840 60 1880
rect 4120 1840 4200 1880
rect 0 1820 40 1840
rect 4160 1820 4200 1840
rect 80 1760 140 1800
rect 4060 1760 4120 1800
rect 80 1740 120 1760
rect 160 1710 200 1760
rect 160 1430 165 1710
rect 195 1430 200 1710
rect 160 1420 200 1430
rect 1120 1710 1160 1720
rect 1120 1430 1125 1710
rect 1155 1430 1160 1710
rect 1120 1420 1160 1430
rect 2080 1710 2120 1720
rect 2080 1430 2085 1710
rect 2115 1430 2120 1710
rect 2080 1400 2120 1430
rect 3040 1710 3080 1720
rect 3040 1430 3045 1710
rect 3075 1430 3080 1710
rect 3040 1420 3080 1430
rect 4000 1710 4040 1760
rect 4000 1430 4005 1710
rect 4035 1430 4040 1710
rect 4000 1420 4040 1430
rect 4080 1740 4120 1760
rect 1120 1360 3080 1400
rect 160 1330 200 1340
rect 160 1050 165 1330
rect 195 1050 200 1330
rect 160 1040 200 1050
rect 1120 1330 1160 1360
rect 1120 1050 1125 1330
rect 1155 1050 1160 1330
rect 1120 1040 1160 1050
rect 2080 1330 2120 1340
rect 2080 1050 2085 1330
rect 2115 1050 2120 1330
rect 2080 1040 2120 1050
rect 3040 1330 3080 1360
rect 3040 1050 3045 1330
rect 3075 1050 3080 1330
rect 3040 1040 3080 1050
rect 4000 1330 4040 1340
rect 4000 1050 4005 1330
rect 4035 1050 4040 1330
rect 4000 1040 4040 1050
rect 260 995 1060 1000
rect 260 965 270 995
rect 1050 965 1060 995
rect 260 960 1060 965
rect 1220 995 2020 1000
rect 1220 965 1230 995
rect 2010 965 2020 995
rect 1220 960 2020 965
rect 2180 995 2980 1000
rect 2180 965 2190 995
rect 2970 965 2980 995
rect 2180 960 2980 965
rect 3140 995 3940 1000
rect 3140 965 3150 995
rect 3930 965 3940 995
rect 3140 960 3940 965
rect 80 920 120 960
rect 4080 920 4120 960
rect 80 880 140 920
rect 4060 880 4120 920
rect 0 840 40 860
rect 4160 840 4200 860
rect 0 800 60 840
rect 4140 800 4200 840
rect 0 520 40 800
rect 80 670 120 760
rect 80 650 90 670
rect 110 650 120 670
rect 80 560 120 650
rect 240 670 280 760
rect 240 650 250 670
rect 270 650 280 670
rect 240 560 280 650
rect 320 670 360 760
rect 320 650 330 670
rect 350 650 360 670
rect 320 560 360 650
rect 400 670 440 760
rect 400 650 410 670
rect 430 650 440 670
rect 400 560 440 650
rect 480 670 520 760
rect 480 650 490 670
rect 510 650 520 670
rect 480 560 520 650
rect 560 670 600 760
rect 560 650 570 670
rect 590 650 600 670
rect 560 560 600 650
rect 720 670 760 760
rect 720 650 730 670
rect 750 650 760 670
rect 720 560 760 650
rect 800 670 840 760
rect 800 650 810 670
rect 830 650 840 670
rect 800 560 840 650
rect 880 670 920 760
rect 880 650 890 670
rect 910 650 920 670
rect 880 560 920 650
rect 960 670 1000 760
rect 960 650 970 670
rect 990 650 1000 670
rect 960 560 1000 650
rect 1040 670 1080 760
rect 1040 650 1050 670
rect 1070 650 1080 670
rect 1040 560 1080 650
rect 1120 670 1160 760
rect 1120 650 1130 670
rect 1150 650 1160 670
rect 1120 560 1160 650
rect 1200 670 1240 760
rect 1200 650 1210 670
rect 1230 650 1240 670
rect 1200 560 1240 650
rect 1280 670 1320 760
rect 1280 650 1290 670
rect 1310 650 1320 670
rect 1280 560 1320 650
rect 1360 670 1400 760
rect 1360 650 1370 670
rect 1390 650 1400 670
rect 1360 560 1400 650
rect 1440 670 1480 760
rect 1440 650 1450 670
rect 1470 650 1480 670
rect 1440 560 1480 650
rect 1520 670 1560 760
rect 1520 650 1530 670
rect 1550 650 1560 670
rect 1520 560 1560 650
rect 1680 670 1720 760
rect 1680 650 1690 670
rect 1710 650 1720 670
rect 1680 560 1720 650
rect 1760 670 1800 760
rect 1760 650 1770 670
rect 1790 650 1800 670
rect 1760 560 1800 650
rect 1840 670 1880 760
rect 1840 650 1850 670
rect 1870 650 1880 670
rect 1840 560 1880 650
rect 1920 670 1960 760
rect 1920 650 1930 670
rect 1950 650 1960 670
rect 1920 560 1960 650
rect 2000 670 2040 760
rect 2000 650 2010 670
rect 2030 650 2040 670
rect 2000 560 2040 650
rect 2160 670 2200 760
rect 2160 650 2170 670
rect 2190 650 2200 670
rect 2160 560 2200 650
rect 2240 670 2280 760
rect 2240 650 2250 670
rect 2270 650 2280 670
rect 2240 560 2280 650
rect 2320 670 2360 760
rect 2320 650 2330 670
rect 2350 650 2360 670
rect 2320 560 2360 650
rect 2400 670 2440 760
rect 2400 650 2410 670
rect 2430 650 2440 670
rect 2400 560 2440 650
rect 2480 670 2520 760
rect 2480 650 2490 670
rect 2510 650 2520 670
rect 2480 560 2520 650
rect 2640 670 2680 760
rect 2640 650 2650 670
rect 2670 650 2680 670
rect 2640 560 2680 650
rect 2720 670 2760 760
rect 2720 650 2730 670
rect 2750 650 2760 670
rect 2720 560 2760 650
rect 2800 670 2840 760
rect 2800 650 2810 670
rect 2830 650 2840 670
rect 2800 560 2840 650
rect 2880 670 2920 760
rect 2880 650 2890 670
rect 2910 650 2920 670
rect 2880 560 2920 650
rect 2960 670 3000 760
rect 2960 650 2970 670
rect 2990 650 3000 670
rect 2960 560 3000 650
rect 3040 670 3080 760
rect 3040 650 3050 670
rect 3070 650 3080 670
rect 3040 560 3080 650
rect 3120 670 3160 760
rect 3120 650 3130 670
rect 3150 650 3160 670
rect 3120 560 3160 650
rect 3200 670 3240 760
rect 3200 650 3210 670
rect 3230 650 3240 670
rect 3200 560 3240 650
rect 3280 670 3320 760
rect 3280 650 3290 670
rect 3310 650 3320 670
rect 3280 560 3320 650
rect 3360 670 3400 760
rect 3360 650 3370 670
rect 3390 650 3400 670
rect 3360 560 3400 650
rect 3440 670 3480 760
rect 3440 650 3450 670
rect 3470 650 3480 670
rect 3440 560 3480 650
rect 3600 670 3640 760
rect 3600 650 3610 670
rect 3630 650 3640 670
rect 3600 560 3640 650
rect 3680 670 3720 760
rect 3680 650 3690 670
rect 3710 650 3720 670
rect 3680 560 3720 650
rect 3760 670 3800 760
rect 3760 650 3770 670
rect 3790 650 3800 670
rect 3760 560 3800 650
rect 3840 670 3880 760
rect 3840 650 3850 670
rect 3870 650 3880 670
rect 3840 560 3880 650
rect 3920 670 3960 760
rect 3920 650 3930 670
rect 3950 650 3960 670
rect 3920 560 3960 650
rect 4080 670 4120 760
rect 4080 650 4090 670
rect 4110 650 4120 670
rect 4080 560 4120 650
rect 4160 520 4200 800
rect 0 480 60 520
rect 4140 480 4200 520
rect 0 460 40 480
rect 4160 460 4200 480
rect 260 435 1060 440
rect 260 405 270 435
rect 1050 405 1060 435
rect 260 400 1060 405
rect 1220 435 2020 440
rect 1220 405 1230 435
rect 2010 405 2020 435
rect 1220 400 2020 405
rect 2180 435 2980 440
rect 2180 405 2190 435
rect 2970 405 2980 435
rect 2180 400 2980 405
rect 3140 435 3940 440
rect 3140 405 3150 435
rect 3930 405 3940 435
rect 3140 400 3940 405
rect 160 370 200 380
rect 160 290 165 370
rect 195 290 200 370
rect 160 280 200 290
rect 1120 370 1160 380
rect 1120 290 1125 370
rect 1155 290 1160 370
rect 1120 240 1160 290
rect 2080 370 2120 380
rect 2080 290 2085 370
rect 2115 290 2120 370
rect 2080 280 2120 290
rect 3040 370 3080 380
rect 3040 290 3045 370
rect 3075 290 3080 370
rect 3040 240 3080 290
rect 4000 370 4040 380
rect 4000 290 4005 370
rect 4035 290 4040 370
rect 4000 280 4040 290
rect 1120 200 3080 240
rect 0 40 40 60
rect 160 170 200 180
rect 160 90 165 170
rect 195 90 200 170
rect 160 40 200 90
rect 1120 170 1160 180
rect 1120 90 1125 170
rect 1155 90 1160 170
rect 1120 80 1160 90
rect 2080 170 2120 200
rect 2080 90 2085 170
rect 2115 90 2120 170
rect 2080 80 2120 90
rect 3040 170 3080 180
rect 3040 90 3045 170
rect 3075 90 3080 170
rect 3040 80 3080 90
rect 4000 170 4040 180
rect 4000 90 4005 170
rect 4035 90 4040 170
rect 4000 40 4040 90
rect 4160 40 4200 60
rect 0 0 60 40
rect 4140 0 4200 40
<< viali >>
rect 165 2550 195 2830
rect 1125 2550 1155 2830
rect 2085 2550 2115 2830
rect 3045 2550 3075 2830
rect 4005 2550 4035 2830
rect 165 2170 195 2450
rect 1125 2170 1155 2450
rect 2085 2170 2115 2450
rect 3045 2170 3075 2450
rect 4005 2170 4035 2450
rect 270 2085 1050 2115
rect 1230 2085 2010 2115
rect 2190 2085 2970 2115
rect 3150 2085 3930 2115
rect 165 1430 195 1710
rect 1125 1430 1155 1710
rect 2085 1430 2115 1710
rect 3045 1430 3075 1710
rect 4005 1430 4035 1710
rect 165 1050 195 1330
rect 1125 1050 1155 1330
rect 2085 1050 2115 1330
rect 3045 1050 3075 1330
rect 4005 1050 4035 1330
rect 270 965 1050 995
rect 1230 965 2010 995
rect 2190 965 2970 995
rect 3150 965 3930 995
rect 90 650 110 670
rect 250 650 270 670
rect 330 650 350 670
rect 410 650 430 670
rect 490 650 510 670
rect 570 650 590 670
rect 730 650 750 670
rect 810 650 830 670
rect 890 650 910 670
rect 970 650 990 670
rect 1050 650 1070 670
rect 1130 650 1150 670
rect 1210 650 1230 670
rect 1290 650 1310 670
rect 1370 650 1390 670
rect 1450 650 1470 670
rect 1530 650 1550 670
rect 1690 650 1710 670
rect 1770 650 1790 670
rect 1850 650 1870 670
rect 1930 650 1950 670
rect 2010 650 2030 670
rect 2170 650 2190 670
rect 2250 650 2270 670
rect 2330 650 2350 670
rect 2410 650 2430 670
rect 2490 650 2510 670
rect 2650 650 2670 670
rect 2730 650 2750 670
rect 2810 650 2830 670
rect 2890 650 2910 670
rect 2970 650 2990 670
rect 3050 650 3070 670
rect 3130 650 3150 670
rect 3210 650 3230 670
rect 3290 650 3310 670
rect 3370 650 3390 670
rect 3450 650 3470 670
rect 3610 650 3630 670
rect 3690 650 3710 670
rect 3770 650 3790 670
rect 3850 650 3870 670
rect 3930 650 3950 670
rect 4090 650 4110 670
rect 270 405 1050 435
rect 1230 405 2010 435
rect 2190 405 2970 435
rect 3150 405 3930 435
rect 165 290 195 370
rect 1125 290 1155 370
rect 2085 290 2115 370
rect 3045 290 3075 370
rect 4005 290 4035 370
rect 165 90 195 170
rect 1125 90 1155 170
rect 2085 90 2115 170
rect 3045 90 3075 170
rect 4005 90 4035 170
<< metal1 >>
rect 160 2830 200 2840
rect 160 2550 165 2830
rect 195 2550 200 2830
rect 160 2450 200 2550
rect 1120 2830 1160 2840
rect 1120 2550 1125 2830
rect 1155 2550 1160 2830
rect 1120 2540 1160 2550
rect 2080 2830 2120 2840
rect 2080 2550 2085 2830
rect 2115 2550 2120 2830
rect 2080 2540 2120 2550
rect 3040 2830 3080 2840
rect 3040 2550 3045 2830
rect 3075 2550 3080 2830
rect 3040 2540 3080 2550
rect 4000 2830 4040 2840
rect 4000 2550 4005 2830
rect 4035 2550 4040 2830
rect 160 2170 165 2450
rect 195 2170 200 2450
rect 0 1995 40 2000
rect 0 1965 5 1995
rect 35 1965 40 1995
rect 0 1835 40 1965
rect 0 1805 5 1835
rect 35 1805 40 1835
rect 0 1800 40 1805
rect 80 1995 120 2000
rect 80 1965 85 1995
rect 115 1965 120 1995
rect 80 1835 120 1965
rect 80 1805 85 1835
rect 115 1805 120 1835
rect 80 1800 120 1805
rect 160 1995 200 2170
rect 1120 2450 1160 2460
rect 1120 2170 1125 2450
rect 1155 2170 1160 2450
rect 1120 2160 1160 2170
rect 2080 2450 2120 2460
rect 2080 2170 2085 2450
rect 2115 2170 2120 2450
rect 260 2115 1060 2120
rect 260 2085 270 2115
rect 1050 2085 1060 2115
rect 260 2080 1060 2085
rect 1220 2115 2020 2120
rect 1220 2085 1230 2115
rect 2010 2085 2020 2115
rect 1220 2080 2020 2085
rect 160 1965 165 1995
rect 195 1965 200 1995
rect 160 1835 200 1965
rect 160 1805 165 1835
rect 195 1805 200 1835
rect 160 1710 200 1805
rect 240 1995 280 2000
rect 240 1965 245 1995
rect 275 1965 280 1995
rect 240 1835 280 1965
rect 240 1805 245 1835
rect 275 1805 280 1835
rect 240 1800 280 1805
rect 320 1995 360 2000
rect 320 1965 325 1995
rect 355 1965 360 1995
rect 320 1835 360 1965
rect 320 1805 325 1835
rect 355 1805 360 1835
rect 320 1800 360 1805
rect 400 1995 440 2000
rect 400 1965 405 1995
rect 435 1965 440 1995
rect 400 1835 440 1965
rect 400 1805 405 1835
rect 435 1805 440 1835
rect 400 1800 440 1805
rect 480 1995 520 2000
rect 480 1965 485 1995
rect 515 1965 520 1995
rect 480 1835 520 1965
rect 480 1805 485 1835
rect 515 1805 520 1835
rect 480 1800 520 1805
rect 560 1995 600 2000
rect 560 1965 565 1995
rect 595 1965 600 1995
rect 560 1835 600 1965
rect 640 1915 680 2080
rect 640 1885 645 1915
rect 675 1885 680 1915
rect 640 1880 680 1885
rect 720 1995 760 2000
rect 720 1965 725 1995
rect 755 1965 760 1995
rect 560 1805 565 1835
rect 595 1805 600 1835
rect 560 1800 600 1805
rect 720 1835 760 1965
rect 720 1805 725 1835
rect 755 1805 760 1835
rect 720 1800 760 1805
rect 800 1995 840 2000
rect 800 1965 805 1995
rect 835 1965 840 1995
rect 800 1835 840 1965
rect 800 1805 805 1835
rect 835 1805 840 1835
rect 800 1800 840 1805
rect 880 1995 920 2000
rect 880 1965 885 1995
rect 915 1965 920 1995
rect 880 1835 920 1965
rect 880 1805 885 1835
rect 915 1805 920 1835
rect 880 1800 920 1805
rect 960 1995 1000 2000
rect 960 1965 965 1995
rect 995 1965 1000 1995
rect 960 1835 1000 1965
rect 960 1805 965 1835
rect 995 1805 1000 1835
rect 960 1800 1000 1805
rect 1040 1995 1080 2000
rect 1040 1965 1045 1995
rect 1075 1965 1080 1995
rect 1040 1835 1080 1965
rect 1040 1805 1045 1835
rect 1075 1805 1080 1835
rect 1040 1800 1080 1805
rect 1120 1995 1160 2000
rect 1120 1965 1125 1995
rect 1155 1965 1160 1995
rect 1120 1835 1160 1965
rect 1120 1805 1125 1835
rect 1155 1805 1160 1835
rect 1120 1800 1160 1805
rect 1200 1995 1240 2000
rect 1200 1965 1205 1995
rect 1235 1965 1240 1995
rect 1200 1835 1240 1965
rect 1200 1805 1205 1835
rect 1235 1805 1240 1835
rect 1200 1800 1240 1805
rect 1280 1995 1320 2000
rect 1280 1965 1285 1995
rect 1315 1965 1320 1995
rect 1280 1835 1320 1965
rect 1280 1805 1285 1835
rect 1315 1805 1320 1835
rect 1280 1800 1320 1805
rect 1360 1995 1400 2000
rect 1360 1965 1365 1995
rect 1395 1965 1400 1995
rect 1360 1835 1400 1965
rect 1360 1805 1365 1835
rect 1395 1805 1400 1835
rect 1360 1800 1400 1805
rect 1440 1995 1480 2000
rect 1440 1965 1445 1995
rect 1475 1965 1480 1995
rect 1440 1835 1480 1965
rect 1440 1805 1445 1835
rect 1475 1805 1480 1835
rect 1440 1800 1480 1805
rect 1520 1995 1560 2000
rect 1520 1965 1525 1995
rect 1555 1965 1560 1995
rect 1520 1835 1560 1965
rect 1600 1915 1640 2080
rect 1600 1885 1605 1915
rect 1635 1885 1640 1915
rect 1600 1880 1640 1885
rect 1680 1995 1720 2000
rect 1680 1965 1685 1995
rect 1715 1965 1720 1995
rect 1520 1805 1525 1835
rect 1555 1805 1560 1835
rect 1520 1800 1560 1805
rect 1680 1835 1720 1965
rect 1680 1805 1685 1835
rect 1715 1805 1720 1835
rect 1680 1800 1720 1805
rect 1760 1995 1800 2000
rect 1760 1965 1765 1995
rect 1795 1965 1800 1995
rect 1760 1835 1800 1965
rect 1760 1805 1765 1835
rect 1795 1805 1800 1835
rect 1760 1800 1800 1805
rect 1840 1995 1880 2000
rect 1840 1965 1845 1995
rect 1875 1965 1880 1995
rect 1840 1835 1880 1965
rect 1840 1805 1845 1835
rect 1875 1805 1880 1835
rect 1840 1800 1880 1805
rect 1920 1995 1960 2000
rect 1920 1965 1925 1995
rect 1955 1965 1960 1995
rect 1920 1835 1960 1965
rect 1920 1805 1925 1835
rect 1955 1805 1960 1835
rect 1920 1800 1960 1805
rect 2000 1995 2040 2000
rect 2000 1965 2005 1995
rect 2035 1965 2040 1995
rect 2000 1835 2040 1965
rect 2000 1805 2005 1835
rect 2035 1805 2040 1835
rect 2000 1800 2040 1805
rect 2080 1995 2120 2170
rect 3040 2450 3080 2460
rect 3040 2170 3045 2450
rect 3075 2170 3080 2450
rect 3040 2160 3080 2170
rect 4000 2450 4040 2550
rect 4000 2170 4005 2450
rect 4035 2170 4040 2450
rect 2180 2115 2980 2120
rect 2180 2085 2190 2115
rect 2970 2085 2980 2115
rect 2180 2080 2980 2085
rect 3140 2115 3940 2120
rect 3140 2085 3150 2115
rect 3930 2085 3940 2115
rect 3140 2080 3940 2085
rect 2080 1965 2085 1995
rect 2115 1965 2120 1995
rect 2080 1835 2120 1965
rect 2080 1805 2085 1835
rect 2115 1805 2120 1835
rect 2080 1800 2120 1805
rect 2160 1995 2200 2000
rect 2160 1965 2165 1995
rect 2195 1965 2200 1995
rect 2160 1835 2200 1965
rect 2160 1805 2165 1835
rect 2195 1805 2200 1835
rect 2160 1800 2200 1805
rect 2240 1995 2280 2000
rect 2240 1965 2245 1995
rect 2275 1965 2280 1995
rect 2240 1835 2280 1965
rect 2240 1805 2245 1835
rect 2275 1805 2280 1835
rect 2240 1800 2280 1805
rect 2320 1995 2360 2000
rect 2320 1965 2325 1995
rect 2355 1965 2360 1995
rect 2320 1835 2360 1965
rect 2320 1805 2325 1835
rect 2355 1805 2360 1835
rect 2320 1800 2360 1805
rect 2400 1995 2440 2000
rect 2400 1965 2405 1995
rect 2435 1965 2440 1995
rect 2400 1835 2440 1965
rect 2400 1805 2405 1835
rect 2435 1805 2440 1835
rect 2400 1800 2440 1805
rect 2480 1995 2520 2000
rect 2480 1965 2485 1995
rect 2515 1965 2520 1995
rect 2480 1835 2520 1965
rect 2560 1915 2600 2080
rect 2560 1885 2565 1915
rect 2595 1885 2600 1915
rect 2560 1880 2600 1885
rect 2640 1995 2680 2000
rect 2640 1965 2645 1995
rect 2675 1965 2680 1995
rect 2480 1805 2485 1835
rect 2515 1805 2520 1835
rect 2480 1800 2520 1805
rect 2640 1835 2680 1965
rect 2640 1805 2645 1835
rect 2675 1805 2680 1835
rect 2640 1800 2680 1805
rect 2720 1995 2760 2000
rect 2720 1965 2725 1995
rect 2755 1965 2760 1995
rect 2720 1835 2760 1965
rect 2720 1805 2725 1835
rect 2755 1805 2760 1835
rect 2720 1800 2760 1805
rect 2800 1995 2840 2000
rect 2800 1965 2805 1995
rect 2835 1965 2840 1995
rect 2800 1835 2840 1965
rect 2800 1805 2805 1835
rect 2835 1805 2840 1835
rect 2800 1800 2840 1805
rect 2880 1995 2920 2000
rect 2880 1965 2885 1995
rect 2915 1965 2920 1995
rect 2880 1835 2920 1965
rect 2880 1805 2885 1835
rect 2915 1805 2920 1835
rect 2880 1800 2920 1805
rect 2960 1995 3000 2000
rect 2960 1965 2965 1995
rect 2995 1965 3000 1995
rect 2960 1835 3000 1965
rect 2960 1805 2965 1835
rect 2995 1805 3000 1835
rect 2960 1800 3000 1805
rect 3040 1995 3080 2000
rect 3040 1965 3045 1995
rect 3075 1965 3080 1995
rect 3040 1835 3080 1965
rect 3040 1805 3045 1835
rect 3075 1805 3080 1835
rect 3040 1800 3080 1805
rect 3120 1995 3160 2000
rect 3120 1965 3125 1995
rect 3155 1965 3160 1995
rect 3120 1835 3160 1965
rect 3120 1805 3125 1835
rect 3155 1805 3160 1835
rect 3120 1800 3160 1805
rect 3200 1995 3240 2000
rect 3200 1965 3205 1995
rect 3235 1965 3240 1995
rect 3200 1835 3240 1965
rect 3200 1805 3205 1835
rect 3235 1805 3240 1835
rect 3200 1800 3240 1805
rect 3280 1995 3320 2000
rect 3280 1965 3285 1995
rect 3315 1965 3320 1995
rect 3280 1835 3320 1965
rect 3280 1805 3285 1835
rect 3315 1805 3320 1835
rect 3280 1800 3320 1805
rect 3360 1995 3400 2000
rect 3360 1965 3365 1995
rect 3395 1965 3400 1995
rect 3360 1835 3400 1965
rect 3360 1805 3365 1835
rect 3395 1805 3400 1835
rect 3360 1800 3400 1805
rect 3440 1995 3480 2000
rect 3440 1965 3445 1995
rect 3475 1965 3480 1995
rect 3440 1835 3480 1965
rect 3520 1915 3560 2080
rect 3520 1885 3525 1915
rect 3555 1885 3560 1915
rect 3520 1880 3560 1885
rect 3600 1995 3640 2000
rect 3600 1965 3605 1995
rect 3635 1965 3640 1995
rect 3440 1805 3445 1835
rect 3475 1805 3480 1835
rect 3440 1800 3480 1805
rect 3600 1835 3640 1965
rect 3600 1805 3605 1835
rect 3635 1805 3640 1835
rect 3600 1800 3640 1805
rect 3680 1995 3720 2000
rect 3680 1965 3685 1995
rect 3715 1965 3720 1995
rect 3680 1835 3720 1965
rect 3680 1805 3685 1835
rect 3715 1805 3720 1835
rect 3680 1800 3720 1805
rect 3760 1995 3800 2000
rect 3760 1965 3765 1995
rect 3795 1965 3800 1995
rect 3760 1835 3800 1965
rect 3760 1805 3765 1835
rect 3795 1805 3800 1835
rect 3760 1800 3800 1805
rect 3840 1995 3880 2000
rect 3840 1965 3845 1995
rect 3875 1965 3880 1995
rect 3840 1835 3880 1965
rect 3840 1805 3845 1835
rect 3875 1805 3880 1835
rect 3840 1800 3880 1805
rect 3920 1995 3960 2000
rect 3920 1965 3925 1995
rect 3955 1965 3960 1995
rect 3920 1835 3960 1965
rect 3920 1805 3925 1835
rect 3955 1805 3960 1835
rect 3920 1800 3960 1805
rect 4000 1995 4040 2170
rect 4000 1965 4005 1995
rect 4035 1965 4040 1995
rect 4000 1835 4040 1965
rect 4000 1805 4005 1835
rect 4035 1805 4040 1835
rect 160 1430 165 1710
rect 195 1430 200 1710
rect 160 1420 200 1430
rect 1120 1710 1160 1720
rect 1120 1430 1125 1710
rect 1155 1430 1160 1710
rect 1120 1420 1160 1430
rect 2080 1710 2120 1720
rect 2080 1430 2085 1710
rect 2115 1430 2120 1710
rect 2080 1400 2120 1430
rect 3040 1710 3080 1720
rect 3040 1430 3045 1710
rect 3075 1430 3080 1710
rect 3040 1420 3080 1430
rect 4000 1710 4040 1805
rect 4080 1995 4120 2000
rect 4080 1965 4085 1995
rect 4115 1965 4120 1995
rect 4080 1835 4120 1965
rect 4080 1805 4085 1835
rect 4115 1805 4120 1835
rect 4080 1800 4120 1805
rect 4160 1995 4200 2000
rect 4160 1965 4165 1995
rect 4195 1965 4200 1995
rect 4160 1835 4200 1965
rect 4160 1805 4165 1835
rect 4195 1805 4200 1835
rect 4160 1800 4200 1805
rect 4000 1430 4005 1710
rect 4035 1430 4040 1710
rect 4000 1420 4040 1430
rect 1120 1395 1160 1400
rect 1120 1365 1125 1395
rect 1155 1365 1160 1395
rect 160 1330 200 1340
rect 160 1050 165 1330
rect 195 1050 200 1330
rect 80 670 120 680
rect 80 650 90 670
rect 110 650 120 670
rect 80 640 120 650
rect 160 595 200 1050
rect 1120 1330 1160 1365
rect 3040 1395 3080 1400
rect 3040 1365 3045 1395
rect 3075 1365 3080 1395
rect 1120 1050 1125 1330
rect 1155 1050 1160 1330
rect 1120 1040 1160 1050
rect 2080 1330 2120 1340
rect 2080 1050 2085 1330
rect 2115 1050 2120 1330
rect 260 995 1060 1000
rect 260 965 270 995
rect 1050 965 1060 995
rect 260 960 1060 965
rect 1220 995 2020 1000
rect 1220 965 1230 995
rect 2010 965 2020 995
rect 1220 960 2020 965
rect 640 755 680 960
rect 640 725 645 755
rect 675 725 680 755
rect 240 670 280 680
rect 240 650 250 670
rect 270 650 280 670
rect 240 640 280 650
rect 320 670 360 680
rect 320 650 330 670
rect 350 650 360 670
rect 320 640 360 650
rect 400 670 440 680
rect 400 650 410 670
rect 430 650 440 670
rect 400 640 440 650
rect 480 670 520 680
rect 480 650 490 670
rect 510 650 520 670
rect 480 640 520 650
rect 560 670 600 680
rect 560 650 570 670
rect 590 650 600 670
rect 560 640 600 650
rect 160 565 165 595
rect 195 565 200 595
rect 160 370 200 565
rect 640 440 680 725
rect 1600 755 1640 960
rect 1600 725 1605 755
rect 1635 725 1640 755
rect 720 670 760 680
rect 720 650 730 670
rect 750 650 760 670
rect 720 640 760 650
rect 800 670 840 680
rect 800 650 810 670
rect 830 650 840 670
rect 800 640 840 650
rect 880 670 920 680
rect 880 650 890 670
rect 910 650 920 670
rect 880 640 920 650
rect 960 670 1000 680
rect 960 650 970 670
rect 990 650 1000 670
rect 960 640 1000 650
rect 1040 670 1080 680
rect 1040 650 1050 670
rect 1070 650 1080 670
rect 1040 640 1080 650
rect 1120 670 1160 680
rect 1120 650 1130 670
rect 1150 650 1160 670
rect 1120 640 1160 650
rect 1200 670 1240 680
rect 1200 650 1210 670
rect 1230 650 1240 670
rect 1200 640 1240 650
rect 1280 670 1320 680
rect 1280 650 1290 670
rect 1310 650 1320 670
rect 1280 640 1320 650
rect 1360 670 1400 680
rect 1360 650 1370 670
rect 1390 650 1400 670
rect 1360 640 1400 650
rect 1440 670 1480 680
rect 1440 650 1450 670
rect 1470 650 1480 670
rect 1440 640 1480 650
rect 1520 670 1560 680
rect 1520 650 1530 670
rect 1550 650 1560 670
rect 1520 640 1560 650
rect 1600 440 1640 725
rect 1680 670 1720 680
rect 1680 650 1690 670
rect 1710 650 1720 670
rect 1680 640 1720 650
rect 1760 670 1800 680
rect 1760 650 1770 670
rect 1790 650 1800 670
rect 1760 640 1800 650
rect 1840 670 1880 680
rect 1840 650 1850 670
rect 1870 650 1880 670
rect 1840 640 1880 650
rect 1920 670 1960 680
rect 1920 650 1930 670
rect 1950 650 1960 670
rect 1920 640 1960 650
rect 2000 670 2040 680
rect 2000 650 2010 670
rect 2030 650 2040 670
rect 2000 640 2040 650
rect 2080 595 2120 1050
rect 3040 1330 3080 1365
rect 3040 1050 3045 1330
rect 3075 1050 3080 1330
rect 3040 1040 3080 1050
rect 4000 1330 4040 1340
rect 4000 1050 4005 1330
rect 4035 1050 4040 1330
rect 2180 995 2980 1000
rect 2180 965 2190 995
rect 2970 965 2980 995
rect 2180 960 2980 965
rect 3140 995 3940 1000
rect 3140 965 3150 995
rect 3930 965 3940 995
rect 3140 960 3940 965
rect 2560 755 2600 960
rect 2560 725 2565 755
rect 2595 725 2600 755
rect 2160 670 2200 680
rect 2160 650 2170 670
rect 2190 650 2200 670
rect 2160 640 2200 650
rect 2240 670 2280 680
rect 2240 650 2250 670
rect 2270 650 2280 670
rect 2240 640 2280 650
rect 2320 670 2360 680
rect 2320 650 2330 670
rect 2350 650 2360 670
rect 2320 640 2360 650
rect 2400 670 2440 680
rect 2400 650 2410 670
rect 2430 650 2440 670
rect 2400 640 2440 650
rect 2480 670 2520 680
rect 2480 650 2490 670
rect 2510 650 2520 670
rect 2480 640 2520 650
rect 2080 565 2085 595
rect 2115 565 2120 595
rect 260 435 1060 440
rect 260 405 270 435
rect 1050 405 1060 435
rect 260 400 1060 405
rect 1220 435 2020 440
rect 1220 405 1230 435
rect 2010 405 2020 435
rect 1220 400 2020 405
rect 160 290 165 370
rect 195 290 200 370
rect 160 280 200 290
rect 1120 370 1160 380
rect 1120 290 1125 370
rect 1155 290 1160 370
rect 1120 275 1160 290
rect 2080 370 2120 565
rect 2560 440 2600 725
rect 3520 755 3560 960
rect 3520 725 3525 755
rect 3555 725 3560 755
rect 2640 670 2680 680
rect 2640 650 2650 670
rect 2670 650 2680 670
rect 2640 640 2680 650
rect 2720 670 2760 680
rect 2720 650 2730 670
rect 2750 650 2760 670
rect 2720 640 2760 650
rect 2800 670 2840 680
rect 2800 650 2810 670
rect 2830 650 2840 670
rect 2800 640 2840 650
rect 2880 670 2920 680
rect 2880 650 2890 670
rect 2910 650 2920 670
rect 2880 640 2920 650
rect 2960 670 3000 680
rect 2960 650 2970 670
rect 2990 650 3000 670
rect 2960 640 3000 650
rect 3040 670 3080 680
rect 3040 650 3050 670
rect 3070 650 3080 670
rect 3040 640 3080 650
rect 3120 670 3160 680
rect 3120 650 3130 670
rect 3150 650 3160 670
rect 3120 640 3160 650
rect 3200 670 3240 680
rect 3200 650 3210 670
rect 3230 650 3240 670
rect 3200 640 3240 650
rect 3280 670 3320 680
rect 3280 650 3290 670
rect 3310 650 3320 670
rect 3280 640 3320 650
rect 3360 670 3400 680
rect 3360 650 3370 670
rect 3390 650 3400 670
rect 3360 640 3400 650
rect 3440 670 3480 680
rect 3440 650 3450 670
rect 3470 650 3480 670
rect 3440 640 3480 650
rect 3520 440 3560 725
rect 3600 670 3640 680
rect 3600 650 3610 670
rect 3630 650 3640 670
rect 3600 640 3640 650
rect 3680 670 3720 680
rect 3680 650 3690 670
rect 3710 650 3720 670
rect 3680 640 3720 650
rect 3760 670 3800 680
rect 3760 650 3770 670
rect 3790 650 3800 670
rect 3760 640 3800 650
rect 3840 670 3880 680
rect 3840 650 3850 670
rect 3870 650 3880 670
rect 3840 640 3880 650
rect 3920 670 3960 680
rect 3920 650 3930 670
rect 3950 650 3960 670
rect 3920 640 3960 650
rect 4000 595 4040 1050
rect 4080 670 4120 680
rect 4080 650 4090 670
rect 4110 650 4120 670
rect 4080 640 4120 650
rect 4000 565 4005 595
rect 4035 565 4040 595
rect 2180 435 2980 440
rect 2180 405 2190 435
rect 2970 405 2980 435
rect 2180 400 2980 405
rect 3140 435 3940 440
rect 3140 405 3150 435
rect 3930 405 3940 435
rect 3140 400 3940 405
rect 2080 290 2085 370
rect 2115 290 2120 370
rect 2080 280 2120 290
rect 3040 370 3080 380
rect 3040 290 3045 370
rect 3075 290 3080 370
rect 1120 245 1125 275
rect 1155 245 1160 275
rect 1120 240 1160 245
rect 3040 275 3080 290
rect 4000 370 4040 565
rect 4000 290 4005 370
rect 4035 290 4040 370
rect 4000 280 4040 290
rect 3040 245 3045 275
rect 3075 245 3080 275
rect 3040 240 3080 245
rect 160 170 200 180
rect 160 90 165 170
rect 195 90 200 170
rect 160 80 200 90
rect 1120 170 1160 180
rect 1120 90 1125 170
rect 1155 90 1160 170
rect 1120 80 1160 90
rect 2080 170 2120 200
rect 2080 90 2085 170
rect 2115 90 2120 170
rect 2080 80 2120 90
rect 3040 170 3080 180
rect 3040 90 3045 170
rect 3075 90 3080 170
rect 3040 80 3080 90
rect 4000 170 4040 180
rect 4000 90 4005 170
rect 4035 90 4040 170
rect 4000 80 4040 90
<< via1 >>
rect 2085 2650 2115 2830
rect 5 1965 35 1995
rect 5 1805 35 1835
rect 85 1965 115 1995
rect 85 1805 115 1835
rect 165 1965 195 1995
rect 165 1805 195 1835
rect 245 1965 275 1995
rect 245 1805 275 1835
rect 325 1965 355 1995
rect 325 1805 355 1835
rect 405 1965 435 1995
rect 405 1805 435 1835
rect 485 1965 515 1995
rect 485 1805 515 1835
rect 565 1965 595 1995
rect 645 1885 675 1915
rect 725 1965 755 1995
rect 565 1805 595 1835
rect 725 1805 755 1835
rect 805 1965 835 1995
rect 805 1805 835 1835
rect 885 1965 915 1995
rect 885 1805 915 1835
rect 965 1965 995 1995
rect 965 1805 995 1835
rect 1045 1965 1075 1995
rect 1045 1805 1075 1835
rect 1125 1965 1155 1995
rect 1125 1805 1155 1835
rect 1205 1965 1235 1995
rect 1205 1805 1235 1835
rect 1285 1965 1315 1995
rect 1285 1805 1315 1835
rect 1365 1965 1395 1995
rect 1365 1805 1395 1835
rect 1445 1965 1475 1995
rect 1445 1805 1475 1835
rect 1525 1965 1555 1995
rect 1605 1885 1635 1915
rect 1685 1965 1715 1995
rect 1525 1805 1555 1835
rect 1685 1805 1715 1835
rect 1765 1965 1795 1995
rect 1765 1805 1795 1835
rect 1845 1965 1875 1995
rect 1845 1805 1875 1835
rect 1925 1965 1955 1995
rect 1925 1805 1955 1835
rect 2005 1965 2035 1995
rect 2005 1805 2035 1835
rect 2085 1965 2115 1995
rect 2085 1805 2115 1835
rect 2165 1965 2195 1995
rect 2165 1805 2195 1835
rect 2245 1965 2275 1995
rect 2245 1805 2275 1835
rect 2325 1965 2355 1995
rect 2325 1805 2355 1835
rect 2405 1965 2435 1995
rect 2405 1805 2435 1835
rect 2485 1965 2515 1995
rect 2565 1885 2595 1915
rect 2645 1965 2675 1995
rect 2485 1805 2515 1835
rect 2645 1805 2675 1835
rect 2725 1965 2755 1995
rect 2725 1805 2755 1835
rect 2805 1965 2835 1995
rect 2805 1805 2835 1835
rect 2885 1965 2915 1995
rect 2885 1805 2915 1835
rect 2965 1965 2995 1995
rect 2965 1805 2995 1835
rect 3045 1965 3075 1995
rect 3045 1805 3075 1835
rect 3125 1965 3155 1995
rect 3125 1805 3155 1835
rect 3205 1965 3235 1995
rect 3205 1805 3235 1835
rect 3285 1965 3315 1995
rect 3285 1805 3315 1835
rect 3365 1965 3395 1995
rect 3365 1805 3395 1835
rect 3445 1965 3475 1995
rect 3525 1885 3555 1915
rect 3605 1965 3635 1995
rect 3445 1805 3475 1835
rect 3605 1805 3635 1835
rect 3685 1965 3715 1995
rect 3685 1805 3715 1835
rect 3765 1965 3795 1995
rect 3765 1805 3795 1835
rect 3845 1965 3875 1995
rect 3845 1805 3875 1835
rect 3925 1965 3955 1995
rect 3925 1805 3955 1835
rect 4005 1965 4035 1995
rect 4005 1805 4035 1835
rect 4085 1965 4115 1995
rect 4085 1805 4115 1835
rect 4165 1965 4195 1995
rect 4165 1805 4195 1835
rect 1125 1365 1155 1395
rect 3045 1365 3075 1395
rect 645 725 675 755
rect 165 565 195 595
rect 1605 725 1635 755
rect 2565 725 2595 755
rect 2085 565 2115 595
rect 3525 725 3555 755
rect 4005 565 4035 595
rect 1125 245 1155 275
rect 3045 245 3075 275
rect 165 90 195 170
rect 4005 90 4035 170
<< metal2 >>
rect 2080 2830 2120 2840
rect 2080 2650 2085 2830
rect 2115 2650 2120 2830
rect 2080 2640 2120 2650
rect 0 1995 4200 2000
rect 0 1965 5 1995
rect 35 1965 85 1995
rect 115 1965 165 1995
rect 195 1965 245 1995
rect 275 1965 325 1995
rect 355 1965 405 1995
rect 435 1965 485 1995
rect 515 1965 565 1995
rect 595 1965 725 1995
rect 755 1965 805 1995
rect 835 1965 885 1995
rect 915 1965 965 1995
rect 995 1965 1045 1995
rect 1075 1965 1125 1995
rect 1155 1965 1205 1995
rect 1235 1965 1285 1995
rect 1315 1965 1365 1995
rect 1395 1965 1445 1995
rect 1475 1965 1525 1995
rect 1555 1965 1685 1995
rect 1715 1965 1765 1995
rect 1795 1965 1845 1995
rect 1875 1965 1925 1995
rect 1955 1965 2005 1995
rect 2035 1965 2085 1995
rect 2115 1965 2165 1995
rect 2195 1965 2245 1995
rect 2275 1965 2325 1995
rect 2355 1965 2405 1995
rect 2435 1965 2485 1995
rect 2515 1965 2645 1995
rect 2675 1965 2725 1995
rect 2755 1965 2805 1995
rect 2835 1965 2885 1995
rect 2915 1965 2965 1995
rect 2995 1965 3045 1995
rect 3075 1965 3125 1995
rect 3155 1965 3205 1995
rect 3235 1965 3285 1995
rect 3315 1965 3365 1995
rect 3395 1965 3445 1995
rect 3475 1965 3605 1995
rect 3635 1965 3685 1995
rect 3715 1965 3765 1995
rect 3795 1965 3845 1995
rect 3875 1965 3925 1995
rect 3955 1965 4005 1995
rect 4035 1965 4085 1995
rect 4115 1965 4165 1995
rect 4195 1965 4200 1995
rect 0 1960 4200 1965
rect 0 1915 4200 1920
rect 0 1885 645 1915
rect 675 1885 1605 1915
rect 1635 1885 2565 1915
rect 2595 1885 3525 1915
rect 3555 1885 4200 1915
rect 0 1880 4200 1885
rect 0 1835 4200 1840
rect 0 1805 5 1835
rect 35 1805 85 1835
rect 115 1805 165 1835
rect 195 1805 245 1835
rect 275 1805 325 1835
rect 355 1805 405 1835
rect 435 1805 485 1835
rect 515 1805 565 1835
rect 595 1805 725 1835
rect 755 1805 805 1835
rect 835 1805 885 1835
rect 915 1805 965 1835
rect 995 1805 1045 1835
rect 1075 1805 1125 1835
rect 1155 1805 1205 1835
rect 1235 1805 1285 1835
rect 1315 1805 1365 1835
rect 1395 1805 1445 1835
rect 1475 1805 1525 1835
rect 1555 1805 1685 1835
rect 1715 1805 1765 1835
rect 1795 1805 1845 1835
rect 1875 1805 1925 1835
rect 1955 1805 2005 1835
rect 2035 1805 2085 1835
rect 2115 1805 2165 1835
rect 2195 1805 2245 1835
rect 2275 1805 2325 1835
rect 2355 1805 2405 1835
rect 2435 1805 2485 1835
rect 2515 1805 2645 1835
rect 2675 1805 2725 1835
rect 2755 1805 2805 1835
rect 2835 1805 2885 1835
rect 2915 1805 2965 1835
rect 2995 1805 3045 1835
rect 3075 1805 3125 1835
rect 3155 1805 3205 1835
rect 3235 1805 3285 1835
rect 3315 1805 3365 1835
rect 3395 1805 3445 1835
rect 3475 1805 3605 1835
rect 3635 1805 3685 1835
rect 3715 1805 3765 1835
rect 3795 1805 3845 1835
rect 3875 1805 3925 1835
rect 3955 1805 4005 1835
rect 4035 1805 4085 1835
rect 4115 1805 4165 1835
rect 4195 1805 4200 1835
rect 0 1800 4200 1805
rect 0 1395 4200 1400
rect 0 1365 1125 1395
rect 1155 1365 3045 1395
rect 3075 1365 4200 1395
rect 0 1360 4200 1365
rect 0 835 4200 840
rect 0 805 85 835
rect 115 805 245 835
rect 275 805 325 835
rect 355 805 405 835
rect 435 805 485 835
rect 515 805 565 835
rect 595 805 725 835
rect 755 805 805 835
rect 835 805 885 835
rect 915 805 965 835
rect 995 805 1045 835
rect 1075 805 1125 835
rect 1155 805 1205 835
rect 1235 805 1285 835
rect 1315 805 1365 835
rect 1395 805 1445 835
rect 1475 805 1525 835
rect 1555 805 1685 835
rect 1715 805 1765 835
rect 1795 805 1845 835
rect 1875 805 1925 835
rect 1955 805 2005 835
rect 2035 805 2165 835
rect 2195 805 2245 835
rect 2275 805 2325 835
rect 2355 805 2405 835
rect 2435 805 2485 835
rect 2515 805 2645 835
rect 2675 805 2725 835
rect 2755 805 2805 835
rect 2835 805 2885 835
rect 2915 805 2965 835
rect 2995 805 3045 835
rect 3075 805 3125 835
rect 3155 805 3205 835
rect 3235 805 3285 835
rect 3315 805 3365 835
rect 3395 805 3445 835
rect 3475 805 3605 835
rect 3635 805 3685 835
rect 3715 805 3765 835
rect 3795 805 3845 835
rect 3875 805 3925 835
rect 3955 805 4085 835
rect 4115 805 4200 835
rect 0 800 4200 805
rect 0 755 4200 760
rect 0 725 645 755
rect 675 725 1605 755
rect 1635 725 2565 755
rect 2595 725 3525 755
rect 3555 725 4200 755
rect 0 720 4200 725
rect 0 675 4200 680
rect 0 645 85 675
rect 115 645 245 675
rect 275 645 325 675
rect 355 645 405 675
rect 435 645 485 675
rect 515 645 565 675
rect 595 645 725 675
rect 755 645 805 675
rect 835 645 885 675
rect 915 645 965 675
rect 995 645 1045 675
rect 1075 645 1125 675
rect 1155 645 1205 675
rect 1235 645 1285 675
rect 1315 645 1365 675
rect 1395 645 1445 675
rect 1475 645 1525 675
rect 1555 645 1685 675
rect 1715 645 1765 675
rect 1795 645 1845 675
rect 1875 645 1925 675
rect 1955 645 2005 675
rect 2035 645 2165 675
rect 2195 645 2245 675
rect 2275 645 2325 675
rect 2355 645 2405 675
rect 2435 645 2485 675
rect 2515 645 2645 675
rect 2675 645 2725 675
rect 2755 645 2805 675
rect 2835 645 2885 675
rect 2915 645 2965 675
rect 2995 645 3045 675
rect 3075 645 3125 675
rect 3155 645 3205 675
rect 3235 645 3285 675
rect 3315 645 3365 675
rect 3395 645 3445 675
rect 3475 645 3605 675
rect 3635 645 3685 675
rect 3715 645 3765 675
rect 3795 645 3845 675
rect 3875 645 3925 675
rect 3955 645 4085 675
rect 4115 645 4200 675
rect 0 640 4200 645
rect 0 595 4200 600
rect 0 565 165 595
rect 195 565 2085 595
rect 2115 565 4005 595
rect 4035 565 4200 595
rect 0 560 4200 565
rect 0 515 4200 520
rect 0 485 85 515
rect 115 485 245 515
rect 275 485 325 515
rect 355 485 405 515
rect 435 485 485 515
rect 515 485 565 515
rect 595 485 725 515
rect 755 485 805 515
rect 835 485 885 515
rect 915 485 965 515
rect 995 485 1045 515
rect 1075 485 1125 515
rect 1155 485 1205 515
rect 1235 485 1285 515
rect 1315 485 1365 515
rect 1395 485 1445 515
rect 1475 485 1525 515
rect 1555 485 1685 515
rect 1715 485 1765 515
rect 1795 485 1845 515
rect 1875 485 1925 515
rect 1955 485 2005 515
rect 2035 485 2165 515
rect 2195 485 2245 515
rect 2275 485 2325 515
rect 2355 485 2405 515
rect 2435 485 2485 515
rect 2515 485 2645 515
rect 2675 485 2725 515
rect 2755 485 2805 515
rect 2835 485 2885 515
rect 2915 485 2965 515
rect 2995 485 3045 515
rect 3075 485 3125 515
rect 3155 485 3205 515
rect 3235 485 3285 515
rect 3315 485 3365 515
rect 3395 485 3445 515
rect 3475 485 3605 515
rect 3635 485 3685 515
rect 3715 485 3765 515
rect 3795 485 3845 515
rect 3875 485 3925 515
rect 3955 485 4085 515
rect 4115 485 4200 515
rect 0 480 4200 485
rect 0 275 4200 280
rect 0 245 1125 275
rect 1155 245 3045 275
rect 3075 245 4200 275
rect 0 240 4200 245
rect 160 170 200 180
rect 160 90 165 170
rect 195 90 200 170
rect 160 80 200 90
rect 4000 170 4040 180
rect 4000 90 4005 170
rect 4035 90 4040 170
rect 4000 80 4040 90
<< via2 >>
rect 2085 2650 2115 2830
rect 5 1965 35 1995
rect 85 1965 115 1995
rect 165 1965 195 1995
rect 245 1965 275 1995
rect 325 1965 355 1995
rect 405 1965 435 1995
rect 485 1965 515 1995
rect 565 1965 595 1995
rect 725 1965 755 1995
rect 805 1965 835 1995
rect 885 1965 915 1995
rect 965 1965 995 1995
rect 1045 1965 1075 1995
rect 1125 1965 1155 1995
rect 1205 1965 1235 1995
rect 1285 1965 1315 1995
rect 1365 1965 1395 1995
rect 1445 1965 1475 1995
rect 1525 1965 1555 1995
rect 1685 1965 1715 1995
rect 1765 1965 1795 1995
rect 1845 1965 1875 1995
rect 1925 1965 1955 1995
rect 2005 1965 2035 1995
rect 2085 1965 2115 1995
rect 2165 1965 2195 1995
rect 2245 1965 2275 1995
rect 2325 1965 2355 1995
rect 2405 1965 2435 1995
rect 2485 1965 2515 1995
rect 2645 1965 2675 1995
rect 2725 1965 2755 1995
rect 2805 1965 2835 1995
rect 2885 1965 2915 1995
rect 2965 1965 2995 1995
rect 3045 1965 3075 1995
rect 3125 1965 3155 1995
rect 3205 1965 3235 1995
rect 3285 1965 3315 1995
rect 3365 1965 3395 1995
rect 3445 1965 3475 1995
rect 3605 1965 3635 1995
rect 3685 1965 3715 1995
rect 3765 1965 3795 1995
rect 3845 1965 3875 1995
rect 3925 1965 3955 1995
rect 4005 1965 4035 1995
rect 4085 1965 4115 1995
rect 4165 1965 4195 1995
rect 5 1805 35 1835
rect 85 1805 115 1835
rect 165 1805 195 1835
rect 245 1805 275 1835
rect 325 1805 355 1835
rect 405 1805 435 1835
rect 485 1805 515 1835
rect 565 1805 595 1835
rect 725 1805 755 1835
rect 805 1805 835 1835
rect 885 1805 915 1835
rect 965 1805 995 1835
rect 1045 1805 1075 1835
rect 1125 1805 1155 1835
rect 1205 1805 1235 1835
rect 1285 1805 1315 1835
rect 1365 1805 1395 1835
rect 1445 1805 1475 1835
rect 1525 1805 1555 1835
rect 1685 1805 1715 1835
rect 1765 1805 1795 1835
rect 1845 1805 1875 1835
rect 1925 1805 1955 1835
rect 2005 1805 2035 1835
rect 2085 1805 2115 1835
rect 2165 1805 2195 1835
rect 2245 1805 2275 1835
rect 2325 1805 2355 1835
rect 2405 1805 2435 1835
rect 2485 1805 2515 1835
rect 2645 1805 2675 1835
rect 2725 1805 2755 1835
rect 2805 1805 2835 1835
rect 2885 1805 2915 1835
rect 2965 1805 2995 1835
rect 3045 1805 3075 1835
rect 3125 1805 3155 1835
rect 3205 1805 3235 1835
rect 3285 1805 3315 1835
rect 3365 1805 3395 1835
rect 3445 1805 3475 1835
rect 3605 1805 3635 1835
rect 3685 1805 3715 1835
rect 3765 1805 3795 1835
rect 3845 1805 3875 1835
rect 3925 1805 3955 1835
rect 4005 1805 4035 1835
rect 4085 1805 4115 1835
rect 4165 1805 4195 1835
rect 85 805 115 835
rect 245 805 275 835
rect 325 805 355 835
rect 405 805 435 835
rect 485 805 515 835
rect 565 805 595 835
rect 725 805 755 835
rect 805 805 835 835
rect 885 805 915 835
rect 965 805 995 835
rect 1045 805 1075 835
rect 1125 805 1155 835
rect 1205 805 1235 835
rect 1285 805 1315 835
rect 1365 805 1395 835
rect 1445 805 1475 835
rect 1525 805 1555 835
rect 1685 805 1715 835
rect 1765 805 1795 835
rect 1845 805 1875 835
rect 1925 805 1955 835
rect 2005 805 2035 835
rect 2165 805 2195 835
rect 2245 805 2275 835
rect 2325 805 2355 835
rect 2405 805 2435 835
rect 2485 805 2515 835
rect 2645 805 2675 835
rect 2725 805 2755 835
rect 2805 805 2835 835
rect 2885 805 2915 835
rect 2965 805 2995 835
rect 3045 805 3075 835
rect 3125 805 3155 835
rect 3205 805 3235 835
rect 3285 805 3315 835
rect 3365 805 3395 835
rect 3445 805 3475 835
rect 3605 805 3635 835
rect 3685 805 3715 835
rect 3765 805 3795 835
rect 3845 805 3875 835
rect 3925 805 3955 835
rect 4085 805 4115 835
rect 85 645 115 675
rect 245 645 275 675
rect 325 645 355 675
rect 405 645 435 675
rect 485 645 515 675
rect 565 645 595 675
rect 725 645 755 675
rect 805 645 835 675
rect 885 645 915 675
rect 965 645 995 675
rect 1045 645 1075 675
rect 1125 645 1155 675
rect 1205 645 1235 675
rect 1285 645 1315 675
rect 1365 645 1395 675
rect 1445 645 1475 675
rect 1525 645 1555 675
rect 1685 645 1715 675
rect 1765 645 1795 675
rect 1845 645 1875 675
rect 1925 645 1955 675
rect 2005 645 2035 675
rect 2165 645 2195 675
rect 2245 645 2275 675
rect 2325 645 2355 675
rect 2405 645 2435 675
rect 2485 645 2515 675
rect 2645 645 2675 675
rect 2725 645 2755 675
rect 2805 645 2835 675
rect 2885 645 2915 675
rect 2965 645 2995 675
rect 3045 645 3075 675
rect 3125 645 3155 675
rect 3205 645 3235 675
rect 3285 645 3315 675
rect 3365 645 3395 675
rect 3445 645 3475 675
rect 3605 645 3635 675
rect 3685 645 3715 675
rect 3765 645 3795 675
rect 3845 645 3875 675
rect 3925 645 3955 675
rect 4085 645 4115 675
rect 85 485 115 515
rect 245 485 275 515
rect 325 485 355 515
rect 405 485 435 515
rect 485 485 515 515
rect 565 485 595 515
rect 725 485 755 515
rect 805 485 835 515
rect 885 485 915 515
rect 965 485 995 515
rect 1045 485 1075 515
rect 1125 485 1155 515
rect 1205 485 1235 515
rect 1285 485 1315 515
rect 1365 485 1395 515
rect 1445 485 1475 515
rect 1525 485 1555 515
rect 1685 485 1715 515
rect 1765 485 1795 515
rect 1845 485 1875 515
rect 1925 485 1955 515
rect 2005 485 2035 515
rect 2165 485 2195 515
rect 2245 485 2275 515
rect 2325 485 2355 515
rect 2405 485 2435 515
rect 2485 485 2515 515
rect 2645 485 2675 515
rect 2725 485 2755 515
rect 2805 485 2835 515
rect 2885 485 2915 515
rect 2965 485 2995 515
rect 3045 485 3075 515
rect 3125 485 3155 515
rect 3205 485 3235 515
rect 3285 485 3315 515
rect 3365 485 3395 515
rect 3445 485 3475 515
rect 3605 485 3635 515
rect 3685 485 3715 515
rect 3765 485 3795 515
rect 3845 485 3875 515
rect 3925 485 3955 515
rect 4085 485 4115 515
rect 165 90 195 170
rect 4005 90 4035 170
<< metal3 >>
rect 2080 2831 2120 2840
rect 2080 2649 2084 2831
rect 2116 2649 2120 2831
rect 2080 2640 2120 2649
rect 0 1996 40 2000
rect 0 1964 4 1996
rect 36 1964 40 1996
rect 0 1836 40 1964
rect 0 1804 4 1836
rect 36 1804 40 1836
rect 0 1800 40 1804
rect 80 1996 120 2000
rect 80 1964 84 1996
rect 116 1964 120 1996
rect 80 1836 120 1964
rect 80 1804 84 1836
rect 116 1804 120 1836
rect 80 1800 120 1804
rect 160 1996 200 2000
rect 160 1964 164 1996
rect 196 1964 200 1996
rect 160 1836 200 1964
rect 160 1804 164 1836
rect 196 1804 200 1836
rect 160 1800 200 1804
rect 240 1996 280 2000
rect 240 1964 244 1996
rect 276 1964 280 1996
rect 240 1836 280 1964
rect 240 1804 244 1836
rect 276 1804 280 1836
rect 240 1800 280 1804
rect 320 1996 360 2000
rect 320 1964 324 1996
rect 356 1964 360 1996
rect 320 1836 360 1964
rect 320 1804 324 1836
rect 356 1804 360 1836
rect 320 1800 360 1804
rect 400 1996 440 2000
rect 400 1964 404 1996
rect 436 1964 440 1996
rect 400 1836 440 1964
rect 400 1804 404 1836
rect 436 1804 440 1836
rect 400 1800 440 1804
rect 480 1996 520 2000
rect 480 1964 484 1996
rect 516 1964 520 1996
rect 480 1836 520 1964
rect 480 1804 484 1836
rect 516 1804 520 1836
rect 480 1800 520 1804
rect 560 1996 600 2000
rect 560 1964 564 1996
rect 596 1964 600 1996
rect 560 1836 600 1964
rect 560 1804 564 1836
rect 596 1804 600 1836
rect 560 1800 600 1804
rect 720 1996 760 2000
rect 720 1964 724 1996
rect 756 1964 760 1996
rect 720 1836 760 1964
rect 720 1804 724 1836
rect 756 1804 760 1836
rect 720 1800 760 1804
rect 800 1996 840 2000
rect 800 1964 804 1996
rect 836 1964 840 1996
rect 800 1836 840 1964
rect 800 1804 804 1836
rect 836 1804 840 1836
rect 800 1800 840 1804
rect 880 1996 920 2000
rect 880 1964 884 1996
rect 916 1964 920 1996
rect 880 1836 920 1964
rect 880 1804 884 1836
rect 916 1804 920 1836
rect 880 1800 920 1804
rect 960 1996 1000 2000
rect 960 1964 964 1996
rect 996 1964 1000 1996
rect 960 1836 1000 1964
rect 960 1804 964 1836
rect 996 1804 1000 1836
rect 960 1800 1000 1804
rect 1040 1996 1080 2000
rect 1040 1964 1044 1996
rect 1076 1964 1080 1996
rect 1040 1836 1080 1964
rect 1040 1804 1044 1836
rect 1076 1804 1080 1836
rect 1040 1800 1080 1804
rect 1120 1996 1160 2000
rect 1120 1964 1124 1996
rect 1156 1964 1160 1996
rect 1120 1836 1160 1964
rect 1120 1804 1124 1836
rect 1156 1804 1160 1836
rect 1120 1800 1160 1804
rect 1200 1996 1240 2000
rect 1200 1964 1204 1996
rect 1236 1964 1240 1996
rect 1200 1836 1240 1964
rect 1200 1804 1204 1836
rect 1236 1804 1240 1836
rect 1200 1800 1240 1804
rect 1280 1996 1320 2000
rect 1280 1964 1284 1996
rect 1316 1964 1320 1996
rect 1280 1836 1320 1964
rect 1280 1804 1284 1836
rect 1316 1804 1320 1836
rect 1280 1800 1320 1804
rect 1360 1996 1400 2000
rect 1360 1964 1364 1996
rect 1396 1964 1400 1996
rect 1360 1836 1400 1964
rect 1360 1804 1364 1836
rect 1396 1804 1400 1836
rect 1360 1800 1400 1804
rect 1440 1996 1480 2000
rect 1440 1964 1444 1996
rect 1476 1964 1480 1996
rect 1440 1836 1480 1964
rect 1440 1804 1444 1836
rect 1476 1804 1480 1836
rect 1440 1800 1480 1804
rect 1520 1996 1560 2000
rect 1520 1964 1524 1996
rect 1556 1964 1560 1996
rect 1520 1836 1560 1964
rect 1520 1804 1524 1836
rect 1556 1804 1560 1836
rect 1520 1800 1560 1804
rect 1680 1996 1720 2000
rect 1680 1964 1684 1996
rect 1716 1964 1720 1996
rect 1680 1836 1720 1964
rect 1680 1804 1684 1836
rect 1716 1804 1720 1836
rect 1680 1800 1720 1804
rect 1760 1996 1800 2000
rect 1760 1964 1764 1996
rect 1796 1964 1800 1996
rect 1760 1836 1800 1964
rect 1760 1804 1764 1836
rect 1796 1804 1800 1836
rect 1760 1800 1800 1804
rect 1840 1996 1880 2000
rect 1840 1964 1844 1996
rect 1876 1964 1880 1996
rect 1840 1836 1880 1964
rect 1840 1804 1844 1836
rect 1876 1804 1880 1836
rect 1840 1800 1880 1804
rect 1920 1996 1960 2000
rect 1920 1964 1924 1996
rect 1956 1964 1960 1996
rect 1920 1836 1960 1964
rect 1920 1804 1924 1836
rect 1956 1804 1960 1836
rect 1920 1800 1960 1804
rect 2000 1996 2040 2000
rect 2000 1964 2004 1996
rect 2036 1964 2040 1996
rect 2000 1836 2040 1964
rect 2000 1804 2004 1836
rect 2036 1804 2040 1836
rect 2000 1800 2040 1804
rect 2080 1996 2120 2000
rect 2080 1964 2084 1996
rect 2116 1964 2120 1996
rect 2080 1836 2120 1964
rect 2080 1804 2084 1836
rect 2116 1804 2120 1836
rect 2080 1800 2120 1804
rect 2160 1996 2200 2000
rect 2160 1964 2164 1996
rect 2196 1964 2200 1996
rect 2160 1836 2200 1964
rect 2160 1804 2164 1836
rect 2196 1804 2200 1836
rect 2160 1800 2200 1804
rect 2240 1996 2280 2000
rect 2240 1964 2244 1996
rect 2276 1964 2280 1996
rect 2240 1836 2280 1964
rect 2240 1804 2244 1836
rect 2276 1804 2280 1836
rect 2240 1800 2280 1804
rect 2320 1996 2360 2000
rect 2320 1964 2324 1996
rect 2356 1964 2360 1996
rect 2320 1836 2360 1964
rect 2320 1804 2324 1836
rect 2356 1804 2360 1836
rect 2320 1800 2360 1804
rect 2400 1996 2440 2000
rect 2400 1964 2404 1996
rect 2436 1964 2440 1996
rect 2400 1836 2440 1964
rect 2400 1804 2404 1836
rect 2436 1804 2440 1836
rect 2400 1800 2440 1804
rect 2480 1996 2520 2000
rect 2480 1964 2484 1996
rect 2516 1964 2520 1996
rect 2480 1836 2520 1964
rect 2480 1804 2484 1836
rect 2516 1804 2520 1836
rect 2480 1800 2520 1804
rect 2640 1996 2680 2000
rect 2640 1964 2644 1996
rect 2676 1964 2680 1996
rect 2640 1836 2680 1964
rect 2640 1804 2644 1836
rect 2676 1804 2680 1836
rect 2640 1800 2680 1804
rect 2720 1996 2760 2000
rect 2720 1964 2724 1996
rect 2756 1964 2760 1996
rect 2720 1836 2760 1964
rect 2720 1804 2724 1836
rect 2756 1804 2760 1836
rect 2720 1800 2760 1804
rect 2800 1996 2840 2000
rect 2800 1964 2804 1996
rect 2836 1964 2840 1996
rect 2800 1836 2840 1964
rect 2800 1804 2804 1836
rect 2836 1804 2840 1836
rect 2800 1800 2840 1804
rect 2880 1996 2920 2000
rect 2880 1964 2884 1996
rect 2916 1964 2920 1996
rect 2880 1836 2920 1964
rect 2880 1804 2884 1836
rect 2916 1804 2920 1836
rect 2880 1800 2920 1804
rect 2960 1996 3000 2000
rect 2960 1964 2964 1996
rect 2996 1964 3000 1996
rect 2960 1836 3000 1964
rect 2960 1804 2964 1836
rect 2996 1804 3000 1836
rect 2960 1800 3000 1804
rect 3040 1996 3080 2000
rect 3040 1964 3044 1996
rect 3076 1964 3080 1996
rect 3040 1836 3080 1964
rect 3040 1804 3044 1836
rect 3076 1804 3080 1836
rect 3040 1800 3080 1804
rect 3120 1996 3160 2000
rect 3120 1964 3124 1996
rect 3156 1964 3160 1996
rect 3120 1836 3160 1964
rect 3120 1804 3124 1836
rect 3156 1804 3160 1836
rect 3120 1800 3160 1804
rect 3200 1996 3240 2000
rect 3200 1964 3204 1996
rect 3236 1964 3240 1996
rect 3200 1836 3240 1964
rect 3200 1804 3204 1836
rect 3236 1804 3240 1836
rect 3200 1800 3240 1804
rect 3280 1996 3320 2000
rect 3280 1964 3284 1996
rect 3316 1964 3320 1996
rect 3280 1836 3320 1964
rect 3280 1804 3284 1836
rect 3316 1804 3320 1836
rect 3280 1800 3320 1804
rect 3360 1996 3400 2000
rect 3360 1964 3364 1996
rect 3396 1964 3400 1996
rect 3360 1836 3400 1964
rect 3360 1804 3364 1836
rect 3396 1804 3400 1836
rect 3360 1800 3400 1804
rect 3440 1996 3480 2000
rect 3440 1964 3444 1996
rect 3476 1964 3480 1996
rect 3440 1836 3480 1964
rect 3440 1804 3444 1836
rect 3476 1804 3480 1836
rect 3440 1800 3480 1804
rect 3600 1996 3640 2000
rect 3600 1964 3604 1996
rect 3636 1964 3640 1996
rect 3600 1836 3640 1964
rect 3600 1804 3604 1836
rect 3636 1804 3640 1836
rect 3600 1800 3640 1804
rect 3680 1996 3720 2000
rect 3680 1964 3684 1996
rect 3716 1964 3720 1996
rect 3680 1836 3720 1964
rect 3680 1804 3684 1836
rect 3716 1804 3720 1836
rect 3680 1800 3720 1804
rect 3760 1996 3800 2000
rect 3760 1964 3764 1996
rect 3796 1964 3800 1996
rect 3760 1836 3800 1964
rect 3760 1804 3764 1836
rect 3796 1804 3800 1836
rect 3760 1800 3800 1804
rect 3840 1996 3880 2000
rect 3840 1964 3844 1996
rect 3876 1964 3880 1996
rect 3840 1836 3880 1964
rect 3840 1804 3844 1836
rect 3876 1804 3880 1836
rect 3840 1800 3880 1804
rect 3920 1996 3960 2000
rect 3920 1964 3924 1996
rect 3956 1964 3960 1996
rect 3920 1836 3960 1964
rect 3920 1804 3924 1836
rect 3956 1804 3960 1836
rect 3920 1800 3960 1804
rect 4000 1996 4040 2000
rect 4000 1964 4004 1996
rect 4036 1964 4040 1996
rect 4000 1836 4040 1964
rect 4000 1804 4004 1836
rect 4036 1804 4040 1836
rect 4000 1800 4040 1804
rect 4080 1996 4120 2000
rect 4080 1964 4084 1996
rect 4116 1964 4120 1996
rect 4080 1836 4120 1964
rect 4080 1804 4084 1836
rect 4116 1804 4120 1836
rect 4080 1800 4120 1804
rect 4160 1996 4200 2000
rect 4160 1964 4164 1996
rect 4196 1964 4200 1996
rect 4160 1836 4200 1964
rect 4160 1804 4164 1836
rect 4196 1804 4200 1836
rect 4160 1800 4200 1804
rect 80 835 120 840
rect 80 805 85 835
rect 115 805 120 835
rect 80 676 120 805
rect 80 644 84 676
rect 116 644 120 676
rect 80 515 120 644
rect 80 485 85 515
rect 115 485 120 515
rect 80 480 120 485
rect 240 835 280 840
rect 240 805 245 835
rect 275 805 280 835
rect 240 675 280 805
rect 240 645 245 675
rect 275 645 280 675
rect 240 515 280 645
rect 240 485 245 515
rect 275 485 280 515
rect 240 480 280 485
rect 320 835 360 840
rect 320 805 325 835
rect 355 805 360 835
rect 320 675 360 805
rect 320 645 325 675
rect 355 645 360 675
rect 320 515 360 645
rect 320 485 325 515
rect 355 485 360 515
rect 320 480 360 485
rect 400 835 440 840
rect 400 805 405 835
rect 435 805 440 835
rect 400 675 440 805
rect 400 645 405 675
rect 435 645 440 675
rect 400 515 440 645
rect 400 485 405 515
rect 435 485 440 515
rect 400 480 440 485
rect 480 835 520 840
rect 480 805 485 835
rect 515 805 520 835
rect 480 675 520 805
rect 480 645 485 675
rect 515 645 520 675
rect 480 515 520 645
rect 480 485 485 515
rect 515 485 520 515
rect 480 480 520 485
rect 560 835 600 840
rect 560 805 565 835
rect 595 805 600 835
rect 560 675 600 805
rect 560 645 565 675
rect 595 645 600 675
rect 560 515 600 645
rect 560 485 565 515
rect 595 485 600 515
rect 560 480 600 485
rect 720 835 760 840
rect 720 805 725 835
rect 755 805 760 835
rect 720 675 760 805
rect 720 645 725 675
rect 755 645 760 675
rect 720 515 760 645
rect 720 485 725 515
rect 755 485 760 515
rect 720 480 760 485
rect 800 835 840 840
rect 800 805 805 835
rect 835 805 840 835
rect 800 675 840 805
rect 800 645 805 675
rect 835 645 840 675
rect 800 515 840 645
rect 800 485 805 515
rect 835 485 840 515
rect 800 480 840 485
rect 880 835 920 840
rect 880 805 885 835
rect 915 805 920 835
rect 880 675 920 805
rect 880 645 885 675
rect 915 645 920 675
rect 880 515 920 645
rect 880 485 885 515
rect 915 485 920 515
rect 880 480 920 485
rect 960 835 1000 840
rect 960 805 965 835
rect 995 805 1000 835
rect 960 675 1000 805
rect 960 645 965 675
rect 995 645 1000 675
rect 960 515 1000 645
rect 960 485 965 515
rect 995 485 1000 515
rect 960 480 1000 485
rect 1040 835 1080 840
rect 1040 805 1045 835
rect 1075 805 1080 835
rect 1040 675 1080 805
rect 1040 645 1045 675
rect 1075 645 1080 675
rect 1040 515 1080 645
rect 1040 485 1045 515
rect 1075 485 1080 515
rect 1040 480 1080 485
rect 1120 835 1160 840
rect 1120 805 1125 835
rect 1155 805 1160 835
rect 1120 675 1160 805
rect 1120 645 1125 675
rect 1155 645 1160 675
rect 1120 515 1160 645
rect 1120 485 1125 515
rect 1155 485 1160 515
rect 1120 480 1160 485
rect 1200 835 1240 840
rect 1200 805 1205 835
rect 1235 805 1240 835
rect 1200 675 1240 805
rect 1200 645 1205 675
rect 1235 645 1240 675
rect 1200 515 1240 645
rect 1200 485 1205 515
rect 1235 485 1240 515
rect 1200 480 1240 485
rect 1280 835 1320 840
rect 1280 805 1285 835
rect 1315 805 1320 835
rect 1280 675 1320 805
rect 1280 645 1285 675
rect 1315 645 1320 675
rect 1280 515 1320 645
rect 1280 485 1285 515
rect 1315 485 1320 515
rect 1280 480 1320 485
rect 1360 835 1400 840
rect 1360 805 1365 835
rect 1395 805 1400 835
rect 1360 675 1400 805
rect 1360 645 1365 675
rect 1395 645 1400 675
rect 1360 515 1400 645
rect 1360 485 1365 515
rect 1395 485 1400 515
rect 1360 480 1400 485
rect 1440 835 1480 840
rect 1440 805 1445 835
rect 1475 805 1480 835
rect 1440 675 1480 805
rect 1440 645 1445 675
rect 1475 645 1480 675
rect 1440 515 1480 645
rect 1440 485 1445 515
rect 1475 485 1480 515
rect 1440 480 1480 485
rect 1520 835 1560 840
rect 1520 805 1525 835
rect 1555 805 1560 835
rect 1520 675 1560 805
rect 1520 645 1525 675
rect 1555 645 1560 675
rect 1520 515 1560 645
rect 1520 485 1525 515
rect 1555 485 1560 515
rect 1520 480 1560 485
rect 1680 835 1720 840
rect 1680 805 1685 835
rect 1715 805 1720 835
rect 1680 675 1720 805
rect 1680 645 1685 675
rect 1715 645 1720 675
rect 1680 515 1720 645
rect 1680 485 1685 515
rect 1715 485 1720 515
rect 1680 480 1720 485
rect 1760 835 1800 840
rect 1760 805 1765 835
rect 1795 805 1800 835
rect 1760 675 1800 805
rect 1760 645 1765 675
rect 1795 645 1800 675
rect 1760 515 1800 645
rect 1760 485 1765 515
rect 1795 485 1800 515
rect 1760 480 1800 485
rect 1840 835 1880 840
rect 1840 805 1845 835
rect 1875 805 1880 835
rect 1840 675 1880 805
rect 1840 645 1845 675
rect 1875 645 1880 675
rect 1840 515 1880 645
rect 1840 485 1845 515
rect 1875 485 1880 515
rect 1840 480 1880 485
rect 1920 835 1960 840
rect 1920 805 1925 835
rect 1955 805 1960 835
rect 1920 675 1960 805
rect 1920 645 1925 675
rect 1955 645 1960 675
rect 1920 515 1960 645
rect 1920 485 1925 515
rect 1955 485 1960 515
rect 1920 480 1960 485
rect 2000 835 2040 840
rect 2000 805 2005 835
rect 2035 805 2040 835
rect 2000 675 2040 805
rect 2000 645 2005 675
rect 2035 645 2040 675
rect 2000 515 2040 645
rect 2000 485 2005 515
rect 2035 485 2040 515
rect 2000 480 2040 485
rect 2160 835 2200 840
rect 2160 805 2165 835
rect 2195 805 2200 835
rect 2160 675 2200 805
rect 2160 645 2165 675
rect 2195 645 2200 675
rect 2160 515 2200 645
rect 2160 485 2165 515
rect 2195 485 2200 515
rect 2160 480 2200 485
rect 2240 835 2280 840
rect 2240 805 2245 835
rect 2275 805 2280 835
rect 2240 675 2280 805
rect 2240 645 2245 675
rect 2275 645 2280 675
rect 2240 515 2280 645
rect 2240 485 2245 515
rect 2275 485 2280 515
rect 2240 480 2280 485
rect 2320 835 2360 840
rect 2320 805 2325 835
rect 2355 805 2360 835
rect 2320 675 2360 805
rect 2320 645 2325 675
rect 2355 645 2360 675
rect 2320 515 2360 645
rect 2320 485 2325 515
rect 2355 485 2360 515
rect 2320 480 2360 485
rect 2400 835 2440 840
rect 2400 805 2405 835
rect 2435 805 2440 835
rect 2400 675 2440 805
rect 2400 645 2405 675
rect 2435 645 2440 675
rect 2400 515 2440 645
rect 2400 485 2405 515
rect 2435 485 2440 515
rect 2400 480 2440 485
rect 2480 835 2520 840
rect 2480 805 2485 835
rect 2515 805 2520 835
rect 2480 675 2520 805
rect 2480 645 2485 675
rect 2515 645 2520 675
rect 2480 515 2520 645
rect 2480 485 2485 515
rect 2515 485 2520 515
rect 2480 480 2520 485
rect 2640 835 2680 840
rect 2640 805 2645 835
rect 2675 805 2680 835
rect 2640 675 2680 805
rect 2640 645 2645 675
rect 2675 645 2680 675
rect 2640 515 2680 645
rect 2640 485 2645 515
rect 2675 485 2680 515
rect 2640 480 2680 485
rect 2720 835 2760 840
rect 2720 805 2725 835
rect 2755 805 2760 835
rect 2720 675 2760 805
rect 2720 645 2725 675
rect 2755 645 2760 675
rect 2720 515 2760 645
rect 2720 485 2725 515
rect 2755 485 2760 515
rect 2720 480 2760 485
rect 2800 835 2840 840
rect 2800 805 2805 835
rect 2835 805 2840 835
rect 2800 675 2840 805
rect 2800 645 2805 675
rect 2835 645 2840 675
rect 2800 515 2840 645
rect 2800 485 2805 515
rect 2835 485 2840 515
rect 2800 480 2840 485
rect 2880 835 2920 840
rect 2880 805 2885 835
rect 2915 805 2920 835
rect 2880 675 2920 805
rect 2880 645 2885 675
rect 2915 645 2920 675
rect 2880 515 2920 645
rect 2880 485 2885 515
rect 2915 485 2920 515
rect 2880 480 2920 485
rect 2960 835 3000 840
rect 2960 805 2965 835
rect 2995 805 3000 835
rect 2960 675 3000 805
rect 2960 645 2965 675
rect 2995 645 3000 675
rect 2960 515 3000 645
rect 2960 485 2965 515
rect 2995 485 3000 515
rect 2960 480 3000 485
rect 3040 835 3080 840
rect 3040 805 3045 835
rect 3075 805 3080 835
rect 3040 675 3080 805
rect 3040 645 3045 675
rect 3075 645 3080 675
rect 3040 515 3080 645
rect 3040 485 3045 515
rect 3075 485 3080 515
rect 3040 480 3080 485
rect 3120 835 3160 840
rect 3120 805 3125 835
rect 3155 805 3160 835
rect 3120 675 3160 805
rect 3120 645 3125 675
rect 3155 645 3160 675
rect 3120 515 3160 645
rect 3120 485 3125 515
rect 3155 485 3160 515
rect 3120 480 3160 485
rect 3200 835 3240 840
rect 3200 805 3205 835
rect 3235 805 3240 835
rect 3200 675 3240 805
rect 3200 645 3205 675
rect 3235 645 3240 675
rect 3200 515 3240 645
rect 3200 485 3205 515
rect 3235 485 3240 515
rect 3200 480 3240 485
rect 3280 835 3320 840
rect 3280 805 3285 835
rect 3315 805 3320 835
rect 3280 675 3320 805
rect 3280 645 3285 675
rect 3315 645 3320 675
rect 3280 515 3320 645
rect 3280 485 3285 515
rect 3315 485 3320 515
rect 3280 480 3320 485
rect 3360 835 3400 840
rect 3360 805 3365 835
rect 3395 805 3400 835
rect 3360 675 3400 805
rect 3360 645 3365 675
rect 3395 645 3400 675
rect 3360 515 3400 645
rect 3360 485 3365 515
rect 3395 485 3400 515
rect 3360 480 3400 485
rect 3440 835 3480 840
rect 3440 805 3445 835
rect 3475 805 3480 835
rect 3440 675 3480 805
rect 3440 645 3445 675
rect 3475 645 3480 675
rect 3440 515 3480 645
rect 3440 485 3445 515
rect 3475 485 3480 515
rect 3440 480 3480 485
rect 3600 835 3640 840
rect 3600 805 3605 835
rect 3635 805 3640 835
rect 3600 675 3640 805
rect 3600 645 3605 675
rect 3635 645 3640 675
rect 3600 515 3640 645
rect 3600 485 3605 515
rect 3635 485 3640 515
rect 3600 480 3640 485
rect 3680 835 3720 840
rect 3680 805 3685 835
rect 3715 805 3720 835
rect 3680 675 3720 805
rect 3680 645 3685 675
rect 3715 645 3720 675
rect 3680 515 3720 645
rect 3680 485 3685 515
rect 3715 485 3720 515
rect 3680 480 3720 485
rect 3760 835 3800 840
rect 3760 805 3765 835
rect 3795 805 3800 835
rect 3760 675 3800 805
rect 3760 645 3765 675
rect 3795 645 3800 675
rect 3760 515 3800 645
rect 3760 485 3765 515
rect 3795 485 3800 515
rect 3760 480 3800 485
rect 3840 835 3880 840
rect 3840 805 3845 835
rect 3875 805 3880 835
rect 3840 675 3880 805
rect 3840 645 3845 675
rect 3875 645 3880 675
rect 3840 515 3880 645
rect 3840 485 3845 515
rect 3875 485 3880 515
rect 3840 480 3880 485
rect 3920 835 3960 840
rect 3920 805 3925 835
rect 3955 805 3960 835
rect 3920 675 3960 805
rect 3920 645 3925 675
rect 3955 645 3960 675
rect 3920 515 3960 645
rect 3920 485 3925 515
rect 3955 485 3960 515
rect 3920 480 3960 485
rect 4080 835 4120 840
rect 4080 805 4085 835
rect 4115 805 4120 835
rect 4080 675 4120 805
rect 4080 645 4085 675
rect 4115 645 4120 675
rect 4080 515 4120 645
rect 4080 485 4085 515
rect 4115 485 4120 515
rect 4080 480 4120 485
rect 160 171 200 180
rect 160 89 164 171
rect 196 89 200 171
rect 160 80 200 89
rect 4000 171 4040 180
rect 4000 89 4004 171
rect 4036 89 4040 171
rect 4000 80 4040 89
<< via3 >>
rect 2084 2830 2116 2831
rect 2084 2650 2085 2830
rect 2085 2650 2115 2830
rect 2115 2650 2116 2830
rect 2084 2649 2116 2650
rect 4 1995 36 1996
rect 4 1965 5 1995
rect 5 1965 35 1995
rect 35 1965 36 1995
rect 4 1964 36 1965
rect 4 1835 36 1836
rect 4 1805 5 1835
rect 5 1805 35 1835
rect 35 1805 36 1835
rect 4 1804 36 1805
rect 84 1995 116 1996
rect 84 1965 85 1995
rect 85 1965 115 1995
rect 115 1965 116 1995
rect 84 1964 116 1965
rect 84 1835 116 1836
rect 84 1805 85 1835
rect 85 1805 115 1835
rect 115 1805 116 1835
rect 84 1804 116 1805
rect 164 1995 196 1996
rect 164 1965 165 1995
rect 165 1965 195 1995
rect 195 1965 196 1995
rect 164 1964 196 1965
rect 164 1835 196 1836
rect 164 1805 165 1835
rect 165 1805 195 1835
rect 195 1805 196 1835
rect 164 1804 196 1805
rect 244 1995 276 1996
rect 244 1965 245 1995
rect 245 1965 275 1995
rect 275 1965 276 1995
rect 244 1964 276 1965
rect 244 1835 276 1836
rect 244 1805 245 1835
rect 245 1805 275 1835
rect 275 1805 276 1835
rect 244 1804 276 1805
rect 324 1995 356 1996
rect 324 1965 325 1995
rect 325 1965 355 1995
rect 355 1965 356 1995
rect 324 1964 356 1965
rect 324 1835 356 1836
rect 324 1805 325 1835
rect 325 1805 355 1835
rect 355 1805 356 1835
rect 324 1804 356 1805
rect 404 1995 436 1996
rect 404 1965 405 1995
rect 405 1965 435 1995
rect 435 1965 436 1995
rect 404 1964 436 1965
rect 404 1835 436 1836
rect 404 1805 405 1835
rect 405 1805 435 1835
rect 435 1805 436 1835
rect 404 1804 436 1805
rect 484 1995 516 1996
rect 484 1965 485 1995
rect 485 1965 515 1995
rect 515 1965 516 1995
rect 484 1964 516 1965
rect 484 1835 516 1836
rect 484 1805 485 1835
rect 485 1805 515 1835
rect 515 1805 516 1835
rect 484 1804 516 1805
rect 564 1995 596 1996
rect 564 1965 565 1995
rect 565 1965 595 1995
rect 595 1965 596 1995
rect 564 1964 596 1965
rect 564 1835 596 1836
rect 564 1805 565 1835
rect 565 1805 595 1835
rect 595 1805 596 1835
rect 564 1804 596 1805
rect 724 1995 756 1996
rect 724 1965 725 1995
rect 725 1965 755 1995
rect 755 1965 756 1995
rect 724 1964 756 1965
rect 724 1835 756 1836
rect 724 1805 725 1835
rect 725 1805 755 1835
rect 755 1805 756 1835
rect 724 1804 756 1805
rect 804 1995 836 1996
rect 804 1965 805 1995
rect 805 1965 835 1995
rect 835 1965 836 1995
rect 804 1964 836 1965
rect 804 1835 836 1836
rect 804 1805 805 1835
rect 805 1805 835 1835
rect 835 1805 836 1835
rect 804 1804 836 1805
rect 884 1995 916 1996
rect 884 1965 885 1995
rect 885 1965 915 1995
rect 915 1965 916 1995
rect 884 1964 916 1965
rect 884 1835 916 1836
rect 884 1805 885 1835
rect 885 1805 915 1835
rect 915 1805 916 1835
rect 884 1804 916 1805
rect 964 1995 996 1996
rect 964 1965 965 1995
rect 965 1965 995 1995
rect 995 1965 996 1995
rect 964 1964 996 1965
rect 964 1835 996 1836
rect 964 1805 965 1835
rect 965 1805 995 1835
rect 995 1805 996 1835
rect 964 1804 996 1805
rect 1044 1995 1076 1996
rect 1044 1965 1045 1995
rect 1045 1965 1075 1995
rect 1075 1965 1076 1995
rect 1044 1964 1076 1965
rect 1044 1835 1076 1836
rect 1044 1805 1045 1835
rect 1045 1805 1075 1835
rect 1075 1805 1076 1835
rect 1044 1804 1076 1805
rect 1124 1995 1156 1996
rect 1124 1965 1125 1995
rect 1125 1965 1155 1995
rect 1155 1965 1156 1995
rect 1124 1964 1156 1965
rect 1124 1835 1156 1836
rect 1124 1805 1125 1835
rect 1125 1805 1155 1835
rect 1155 1805 1156 1835
rect 1124 1804 1156 1805
rect 1204 1995 1236 1996
rect 1204 1965 1205 1995
rect 1205 1965 1235 1995
rect 1235 1965 1236 1995
rect 1204 1964 1236 1965
rect 1204 1835 1236 1836
rect 1204 1805 1205 1835
rect 1205 1805 1235 1835
rect 1235 1805 1236 1835
rect 1204 1804 1236 1805
rect 1284 1995 1316 1996
rect 1284 1965 1285 1995
rect 1285 1965 1315 1995
rect 1315 1965 1316 1995
rect 1284 1964 1316 1965
rect 1284 1835 1316 1836
rect 1284 1805 1285 1835
rect 1285 1805 1315 1835
rect 1315 1805 1316 1835
rect 1284 1804 1316 1805
rect 1364 1995 1396 1996
rect 1364 1965 1365 1995
rect 1365 1965 1395 1995
rect 1395 1965 1396 1995
rect 1364 1964 1396 1965
rect 1364 1835 1396 1836
rect 1364 1805 1365 1835
rect 1365 1805 1395 1835
rect 1395 1805 1396 1835
rect 1364 1804 1396 1805
rect 1444 1995 1476 1996
rect 1444 1965 1445 1995
rect 1445 1965 1475 1995
rect 1475 1965 1476 1995
rect 1444 1964 1476 1965
rect 1444 1835 1476 1836
rect 1444 1805 1445 1835
rect 1445 1805 1475 1835
rect 1475 1805 1476 1835
rect 1444 1804 1476 1805
rect 1524 1995 1556 1996
rect 1524 1965 1525 1995
rect 1525 1965 1555 1995
rect 1555 1965 1556 1995
rect 1524 1964 1556 1965
rect 1524 1835 1556 1836
rect 1524 1805 1525 1835
rect 1525 1805 1555 1835
rect 1555 1805 1556 1835
rect 1524 1804 1556 1805
rect 1684 1995 1716 1996
rect 1684 1965 1685 1995
rect 1685 1965 1715 1995
rect 1715 1965 1716 1995
rect 1684 1964 1716 1965
rect 1684 1835 1716 1836
rect 1684 1805 1685 1835
rect 1685 1805 1715 1835
rect 1715 1805 1716 1835
rect 1684 1804 1716 1805
rect 1764 1995 1796 1996
rect 1764 1965 1765 1995
rect 1765 1965 1795 1995
rect 1795 1965 1796 1995
rect 1764 1964 1796 1965
rect 1764 1835 1796 1836
rect 1764 1805 1765 1835
rect 1765 1805 1795 1835
rect 1795 1805 1796 1835
rect 1764 1804 1796 1805
rect 1844 1995 1876 1996
rect 1844 1965 1845 1995
rect 1845 1965 1875 1995
rect 1875 1965 1876 1995
rect 1844 1964 1876 1965
rect 1844 1835 1876 1836
rect 1844 1805 1845 1835
rect 1845 1805 1875 1835
rect 1875 1805 1876 1835
rect 1844 1804 1876 1805
rect 1924 1995 1956 1996
rect 1924 1965 1925 1995
rect 1925 1965 1955 1995
rect 1955 1965 1956 1995
rect 1924 1964 1956 1965
rect 1924 1835 1956 1836
rect 1924 1805 1925 1835
rect 1925 1805 1955 1835
rect 1955 1805 1956 1835
rect 1924 1804 1956 1805
rect 2004 1995 2036 1996
rect 2004 1965 2005 1995
rect 2005 1965 2035 1995
rect 2035 1965 2036 1995
rect 2004 1964 2036 1965
rect 2004 1835 2036 1836
rect 2004 1805 2005 1835
rect 2005 1805 2035 1835
rect 2035 1805 2036 1835
rect 2004 1804 2036 1805
rect 2084 1995 2116 1996
rect 2084 1965 2085 1995
rect 2085 1965 2115 1995
rect 2115 1965 2116 1995
rect 2084 1964 2116 1965
rect 2084 1835 2116 1836
rect 2084 1805 2085 1835
rect 2085 1805 2115 1835
rect 2115 1805 2116 1835
rect 2084 1804 2116 1805
rect 2164 1995 2196 1996
rect 2164 1965 2165 1995
rect 2165 1965 2195 1995
rect 2195 1965 2196 1995
rect 2164 1964 2196 1965
rect 2164 1835 2196 1836
rect 2164 1805 2165 1835
rect 2165 1805 2195 1835
rect 2195 1805 2196 1835
rect 2164 1804 2196 1805
rect 2244 1995 2276 1996
rect 2244 1965 2245 1995
rect 2245 1965 2275 1995
rect 2275 1965 2276 1995
rect 2244 1964 2276 1965
rect 2244 1835 2276 1836
rect 2244 1805 2245 1835
rect 2245 1805 2275 1835
rect 2275 1805 2276 1835
rect 2244 1804 2276 1805
rect 2324 1995 2356 1996
rect 2324 1965 2325 1995
rect 2325 1965 2355 1995
rect 2355 1965 2356 1995
rect 2324 1964 2356 1965
rect 2324 1835 2356 1836
rect 2324 1805 2325 1835
rect 2325 1805 2355 1835
rect 2355 1805 2356 1835
rect 2324 1804 2356 1805
rect 2404 1995 2436 1996
rect 2404 1965 2405 1995
rect 2405 1965 2435 1995
rect 2435 1965 2436 1995
rect 2404 1964 2436 1965
rect 2404 1835 2436 1836
rect 2404 1805 2405 1835
rect 2405 1805 2435 1835
rect 2435 1805 2436 1835
rect 2404 1804 2436 1805
rect 2484 1995 2516 1996
rect 2484 1965 2485 1995
rect 2485 1965 2515 1995
rect 2515 1965 2516 1995
rect 2484 1964 2516 1965
rect 2484 1835 2516 1836
rect 2484 1805 2485 1835
rect 2485 1805 2515 1835
rect 2515 1805 2516 1835
rect 2484 1804 2516 1805
rect 2644 1995 2676 1996
rect 2644 1965 2645 1995
rect 2645 1965 2675 1995
rect 2675 1965 2676 1995
rect 2644 1964 2676 1965
rect 2644 1835 2676 1836
rect 2644 1805 2645 1835
rect 2645 1805 2675 1835
rect 2675 1805 2676 1835
rect 2644 1804 2676 1805
rect 2724 1995 2756 1996
rect 2724 1965 2725 1995
rect 2725 1965 2755 1995
rect 2755 1965 2756 1995
rect 2724 1964 2756 1965
rect 2724 1835 2756 1836
rect 2724 1805 2725 1835
rect 2725 1805 2755 1835
rect 2755 1805 2756 1835
rect 2724 1804 2756 1805
rect 2804 1995 2836 1996
rect 2804 1965 2805 1995
rect 2805 1965 2835 1995
rect 2835 1965 2836 1995
rect 2804 1964 2836 1965
rect 2804 1835 2836 1836
rect 2804 1805 2805 1835
rect 2805 1805 2835 1835
rect 2835 1805 2836 1835
rect 2804 1804 2836 1805
rect 2884 1995 2916 1996
rect 2884 1965 2885 1995
rect 2885 1965 2915 1995
rect 2915 1965 2916 1995
rect 2884 1964 2916 1965
rect 2884 1835 2916 1836
rect 2884 1805 2885 1835
rect 2885 1805 2915 1835
rect 2915 1805 2916 1835
rect 2884 1804 2916 1805
rect 2964 1995 2996 1996
rect 2964 1965 2965 1995
rect 2965 1965 2995 1995
rect 2995 1965 2996 1995
rect 2964 1964 2996 1965
rect 2964 1835 2996 1836
rect 2964 1805 2965 1835
rect 2965 1805 2995 1835
rect 2995 1805 2996 1835
rect 2964 1804 2996 1805
rect 3044 1995 3076 1996
rect 3044 1965 3045 1995
rect 3045 1965 3075 1995
rect 3075 1965 3076 1995
rect 3044 1964 3076 1965
rect 3044 1835 3076 1836
rect 3044 1805 3045 1835
rect 3045 1805 3075 1835
rect 3075 1805 3076 1835
rect 3044 1804 3076 1805
rect 3124 1995 3156 1996
rect 3124 1965 3125 1995
rect 3125 1965 3155 1995
rect 3155 1965 3156 1995
rect 3124 1964 3156 1965
rect 3124 1835 3156 1836
rect 3124 1805 3125 1835
rect 3125 1805 3155 1835
rect 3155 1805 3156 1835
rect 3124 1804 3156 1805
rect 3204 1995 3236 1996
rect 3204 1965 3205 1995
rect 3205 1965 3235 1995
rect 3235 1965 3236 1995
rect 3204 1964 3236 1965
rect 3204 1835 3236 1836
rect 3204 1805 3205 1835
rect 3205 1805 3235 1835
rect 3235 1805 3236 1835
rect 3204 1804 3236 1805
rect 3284 1995 3316 1996
rect 3284 1965 3285 1995
rect 3285 1965 3315 1995
rect 3315 1965 3316 1995
rect 3284 1964 3316 1965
rect 3284 1835 3316 1836
rect 3284 1805 3285 1835
rect 3285 1805 3315 1835
rect 3315 1805 3316 1835
rect 3284 1804 3316 1805
rect 3364 1995 3396 1996
rect 3364 1965 3365 1995
rect 3365 1965 3395 1995
rect 3395 1965 3396 1995
rect 3364 1964 3396 1965
rect 3364 1835 3396 1836
rect 3364 1805 3365 1835
rect 3365 1805 3395 1835
rect 3395 1805 3396 1835
rect 3364 1804 3396 1805
rect 3444 1995 3476 1996
rect 3444 1965 3445 1995
rect 3445 1965 3475 1995
rect 3475 1965 3476 1995
rect 3444 1964 3476 1965
rect 3444 1835 3476 1836
rect 3444 1805 3445 1835
rect 3445 1805 3475 1835
rect 3475 1805 3476 1835
rect 3444 1804 3476 1805
rect 3604 1995 3636 1996
rect 3604 1965 3605 1995
rect 3605 1965 3635 1995
rect 3635 1965 3636 1995
rect 3604 1964 3636 1965
rect 3604 1835 3636 1836
rect 3604 1805 3605 1835
rect 3605 1805 3635 1835
rect 3635 1805 3636 1835
rect 3604 1804 3636 1805
rect 3684 1995 3716 1996
rect 3684 1965 3685 1995
rect 3685 1965 3715 1995
rect 3715 1965 3716 1995
rect 3684 1964 3716 1965
rect 3684 1835 3716 1836
rect 3684 1805 3685 1835
rect 3685 1805 3715 1835
rect 3715 1805 3716 1835
rect 3684 1804 3716 1805
rect 3764 1995 3796 1996
rect 3764 1965 3765 1995
rect 3765 1965 3795 1995
rect 3795 1965 3796 1995
rect 3764 1964 3796 1965
rect 3764 1835 3796 1836
rect 3764 1805 3765 1835
rect 3765 1805 3795 1835
rect 3795 1805 3796 1835
rect 3764 1804 3796 1805
rect 3844 1995 3876 1996
rect 3844 1965 3845 1995
rect 3845 1965 3875 1995
rect 3875 1965 3876 1995
rect 3844 1964 3876 1965
rect 3844 1835 3876 1836
rect 3844 1805 3845 1835
rect 3845 1805 3875 1835
rect 3875 1805 3876 1835
rect 3844 1804 3876 1805
rect 3924 1995 3956 1996
rect 3924 1965 3925 1995
rect 3925 1965 3955 1995
rect 3955 1965 3956 1995
rect 3924 1964 3956 1965
rect 3924 1835 3956 1836
rect 3924 1805 3925 1835
rect 3925 1805 3955 1835
rect 3955 1805 3956 1835
rect 3924 1804 3956 1805
rect 4004 1995 4036 1996
rect 4004 1965 4005 1995
rect 4005 1965 4035 1995
rect 4035 1965 4036 1995
rect 4004 1964 4036 1965
rect 4004 1835 4036 1836
rect 4004 1805 4005 1835
rect 4005 1805 4035 1835
rect 4035 1805 4036 1835
rect 4004 1804 4036 1805
rect 4084 1995 4116 1996
rect 4084 1965 4085 1995
rect 4085 1965 4115 1995
rect 4115 1965 4116 1995
rect 4084 1964 4116 1965
rect 4084 1835 4116 1836
rect 4084 1805 4085 1835
rect 4085 1805 4115 1835
rect 4115 1805 4116 1835
rect 4084 1804 4116 1805
rect 4164 1995 4196 1996
rect 4164 1965 4165 1995
rect 4165 1965 4195 1995
rect 4195 1965 4196 1995
rect 4164 1964 4196 1965
rect 4164 1835 4196 1836
rect 4164 1805 4165 1835
rect 4165 1805 4195 1835
rect 4195 1805 4196 1835
rect 4164 1804 4196 1805
rect 84 675 116 676
rect 84 645 85 675
rect 85 645 115 675
rect 115 645 116 675
rect 84 644 116 645
rect 164 170 196 171
rect 164 90 165 170
rect 165 90 195 170
rect 195 90 196 170
rect 164 89 196 90
rect 4004 170 4036 171
rect 4004 90 4005 170
rect 4005 90 4035 170
rect 4035 90 4036 170
rect 4004 89 4036 90
<< metal4 >>
rect 0 2831 4200 2840
rect 0 2800 2084 2831
rect 0 2680 120 2800
rect 240 2680 2084 2800
rect 0 2649 2084 2680
rect 2116 2800 4200 2831
rect 2116 2680 3960 2800
rect 4080 2680 4200 2800
rect 2116 2649 4200 2680
rect 0 2640 4200 2649
rect 0 1996 4200 2000
rect 0 1964 4 1996
rect 36 1964 84 1996
rect 116 1964 164 1996
rect 196 1964 244 1996
rect 276 1964 324 1996
rect 356 1964 404 1996
rect 436 1964 484 1996
rect 516 1964 564 1996
rect 596 1964 724 1996
rect 756 1964 804 1996
rect 836 1964 884 1996
rect 916 1964 964 1996
rect 996 1964 1044 1996
rect 1076 1964 1124 1996
rect 1156 1964 1204 1996
rect 1236 1964 1284 1996
rect 1316 1964 1364 1996
rect 1396 1964 1444 1996
rect 1476 1964 1524 1996
rect 1556 1964 1684 1996
rect 1716 1964 1764 1996
rect 1796 1964 1844 1996
rect 1876 1964 1924 1996
rect 1956 1964 2004 1996
rect 2036 1964 2084 1996
rect 2116 1964 2164 1996
rect 2196 1964 2244 1996
rect 2276 1964 2324 1996
rect 2356 1964 2404 1996
rect 2436 1964 2484 1996
rect 2516 1964 2644 1996
rect 2676 1964 2724 1996
rect 2756 1964 2804 1996
rect 2836 1964 2884 1996
rect 2916 1964 2964 1996
rect 2996 1964 3044 1996
rect 3076 1964 3124 1996
rect 3156 1964 3204 1996
rect 3236 1964 3284 1996
rect 3316 1964 3364 1996
rect 3396 1964 3444 1996
rect 3476 1964 3604 1996
rect 3636 1964 3684 1996
rect 3716 1964 3764 1996
rect 3796 1964 3844 1996
rect 3876 1964 3924 1996
rect 3956 1964 4004 1996
rect 4036 1964 4084 1996
rect 4116 1964 4164 1996
rect 4196 1964 4200 1996
rect 0 1960 4200 1964
rect 0 1840 600 1960
rect 720 1840 3480 1960
rect 3600 1840 4200 1960
rect 0 1836 4200 1840
rect 0 1804 4 1836
rect 36 1804 84 1836
rect 116 1804 164 1836
rect 196 1804 244 1836
rect 276 1804 324 1836
rect 356 1804 404 1836
rect 436 1804 484 1836
rect 516 1804 564 1836
rect 596 1804 724 1836
rect 756 1804 804 1836
rect 836 1804 884 1836
rect 916 1804 964 1836
rect 996 1804 1044 1836
rect 1076 1804 1124 1836
rect 1156 1804 1204 1836
rect 1236 1804 1284 1836
rect 1316 1804 1364 1836
rect 1396 1804 1444 1836
rect 1476 1804 1524 1836
rect 1556 1804 1684 1836
rect 1716 1804 1764 1836
rect 1796 1804 1844 1836
rect 1876 1804 1924 1836
rect 1956 1804 2004 1836
rect 2036 1804 2084 1836
rect 2116 1804 2164 1836
rect 2196 1804 2244 1836
rect 2276 1804 2324 1836
rect 2356 1804 2404 1836
rect 2436 1804 2484 1836
rect 2516 1804 2644 1836
rect 2676 1804 2724 1836
rect 2756 1804 2804 1836
rect 2836 1804 2884 1836
rect 2916 1804 2964 1836
rect 2996 1804 3044 1836
rect 3076 1804 3124 1836
rect 3156 1804 3204 1836
rect 3236 1804 3284 1836
rect 3316 1804 3364 1836
rect 3396 1804 3444 1836
rect 3476 1804 3604 1836
rect 3636 1804 3684 1836
rect 3716 1804 3764 1836
rect 3796 1804 3844 1836
rect 3876 1804 3924 1836
rect 3956 1804 4004 1836
rect 4036 1804 4084 1836
rect 4116 1804 4164 1836
rect 4196 1804 4200 1836
rect 0 1800 4200 1804
rect 0 760 40 840
rect 4160 760 4200 840
rect 0 720 4200 760
rect 0 676 1080 720
rect 0 644 84 676
rect 116 644 1080 676
rect 0 600 1080 644
rect 1200 600 2040 720
rect 2160 600 3000 720
rect 3120 600 4200 720
rect 0 560 4200 600
rect 0 171 4200 200
rect 0 89 164 171
rect 196 160 4004 171
rect 196 89 1560 160
rect 0 40 1560 89
rect 1680 40 2520 160
rect 2640 89 4004 160
rect 4036 89 4200 171
rect 2640 40 4200 89
rect 0 0 4200 40
<< via4 >>
rect 120 2680 240 2800
rect 3960 2680 4080 2800
rect 600 1840 720 1960
rect 3480 1840 3600 1960
rect 1080 600 1200 720
rect 2040 600 2160 720
rect 3000 600 3120 720
rect 1560 40 1680 160
rect 2520 40 2640 160
<< metal5 >>
rect 60 2800 280 3000
rect 60 2680 120 2800
rect 240 2680 280 2800
rect 60 1540 280 2680
rect 80 0 280 1540
rect 560 1960 760 3000
rect 560 1840 600 1960
rect 720 1840 760 1960
rect 560 0 760 1840
rect 1040 720 1240 3000
rect 1040 600 1080 720
rect 1200 600 1240 720
rect 1040 0 1240 600
rect 1520 160 1720 3000
rect 1520 40 1560 160
rect 1680 40 1720 160
rect 1520 0 1720 40
rect 2000 720 2200 3000
rect 2000 600 2040 720
rect 2160 600 2200 720
rect 2000 0 2200 600
rect 2480 160 2680 3000
rect 2480 40 2520 160
rect 2640 40 2680 160
rect 2480 0 2680 40
rect 2960 720 3160 3000
rect 2960 600 3000 720
rect 3120 600 3160 720
rect 2960 0 3160 600
rect 3440 1960 3640 3000
rect 3440 1840 3480 1960
rect 3600 1840 3640 1960
rect 3440 0 3640 1840
rect 3920 2800 4120 3000
rect 3920 2680 3960 2800
rect 4080 2680 4120 2800
rect 3920 0 4120 2680
<< labels >>
rlabel metal2 0 720 4200 760 0 in
port 0 nsew
rlabel metal2 0 560 4200 600 0 out
port 1 nsew
rlabel locali 2080 2480 2120 2520 0 xpa
rlabel metal2 0 1360 4200 1400 0 xpb
port 2 nsew
rlabel metal2 0 240 4200 280 0 xn
port 3 nsew
rlabel metal5 80 0 280 2000 0 vdda
port 4 nsew
rlabel metal5 560 0 760 2000 0 vddx
port 5 nsew
rlabel metal2 0 1880 4200 1920 0 bp
port 6 nsew
rlabel metal5 1040 0 1240 2000 0 gnda
port 7 nsew
rlabel metal5 1520 0 1720 2000 0 vssa
port 8 nsew
rlabel metal1 1120 80 1160 180 0 n1
rlabel metal1 3040 80 3080 180 0 n2
rlabel metal1 3040 1420 3080 1720 0 pb2
rlabel metal1 1120 1420 1160 1720 0 pb1
rlabel metal1 3040 2540 3080 2840 0 pa2
rlabel metal1 1120 2540 1160 2840 0 pa1
<< end >>
