magic
tech sky130A
timestamp 1638390070
<< nwell >>
rect 60 4420 4140 4980
rect 60 2100 4140 2660
rect 60 1380 4140 1940
rect 60 660 4140 1220
<< nmos >>
rect 260 3760 1060 3860
rect 1220 3760 2020 3860
rect 2180 3760 2980 3860
rect 3140 3760 3940 3860
rect 260 3460 1060 3560
rect 1220 3460 2020 3560
rect 2180 3460 2980 3560
rect 3140 3460 3940 3560
rect 260 80 1060 180
rect 1220 80 2020 180
rect 2180 80 2980 180
rect 3140 80 3940 180
rect 260 -440 1060 -340
rect 1220 -440 2020 -340
rect 2180 -440 2980 -340
rect 3140 -440 3940 -340
<< pmoslvt >>
rect 260 4580 1060 4880
rect 1220 4580 2020 4880
rect 2180 4580 2980 4880
rect 3140 4580 3940 4880
rect 260 2200 1060 2500
rect 1220 2200 2020 2500
rect 2180 2200 2980 2500
rect 3140 2200 3940 2500
rect 260 1540 1060 1840
rect 1220 1540 2020 1840
rect 2180 1540 2980 1840
rect 3140 1540 3940 1840
rect 260 820 1060 1120
rect 1220 820 2020 1120
rect 2180 820 2980 1120
rect 3140 820 3940 1120
<< ndiff >>
rect 160 3850 260 3860
rect 160 3770 165 3850
rect 195 3770 260 3850
rect 160 3760 260 3770
rect 1060 3850 1220 3860
rect 1060 3770 1125 3850
rect 1155 3770 1220 3850
rect 1060 3760 1220 3770
rect 2020 3850 2180 3860
rect 2020 3770 2085 3850
rect 2115 3770 2180 3850
rect 2020 3760 2180 3770
rect 2980 3850 3140 3860
rect 2980 3770 3045 3850
rect 3075 3770 3140 3850
rect 2980 3760 3140 3770
rect 3940 3850 4040 3860
rect 3940 3770 4005 3850
rect 4035 3770 4040 3850
rect 3940 3760 4040 3770
rect 160 3550 260 3560
rect 160 3470 165 3550
rect 195 3470 260 3550
rect 160 3460 260 3470
rect 1060 3550 1220 3560
rect 1060 3470 1125 3550
rect 1155 3470 1220 3550
rect 1060 3460 1220 3470
rect 2020 3550 2180 3560
rect 2020 3470 2085 3550
rect 2115 3470 2180 3550
rect 2020 3460 2180 3470
rect 2980 3550 3140 3560
rect 2980 3470 3045 3550
rect 3075 3470 3140 3550
rect 2980 3460 3140 3470
rect 3940 3550 4040 3560
rect 3940 3470 4005 3550
rect 4035 3470 4040 3550
rect 3940 3460 4040 3470
rect 160 170 260 180
rect 160 90 165 170
rect 195 90 260 170
rect 160 80 260 90
rect 1060 170 1220 180
rect 1060 90 1125 170
rect 1155 90 1220 170
rect 1060 80 1220 90
rect 2020 170 2180 180
rect 2020 90 2085 170
rect 2115 90 2180 170
rect 2020 80 2180 90
rect 2980 170 3140 180
rect 2980 90 3045 170
rect 3075 90 3140 170
rect 2980 80 3140 90
rect 3940 170 4040 180
rect 3940 90 4005 170
rect 4035 90 4040 170
rect 3940 80 4040 90
rect 160 -350 260 -340
rect 160 -430 165 -350
rect 195 -430 260 -350
rect 160 -440 260 -430
rect 1060 -350 1220 -340
rect 1060 -430 1125 -350
rect 1155 -430 1220 -350
rect 1060 -440 1220 -430
rect 2020 -350 2180 -340
rect 2020 -430 2085 -350
rect 2115 -430 2180 -350
rect 2020 -440 2180 -430
rect 2980 -350 3140 -340
rect 2980 -430 3045 -350
rect 3075 -430 3140 -350
rect 2980 -440 3140 -430
rect 3940 -350 4040 -340
rect 3940 -430 4005 -350
rect 4035 -430 4040 -350
rect 3940 -440 4040 -430
<< pdiff >>
rect 160 4870 260 4880
rect 160 4590 165 4870
rect 195 4590 260 4870
rect 160 4580 260 4590
rect 1060 4870 1220 4880
rect 1060 4590 1125 4870
rect 1155 4590 1220 4870
rect 1060 4580 1220 4590
rect 2020 4870 2180 4880
rect 2020 4590 2085 4870
rect 2115 4590 2180 4870
rect 2020 4580 2180 4590
rect 2980 4870 3140 4880
rect 2980 4590 3045 4870
rect 3075 4590 3140 4870
rect 2980 4580 3140 4590
rect 3940 4870 4040 4880
rect 3940 4590 4005 4870
rect 4035 4590 4040 4870
rect 3940 4580 4040 4590
rect 160 2490 260 2500
rect 160 2210 165 2490
rect 195 2210 260 2490
rect 160 2200 260 2210
rect 1060 2490 1220 2500
rect 1060 2210 1125 2490
rect 1155 2210 1220 2490
rect 1060 2200 1220 2210
rect 2020 2490 2180 2500
rect 2020 2210 2085 2490
rect 2115 2210 2180 2490
rect 2020 2200 2180 2210
rect 2980 2490 3140 2500
rect 2980 2210 3045 2490
rect 3075 2210 3140 2490
rect 2980 2200 3140 2210
rect 3940 2490 4040 2500
rect 3940 2210 4005 2490
rect 4035 2210 4040 2490
rect 3940 2200 4040 2210
rect 160 1830 260 1840
rect 160 1550 165 1830
rect 195 1550 260 1830
rect 160 1540 260 1550
rect 1060 1830 1220 1840
rect 1060 1550 1125 1830
rect 1155 1550 1220 1830
rect 1060 1540 1220 1550
rect 2020 1830 2180 1840
rect 2020 1550 2085 1830
rect 2115 1550 2180 1830
rect 2020 1540 2180 1550
rect 2980 1830 3140 1840
rect 2980 1550 3045 1830
rect 3075 1550 3140 1830
rect 2980 1540 3140 1550
rect 3940 1830 4040 1840
rect 3940 1550 4005 1830
rect 4035 1550 4040 1830
rect 3940 1540 4040 1550
rect 160 1110 260 1120
rect 160 830 165 1110
rect 195 830 260 1110
rect 160 820 260 830
rect 1060 1110 1220 1120
rect 1060 830 1125 1110
rect 1155 830 1220 1110
rect 1060 820 1220 830
rect 2020 1110 2180 1120
rect 2020 830 2085 1110
rect 2115 830 2180 1110
rect 2020 820 2180 830
rect 2980 1110 3140 1120
rect 2980 830 3045 1110
rect 3075 830 3140 1110
rect 2980 820 3140 830
rect 3940 1110 4040 1120
rect 3940 830 4005 1110
rect 4035 830 4040 1110
rect 3940 820 4040 830
<< ndiffc >>
rect 165 3770 195 3850
rect 1125 3770 1155 3850
rect 2085 3770 2115 3850
rect 3045 3770 3075 3850
rect 4005 3770 4035 3850
rect 165 3470 195 3550
rect 1125 3470 1155 3550
rect 2085 3470 2115 3550
rect 3045 3470 3075 3550
rect 4005 3470 4035 3550
rect 165 90 195 170
rect 1125 90 1155 170
rect 2085 90 2115 170
rect 3045 90 3075 170
rect 4005 90 4035 170
rect 165 -430 195 -350
rect 1125 -430 1155 -350
rect 2085 -430 2115 -350
rect 3045 -430 3075 -350
rect 4005 -430 4035 -350
<< pdiffc >>
rect 165 4590 195 4870
rect 1125 4590 1155 4870
rect 2085 4590 2115 4870
rect 3045 4590 3075 4870
rect 4005 4590 4035 4870
rect 165 2210 195 2490
rect 1125 2210 1155 2490
rect 2085 2210 2115 2490
rect 3045 2210 3075 2490
rect 4005 2210 4035 2490
rect 165 1550 195 1830
rect 1125 1550 1155 1830
rect 2085 1550 2115 1830
rect 3045 1550 3075 1830
rect 4005 1550 4035 1830
rect 165 830 195 1110
rect 1125 830 1155 1110
rect 2085 830 2115 1110
rect 3045 830 3075 1110
rect 4005 830 4035 1110
<< psubdiff >>
rect 0 5000 60 5040
rect 4140 5000 4200 5040
rect 0 4980 40 5000
rect 4160 4980 4200 5000
rect 0 4400 40 4420
rect 4160 4400 4200 4420
rect 0 4360 60 4400
rect 4140 4360 4200 4400
rect 0 4000 40 4360
rect 4160 4000 4200 4360
rect 0 3960 60 4000
rect 4140 3960 4200 4000
rect 0 3940 40 3960
rect 0 3720 40 3740
rect 4160 3720 4200 3960
rect 0 3680 60 3720
rect 4140 3680 4200 3720
rect 0 3600 60 3640
rect 4140 3600 4200 3640
rect 0 3580 40 3600
rect 0 3360 40 3380
rect 4160 3360 4200 3600
rect 0 3320 60 3360
rect 4140 3320 4200 3360
rect 0 2720 40 3320
rect 4160 2720 4200 3320
rect 0 2680 60 2720
rect 4140 2680 4200 2720
rect 0 2660 40 2680
rect 4160 2660 4200 2680
rect 0 2080 40 2100
rect 4160 2080 4200 2100
rect 0 2040 60 2080
rect 4140 2040 4200 2080
rect 0 1960 60 2000
rect 4140 1960 4200 2000
rect 0 1940 40 1960
rect 4160 1940 4200 1960
rect 0 1360 40 1380
rect 4160 1360 4200 1380
rect 0 1320 60 1360
rect 4120 1320 4200 1360
rect 0 1240 60 1280
rect 4120 1240 4200 1280
rect 0 1220 40 1240
rect 4160 1220 4200 1240
rect 0 640 40 660
rect 0 600 60 640
rect 4140 600 4160 640
rect 0 280 60 320
rect 4140 280 4160 320
rect 0 260 40 280
rect 0 40 40 60
rect 4160 40 4200 60
rect 0 0 60 40
rect 4140 0 4200 40
rect 0 -240 60 -200
rect 4140 -240 4200 -200
rect 0 -260 40 -240
rect 4160 -260 4200 -240
rect 0 -480 40 -460
rect 4160 -480 4200 -460
rect 0 -520 60 -480
rect 4140 -520 4200 -480
<< nsubdiff >>
rect 80 4920 140 4960
rect 4060 4920 4120 4960
rect 80 4900 120 4920
rect 4080 4900 4120 4920
rect 80 4480 120 4500
rect 4080 4480 4120 4500
rect 80 4440 140 4480
rect 4060 4440 4120 4480
rect 80 2600 140 2640
rect 4060 2600 4120 2640
rect 80 2580 120 2600
rect 4080 2580 4120 2600
rect 80 2160 120 2180
rect 4080 2160 4120 2180
rect 80 2120 140 2160
rect 4060 2120 4120 2160
rect 80 1880 140 1920
rect 4060 1880 4120 1920
rect 80 1860 120 1880
rect 4080 1860 4120 1880
rect 80 1440 120 1460
rect 4080 1440 4120 1460
rect 80 1400 140 1440
rect 4060 1400 4120 1440
rect 80 1160 140 1200
rect 4060 1160 4120 1200
rect 80 1140 120 1160
rect 4080 1140 4120 1160
rect 80 720 120 740
rect 4080 720 4120 740
rect 80 680 140 720
rect 4060 680 4120 720
<< psubdiffcont >>
rect 60 5000 4140 5040
rect 0 4420 40 4980
rect 4160 4420 4200 4980
rect 60 4360 4140 4400
rect 60 3960 4140 4000
rect 0 3740 40 3940
rect 60 3680 4140 3720
rect 60 3600 4140 3640
rect 0 3380 40 3580
rect 60 3320 4140 3360
rect 60 2680 4140 2720
rect 0 2100 40 2660
rect 4160 2100 4200 2660
rect 60 2040 4140 2080
rect 60 1960 4140 2000
rect 0 1380 40 1940
rect 4160 1380 4200 1940
rect 60 1320 4120 1360
rect 60 1240 4120 1280
rect 0 660 40 1220
rect 60 600 4140 640
rect 60 280 4140 320
rect 0 60 40 260
rect 4160 60 4200 1220
rect 60 0 4140 40
rect 60 -240 4140 -200
rect 0 -460 40 -260
rect 4160 -460 4200 -260
rect 60 -520 4140 -480
<< nsubdiffcont >>
rect 140 4920 4060 4960
rect 80 4500 120 4900
rect 4080 4500 4120 4900
rect 140 4440 4060 4480
rect 140 2600 4060 2640
rect 80 2180 120 2580
rect 4080 2180 4120 2580
rect 140 2120 4060 2160
rect 140 1880 4060 1920
rect 80 1460 120 1860
rect 4080 1460 4120 1860
rect 140 1400 4060 1440
rect 140 1160 4060 1200
rect 80 740 120 1140
rect 4080 740 4120 1140
rect 140 680 4060 720
<< poly >>
rect 260 4880 1060 4900
rect 1220 4880 2020 4900
rect 2180 4880 2980 4900
rect 3140 4880 3940 4900
rect 260 4555 1060 4580
rect 260 4525 270 4555
rect 1050 4525 1060 4555
rect 260 4520 1060 4525
rect 1220 4555 2020 4580
rect 1220 4525 1230 4555
rect 2010 4525 2020 4555
rect 1220 4520 2020 4525
rect 2180 4555 2980 4580
rect 2180 4525 2190 4555
rect 2970 4525 2980 4555
rect 2180 4520 2980 4525
rect 3140 4555 3940 4580
rect 3140 4525 3150 4555
rect 3930 4525 3940 4555
rect 3140 4520 3940 4525
rect 260 3915 1060 3920
rect 260 3885 270 3915
rect 1050 3885 1060 3915
rect 260 3860 1060 3885
rect 1220 3915 2020 3920
rect 1220 3885 1230 3915
rect 2010 3885 2020 3915
rect 1220 3860 2020 3885
rect 2180 3915 2980 3920
rect 2180 3885 2190 3915
rect 2970 3885 2980 3915
rect 2180 3860 2980 3885
rect 3140 3915 3940 3920
rect 3140 3885 3150 3915
rect 3930 3885 3940 3915
rect 3140 3860 3940 3885
rect 260 3740 1060 3760
rect 1220 3740 2020 3760
rect 2180 3740 2980 3760
rect 3140 3740 3940 3760
rect 260 3560 1060 3580
rect 1220 3560 2020 3580
rect 2180 3560 2980 3580
rect 3140 3560 3940 3580
rect 260 3435 1060 3460
rect 260 3405 270 3435
rect 1050 3405 1060 3435
rect 260 3400 1060 3405
rect 1220 3435 2020 3460
rect 1220 3405 1230 3435
rect 2010 3405 2020 3435
rect 1220 3400 2020 3405
rect 2180 3435 2980 3460
rect 2180 3405 2190 3435
rect 2970 3405 2980 3435
rect 2180 3400 2980 3405
rect 3140 3435 3940 3460
rect 3140 3405 3150 3435
rect 3930 3405 3940 3435
rect 3140 3400 3940 3405
rect 260 2555 1060 2560
rect 260 2525 270 2555
rect 1050 2525 1060 2555
rect 260 2500 1060 2525
rect 1220 2555 2020 2560
rect 1220 2525 1230 2555
rect 2010 2525 2020 2555
rect 1220 2500 2020 2525
rect 2180 2555 2980 2560
rect 2180 2525 2190 2555
rect 2970 2525 2980 2555
rect 2180 2500 2980 2525
rect 3140 2555 3940 2560
rect 3140 2525 3150 2555
rect 3930 2525 3940 2555
rect 3140 2500 3940 2525
rect 260 2180 1060 2200
rect 1220 2180 2020 2200
rect 2180 2180 2980 2200
rect 3140 2180 3940 2200
rect 260 1840 1060 1860
rect 1220 1840 2020 1860
rect 2180 1840 2980 1860
rect 3140 1840 3940 1860
rect 260 1515 1060 1540
rect 260 1485 270 1515
rect 1050 1485 1060 1515
rect 260 1480 1060 1485
rect 1220 1515 2020 1540
rect 1220 1485 1230 1515
rect 2010 1485 2020 1515
rect 1220 1480 2020 1485
rect 2180 1515 2980 1540
rect 2180 1485 2190 1515
rect 2970 1485 2980 1515
rect 2180 1480 2980 1485
rect 3140 1515 3940 1540
rect 3140 1485 3150 1515
rect 3930 1485 3940 1515
rect 3140 1480 3940 1485
rect 260 1120 1060 1140
rect 1220 1120 2020 1140
rect 2180 1120 2980 1140
rect 3140 1120 3940 1140
rect 260 795 1060 820
rect 260 765 270 795
rect 1050 765 1060 795
rect 260 760 1060 765
rect 1220 795 2020 820
rect 1220 765 1230 795
rect 2010 765 2020 795
rect 1220 760 2020 765
rect 2180 795 2980 820
rect 2180 765 2190 795
rect 2970 765 2980 795
rect 2180 760 2980 765
rect 3140 795 3940 820
rect 3140 765 3150 795
rect 3930 765 3940 795
rect 3140 760 3940 765
rect 260 235 1060 240
rect 260 205 270 235
rect 1050 205 1060 235
rect 260 180 1060 205
rect 1220 235 2020 240
rect 1220 205 1230 235
rect 2010 205 2020 235
rect 1220 180 2020 205
rect 2180 235 2980 240
rect 2180 205 2190 235
rect 2970 205 2980 235
rect 2180 180 2980 205
rect 3140 235 3940 240
rect 3140 205 3150 235
rect 3930 205 3940 235
rect 3140 180 3940 205
rect 260 60 1060 80
rect 1220 60 2020 80
rect 2180 60 2980 80
rect 3140 60 3940 80
rect 260 -285 1060 -280
rect 260 -315 270 -285
rect 1050 -315 1060 -285
rect 260 -340 1060 -315
rect 1220 -285 2020 -280
rect 1220 -315 1230 -285
rect 2010 -315 2020 -285
rect 1220 -340 2020 -315
rect 2180 -285 2980 -280
rect 2180 -315 2190 -285
rect 2970 -315 2980 -285
rect 2180 -340 2980 -315
rect 3140 -285 3940 -280
rect 3140 -315 3150 -285
rect 3930 -315 3940 -285
rect 3140 -340 3940 -315
rect 260 -460 1060 -440
rect 1220 -460 2020 -440
rect 2180 -460 2980 -440
rect 3140 -460 3940 -440
<< polycont >>
rect 270 4525 1050 4555
rect 1230 4525 2010 4555
rect 2190 4525 2970 4555
rect 3150 4525 3930 4555
rect 270 3885 1050 3915
rect 1230 3885 2010 3915
rect 2190 3885 2970 3915
rect 3150 3885 3930 3915
rect 270 3405 1050 3435
rect 1230 3405 2010 3435
rect 2190 3405 2970 3435
rect 3150 3405 3930 3435
rect 270 2525 1050 2555
rect 1230 2525 2010 2555
rect 2190 2525 2970 2555
rect 3150 2525 3930 2555
rect 270 1485 1050 1515
rect 1230 1485 2010 1515
rect 2190 1485 2970 1515
rect 3150 1485 3930 1515
rect 270 765 1050 795
rect 1230 765 2010 795
rect 2190 765 2970 795
rect 3150 765 3930 795
rect 270 205 1050 235
rect 1230 205 2010 235
rect 2190 205 2970 235
rect 3150 205 3930 235
rect 270 -315 1050 -285
rect 1230 -315 2010 -285
rect 2190 -315 2970 -285
rect 3150 -315 3930 -285
<< locali >>
rect 0 5000 60 5040
rect 4140 5000 4200 5040
rect 0 4980 40 5000
rect 4160 4980 4200 5000
rect 80 4920 140 4960
rect 4060 4920 4120 4960
rect 80 4900 120 4920
rect 160 4870 200 4920
rect 4080 4900 4120 4920
rect 160 4590 165 4870
rect 195 4590 200 4870
rect 160 4580 200 4590
rect 1120 4870 1160 4880
rect 1120 4590 1125 4870
rect 1155 4590 1160 4870
rect 1120 4580 1160 4590
rect 2080 4870 2120 4880
rect 2080 4590 2085 4870
rect 2115 4590 2120 4870
rect 2080 4580 2120 4590
rect 3040 4870 3080 4880
rect 3040 4590 3045 4870
rect 3075 4590 3080 4870
rect 3040 4580 3080 4590
rect 4000 4870 4040 4880
rect 4000 4590 4005 4870
rect 4035 4590 4040 4870
rect 4000 4580 4040 4590
rect 260 4555 1060 4560
rect 260 4525 270 4555
rect 1050 4525 1060 4555
rect 260 4520 1060 4525
rect 1220 4555 2020 4560
rect 1220 4525 1230 4555
rect 2010 4525 2020 4555
rect 1220 4520 2020 4525
rect 2180 4555 2980 4560
rect 2180 4525 2190 4555
rect 2970 4525 2980 4555
rect 2180 4520 2980 4525
rect 3140 4555 3940 4560
rect 3140 4525 3150 4555
rect 3930 4525 3940 4555
rect 3140 4520 3940 4525
rect 80 4480 120 4500
rect 4080 4480 4120 4500
rect 80 4440 140 4480
rect 4060 4440 4120 4480
rect 0 4400 40 4420
rect 4160 4400 4200 4420
rect 0 4360 60 4400
rect 4140 4360 4200 4400
rect 0 4000 40 4360
rect 80 4230 4120 4320
rect 80 4210 90 4230
rect 110 4210 4090 4230
rect 4110 4210 4120 4230
rect 80 4200 4120 4210
rect 80 4150 4120 4160
rect 80 4130 90 4150
rect 110 4130 4090 4150
rect 4110 4130 4120 4150
rect 80 4040 4120 4130
rect 4160 4000 4200 4360
rect 0 3960 60 4000
rect 4140 3960 4200 4000
rect 0 3940 40 3960
rect 260 3915 1060 3920
rect 260 3885 270 3915
rect 1050 3885 1060 3915
rect 260 3880 1060 3885
rect 1220 3915 2020 3920
rect 1220 3885 1230 3915
rect 2010 3885 2020 3915
rect 1220 3880 2020 3885
rect 2180 3915 2980 3920
rect 2180 3885 2190 3915
rect 2970 3885 2980 3915
rect 2180 3880 2980 3885
rect 3140 3915 3940 3920
rect 3140 3885 3150 3915
rect 3930 3885 3940 3915
rect 3140 3880 3940 3885
rect 0 3720 40 3740
rect 160 3850 200 3860
rect 160 3770 165 3850
rect 195 3770 200 3850
rect 160 3720 200 3770
rect 1120 3850 1160 3860
rect 1120 3770 1125 3850
rect 1155 3770 1160 3850
rect 1120 3760 1160 3770
rect 2080 3850 2120 3860
rect 2080 3770 2085 3850
rect 2115 3770 2120 3850
rect 2080 3760 2120 3770
rect 3040 3850 3080 3860
rect 3040 3770 3045 3850
rect 3075 3770 3080 3850
rect 3040 3760 3080 3770
rect 4000 3850 4040 3860
rect 4000 3770 4005 3850
rect 4035 3770 4040 3850
rect 4000 3760 4040 3770
rect 4160 3720 4200 3960
rect 0 3680 60 3720
rect 4140 3680 4200 3720
rect 0 3640 40 3680
rect 4160 3640 4200 3680
rect 0 3600 60 3640
rect 4140 3600 4200 3640
rect 0 3580 40 3600
rect 160 3550 200 3600
rect 160 3470 165 3550
rect 195 3470 200 3550
rect 160 3460 200 3470
rect 1120 3550 1160 3560
rect 1120 3470 1125 3550
rect 1155 3470 1160 3550
rect 1120 3460 1160 3470
rect 2080 3550 2120 3560
rect 2080 3470 2085 3550
rect 2115 3470 2120 3550
rect 2080 3460 2120 3470
rect 3040 3550 3080 3560
rect 3040 3470 3045 3550
rect 3075 3470 3080 3550
rect 3040 3460 3080 3470
rect 4000 3550 4040 3560
rect 4000 3470 4005 3550
rect 4035 3470 4040 3550
rect 4000 3460 4040 3470
rect 260 3435 1060 3440
rect 260 3405 270 3435
rect 1050 3405 1060 3435
rect 260 3400 1060 3405
rect 1220 3435 2020 3440
rect 1220 3405 1230 3435
rect 2010 3405 2020 3435
rect 1220 3400 2020 3405
rect 2180 3435 2980 3440
rect 2180 3405 2190 3435
rect 2970 3405 2980 3435
rect 2180 3400 2980 3405
rect 3140 3435 3940 3440
rect 3140 3405 3150 3435
rect 3930 3405 3940 3435
rect 3140 3400 3940 3405
rect 0 3360 40 3380
rect 4160 3360 4200 3600
rect 0 3320 60 3360
rect 4140 3320 4200 3360
rect 0 2720 40 3320
rect 80 3190 4120 3280
rect 80 3170 90 3190
rect 110 3170 4090 3190
rect 4110 3170 4120 3190
rect 80 3160 4120 3170
rect 80 3110 4120 3120
rect 80 3090 90 3110
rect 110 3090 4090 3110
rect 4110 3090 4120 3110
rect 80 2950 4120 3090
rect 80 2930 90 2950
rect 110 2930 4090 2950
rect 4110 2930 4120 2950
rect 80 2920 4120 2930
rect 80 2870 4120 2880
rect 80 2850 90 2870
rect 110 2850 4090 2870
rect 4110 2850 4120 2870
rect 80 2760 4120 2850
rect 4160 2720 4200 3320
rect 0 2680 60 2720
rect 4140 2680 4200 2720
rect 0 2660 40 2680
rect 4160 2660 4200 2680
rect 80 2600 140 2640
rect 4060 2600 4120 2640
rect 80 2580 120 2600
rect 4080 2580 4120 2600
rect 260 2555 1060 2560
rect 260 2525 270 2555
rect 1050 2525 1060 2555
rect 260 2520 1060 2525
rect 1220 2555 2020 2560
rect 1220 2525 1230 2555
rect 2010 2525 2020 2555
rect 1220 2520 2020 2525
rect 2180 2555 2980 2560
rect 2180 2525 2190 2555
rect 2970 2525 2980 2555
rect 2180 2520 2980 2525
rect 3140 2555 3940 2560
rect 3140 2525 3150 2555
rect 3930 2525 3940 2555
rect 3140 2520 3940 2525
rect 80 2160 120 2180
rect 160 2490 200 2500
rect 160 2210 165 2490
rect 195 2210 200 2490
rect 160 2160 200 2210
rect 1120 2490 1160 2500
rect 1120 2210 1125 2490
rect 1155 2210 1160 2490
rect 1120 2200 1160 2210
rect 2080 2490 2120 2500
rect 2080 2210 2085 2490
rect 2115 2210 2120 2490
rect 2080 2200 2120 2210
rect 3040 2490 3080 2500
rect 3040 2210 3045 2490
rect 3075 2210 3080 2490
rect 3040 2200 3080 2210
rect 4000 2490 4040 2500
rect 4000 2210 4005 2490
rect 4035 2210 4040 2490
rect 4000 2200 4040 2210
rect 4080 2160 4120 2180
rect 80 2120 140 2160
rect 4060 2120 4120 2160
rect 0 2080 40 2100
rect 4160 2080 4200 2100
rect 0 2040 60 2080
rect 4140 2040 4200 2080
rect 0 2000 40 2040
rect 4160 2000 4200 2040
rect 0 1960 60 2000
rect 4140 1960 4200 2000
rect 0 1940 40 1960
rect 4160 1940 4200 1960
rect 80 1880 140 1920
rect 4060 1880 4120 1920
rect 80 1860 120 1880
rect 160 1830 200 1840
rect 160 1550 165 1830
rect 195 1550 200 1830
rect 160 1540 200 1550
rect 1120 1830 1160 1840
rect 1120 1550 1125 1830
rect 1155 1550 1160 1830
rect 1120 1540 1160 1550
rect 2080 1830 2120 1840
rect 2080 1550 2085 1830
rect 2115 1550 2120 1830
rect 2080 1540 2120 1550
rect 3040 1830 3080 1840
rect 3040 1550 3045 1830
rect 3075 1550 3080 1830
rect 3040 1540 3080 1550
rect 4000 1830 4040 1880
rect 4000 1550 4005 1830
rect 4035 1550 4040 1830
rect 4000 1540 4040 1550
rect 4080 1860 4120 1880
rect 260 1515 1060 1520
rect 260 1485 270 1515
rect 1050 1485 1060 1515
rect 260 1480 1060 1485
rect 1220 1515 2020 1520
rect 1220 1485 1230 1515
rect 2010 1485 2020 1515
rect 1220 1480 2020 1485
rect 2180 1515 2980 1520
rect 2180 1485 2190 1515
rect 2970 1485 2980 1515
rect 2180 1480 2980 1485
rect 3140 1515 3940 1520
rect 3140 1485 3150 1515
rect 3930 1485 3940 1515
rect 3140 1480 3940 1485
rect 80 1440 120 1460
rect 4080 1440 4120 1460
rect 80 1400 140 1440
rect 4060 1400 4120 1440
rect 0 1360 40 1380
rect 4160 1360 4200 1380
rect 0 1320 60 1360
rect 4120 1320 4200 1360
rect 0 1280 40 1320
rect 4160 1280 4200 1320
rect 0 1240 60 1280
rect 4120 1240 4200 1280
rect 0 1220 40 1240
rect 4160 1220 4200 1240
rect 80 1160 140 1200
rect 4060 1160 4120 1200
rect 80 1140 120 1160
rect 160 1110 200 1160
rect 4080 1140 4120 1160
rect 160 830 165 1110
rect 195 830 200 1110
rect 160 820 200 830
rect 1120 1110 1160 1120
rect 1120 830 1125 1110
rect 1155 830 1160 1110
rect 1120 820 1160 830
rect 2080 1110 2120 1120
rect 2080 830 2085 1110
rect 2115 830 2120 1110
rect 2080 820 2120 830
rect 3040 1110 3080 1120
rect 3040 830 3045 1110
rect 3075 830 3080 1110
rect 3040 820 3080 830
rect 4000 1110 4040 1120
rect 4000 830 4005 1110
rect 4035 830 4040 1110
rect 4000 820 4040 830
rect 260 795 1060 800
rect 260 765 270 795
rect 1050 765 1060 795
rect 260 760 1060 765
rect 1220 795 2020 800
rect 1220 765 1230 795
rect 2010 765 2020 795
rect 1220 760 2020 765
rect 2180 795 2980 800
rect 2180 765 2190 795
rect 2970 765 2980 795
rect 2180 760 2980 765
rect 3140 795 3940 800
rect 3140 765 3150 795
rect 3930 765 3940 795
rect 3140 760 3940 765
rect 80 720 120 740
rect 4080 720 4120 740
rect 80 680 140 720
rect 4060 680 4120 720
rect 0 640 40 660
rect 0 600 60 640
rect 4140 600 4160 640
rect 0 320 40 600
rect 80 470 4120 560
rect 80 450 90 470
rect 110 450 170 470
rect 190 450 250 470
rect 270 450 330 470
rect 350 450 410 470
rect 430 450 490 470
rect 510 450 570 470
rect 590 450 730 470
rect 750 450 810 470
rect 830 450 890 470
rect 910 450 970 470
rect 990 450 1050 470
rect 1070 450 1130 470
rect 1150 450 1210 470
rect 1230 450 1290 470
rect 1310 450 1370 470
rect 1390 450 1450 470
rect 1470 450 1530 470
rect 1550 450 1690 470
rect 1710 450 1770 470
rect 1790 450 1850 470
rect 1870 450 1930 470
rect 1950 450 2010 470
rect 2030 450 2090 470
rect 2110 450 2170 470
rect 2190 450 2250 470
rect 2270 450 2330 470
rect 2350 450 2410 470
rect 2430 450 2490 470
rect 2510 450 2650 470
rect 2670 450 2730 470
rect 2750 450 2810 470
rect 2830 450 2890 470
rect 2910 450 2970 470
rect 2990 450 3050 470
rect 3070 450 3130 470
rect 3150 450 3210 470
rect 3230 450 3290 470
rect 3310 450 3370 470
rect 3390 450 3450 470
rect 3470 450 3610 470
rect 3630 450 3690 470
rect 3710 450 3770 470
rect 3790 450 3850 470
rect 3870 450 3930 470
rect 3950 450 4090 470
rect 4110 450 4120 470
rect 80 360 4120 450
rect 0 280 60 320
rect 4140 280 4160 320
rect 0 260 40 280
rect 260 235 1060 240
rect 260 205 270 235
rect 1050 205 1060 235
rect 260 200 1060 205
rect 1220 235 2020 240
rect 1220 205 1230 235
rect 2010 205 2020 235
rect 1220 200 2020 205
rect 2180 235 2980 240
rect 2180 205 2190 235
rect 2970 205 2980 235
rect 2180 200 2980 205
rect 3140 235 3940 240
rect 3140 205 3150 235
rect 3930 205 3940 235
rect 3140 200 3940 205
rect 0 40 40 60
rect 160 170 200 180
rect 160 90 165 170
rect 195 90 200 170
rect 160 40 200 90
rect 1120 170 1160 180
rect 1120 90 1125 170
rect 1155 90 1160 170
rect 1120 80 1160 90
rect 2080 170 2120 180
rect 2080 90 2085 170
rect 2115 90 2120 170
rect 2080 80 2120 90
rect 3040 170 3080 180
rect 3040 90 3045 170
rect 3075 90 3080 170
rect 3040 80 3080 90
rect 4000 170 4040 180
rect 4000 90 4005 170
rect 4035 90 4040 170
rect 4000 80 4040 90
rect 4160 40 4200 60
rect 0 0 60 40
rect 4140 0 4200 40
rect 0 -200 40 0
rect 80 -50 4120 -40
rect 80 -70 90 -50
rect 110 -70 170 -50
rect 190 -70 250 -50
rect 270 -70 330 -50
rect 350 -70 410 -50
rect 430 -70 490 -50
rect 510 -70 570 -50
rect 590 -70 730 -50
rect 750 -70 810 -50
rect 830 -70 890 -50
rect 910 -70 970 -50
rect 990 -70 1050 -50
rect 1070 -70 1130 -50
rect 1150 -70 1210 -50
rect 1230 -70 1290 -50
rect 1310 -70 1370 -50
rect 1390 -70 1450 -50
rect 1470 -70 1530 -50
rect 1550 -70 1690 -50
rect 1710 -70 1770 -50
rect 1790 -70 1850 -50
rect 1870 -70 1930 -50
rect 1950 -70 2010 -50
rect 2030 -70 2090 -50
rect 2110 -70 2170 -50
rect 2190 -70 2250 -50
rect 2270 -70 2330 -50
rect 2350 -70 2410 -50
rect 2430 -70 2490 -50
rect 2510 -70 2650 -50
rect 2670 -70 2730 -50
rect 2750 -70 2810 -50
rect 2830 -70 2890 -50
rect 2910 -70 2970 -50
rect 2990 -70 3050 -50
rect 3070 -70 3130 -50
rect 3150 -70 3210 -50
rect 3230 -70 3290 -50
rect 3310 -70 3370 -50
rect 3390 -70 3450 -50
rect 3470 -70 3610 -50
rect 3630 -70 3690 -50
rect 3710 -70 3770 -50
rect 3790 -70 3850 -50
rect 3870 -70 3930 -50
rect 3950 -70 4090 -50
rect 4110 -70 4120 -50
rect 80 -160 4120 -70
rect 4160 -200 4200 0
rect 0 -240 60 -200
rect 4140 -240 4200 -200
rect 0 -260 40 -240
rect 4160 -260 4200 -240
rect 260 -285 1060 -280
rect 260 -315 270 -285
rect 1050 -315 1060 -285
rect 260 -320 1060 -315
rect 1220 -285 2020 -280
rect 1220 -315 1230 -285
rect 2010 -315 2020 -285
rect 1220 -320 2020 -315
rect 2180 -285 2980 -280
rect 2180 -315 2190 -285
rect 2970 -315 2980 -285
rect 2180 -320 2980 -315
rect 3140 -285 3940 -280
rect 3140 -315 3150 -285
rect 3930 -315 3940 -285
rect 3140 -320 3940 -315
rect 0 -480 40 -460
rect 160 -350 200 -340
rect 160 -430 165 -350
rect 195 -430 200 -350
rect 160 -480 200 -430
rect 1120 -350 1160 -340
rect 1120 -430 1125 -350
rect 1155 -430 1160 -350
rect 1120 -440 1160 -430
rect 2080 -350 2120 -340
rect 2080 -430 2085 -350
rect 2115 -430 2120 -350
rect 2080 -440 2120 -430
rect 3040 -350 3080 -340
rect 3040 -430 3045 -350
rect 3075 -430 3080 -350
rect 3040 -440 3080 -430
rect 4000 -350 4040 -340
rect 4000 -430 4005 -350
rect 4035 -430 4040 -350
rect 4000 -440 4040 -430
rect 4160 -480 4200 -460
rect 0 -520 60 -480
rect 4140 -520 4200 -480
<< viali >>
rect 165 4590 195 4870
rect 1125 4590 1155 4870
rect 2085 4590 2115 4870
rect 3045 4590 3075 4870
rect 4005 4590 4035 4870
rect 270 4525 1050 4555
rect 1230 4525 2010 4555
rect 2190 4525 2970 4555
rect 3150 4525 3930 4555
rect 90 4210 110 4230
rect 4090 4210 4110 4230
rect 90 4130 110 4150
rect 4090 4130 4110 4150
rect 270 3885 1050 3915
rect 1230 3885 2010 3915
rect 2190 3885 2970 3915
rect 3150 3885 3930 3915
rect 165 3770 195 3850
rect 1125 3770 1155 3850
rect 2085 3770 2115 3850
rect 3045 3770 3075 3850
rect 4005 3770 4035 3850
rect 165 3470 195 3550
rect 1125 3470 1155 3550
rect 2085 3470 2115 3550
rect 3045 3470 3075 3550
rect 4005 3470 4035 3550
rect 270 3405 1050 3435
rect 1230 3405 2010 3435
rect 2190 3405 2970 3435
rect 3150 3405 3930 3435
rect 90 3170 110 3190
rect 4090 3170 4110 3190
rect 90 3090 110 3110
rect 4090 3090 4110 3110
rect 90 2930 110 2950
rect 4090 2930 4110 2950
rect 90 2850 110 2870
rect 4090 2850 4110 2870
rect 270 2525 1050 2555
rect 1230 2525 2010 2555
rect 2190 2525 2970 2555
rect 3150 2525 3930 2555
rect 165 2210 195 2490
rect 1125 2210 1155 2490
rect 2085 2210 2115 2490
rect 3045 2210 3075 2490
rect 4005 2210 4035 2490
rect 165 1550 195 1830
rect 1125 1550 1155 1830
rect 2085 1550 2115 1830
rect 3045 1550 3075 1830
rect 4005 1550 4035 1830
rect 270 1485 1050 1515
rect 1230 1485 2010 1515
rect 2190 1485 2970 1515
rect 3150 1485 3930 1515
rect 165 830 195 1110
rect 1125 830 1155 1110
rect 2085 830 2115 1110
rect 3045 830 3075 1110
rect 4005 830 4035 1110
rect 270 765 1050 795
rect 1230 765 2010 795
rect 2190 765 2970 795
rect 3150 765 3930 795
rect 90 450 110 470
rect 170 450 190 470
rect 250 450 270 470
rect 330 450 350 470
rect 410 450 430 470
rect 490 450 510 470
rect 570 450 590 470
rect 730 450 750 470
rect 810 450 830 470
rect 890 450 910 470
rect 970 450 990 470
rect 1050 450 1070 470
rect 1130 450 1150 470
rect 1210 450 1230 470
rect 1290 450 1310 470
rect 1370 450 1390 470
rect 1450 450 1470 470
rect 1530 450 1550 470
rect 1690 450 1710 470
rect 1770 450 1790 470
rect 1850 450 1870 470
rect 1930 450 1950 470
rect 2010 450 2030 470
rect 2090 450 2110 470
rect 2170 450 2190 470
rect 2250 450 2270 470
rect 2330 450 2350 470
rect 2410 450 2430 470
rect 2490 450 2510 470
rect 2650 450 2670 470
rect 2730 450 2750 470
rect 2810 450 2830 470
rect 2890 450 2910 470
rect 2970 450 2990 470
rect 3050 450 3070 470
rect 3130 450 3150 470
rect 3210 450 3230 470
rect 3290 450 3310 470
rect 3370 450 3390 470
rect 3450 450 3470 470
rect 3610 450 3630 470
rect 3690 450 3710 470
rect 3770 450 3790 470
rect 3850 450 3870 470
rect 3930 450 3950 470
rect 4090 450 4110 470
rect 270 205 1050 235
rect 1230 205 2010 235
rect 2190 205 2970 235
rect 3150 205 3930 235
rect 165 90 195 170
rect 1125 90 1155 170
rect 2085 90 2115 170
rect 3045 90 3075 170
rect 4005 90 4035 170
rect 90 -70 110 -50
rect 170 -70 190 -50
rect 250 -70 270 -50
rect 330 -70 350 -50
rect 410 -70 430 -50
rect 490 -70 510 -50
rect 570 -70 590 -50
rect 730 -70 750 -50
rect 810 -70 830 -50
rect 890 -70 910 -50
rect 970 -70 990 -50
rect 1050 -70 1070 -50
rect 1130 -70 1150 -50
rect 1210 -70 1230 -50
rect 1290 -70 1310 -50
rect 1370 -70 1390 -50
rect 1450 -70 1470 -50
rect 1530 -70 1550 -50
rect 1690 -70 1710 -50
rect 1770 -70 1790 -50
rect 1850 -70 1870 -50
rect 1930 -70 1950 -50
rect 2010 -70 2030 -50
rect 2090 -70 2110 -50
rect 2170 -70 2190 -50
rect 2250 -70 2270 -50
rect 2330 -70 2350 -50
rect 2410 -70 2430 -50
rect 2490 -70 2510 -50
rect 2650 -70 2670 -50
rect 2730 -70 2750 -50
rect 2810 -70 2830 -50
rect 2890 -70 2910 -50
rect 2970 -70 2990 -50
rect 3050 -70 3070 -50
rect 3130 -70 3150 -50
rect 3210 -70 3230 -50
rect 3290 -70 3310 -50
rect 3370 -70 3390 -50
rect 3450 -70 3470 -50
rect 3610 -70 3630 -50
rect 3690 -70 3710 -50
rect 3770 -70 3790 -50
rect 3850 -70 3870 -50
rect 3930 -70 3950 -50
rect 4090 -70 4110 -50
rect 270 -315 1050 -285
rect 1230 -315 2010 -285
rect 2190 -315 2970 -285
rect 3150 -315 3930 -285
rect 165 -430 195 -350
rect 1125 -430 1155 -350
rect 2085 -430 2115 -350
rect 3045 -430 3075 -350
rect 4005 -430 4035 -350
<< metal1 >>
rect 160 4870 200 4880
rect 160 4590 165 4870
rect 195 4590 200 4870
rect 160 4580 200 4590
rect 1120 4870 1160 4880
rect 1120 4590 1125 4870
rect 1155 4590 1160 4870
rect 1120 4580 1160 4590
rect 2080 4870 2120 4880
rect 2080 4590 2085 4870
rect 2115 4590 2120 4870
rect 2080 4580 2120 4590
rect 3040 4870 3080 4880
rect 3040 4590 3045 4870
rect 3075 4590 3080 4870
rect 3040 4580 3080 4590
rect 4000 4870 4040 4880
rect 4000 4590 4005 4870
rect 4035 4590 4040 4870
rect 260 4555 1060 4560
rect 260 4525 270 4555
rect 1050 4525 1060 4555
rect 260 4520 1060 4525
rect 1220 4555 2020 4560
rect 1220 4525 1230 4555
rect 2010 4525 2020 4555
rect 1220 4520 2020 4525
rect 2180 4555 2980 4560
rect 2180 4525 2190 4555
rect 2970 4525 2980 4555
rect 2180 4520 2980 4525
rect 3140 4555 3940 4560
rect 3140 4525 3150 4555
rect 3930 4525 3940 4555
rect 3140 4520 3940 4525
rect 640 4315 680 4520
rect 640 4285 645 4315
rect 675 4285 680 4315
rect 640 4280 680 4285
rect 1600 4315 1640 4520
rect 1600 4285 1605 4315
rect 1635 4285 1640 4315
rect 1600 4280 1640 4285
rect 2560 4315 2600 4520
rect 2560 4285 2565 4315
rect 2595 4285 2600 4315
rect 2560 4280 2600 4285
rect 3520 4315 3560 4520
rect 3520 4285 3525 4315
rect 3555 4285 3560 4315
rect 3520 4280 3560 4285
rect 4000 4315 4040 4590
rect 4000 4285 4005 4315
rect 4035 4285 4040 4315
rect 80 4235 120 4240
rect 80 4205 85 4235
rect 115 4205 120 4235
rect 80 4200 120 4205
rect 80 4155 120 4160
rect 80 4125 85 4155
rect 115 4125 120 4155
rect 80 4120 120 4125
rect 640 4075 680 4080
rect 640 4045 645 4075
rect 675 4045 680 4075
rect 640 3920 680 4045
rect 1600 4075 1640 4080
rect 1600 4045 1605 4075
rect 1635 4045 1640 4075
rect 1600 3920 1640 4045
rect 2560 4075 2600 4080
rect 2560 4045 2565 4075
rect 2595 4045 2600 4075
rect 2560 3920 2600 4045
rect 3520 4075 3560 4080
rect 3520 4045 3525 4075
rect 3555 4045 3560 4075
rect 3520 3920 3560 4045
rect 260 3915 1060 3920
rect 260 3885 270 3915
rect 1050 3885 1060 3915
rect 260 3880 1060 3885
rect 1220 3915 2020 3920
rect 1220 3885 1230 3915
rect 2010 3885 2020 3915
rect 1220 3880 2020 3885
rect 2180 3915 2980 3920
rect 2180 3885 2190 3915
rect 2970 3885 2980 3915
rect 2180 3880 2980 3885
rect 3140 3915 3940 3920
rect 3140 3885 3150 3915
rect 3930 3885 3940 3915
rect 3140 3880 3940 3885
rect 160 3850 200 3860
rect 160 3770 165 3850
rect 195 3770 200 3850
rect 160 3760 200 3770
rect 1120 3850 1160 3860
rect 1120 3770 1125 3850
rect 1155 3770 1160 3850
rect 1120 3760 1160 3770
rect 2080 3850 2120 3860
rect 2080 3770 2085 3850
rect 2115 3770 2120 3850
rect 2080 3760 2120 3770
rect 3040 3850 3080 3860
rect 3040 3770 3045 3850
rect 3075 3770 3080 3850
rect 3040 3760 3080 3770
rect 4000 3850 4040 4285
rect 4080 4235 4120 4240
rect 4080 4205 4085 4235
rect 4115 4205 4120 4235
rect 4080 4200 4120 4205
rect 4080 4155 4120 4160
rect 4080 4125 4085 4155
rect 4115 4125 4120 4155
rect 4080 4120 4120 4125
rect 4000 3770 4005 3850
rect 4035 3770 4040 3850
rect 4000 3760 4040 3770
rect 160 3550 200 3560
rect 160 3470 165 3550
rect 195 3470 200 3550
rect 160 3460 200 3470
rect 1120 3550 1160 3560
rect 1120 3470 1125 3550
rect 1155 3470 1160 3550
rect 1120 3460 1160 3470
rect 2080 3550 2120 3560
rect 2080 3470 2085 3550
rect 2115 3470 2120 3550
rect 2080 3460 2120 3470
rect 3040 3550 3080 3560
rect 3040 3470 3045 3550
rect 3075 3470 3080 3550
rect 3040 3460 3080 3470
rect 4000 3550 4040 3560
rect 4000 3470 4005 3550
rect 4035 3470 4040 3550
rect 260 3435 1060 3440
rect 260 3405 270 3435
rect 1050 3405 1060 3435
rect 260 3400 1060 3405
rect 1220 3435 2020 3440
rect 1220 3405 1230 3435
rect 2010 3405 2020 3435
rect 1220 3400 2020 3405
rect 2180 3435 2980 3440
rect 2180 3405 2190 3435
rect 2970 3405 2980 3435
rect 2180 3400 2980 3405
rect 3140 3435 3940 3440
rect 3140 3405 3150 3435
rect 3930 3405 3940 3435
rect 3140 3400 3940 3405
rect 640 3275 680 3400
rect 640 3245 645 3275
rect 675 3245 680 3275
rect 640 3240 680 3245
rect 1600 3275 1640 3400
rect 1600 3245 1605 3275
rect 1635 3245 1640 3275
rect 1600 3240 1640 3245
rect 2560 3275 2600 3400
rect 2560 3245 2565 3275
rect 2595 3245 2600 3275
rect 2560 3240 2600 3245
rect 3520 3275 3560 3400
rect 3520 3245 3525 3275
rect 3555 3245 3560 3275
rect 3520 3240 3560 3245
rect 80 3195 120 3200
rect 80 3165 85 3195
rect 115 3165 120 3195
rect 80 3160 120 3165
rect 80 3115 120 3120
rect 80 3085 85 3115
rect 115 3085 120 3115
rect 80 3080 120 3085
rect 4000 3035 4040 3470
rect 4080 3195 4120 3200
rect 4080 3165 4085 3195
rect 4115 3165 4120 3195
rect 4080 3160 4120 3165
rect 4080 3115 4120 3120
rect 4080 3085 4085 3115
rect 4115 3085 4120 3115
rect 4080 3080 4120 3085
rect 4000 3005 4005 3035
rect 4035 3005 4040 3035
rect 80 2955 120 2960
rect 80 2925 85 2955
rect 115 2925 120 2955
rect 80 2920 120 2925
rect 80 2875 120 2880
rect 80 2845 85 2875
rect 115 2845 120 2875
rect 80 2840 120 2845
rect 640 2795 680 2800
rect 640 2765 645 2795
rect 675 2765 680 2795
rect 640 2560 680 2765
rect 1600 2795 1640 2800
rect 1600 2765 1605 2795
rect 1635 2765 1640 2795
rect 1600 2560 1640 2765
rect 2560 2795 2600 2800
rect 2560 2765 2565 2795
rect 2595 2765 2600 2795
rect 2560 2560 2600 2765
rect 3520 2795 3560 2800
rect 3520 2765 3525 2795
rect 3555 2765 3560 2795
rect 3520 2560 3560 2765
rect 260 2555 1060 2560
rect 260 2525 270 2555
rect 1050 2525 1060 2555
rect 260 2520 1060 2525
rect 1220 2555 2020 2560
rect 1220 2525 1230 2555
rect 2010 2525 2020 2555
rect 1220 2520 2020 2525
rect 2180 2555 2980 2560
rect 2180 2525 2190 2555
rect 2970 2525 2980 2555
rect 2180 2520 2980 2525
rect 3140 2555 3940 2560
rect 3140 2525 3150 2555
rect 3930 2525 3940 2555
rect 3140 2520 3940 2525
rect 160 2490 200 2500
rect 160 2210 165 2490
rect 195 2210 200 2490
rect 160 2200 200 2210
rect 1120 2490 1160 2500
rect 1120 2210 1125 2490
rect 1155 2210 1160 2490
rect 1120 2200 1160 2210
rect 2080 2490 2120 2500
rect 2080 2210 2085 2490
rect 2115 2210 2120 2490
rect 2080 2200 2120 2210
rect 3040 2490 3080 2500
rect 3040 2210 3045 2490
rect 3075 2210 3080 2490
rect 3040 2200 3080 2210
rect 4000 2490 4040 3005
rect 4080 2955 4120 2960
rect 4080 2925 4085 2955
rect 4115 2925 4120 2955
rect 4080 2920 4120 2925
rect 4080 2875 4120 2880
rect 4080 2845 4085 2875
rect 4115 2845 4120 2875
rect 4080 2840 4120 2845
rect 4000 2210 4005 2490
rect 4035 2210 4040 2490
rect 4000 2200 4040 2210
rect 160 1830 200 1840
rect 160 1550 165 1830
rect 195 1550 200 1830
rect 0 1395 40 1400
rect 0 1365 5 1395
rect 35 1365 40 1395
rect 0 1235 40 1365
rect 0 1205 5 1235
rect 35 1205 40 1235
rect 0 1200 40 1205
rect 80 1395 120 1400
rect 80 1365 85 1395
rect 115 1365 120 1395
rect 80 1235 120 1365
rect 80 1205 85 1235
rect 115 1205 120 1235
rect 80 1200 120 1205
rect 160 1395 200 1550
rect 1120 1830 1160 1840
rect 1120 1550 1125 1830
rect 1155 1550 1160 1830
rect 1120 1540 1160 1550
rect 2080 1830 2120 1840
rect 2080 1550 2085 1830
rect 2115 1550 2120 1830
rect 2080 1540 2120 1550
rect 3040 1830 3080 1840
rect 3040 1550 3045 1830
rect 3075 1550 3080 1830
rect 3040 1540 3080 1550
rect 4000 1830 4040 1840
rect 4000 1550 4005 1830
rect 4035 1550 4040 1830
rect 4000 1540 4040 1550
rect 260 1515 1060 1520
rect 260 1485 270 1515
rect 1050 1485 1060 1515
rect 260 1480 1060 1485
rect 1220 1515 2020 1520
rect 1220 1485 1230 1515
rect 2010 1485 2020 1515
rect 1220 1480 2020 1485
rect 2180 1515 2980 1520
rect 2180 1485 2190 1515
rect 2970 1485 2980 1515
rect 2180 1480 2980 1485
rect 3140 1515 3940 1520
rect 3140 1485 3150 1515
rect 3930 1485 3940 1515
rect 3140 1480 3940 1485
rect 160 1365 165 1395
rect 195 1365 200 1395
rect 160 1235 200 1365
rect 160 1205 165 1235
rect 195 1205 200 1235
rect 160 1110 200 1205
rect 240 1395 280 1400
rect 240 1365 245 1395
rect 275 1365 280 1395
rect 240 1235 280 1365
rect 240 1205 245 1235
rect 275 1205 280 1235
rect 240 1200 280 1205
rect 320 1395 360 1400
rect 320 1365 325 1395
rect 355 1365 360 1395
rect 320 1235 360 1365
rect 320 1205 325 1235
rect 355 1205 360 1235
rect 320 1200 360 1205
rect 400 1395 440 1400
rect 400 1365 405 1395
rect 435 1365 440 1395
rect 400 1235 440 1365
rect 400 1205 405 1235
rect 435 1205 440 1235
rect 400 1200 440 1205
rect 480 1395 520 1400
rect 480 1365 485 1395
rect 515 1365 520 1395
rect 480 1235 520 1365
rect 480 1205 485 1235
rect 515 1205 520 1235
rect 480 1200 520 1205
rect 560 1395 600 1400
rect 560 1365 565 1395
rect 595 1365 600 1395
rect 560 1235 600 1365
rect 640 1315 680 1480
rect 640 1285 645 1315
rect 675 1285 680 1315
rect 640 1280 680 1285
rect 720 1395 760 1400
rect 720 1365 725 1395
rect 755 1365 760 1395
rect 560 1205 565 1235
rect 595 1205 600 1235
rect 560 1200 600 1205
rect 720 1235 760 1365
rect 720 1205 725 1235
rect 755 1205 760 1235
rect 720 1200 760 1205
rect 800 1395 840 1400
rect 800 1365 805 1395
rect 835 1365 840 1395
rect 800 1235 840 1365
rect 800 1205 805 1235
rect 835 1205 840 1235
rect 800 1200 840 1205
rect 880 1395 920 1400
rect 880 1365 885 1395
rect 915 1365 920 1395
rect 880 1235 920 1365
rect 880 1205 885 1235
rect 915 1205 920 1235
rect 880 1200 920 1205
rect 960 1395 1000 1400
rect 960 1365 965 1395
rect 995 1365 1000 1395
rect 960 1235 1000 1365
rect 960 1205 965 1235
rect 995 1205 1000 1235
rect 960 1200 1000 1205
rect 1040 1395 1080 1400
rect 1040 1365 1045 1395
rect 1075 1365 1080 1395
rect 1040 1235 1080 1365
rect 1040 1205 1045 1235
rect 1075 1205 1080 1235
rect 1040 1200 1080 1205
rect 1120 1395 1160 1400
rect 1120 1365 1125 1395
rect 1155 1365 1160 1395
rect 1120 1235 1160 1365
rect 1120 1205 1125 1235
rect 1155 1205 1160 1235
rect 1120 1200 1160 1205
rect 1200 1395 1240 1400
rect 1200 1365 1205 1395
rect 1235 1365 1240 1395
rect 1200 1235 1240 1365
rect 1200 1205 1205 1235
rect 1235 1205 1240 1235
rect 1200 1200 1240 1205
rect 1280 1395 1320 1400
rect 1280 1365 1285 1395
rect 1315 1365 1320 1395
rect 1280 1235 1320 1365
rect 1280 1205 1285 1235
rect 1315 1205 1320 1235
rect 1280 1200 1320 1205
rect 1360 1395 1400 1400
rect 1360 1365 1365 1395
rect 1395 1365 1400 1395
rect 1360 1235 1400 1365
rect 1360 1205 1365 1235
rect 1395 1205 1400 1235
rect 1360 1200 1400 1205
rect 1440 1395 1480 1400
rect 1440 1365 1445 1395
rect 1475 1365 1480 1395
rect 1440 1235 1480 1365
rect 1440 1205 1445 1235
rect 1475 1205 1480 1235
rect 1440 1200 1480 1205
rect 1520 1395 1560 1400
rect 1520 1365 1525 1395
rect 1555 1365 1560 1395
rect 1520 1235 1560 1365
rect 1600 1315 1640 1480
rect 1600 1285 1605 1315
rect 1635 1285 1640 1315
rect 1600 1280 1640 1285
rect 1680 1395 1720 1400
rect 1680 1365 1685 1395
rect 1715 1365 1720 1395
rect 1520 1205 1525 1235
rect 1555 1205 1560 1235
rect 1520 1200 1560 1205
rect 1680 1235 1720 1365
rect 1680 1205 1685 1235
rect 1715 1205 1720 1235
rect 1680 1200 1720 1205
rect 1760 1395 1800 1400
rect 1760 1365 1765 1395
rect 1795 1365 1800 1395
rect 1760 1235 1800 1365
rect 1760 1205 1765 1235
rect 1795 1205 1800 1235
rect 1760 1200 1800 1205
rect 1840 1395 1880 1400
rect 1840 1365 1845 1395
rect 1875 1365 1880 1395
rect 1840 1235 1880 1365
rect 1840 1205 1845 1235
rect 1875 1205 1880 1235
rect 1840 1200 1880 1205
rect 1920 1395 1960 1400
rect 1920 1365 1925 1395
rect 1955 1365 1960 1395
rect 1920 1235 1960 1365
rect 1920 1205 1925 1235
rect 1955 1205 1960 1235
rect 1920 1200 1960 1205
rect 2000 1395 2040 1400
rect 2000 1365 2005 1395
rect 2035 1365 2040 1395
rect 2000 1235 2040 1365
rect 2000 1205 2005 1235
rect 2035 1205 2040 1235
rect 2000 1200 2040 1205
rect 2080 1395 2120 1400
rect 2080 1365 2085 1395
rect 2115 1365 2120 1395
rect 2080 1235 2120 1365
rect 2080 1205 2085 1235
rect 2115 1205 2120 1235
rect 2080 1200 2120 1205
rect 2160 1395 2200 1400
rect 2160 1365 2165 1395
rect 2195 1365 2200 1395
rect 2160 1235 2200 1365
rect 2160 1205 2165 1235
rect 2195 1205 2200 1235
rect 2160 1200 2200 1205
rect 2240 1395 2280 1400
rect 2240 1365 2245 1395
rect 2275 1365 2280 1395
rect 2240 1235 2280 1365
rect 2240 1205 2245 1235
rect 2275 1205 2280 1235
rect 2240 1200 2280 1205
rect 2320 1395 2360 1400
rect 2320 1365 2325 1395
rect 2355 1365 2360 1395
rect 2320 1235 2360 1365
rect 2320 1205 2325 1235
rect 2355 1205 2360 1235
rect 2320 1200 2360 1205
rect 2400 1395 2440 1400
rect 2400 1365 2405 1395
rect 2435 1365 2440 1395
rect 2400 1235 2440 1365
rect 2400 1205 2405 1235
rect 2435 1205 2440 1235
rect 2400 1200 2440 1205
rect 2480 1395 2520 1400
rect 2480 1365 2485 1395
rect 2515 1365 2520 1395
rect 2480 1235 2520 1365
rect 2560 1315 2600 1480
rect 2560 1285 2565 1315
rect 2595 1285 2600 1315
rect 2560 1280 2600 1285
rect 2640 1395 2680 1400
rect 2640 1365 2645 1395
rect 2675 1365 2680 1395
rect 2480 1205 2485 1235
rect 2515 1205 2520 1235
rect 2480 1200 2520 1205
rect 2640 1235 2680 1365
rect 2640 1205 2645 1235
rect 2675 1205 2680 1235
rect 2640 1200 2680 1205
rect 2720 1395 2760 1400
rect 2720 1365 2725 1395
rect 2755 1365 2760 1395
rect 2720 1235 2760 1365
rect 2720 1205 2725 1235
rect 2755 1205 2760 1235
rect 2720 1200 2760 1205
rect 2800 1395 2840 1400
rect 2800 1365 2805 1395
rect 2835 1365 2840 1395
rect 2800 1235 2840 1365
rect 2800 1205 2805 1235
rect 2835 1205 2840 1235
rect 2800 1200 2840 1205
rect 2880 1395 2920 1400
rect 2880 1365 2885 1395
rect 2915 1365 2920 1395
rect 2880 1235 2920 1365
rect 2880 1205 2885 1235
rect 2915 1205 2920 1235
rect 2880 1200 2920 1205
rect 2960 1395 3000 1400
rect 2960 1365 2965 1395
rect 2995 1365 3000 1395
rect 2960 1235 3000 1365
rect 2960 1205 2965 1235
rect 2995 1205 3000 1235
rect 2960 1200 3000 1205
rect 3040 1395 3080 1400
rect 3040 1365 3045 1395
rect 3075 1365 3080 1395
rect 3040 1235 3080 1365
rect 3040 1205 3045 1235
rect 3075 1205 3080 1235
rect 3040 1200 3080 1205
rect 3120 1395 3160 1400
rect 3120 1365 3125 1395
rect 3155 1365 3160 1395
rect 3120 1235 3160 1365
rect 3120 1205 3125 1235
rect 3155 1205 3160 1235
rect 3120 1200 3160 1205
rect 3200 1395 3240 1400
rect 3200 1365 3205 1395
rect 3235 1365 3240 1395
rect 3200 1235 3240 1365
rect 3200 1205 3205 1235
rect 3235 1205 3240 1235
rect 3200 1200 3240 1205
rect 3280 1395 3320 1400
rect 3280 1365 3285 1395
rect 3315 1365 3320 1395
rect 3280 1235 3320 1365
rect 3280 1205 3285 1235
rect 3315 1205 3320 1235
rect 3280 1200 3320 1205
rect 3360 1395 3400 1400
rect 3360 1365 3365 1395
rect 3395 1365 3400 1395
rect 3360 1235 3400 1365
rect 3360 1205 3365 1235
rect 3395 1205 3400 1235
rect 3360 1200 3400 1205
rect 3440 1395 3480 1400
rect 3440 1365 3445 1395
rect 3475 1365 3480 1395
rect 3440 1235 3480 1365
rect 3520 1315 3560 1480
rect 3520 1285 3525 1315
rect 3555 1285 3560 1315
rect 3520 1280 3560 1285
rect 3600 1395 3640 1400
rect 3600 1365 3605 1395
rect 3635 1365 3640 1395
rect 3440 1205 3445 1235
rect 3475 1205 3480 1235
rect 3440 1200 3480 1205
rect 3600 1235 3640 1365
rect 3600 1205 3605 1235
rect 3635 1205 3640 1235
rect 3600 1200 3640 1205
rect 3680 1395 3720 1400
rect 3680 1365 3685 1395
rect 3715 1365 3720 1395
rect 3680 1235 3720 1365
rect 3680 1205 3685 1235
rect 3715 1205 3720 1235
rect 3680 1200 3720 1205
rect 3760 1395 3800 1400
rect 3760 1365 3765 1395
rect 3795 1365 3800 1395
rect 3760 1235 3800 1365
rect 3760 1205 3765 1235
rect 3795 1205 3800 1235
rect 3760 1200 3800 1205
rect 3840 1395 3880 1400
rect 3840 1365 3845 1395
rect 3875 1365 3880 1395
rect 3840 1235 3880 1365
rect 3840 1205 3845 1235
rect 3875 1205 3880 1235
rect 3840 1200 3880 1205
rect 3920 1395 3960 1400
rect 3920 1365 3925 1395
rect 3955 1365 3960 1395
rect 3920 1235 3960 1365
rect 3920 1205 3925 1235
rect 3955 1205 3960 1235
rect 3920 1200 3960 1205
rect 4000 1395 4040 1400
rect 4000 1365 4005 1395
rect 4035 1365 4040 1395
rect 4000 1235 4040 1365
rect 4000 1205 4005 1235
rect 4035 1205 4040 1235
rect 4000 1200 4040 1205
rect 4080 1395 4120 1400
rect 4080 1365 4085 1395
rect 4115 1365 4120 1395
rect 4080 1235 4120 1365
rect 4080 1205 4085 1235
rect 4115 1205 4120 1235
rect 4080 1200 4120 1205
rect 4160 1395 4200 1400
rect 4160 1365 4165 1395
rect 4195 1365 4200 1395
rect 4160 1235 4200 1365
rect 4160 1205 4165 1235
rect 4195 1205 4200 1235
rect 4160 1200 4200 1205
rect 160 830 165 1110
rect 195 830 200 1110
rect 160 820 200 830
rect 1120 1110 1160 1120
rect 1120 830 1125 1110
rect 1155 830 1160 1110
rect 1120 820 1160 830
rect 2080 1110 2120 1120
rect 2080 830 2085 1110
rect 2115 830 2120 1110
rect 2080 820 2120 830
rect 3040 1110 3080 1120
rect 3040 830 3045 1110
rect 3075 830 3080 1110
rect 3040 820 3080 830
rect 4000 1110 4040 1120
rect 4000 830 4005 1110
rect 4035 830 4040 1110
rect 260 795 1060 800
rect 260 765 270 795
rect 1050 765 1060 795
rect 260 760 1060 765
rect 1220 795 2020 800
rect 1220 765 1230 795
rect 2010 765 2020 795
rect 1220 760 2020 765
rect 2180 795 2980 800
rect 2180 765 2190 795
rect 2970 765 2980 795
rect 2180 760 2980 765
rect 3140 795 3940 800
rect 3140 765 3150 795
rect 3930 765 3940 795
rect 3140 760 3940 765
rect 640 555 680 760
rect 640 525 645 555
rect 675 525 680 555
rect 80 475 120 480
rect 80 445 85 475
rect 115 445 120 475
rect 80 440 120 445
rect 160 470 200 480
rect 160 450 170 470
rect 190 450 200 470
rect 160 440 200 450
rect 240 470 280 480
rect 240 450 250 470
rect 270 450 280 470
rect 240 440 280 450
rect 320 470 360 480
rect 320 450 330 470
rect 350 450 360 470
rect 320 440 360 450
rect 400 470 440 480
rect 400 450 410 470
rect 430 450 440 470
rect 400 440 440 450
rect 480 470 520 480
rect 480 450 490 470
rect 510 450 520 470
rect 480 440 520 450
rect 560 470 600 480
rect 560 450 570 470
rect 590 450 600 470
rect 560 440 600 450
rect 640 240 680 525
rect 1600 555 1640 760
rect 1600 525 1605 555
rect 1635 525 1640 555
rect 720 470 760 480
rect 720 450 730 470
rect 750 450 760 470
rect 720 440 760 450
rect 800 470 840 480
rect 800 450 810 470
rect 830 450 840 470
rect 800 440 840 450
rect 880 470 920 480
rect 880 450 890 470
rect 910 450 920 470
rect 880 440 920 450
rect 960 470 1000 480
rect 960 450 970 470
rect 990 450 1000 470
rect 960 440 1000 450
rect 1040 470 1080 480
rect 1040 450 1050 470
rect 1070 450 1080 470
rect 1040 440 1080 450
rect 1120 470 1160 480
rect 1120 450 1130 470
rect 1150 450 1160 470
rect 1120 440 1160 450
rect 1200 470 1240 480
rect 1200 450 1210 470
rect 1230 450 1240 470
rect 1200 440 1240 450
rect 1280 470 1320 480
rect 1280 450 1290 470
rect 1310 450 1320 470
rect 1280 440 1320 450
rect 1360 470 1400 480
rect 1360 450 1370 470
rect 1390 450 1400 470
rect 1360 440 1400 450
rect 1440 470 1480 480
rect 1440 450 1450 470
rect 1470 450 1480 470
rect 1440 440 1480 450
rect 1520 470 1560 480
rect 1520 450 1530 470
rect 1550 450 1560 470
rect 1520 440 1560 450
rect 1600 240 1640 525
rect 2560 555 2600 760
rect 2560 525 2565 555
rect 2595 525 2600 555
rect 1680 470 1720 480
rect 1680 450 1690 470
rect 1710 450 1720 470
rect 1680 440 1720 450
rect 1760 470 1800 480
rect 1760 450 1770 470
rect 1790 450 1800 470
rect 1760 440 1800 450
rect 1840 470 1880 480
rect 1840 450 1850 470
rect 1870 450 1880 470
rect 1840 440 1880 450
rect 1920 470 1960 480
rect 1920 450 1930 470
rect 1950 450 1960 470
rect 1920 440 1960 450
rect 2000 470 2040 480
rect 2000 450 2010 470
rect 2030 450 2040 470
rect 2000 440 2040 450
rect 2080 470 2120 480
rect 2080 450 2090 470
rect 2110 450 2120 470
rect 2080 440 2120 450
rect 2160 470 2200 480
rect 2160 450 2170 470
rect 2190 450 2200 470
rect 2160 440 2200 450
rect 2240 470 2280 480
rect 2240 450 2250 470
rect 2270 450 2280 470
rect 2240 440 2280 450
rect 2320 470 2360 480
rect 2320 450 2330 470
rect 2350 450 2360 470
rect 2320 440 2360 450
rect 2400 470 2440 480
rect 2400 450 2410 470
rect 2430 450 2440 470
rect 2400 440 2440 450
rect 2480 470 2520 480
rect 2480 450 2490 470
rect 2510 450 2520 470
rect 2480 440 2520 450
rect 2560 240 2600 525
rect 3520 555 3560 760
rect 3520 525 3525 555
rect 3555 525 3560 555
rect 2640 470 2680 480
rect 2640 450 2650 470
rect 2670 450 2680 470
rect 2640 440 2680 450
rect 2720 470 2760 480
rect 2720 450 2730 470
rect 2750 450 2760 470
rect 2720 440 2760 450
rect 2800 470 2840 480
rect 2800 450 2810 470
rect 2830 450 2840 470
rect 2800 440 2840 450
rect 2880 470 2920 480
rect 2880 450 2890 470
rect 2910 450 2920 470
rect 2880 440 2920 450
rect 2960 470 3000 480
rect 2960 450 2970 470
rect 2990 450 3000 470
rect 2960 440 3000 450
rect 3040 470 3080 480
rect 3040 450 3050 470
rect 3070 450 3080 470
rect 3040 440 3080 450
rect 3120 470 3160 480
rect 3120 450 3130 470
rect 3150 450 3160 470
rect 3120 440 3160 450
rect 3200 470 3240 480
rect 3200 450 3210 470
rect 3230 450 3240 470
rect 3200 440 3240 450
rect 3280 470 3320 480
rect 3280 450 3290 470
rect 3310 450 3320 470
rect 3280 440 3320 450
rect 3360 470 3400 480
rect 3360 450 3370 470
rect 3390 450 3400 470
rect 3360 440 3400 450
rect 3440 470 3480 480
rect 3440 450 3450 470
rect 3470 450 3480 470
rect 3440 440 3480 450
rect 3520 240 3560 525
rect 4000 555 4040 830
rect 4000 525 4005 555
rect 4035 525 4040 555
rect 3600 470 3640 480
rect 3600 450 3610 470
rect 3630 450 3640 470
rect 3600 440 3640 450
rect 3680 470 3720 480
rect 3680 450 3690 470
rect 3710 450 3720 470
rect 3680 440 3720 450
rect 3760 470 3800 480
rect 3760 450 3770 470
rect 3790 450 3800 470
rect 3760 440 3800 450
rect 3840 470 3880 480
rect 3840 450 3850 470
rect 3870 450 3880 470
rect 3840 440 3880 450
rect 3920 470 3960 480
rect 3920 450 3930 470
rect 3950 450 3960 470
rect 3920 440 3960 450
rect 4000 395 4040 525
rect 4080 470 4120 480
rect 4080 450 4090 470
rect 4110 450 4120 470
rect 4080 440 4120 450
rect 4000 365 4005 395
rect 4035 365 4040 395
rect 260 235 1060 240
rect 260 205 270 235
rect 1050 205 1060 235
rect 260 200 1060 205
rect 1220 235 2020 240
rect 1220 205 1230 235
rect 2010 205 2020 235
rect 1220 200 2020 205
rect 2180 235 2980 240
rect 2180 205 2190 235
rect 2970 205 2980 235
rect 2180 200 2980 205
rect 3140 235 3940 240
rect 3140 205 3150 235
rect 3930 205 3940 235
rect 3140 200 3940 205
rect 160 170 200 180
rect 160 90 165 170
rect 195 90 200 170
rect 160 80 200 90
rect 1120 170 1160 180
rect 1120 90 1125 170
rect 1155 90 1160 170
rect 1120 80 1160 90
rect 2080 170 2120 180
rect 2080 90 2085 170
rect 2115 90 2120 170
rect 2080 80 2120 90
rect 3040 170 3080 180
rect 3040 90 3045 170
rect 3075 90 3080 170
rect 3040 80 3080 90
rect 4000 170 4040 365
rect 4000 90 4005 170
rect 4035 90 4040 170
rect 4000 80 4040 90
rect 80 -45 120 -40
rect 80 -75 85 -45
rect 115 -75 120 -45
rect 80 -80 120 -75
rect 160 -45 200 -40
rect 160 -75 165 -45
rect 195 -75 200 -45
rect 160 -80 200 -75
rect 240 -45 280 -40
rect 240 -75 245 -45
rect 275 -75 280 -45
rect 240 -80 280 -75
rect 320 -45 360 -40
rect 320 -75 325 -45
rect 355 -75 360 -45
rect 320 -80 360 -75
rect 400 -45 440 -40
rect 400 -75 405 -45
rect 435 -75 440 -45
rect 400 -80 440 -75
rect 480 -45 520 -40
rect 480 -75 485 -45
rect 515 -75 520 -45
rect 480 -80 520 -75
rect 560 -45 600 -40
rect 560 -75 565 -45
rect 595 -75 600 -45
rect 560 -80 600 -75
rect 720 -45 760 -40
rect 720 -75 725 -45
rect 755 -75 760 -45
rect 720 -80 760 -75
rect 800 -45 840 -40
rect 800 -75 805 -45
rect 835 -75 840 -45
rect 800 -80 840 -75
rect 880 -45 920 -40
rect 880 -75 885 -45
rect 915 -75 920 -45
rect 880 -80 920 -75
rect 960 -45 1000 -40
rect 960 -75 965 -45
rect 995 -75 1000 -45
rect 960 -80 1000 -75
rect 1040 -45 1080 -40
rect 1040 -75 1045 -45
rect 1075 -75 1080 -45
rect 1040 -80 1080 -75
rect 1120 -45 1160 -40
rect 1120 -75 1125 -45
rect 1155 -75 1160 -45
rect 1120 -80 1160 -75
rect 1200 -45 1240 -40
rect 1200 -75 1205 -45
rect 1235 -75 1240 -45
rect 1200 -80 1240 -75
rect 1280 -45 1320 -40
rect 1280 -75 1285 -45
rect 1315 -75 1320 -45
rect 1280 -80 1320 -75
rect 1360 -45 1400 -40
rect 1360 -75 1365 -45
rect 1395 -75 1400 -45
rect 1360 -80 1400 -75
rect 1440 -45 1480 -40
rect 1440 -75 1445 -45
rect 1475 -75 1480 -45
rect 1440 -80 1480 -75
rect 1520 -45 1560 -40
rect 1520 -75 1525 -45
rect 1555 -75 1560 -45
rect 1520 -80 1560 -75
rect 1680 -45 1720 -40
rect 1680 -75 1685 -45
rect 1715 -75 1720 -45
rect 1680 -80 1720 -75
rect 1760 -45 1800 -40
rect 1760 -75 1765 -45
rect 1795 -75 1800 -45
rect 1760 -80 1800 -75
rect 1840 -45 1880 -40
rect 1840 -75 1845 -45
rect 1875 -75 1880 -45
rect 1840 -80 1880 -75
rect 1920 -45 1960 -40
rect 1920 -75 1925 -45
rect 1955 -75 1960 -45
rect 1920 -80 1960 -75
rect 2000 -45 2040 -40
rect 2000 -75 2005 -45
rect 2035 -75 2040 -45
rect 2000 -80 2040 -75
rect 2080 -45 2120 -40
rect 2080 -75 2085 -45
rect 2115 -75 2120 -45
rect 2080 -80 2120 -75
rect 2160 -45 2200 -40
rect 2160 -75 2165 -45
rect 2195 -75 2200 -45
rect 2160 -80 2200 -75
rect 2240 -45 2280 -40
rect 2240 -75 2245 -45
rect 2275 -75 2280 -45
rect 2240 -80 2280 -75
rect 2320 -45 2360 -40
rect 2320 -75 2325 -45
rect 2355 -75 2360 -45
rect 2320 -80 2360 -75
rect 2400 -45 2440 -40
rect 2400 -75 2405 -45
rect 2435 -75 2440 -45
rect 2400 -80 2440 -75
rect 2480 -45 2520 -40
rect 2480 -75 2485 -45
rect 2515 -75 2520 -45
rect 2480 -80 2520 -75
rect 2640 -45 2680 -40
rect 2640 -75 2645 -45
rect 2675 -75 2680 -45
rect 2640 -80 2680 -75
rect 2720 -45 2760 -40
rect 2720 -75 2725 -45
rect 2755 -75 2760 -45
rect 2720 -80 2760 -75
rect 2800 -45 2840 -40
rect 2800 -75 2805 -45
rect 2835 -75 2840 -45
rect 2800 -80 2840 -75
rect 2880 -45 2920 -40
rect 2880 -75 2885 -45
rect 2915 -75 2920 -45
rect 2880 -80 2920 -75
rect 2960 -45 3000 -40
rect 2960 -75 2965 -45
rect 2995 -75 3000 -45
rect 2960 -80 3000 -75
rect 3040 -45 3080 -40
rect 3040 -75 3045 -45
rect 3075 -75 3080 -45
rect 3040 -80 3080 -75
rect 3120 -45 3160 -40
rect 3120 -75 3125 -45
rect 3155 -75 3160 -45
rect 3120 -80 3160 -75
rect 3200 -45 3240 -40
rect 3200 -75 3205 -45
rect 3235 -75 3240 -45
rect 3200 -80 3240 -75
rect 3280 -45 3320 -40
rect 3280 -75 3285 -45
rect 3315 -75 3320 -45
rect 3280 -80 3320 -75
rect 3360 -45 3400 -40
rect 3360 -75 3365 -45
rect 3395 -75 3400 -45
rect 3360 -80 3400 -75
rect 3440 -45 3480 -40
rect 3440 -75 3445 -45
rect 3475 -75 3480 -45
rect 3440 -80 3480 -75
rect 3600 -45 3640 -40
rect 3600 -75 3605 -45
rect 3635 -75 3640 -45
rect 3600 -80 3640 -75
rect 3680 -45 3720 -40
rect 3680 -75 3685 -45
rect 3715 -75 3720 -45
rect 3680 -80 3720 -75
rect 3760 -45 3800 -40
rect 3760 -75 3765 -45
rect 3795 -75 3800 -45
rect 3760 -80 3800 -75
rect 3840 -45 3880 -40
rect 3840 -75 3845 -45
rect 3875 -75 3880 -45
rect 3840 -80 3880 -75
rect 3920 -45 3960 -40
rect 3920 -75 3925 -45
rect 3955 -75 3960 -45
rect 3920 -80 3960 -75
rect 4080 -45 4120 -40
rect 4080 -75 4085 -45
rect 4115 -75 4120 -45
rect 4080 -80 4120 -75
rect 640 -125 680 -120
rect 640 -155 645 -125
rect 675 -155 680 -125
rect 640 -280 680 -155
rect 1600 -125 1640 -120
rect 1600 -155 1605 -125
rect 1635 -155 1640 -125
rect 1600 -280 1640 -155
rect 2560 -125 2600 -120
rect 2560 -155 2565 -125
rect 2595 -155 2600 -125
rect 2560 -280 2600 -155
rect 3520 -125 3560 -120
rect 3520 -155 3525 -125
rect 3555 -155 3560 -125
rect 3520 -280 3560 -155
rect 4000 -125 4040 -120
rect 4000 -155 4005 -125
rect 4035 -155 4040 -125
rect 260 -285 1060 -280
rect 260 -315 270 -285
rect 1050 -315 1060 -285
rect 260 -320 1060 -315
rect 1220 -285 2020 -280
rect 1220 -315 1230 -285
rect 2010 -315 2020 -285
rect 1220 -320 2020 -315
rect 2180 -285 2980 -280
rect 2180 -315 2190 -285
rect 2970 -315 2980 -285
rect 2180 -320 2980 -315
rect 3140 -285 3940 -280
rect 3140 -315 3150 -285
rect 3930 -315 3940 -285
rect 3140 -320 3940 -315
rect 160 -350 200 -340
rect 160 -430 165 -350
rect 195 -430 200 -350
rect 160 -440 200 -430
rect 1120 -350 1160 -340
rect 1120 -430 1125 -350
rect 1155 -430 1160 -350
rect 1120 -440 1160 -430
rect 2080 -350 2120 -340
rect 2080 -430 2085 -350
rect 2115 -430 2120 -350
rect 2080 -440 2120 -430
rect 3040 -350 3080 -340
rect 3040 -430 3045 -350
rect 3075 -430 3080 -350
rect 3040 -440 3080 -430
rect 4000 -350 4040 -155
rect 4000 -430 4005 -350
rect 4035 -430 4040 -350
rect 4000 -440 4040 -430
<< via1 >>
rect 165 4690 195 4870
rect 645 4285 675 4315
rect 1605 4285 1635 4315
rect 2565 4285 2595 4315
rect 3525 4285 3555 4315
rect 4005 4285 4035 4315
rect 85 4230 115 4235
rect 85 4210 90 4230
rect 90 4210 110 4230
rect 110 4210 115 4230
rect 85 4205 115 4210
rect 85 4150 115 4155
rect 85 4130 90 4150
rect 90 4130 110 4150
rect 110 4130 115 4150
rect 85 4125 115 4130
rect 645 4045 675 4075
rect 1605 4045 1635 4075
rect 2565 4045 2595 4075
rect 3525 4045 3555 4075
rect 165 3770 195 3850
rect 4085 4230 4115 4235
rect 4085 4210 4090 4230
rect 4090 4210 4110 4230
rect 4110 4210 4115 4230
rect 4085 4205 4115 4210
rect 4085 4150 4115 4155
rect 4085 4130 4090 4150
rect 4090 4130 4110 4150
rect 4110 4130 4115 4150
rect 4085 4125 4115 4130
rect 165 3470 195 3550
rect 645 3245 675 3275
rect 1605 3245 1635 3275
rect 2565 3245 2595 3275
rect 3525 3245 3555 3275
rect 85 3190 115 3195
rect 85 3170 90 3190
rect 90 3170 110 3190
rect 110 3170 115 3190
rect 85 3165 115 3170
rect 85 3110 115 3115
rect 85 3090 90 3110
rect 90 3090 110 3110
rect 110 3090 115 3110
rect 85 3085 115 3090
rect 4085 3190 4115 3195
rect 4085 3170 4090 3190
rect 4090 3170 4110 3190
rect 4110 3170 4115 3190
rect 4085 3165 4115 3170
rect 4085 3110 4115 3115
rect 4085 3090 4090 3110
rect 4090 3090 4110 3110
rect 4110 3090 4115 3110
rect 4085 3085 4115 3090
rect 4005 3005 4035 3035
rect 85 2950 115 2955
rect 85 2930 90 2950
rect 90 2930 110 2950
rect 110 2930 115 2950
rect 85 2925 115 2930
rect 85 2870 115 2875
rect 85 2850 90 2870
rect 90 2850 110 2870
rect 110 2850 115 2870
rect 85 2845 115 2850
rect 645 2765 675 2795
rect 1605 2765 1635 2795
rect 2565 2765 2595 2795
rect 3525 2765 3555 2795
rect 165 2210 195 2390
rect 4085 2950 4115 2955
rect 4085 2930 4090 2950
rect 4090 2930 4110 2950
rect 4110 2930 4115 2950
rect 4085 2925 4115 2930
rect 4085 2870 4115 2875
rect 4085 2850 4090 2870
rect 4090 2850 4110 2870
rect 4110 2850 4115 2870
rect 4085 2845 4115 2850
rect 5 1365 35 1395
rect 5 1205 35 1235
rect 85 1365 115 1395
rect 85 1205 115 1235
rect 4005 1650 4035 1830
rect 165 1365 195 1395
rect 165 1205 195 1235
rect 245 1365 275 1395
rect 245 1205 275 1235
rect 325 1365 355 1395
rect 325 1205 355 1235
rect 405 1365 435 1395
rect 405 1205 435 1235
rect 485 1365 515 1395
rect 485 1205 515 1235
rect 565 1365 595 1395
rect 645 1285 675 1315
rect 725 1365 755 1395
rect 565 1205 595 1235
rect 725 1205 755 1235
rect 805 1365 835 1395
rect 805 1205 835 1235
rect 885 1365 915 1395
rect 885 1205 915 1235
rect 965 1365 995 1395
rect 965 1205 995 1235
rect 1045 1365 1075 1395
rect 1045 1205 1075 1235
rect 1125 1365 1155 1395
rect 1125 1205 1155 1235
rect 1205 1365 1235 1395
rect 1205 1205 1235 1235
rect 1285 1365 1315 1395
rect 1285 1205 1315 1235
rect 1365 1365 1395 1395
rect 1365 1205 1395 1235
rect 1445 1365 1475 1395
rect 1445 1205 1475 1235
rect 1525 1365 1555 1395
rect 1605 1285 1635 1315
rect 1685 1365 1715 1395
rect 1525 1205 1555 1235
rect 1685 1205 1715 1235
rect 1765 1365 1795 1395
rect 1765 1205 1795 1235
rect 1845 1365 1875 1395
rect 1845 1205 1875 1235
rect 1925 1365 1955 1395
rect 1925 1205 1955 1235
rect 2005 1365 2035 1395
rect 2005 1205 2035 1235
rect 2085 1365 2115 1395
rect 2085 1205 2115 1235
rect 2165 1365 2195 1395
rect 2165 1205 2195 1235
rect 2245 1365 2275 1395
rect 2245 1205 2275 1235
rect 2325 1365 2355 1395
rect 2325 1205 2355 1235
rect 2405 1365 2435 1395
rect 2405 1205 2435 1235
rect 2485 1365 2515 1395
rect 2565 1285 2595 1315
rect 2645 1365 2675 1395
rect 2485 1205 2515 1235
rect 2645 1205 2675 1235
rect 2725 1365 2755 1395
rect 2725 1205 2755 1235
rect 2805 1365 2835 1395
rect 2805 1205 2835 1235
rect 2885 1365 2915 1395
rect 2885 1205 2915 1235
rect 2965 1365 2995 1395
rect 2965 1205 2995 1235
rect 3045 1365 3075 1395
rect 3045 1205 3075 1235
rect 3125 1365 3155 1395
rect 3125 1205 3155 1235
rect 3205 1365 3235 1395
rect 3205 1205 3235 1235
rect 3285 1365 3315 1395
rect 3285 1205 3315 1235
rect 3365 1365 3395 1395
rect 3365 1205 3395 1235
rect 3445 1365 3475 1395
rect 3525 1285 3555 1315
rect 3605 1365 3635 1395
rect 3445 1205 3475 1235
rect 3605 1205 3635 1235
rect 3685 1365 3715 1395
rect 3685 1205 3715 1235
rect 3765 1365 3795 1395
rect 3765 1205 3795 1235
rect 3845 1365 3875 1395
rect 3845 1205 3875 1235
rect 3925 1365 3955 1395
rect 3925 1205 3955 1235
rect 4005 1365 4035 1395
rect 4005 1205 4035 1235
rect 4085 1365 4115 1395
rect 4085 1205 4115 1235
rect 4165 1365 4195 1395
rect 4165 1205 4195 1235
rect 645 525 675 555
rect 85 470 115 475
rect 85 450 90 470
rect 90 450 110 470
rect 110 450 115 470
rect 85 445 115 450
rect 1605 525 1635 555
rect 2565 525 2595 555
rect 3525 525 3555 555
rect 4005 525 4035 555
rect 4005 365 4035 395
rect 165 90 195 170
rect 85 -50 115 -45
rect 85 -70 90 -50
rect 90 -70 110 -50
rect 110 -70 115 -50
rect 85 -75 115 -70
rect 165 -50 195 -45
rect 165 -70 170 -50
rect 170 -70 190 -50
rect 190 -70 195 -50
rect 165 -75 195 -70
rect 245 -50 275 -45
rect 245 -70 250 -50
rect 250 -70 270 -50
rect 270 -70 275 -50
rect 245 -75 275 -70
rect 325 -50 355 -45
rect 325 -70 330 -50
rect 330 -70 350 -50
rect 350 -70 355 -50
rect 325 -75 355 -70
rect 405 -50 435 -45
rect 405 -70 410 -50
rect 410 -70 430 -50
rect 430 -70 435 -50
rect 405 -75 435 -70
rect 485 -50 515 -45
rect 485 -70 490 -50
rect 490 -70 510 -50
rect 510 -70 515 -50
rect 485 -75 515 -70
rect 565 -50 595 -45
rect 565 -70 570 -50
rect 570 -70 590 -50
rect 590 -70 595 -50
rect 565 -75 595 -70
rect 725 -50 755 -45
rect 725 -70 730 -50
rect 730 -70 750 -50
rect 750 -70 755 -50
rect 725 -75 755 -70
rect 805 -50 835 -45
rect 805 -70 810 -50
rect 810 -70 830 -50
rect 830 -70 835 -50
rect 805 -75 835 -70
rect 885 -50 915 -45
rect 885 -70 890 -50
rect 890 -70 910 -50
rect 910 -70 915 -50
rect 885 -75 915 -70
rect 965 -50 995 -45
rect 965 -70 970 -50
rect 970 -70 990 -50
rect 990 -70 995 -50
rect 965 -75 995 -70
rect 1045 -50 1075 -45
rect 1045 -70 1050 -50
rect 1050 -70 1070 -50
rect 1070 -70 1075 -50
rect 1045 -75 1075 -70
rect 1125 -50 1155 -45
rect 1125 -70 1130 -50
rect 1130 -70 1150 -50
rect 1150 -70 1155 -50
rect 1125 -75 1155 -70
rect 1205 -50 1235 -45
rect 1205 -70 1210 -50
rect 1210 -70 1230 -50
rect 1230 -70 1235 -50
rect 1205 -75 1235 -70
rect 1285 -50 1315 -45
rect 1285 -70 1290 -50
rect 1290 -70 1310 -50
rect 1310 -70 1315 -50
rect 1285 -75 1315 -70
rect 1365 -50 1395 -45
rect 1365 -70 1370 -50
rect 1370 -70 1390 -50
rect 1390 -70 1395 -50
rect 1365 -75 1395 -70
rect 1445 -50 1475 -45
rect 1445 -70 1450 -50
rect 1450 -70 1470 -50
rect 1470 -70 1475 -50
rect 1445 -75 1475 -70
rect 1525 -50 1555 -45
rect 1525 -70 1530 -50
rect 1530 -70 1550 -50
rect 1550 -70 1555 -50
rect 1525 -75 1555 -70
rect 1685 -50 1715 -45
rect 1685 -70 1690 -50
rect 1690 -70 1710 -50
rect 1710 -70 1715 -50
rect 1685 -75 1715 -70
rect 1765 -50 1795 -45
rect 1765 -70 1770 -50
rect 1770 -70 1790 -50
rect 1790 -70 1795 -50
rect 1765 -75 1795 -70
rect 1845 -50 1875 -45
rect 1845 -70 1850 -50
rect 1850 -70 1870 -50
rect 1870 -70 1875 -50
rect 1845 -75 1875 -70
rect 1925 -50 1955 -45
rect 1925 -70 1930 -50
rect 1930 -70 1950 -50
rect 1950 -70 1955 -50
rect 1925 -75 1955 -70
rect 2005 -50 2035 -45
rect 2005 -70 2010 -50
rect 2010 -70 2030 -50
rect 2030 -70 2035 -50
rect 2005 -75 2035 -70
rect 2085 -50 2115 -45
rect 2085 -70 2090 -50
rect 2090 -70 2110 -50
rect 2110 -70 2115 -50
rect 2085 -75 2115 -70
rect 2165 -50 2195 -45
rect 2165 -70 2170 -50
rect 2170 -70 2190 -50
rect 2190 -70 2195 -50
rect 2165 -75 2195 -70
rect 2245 -50 2275 -45
rect 2245 -70 2250 -50
rect 2250 -70 2270 -50
rect 2270 -70 2275 -50
rect 2245 -75 2275 -70
rect 2325 -50 2355 -45
rect 2325 -70 2330 -50
rect 2330 -70 2350 -50
rect 2350 -70 2355 -50
rect 2325 -75 2355 -70
rect 2405 -50 2435 -45
rect 2405 -70 2410 -50
rect 2410 -70 2430 -50
rect 2430 -70 2435 -50
rect 2405 -75 2435 -70
rect 2485 -50 2515 -45
rect 2485 -70 2490 -50
rect 2490 -70 2510 -50
rect 2510 -70 2515 -50
rect 2485 -75 2515 -70
rect 2645 -50 2675 -45
rect 2645 -70 2650 -50
rect 2650 -70 2670 -50
rect 2670 -70 2675 -50
rect 2645 -75 2675 -70
rect 2725 -50 2755 -45
rect 2725 -70 2730 -50
rect 2730 -70 2750 -50
rect 2750 -70 2755 -50
rect 2725 -75 2755 -70
rect 2805 -50 2835 -45
rect 2805 -70 2810 -50
rect 2810 -70 2830 -50
rect 2830 -70 2835 -50
rect 2805 -75 2835 -70
rect 2885 -50 2915 -45
rect 2885 -70 2890 -50
rect 2890 -70 2910 -50
rect 2910 -70 2915 -50
rect 2885 -75 2915 -70
rect 2965 -50 2995 -45
rect 2965 -70 2970 -50
rect 2970 -70 2990 -50
rect 2990 -70 2995 -50
rect 2965 -75 2995 -70
rect 3045 -50 3075 -45
rect 3045 -70 3050 -50
rect 3050 -70 3070 -50
rect 3070 -70 3075 -50
rect 3045 -75 3075 -70
rect 3125 -50 3155 -45
rect 3125 -70 3130 -50
rect 3130 -70 3150 -50
rect 3150 -70 3155 -50
rect 3125 -75 3155 -70
rect 3205 -50 3235 -45
rect 3205 -70 3210 -50
rect 3210 -70 3230 -50
rect 3230 -70 3235 -50
rect 3205 -75 3235 -70
rect 3285 -50 3315 -45
rect 3285 -70 3290 -50
rect 3290 -70 3310 -50
rect 3310 -70 3315 -50
rect 3285 -75 3315 -70
rect 3365 -50 3395 -45
rect 3365 -70 3370 -50
rect 3370 -70 3390 -50
rect 3390 -70 3395 -50
rect 3365 -75 3395 -70
rect 3445 -50 3475 -45
rect 3445 -70 3450 -50
rect 3450 -70 3470 -50
rect 3470 -70 3475 -50
rect 3445 -75 3475 -70
rect 3605 -50 3635 -45
rect 3605 -70 3610 -50
rect 3610 -70 3630 -50
rect 3630 -70 3635 -50
rect 3605 -75 3635 -70
rect 3685 -50 3715 -45
rect 3685 -70 3690 -50
rect 3690 -70 3710 -50
rect 3710 -70 3715 -50
rect 3685 -75 3715 -70
rect 3765 -50 3795 -45
rect 3765 -70 3770 -50
rect 3770 -70 3790 -50
rect 3790 -70 3795 -50
rect 3765 -75 3795 -70
rect 3845 -50 3875 -45
rect 3845 -70 3850 -50
rect 3850 -70 3870 -50
rect 3870 -70 3875 -50
rect 3845 -75 3875 -70
rect 3925 -50 3955 -45
rect 3925 -70 3930 -50
rect 3930 -70 3950 -50
rect 3950 -70 3955 -50
rect 3925 -75 3955 -70
rect 4085 -50 4115 -45
rect 4085 -70 4090 -50
rect 4090 -70 4110 -50
rect 4110 -70 4115 -50
rect 4085 -75 4115 -70
rect 645 -155 675 -125
rect 1605 -155 1635 -125
rect 2565 -155 2595 -125
rect 3525 -155 3555 -125
rect 4005 -155 4035 -125
rect 165 -430 195 -350
<< metal2 >>
rect 160 4870 200 4880
rect 160 4690 165 4870
rect 195 4690 200 4870
rect 160 4680 200 4690
rect 0 4395 4200 4400
rect 0 4365 85 4395
rect 115 4365 165 4395
rect 195 4365 245 4395
rect 275 4365 325 4395
rect 355 4365 405 4395
rect 435 4365 485 4395
rect 515 4365 565 4395
rect 595 4365 725 4395
rect 755 4365 805 4395
rect 835 4365 885 4395
rect 915 4365 965 4395
rect 995 4365 1045 4395
rect 1075 4365 1125 4395
rect 1155 4365 1205 4395
rect 1235 4365 1285 4395
rect 1315 4365 1365 4395
rect 1395 4365 1445 4395
rect 1475 4365 1525 4395
rect 1555 4365 1685 4395
rect 1715 4365 1765 4395
rect 1795 4365 1845 4395
rect 1875 4365 1925 4395
rect 1955 4365 2005 4395
rect 2035 4365 2085 4395
rect 2115 4365 2165 4395
rect 2195 4365 2245 4395
rect 2275 4365 2325 4395
rect 2355 4365 2405 4395
rect 2435 4365 2485 4395
rect 2515 4365 2645 4395
rect 2675 4365 2725 4395
rect 2755 4365 2805 4395
rect 2835 4365 2885 4395
rect 2915 4365 2965 4395
rect 2995 4365 3045 4395
rect 3075 4365 3125 4395
rect 3155 4365 3205 4395
rect 3235 4365 3285 4395
rect 3315 4365 3365 4395
rect 3395 4365 3445 4395
rect 3475 4365 3605 4395
rect 3635 4365 3685 4395
rect 3715 4365 3765 4395
rect 3795 4365 3845 4395
rect 3875 4365 3925 4395
rect 3955 4365 4005 4395
rect 4035 4365 4085 4395
rect 4115 4365 4200 4395
rect 0 4360 4200 4365
rect 0 4315 4200 4320
rect 0 4285 645 4315
rect 675 4285 1605 4315
rect 1635 4285 2565 4315
rect 2595 4285 3525 4315
rect 3555 4285 4005 4315
rect 4035 4285 4200 4315
rect 0 4280 4200 4285
rect 0 4235 4200 4240
rect 0 4205 85 4235
rect 115 4205 165 4235
rect 195 4205 245 4235
rect 275 4205 325 4235
rect 355 4205 405 4235
rect 435 4205 485 4235
rect 515 4205 565 4235
rect 595 4205 725 4235
rect 755 4205 805 4235
rect 835 4205 885 4235
rect 915 4205 965 4235
rect 995 4205 1045 4235
rect 1075 4205 1125 4235
rect 1155 4205 1205 4235
rect 1235 4205 1285 4235
rect 1315 4205 1365 4235
rect 1395 4205 1445 4235
rect 1475 4205 1525 4235
rect 1555 4205 1685 4235
rect 1715 4205 1765 4235
rect 1795 4205 1845 4235
rect 1875 4205 1925 4235
rect 1955 4205 2005 4235
rect 2035 4205 2085 4235
rect 2115 4205 2165 4235
rect 2195 4205 2245 4235
rect 2275 4205 2325 4235
rect 2355 4205 2405 4235
rect 2435 4205 2485 4235
rect 2515 4205 2645 4235
rect 2675 4205 2725 4235
rect 2755 4205 2805 4235
rect 2835 4205 2885 4235
rect 2915 4205 2965 4235
rect 2995 4205 3045 4235
rect 3075 4205 3125 4235
rect 3155 4205 3205 4235
rect 3235 4205 3285 4235
rect 3315 4205 3365 4235
rect 3395 4205 3445 4235
rect 3475 4205 3605 4235
rect 3635 4205 3685 4235
rect 3715 4205 3765 4235
rect 3795 4205 3845 4235
rect 3875 4205 3925 4235
rect 3955 4205 4005 4235
rect 4035 4205 4085 4235
rect 4115 4205 4200 4235
rect 0 4200 4200 4205
rect 0 4155 4200 4160
rect 0 4125 85 4155
rect 115 4125 165 4155
rect 195 4125 245 4155
rect 275 4125 325 4155
rect 355 4125 405 4155
rect 435 4125 485 4155
rect 515 4125 565 4155
rect 595 4125 725 4155
rect 755 4125 805 4155
rect 835 4125 885 4155
rect 915 4125 965 4155
rect 995 4125 1045 4155
rect 1075 4125 1125 4155
rect 1155 4125 1205 4155
rect 1235 4125 1285 4155
rect 1315 4125 1365 4155
rect 1395 4125 1445 4155
rect 1475 4125 1525 4155
rect 1555 4125 1685 4155
rect 1715 4125 1765 4155
rect 1795 4125 1845 4155
rect 1875 4125 1925 4155
rect 1955 4125 2005 4155
rect 2035 4125 2085 4155
rect 2115 4125 2165 4155
rect 2195 4125 2245 4155
rect 2275 4125 2325 4155
rect 2355 4125 2405 4155
rect 2435 4125 2485 4155
rect 2515 4125 2645 4155
rect 2675 4125 2725 4155
rect 2755 4125 2805 4155
rect 2835 4125 2885 4155
rect 2915 4125 2965 4155
rect 2995 4125 3045 4155
rect 3075 4125 3125 4155
rect 3155 4125 3205 4155
rect 3235 4125 3285 4155
rect 3315 4125 3365 4155
rect 3395 4125 3445 4155
rect 3475 4125 3605 4155
rect 3635 4125 3685 4155
rect 3715 4125 3765 4155
rect 3795 4125 3845 4155
rect 3875 4125 3925 4155
rect 3955 4125 4005 4155
rect 4035 4125 4085 4155
rect 4115 4125 4200 4155
rect 0 4120 4200 4125
rect 0 4075 4200 4080
rect 0 4045 645 4075
rect 675 4045 1605 4075
rect 1635 4045 2565 4075
rect 2595 4045 3525 4075
rect 3555 4045 4200 4075
rect 0 4040 4200 4045
rect 0 3995 4200 4000
rect 0 3965 85 3995
rect 115 3965 165 3995
rect 195 3965 245 3995
rect 275 3965 325 3995
rect 355 3965 405 3995
rect 435 3965 485 3995
rect 515 3965 565 3995
rect 595 3965 725 3995
rect 755 3965 805 3995
rect 835 3965 885 3995
rect 915 3965 965 3995
rect 995 3965 1045 3995
rect 1075 3965 1125 3995
rect 1155 3965 1205 3995
rect 1235 3965 1285 3995
rect 1315 3965 1365 3995
rect 1395 3965 1445 3995
rect 1475 3965 1525 3995
rect 1555 3965 1685 3995
rect 1715 3965 1765 3995
rect 1795 3965 1845 3995
rect 1875 3965 1925 3995
rect 1955 3965 2005 3995
rect 2035 3965 2085 3995
rect 2115 3965 2165 3995
rect 2195 3965 2245 3995
rect 2275 3965 2325 3995
rect 2355 3965 2405 3995
rect 2435 3965 2485 3995
rect 2515 3965 2645 3995
rect 2675 3965 2725 3995
rect 2755 3965 2805 3995
rect 2835 3965 2885 3995
rect 2915 3965 2965 3995
rect 2995 3965 3045 3995
rect 3075 3965 3125 3995
rect 3155 3965 3205 3995
rect 3235 3965 3285 3995
rect 3315 3965 3365 3995
rect 3395 3965 3445 3995
rect 3475 3965 3605 3995
rect 3635 3965 3685 3995
rect 3715 3965 3765 3995
rect 3795 3965 3845 3995
rect 3875 3965 3925 3995
rect 3955 3965 4005 3995
rect 4035 3965 4085 3995
rect 4115 3965 4200 3995
rect 0 3960 4200 3965
rect 160 3850 200 3860
rect 160 3770 165 3850
rect 195 3770 200 3850
rect 160 3760 200 3770
rect 160 3550 200 3560
rect 160 3470 165 3550
rect 195 3470 200 3550
rect 160 3460 200 3470
rect 0 3355 4200 3360
rect 0 3325 85 3355
rect 115 3325 165 3355
rect 195 3325 245 3355
rect 275 3325 325 3355
rect 355 3325 405 3355
rect 435 3325 485 3355
rect 515 3325 565 3355
rect 595 3325 725 3355
rect 755 3325 805 3355
rect 835 3325 885 3355
rect 915 3325 965 3355
rect 995 3325 1045 3355
rect 1075 3325 1125 3355
rect 1155 3325 1205 3355
rect 1235 3325 1285 3355
rect 1315 3325 1365 3355
rect 1395 3325 1445 3355
rect 1475 3325 1525 3355
rect 1555 3325 1685 3355
rect 1715 3325 1765 3355
rect 1795 3325 1845 3355
rect 1875 3325 1925 3355
rect 1955 3325 2005 3355
rect 2035 3325 2085 3355
rect 2115 3325 2165 3355
rect 2195 3325 2245 3355
rect 2275 3325 2325 3355
rect 2355 3325 2405 3355
rect 2435 3325 2485 3355
rect 2515 3325 2645 3355
rect 2675 3325 2725 3355
rect 2755 3325 2805 3355
rect 2835 3325 2885 3355
rect 2915 3325 2965 3355
rect 2995 3325 3045 3355
rect 3075 3325 3125 3355
rect 3155 3325 3205 3355
rect 3235 3325 3285 3355
rect 3315 3325 3365 3355
rect 3395 3325 3445 3355
rect 3475 3325 3605 3355
rect 3635 3325 3685 3355
rect 3715 3325 3765 3355
rect 3795 3325 3845 3355
rect 3875 3325 3925 3355
rect 3955 3325 4085 3355
rect 4115 3325 4200 3355
rect 0 3320 4200 3325
rect 0 3275 4200 3280
rect 0 3245 645 3275
rect 675 3245 1605 3275
rect 1635 3245 2565 3275
rect 2595 3245 3525 3275
rect 3555 3245 4200 3275
rect 0 3240 4200 3245
rect 0 3195 4200 3200
rect 0 3165 85 3195
rect 115 3165 165 3195
rect 195 3165 245 3195
rect 275 3165 325 3195
rect 355 3165 405 3195
rect 435 3165 485 3195
rect 515 3165 565 3195
rect 595 3165 725 3195
rect 755 3165 805 3195
rect 835 3165 885 3195
rect 915 3165 965 3195
rect 995 3165 1045 3195
rect 1075 3165 1125 3195
rect 1155 3165 1205 3195
rect 1235 3165 1285 3195
rect 1315 3165 1365 3195
rect 1395 3165 1445 3195
rect 1475 3165 1525 3195
rect 1555 3165 1685 3195
rect 1715 3165 1765 3195
rect 1795 3165 1845 3195
rect 1875 3165 1925 3195
rect 1955 3165 2005 3195
rect 2035 3165 2085 3195
rect 2115 3165 2165 3195
rect 2195 3165 2245 3195
rect 2275 3165 2325 3195
rect 2355 3165 2405 3195
rect 2435 3165 2485 3195
rect 2515 3165 2645 3195
rect 2675 3165 2725 3195
rect 2755 3165 2805 3195
rect 2835 3165 2885 3195
rect 2915 3165 2965 3195
rect 2995 3165 3045 3195
rect 3075 3165 3125 3195
rect 3155 3165 3205 3195
rect 3235 3165 3285 3195
rect 3315 3165 3365 3195
rect 3395 3165 3445 3195
rect 3475 3165 3605 3195
rect 3635 3165 3685 3195
rect 3715 3165 3765 3195
rect 3795 3165 3845 3195
rect 3875 3165 3925 3195
rect 3955 3165 4085 3195
rect 4115 3165 4200 3195
rect 0 3160 4200 3165
rect 0 3115 4200 3120
rect 0 3085 85 3115
rect 115 3085 165 3115
rect 195 3085 245 3115
rect 275 3085 325 3115
rect 355 3085 405 3115
rect 435 3085 485 3115
rect 515 3085 565 3115
rect 595 3085 645 3115
rect 675 3085 725 3115
rect 755 3085 805 3115
rect 835 3085 885 3115
rect 915 3085 965 3115
rect 995 3085 1045 3115
rect 1075 3085 1125 3115
rect 1155 3085 1205 3115
rect 1235 3085 1285 3115
rect 1315 3085 1365 3115
rect 1395 3085 1445 3115
rect 1475 3085 1525 3115
rect 1555 3085 1605 3115
rect 1635 3085 1685 3115
rect 1715 3085 1765 3115
rect 1795 3085 1845 3115
rect 1875 3085 1925 3115
rect 1955 3085 2005 3115
rect 2035 3085 2085 3115
rect 2115 3085 2165 3115
rect 2195 3085 2245 3115
rect 2275 3085 2325 3115
rect 2355 3085 2405 3115
rect 2435 3085 2485 3115
rect 2515 3085 2565 3115
rect 2595 3085 2645 3115
rect 2675 3085 2725 3115
rect 2755 3085 2805 3115
rect 2835 3085 2885 3115
rect 2915 3085 2965 3115
rect 2995 3085 3045 3115
rect 3075 3085 3125 3115
rect 3155 3085 3205 3115
rect 3235 3085 3285 3115
rect 3315 3085 3365 3115
rect 3395 3085 3445 3115
rect 3475 3085 3525 3115
rect 3555 3085 3605 3115
rect 3635 3085 3685 3115
rect 3715 3085 3765 3115
rect 3795 3085 3845 3115
rect 3875 3085 3925 3115
rect 3955 3085 4085 3115
rect 4115 3085 4200 3115
rect 0 3080 4200 3085
rect 0 3035 4200 3040
rect 0 3005 4005 3035
rect 4035 3005 4200 3035
rect 0 3000 4200 3005
rect 0 2955 4200 2960
rect 0 2925 85 2955
rect 115 2925 165 2955
rect 195 2925 245 2955
rect 275 2925 325 2955
rect 355 2925 405 2955
rect 435 2925 485 2955
rect 515 2925 565 2955
rect 595 2925 645 2955
rect 675 2925 725 2955
rect 755 2925 805 2955
rect 835 2925 885 2955
rect 915 2925 965 2955
rect 995 2925 1045 2955
rect 1075 2925 1125 2955
rect 1155 2925 1205 2955
rect 1235 2925 1285 2955
rect 1315 2925 1365 2955
rect 1395 2925 1445 2955
rect 1475 2925 1525 2955
rect 1555 2925 1605 2955
rect 1635 2925 1685 2955
rect 1715 2925 1765 2955
rect 1795 2925 1845 2955
rect 1875 2925 1925 2955
rect 1955 2925 2005 2955
rect 2035 2925 2085 2955
rect 2115 2925 2165 2955
rect 2195 2925 2245 2955
rect 2275 2925 2325 2955
rect 2355 2925 2405 2955
rect 2435 2925 2485 2955
rect 2515 2925 2565 2955
rect 2595 2925 2645 2955
rect 2675 2925 2725 2955
rect 2755 2925 2805 2955
rect 2835 2925 2885 2955
rect 2915 2925 2965 2955
rect 2995 2925 3045 2955
rect 3075 2925 3125 2955
rect 3155 2925 3205 2955
rect 3235 2925 3285 2955
rect 3315 2925 3365 2955
rect 3395 2925 3445 2955
rect 3475 2925 3525 2955
rect 3555 2925 3605 2955
rect 3635 2925 3685 2955
rect 3715 2925 3765 2955
rect 3795 2925 3845 2955
rect 3875 2925 3925 2955
rect 3955 2925 4085 2955
rect 4115 2925 4200 2955
rect 0 2920 4200 2925
rect 0 2875 4200 2880
rect 0 2845 85 2875
rect 115 2845 165 2875
rect 195 2845 245 2875
rect 275 2845 325 2875
rect 355 2845 405 2875
rect 435 2845 485 2875
rect 515 2845 565 2875
rect 595 2845 725 2875
rect 755 2845 805 2875
rect 835 2845 885 2875
rect 915 2845 965 2875
rect 995 2845 1045 2875
rect 1075 2845 1125 2875
rect 1155 2845 1205 2875
rect 1235 2845 1285 2875
rect 1315 2845 1365 2875
rect 1395 2845 1445 2875
rect 1475 2845 1525 2875
rect 1555 2845 1685 2875
rect 1715 2845 1765 2875
rect 1795 2845 1845 2875
rect 1875 2845 1925 2875
rect 1955 2845 2005 2875
rect 2035 2845 2085 2875
rect 2115 2845 2165 2875
rect 2195 2845 2245 2875
rect 2275 2845 2325 2875
rect 2355 2845 2405 2875
rect 2435 2845 2485 2875
rect 2515 2845 2645 2875
rect 2675 2845 2725 2875
rect 2755 2845 2805 2875
rect 2835 2845 2885 2875
rect 2915 2845 2965 2875
rect 2995 2845 3045 2875
rect 3075 2845 3125 2875
rect 3155 2845 3205 2875
rect 3235 2845 3285 2875
rect 3315 2845 3365 2875
rect 3395 2845 3445 2875
rect 3475 2845 3605 2875
rect 3635 2845 3685 2875
rect 3715 2845 3765 2875
rect 3795 2845 3845 2875
rect 3875 2845 3925 2875
rect 3955 2845 4085 2875
rect 4115 2845 4200 2875
rect 0 2840 4200 2845
rect 0 2795 4200 2800
rect 0 2765 645 2795
rect 675 2765 1605 2795
rect 1635 2765 2565 2795
rect 2595 2765 3525 2795
rect 3555 2765 4200 2795
rect 0 2760 4200 2765
rect 0 2715 4200 2720
rect 0 2685 85 2715
rect 115 2685 165 2715
rect 195 2685 245 2715
rect 275 2685 325 2715
rect 355 2685 405 2715
rect 435 2685 485 2715
rect 515 2685 565 2715
rect 595 2685 725 2715
rect 755 2685 805 2715
rect 835 2685 885 2715
rect 915 2685 965 2715
rect 995 2685 1045 2715
rect 1075 2685 1125 2715
rect 1155 2685 1205 2715
rect 1235 2685 1285 2715
rect 1315 2685 1365 2715
rect 1395 2685 1445 2715
rect 1475 2685 1525 2715
rect 1555 2685 1685 2715
rect 1715 2685 1765 2715
rect 1795 2685 1845 2715
rect 1875 2685 1925 2715
rect 1955 2685 2005 2715
rect 2035 2685 2085 2715
rect 2115 2685 2165 2715
rect 2195 2685 2245 2715
rect 2275 2685 2325 2715
rect 2355 2685 2405 2715
rect 2435 2685 2485 2715
rect 2515 2685 2645 2715
rect 2675 2685 2725 2715
rect 2755 2685 2805 2715
rect 2835 2685 2885 2715
rect 2915 2685 2965 2715
rect 2995 2685 3045 2715
rect 3075 2685 3125 2715
rect 3155 2685 3205 2715
rect 3235 2685 3285 2715
rect 3315 2685 3365 2715
rect 3395 2685 3445 2715
rect 3475 2685 3605 2715
rect 3635 2685 3685 2715
rect 3715 2685 3765 2715
rect 3795 2685 3845 2715
rect 3875 2685 3925 2715
rect 3955 2685 4085 2715
rect 4115 2685 4200 2715
rect 0 2680 4200 2685
rect 160 2390 200 2400
rect 160 2210 165 2390
rect 195 2210 200 2390
rect 160 2200 200 2210
rect 4000 1830 4040 1840
rect 4000 1650 4005 1830
rect 4035 1650 4040 1830
rect 4000 1640 4040 1650
rect 0 1395 4200 1400
rect 0 1365 5 1395
rect 35 1365 85 1395
rect 115 1365 165 1395
rect 195 1365 245 1395
rect 275 1365 325 1395
rect 355 1365 405 1395
rect 435 1365 485 1395
rect 515 1365 565 1395
rect 595 1365 725 1395
rect 755 1365 805 1395
rect 835 1365 885 1395
rect 915 1365 965 1395
rect 995 1365 1045 1395
rect 1075 1365 1125 1395
rect 1155 1365 1205 1395
rect 1235 1365 1285 1395
rect 1315 1365 1365 1395
rect 1395 1365 1445 1395
rect 1475 1365 1525 1395
rect 1555 1365 1685 1395
rect 1715 1365 1765 1395
rect 1795 1365 1845 1395
rect 1875 1365 1925 1395
rect 1955 1365 2005 1395
rect 2035 1365 2085 1395
rect 2115 1365 2165 1395
rect 2195 1365 2245 1395
rect 2275 1365 2325 1395
rect 2355 1365 2405 1395
rect 2435 1365 2485 1395
rect 2515 1365 2645 1395
rect 2675 1365 2725 1395
rect 2755 1365 2805 1395
rect 2835 1365 2885 1395
rect 2915 1365 2965 1395
rect 2995 1365 3045 1395
rect 3075 1365 3125 1395
rect 3155 1365 3205 1395
rect 3235 1365 3285 1395
rect 3315 1365 3365 1395
rect 3395 1365 3445 1395
rect 3475 1365 3605 1395
rect 3635 1365 3685 1395
rect 3715 1365 3765 1395
rect 3795 1365 3845 1395
rect 3875 1365 3925 1395
rect 3955 1365 4005 1395
rect 4035 1365 4085 1395
rect 4115 1365 4165 1395
rect 4195 1365 4200 1395
rect 0 1360 4200 1365
rect 0 1315 4200 1320
rect 0 1285 645 1315
rect 675 1285 1605 1315
rect 1635 1285 2565 1315
rect 2595 1285 3525 1315
rect 3555 1285 4200 1315
rect 0 1280 4200 1285
rect 0 1235 4200 1240
rect 0 1205 5 1235
rect 35 1205 85 1235
rect 115 1205 165 1235
rect 195 1205 245 1235
rect 275 1205 325 1235
rect 355 1205 405 1235
rect 435 1205 485 1235
rect 515 1205 565 1235
rect 595 1205 725 1235
rect 755 1205 805 1235
rect 835 1205 885 1235
rect 915 1205 965 1235
rect 995 1205 1045 1235
rect 1075 1205 1125 1235
rect 1155 1205 1205 1235
rect 1235 1205 1285 1235
rect 1315 1205 1365 1235
rect 1395 1205 1445 1235
rect 1475 1205 1525 1235
rect 1555 1205 1685 1235
rect 1715 1205 1765 1235
rect 1795 1205 1845 1235
rect 1875 1205 1925 1235
rect 1955 1205 2005 1235
rect 2035 1205 2085 1235
rect 2115 1205 2165 1235
rect 2195 1205 2245 1235
rect 2275 1205 2325 1235
rect 2355 1205 2405 1235
rect 2435 1205 2485 1235
rect 2515 1205 2645 1235
rect 2675 1205 2725 1235
rect 2755 1205 2805 1235
rect 2835 1205 2885 1235
rect 2915 1205 2965 1235
rect 2995 1205 3045 1235
rect 3075 1205 3125 1235
rect 3155 1205 3205 1235
rect 3235 1205 3285 1235
rect 3315 1205 3365 1235
rect 3395 1205 3445 1235
rect 3475 1205 3605 1235
rect 3635 1205 3685 1235
rect 3715 1205 3765 1235
rect 3795 1205 3845 1235
rect 3875 1205 3925 1235
rect 3955 1205 4005 1235
rect 4035 1205 4085 1235
rect 4115 1205 4165 1235
rect 4195 1205 4200 1235
rect 0 1200 4200 1205
rect 0 635 4200 640
rect 0 605 85 635
rect 115 605 165 635
rect 195 605 245 635
rect 275 605 325 635
rect 355 605 405 635
rect 435 605 485 635
rect 515 605 565 635
rect 595 605 725 635
rect 755 605 805 635
rect 835 605 885 635
rect 915 605 965 635
rect 995 605 1045 635
rect 1075 605 1125 635
rect 1155 605 1205 635
rect 1235 605 1285 635
rect 1315 605 1365 635
rect 1395 605 1445 635
rect 1475 605 1525 635
rect 1555 605 1685 635
rect 1715 605 1765 635
rect 1795 605 1845 635
rect 1875 605 1925 635
rect 1955 605 2005 635
rect 2035 605 2085 635
rect 2115 605 2165 635
rect 2195 605 2245 635
rect 2275 605 2325 635
rect 2355 605 2405 635
rect 2435 605 2485 635
rect 2515 605 2645 635
rect 2675 605 2725 635
rect 2755 605 2805 635
rect 2835 605 2885 635
rect 2915 605 2965 635
rect 2995 605 3045 635
rect 3075 605 3125 635
rect 3155 605 3205 635
rect 3235 605 3285 635
rect 3315 605 3365 635
rect 3395 605 3445 635
rect 3475 605 3605 635
rect 3635 605 3685 635
rect 3715 605 3765 635
rect 3795 605 3845 635
rect 3875 605 3925 635
rect 3955 605 4005 635
rect 4035 605 4085 635
rect 4115 605 4200 635
rect 0 600 4200 605
rect 0 555 4200 560
rect 0 525 645 555
rect 675 525 1605 555
rect 1635 525 2565 555
rect 2595 525 3525 555
rect 3555 525 4005 555
rect 4035 525 4200 555
rect 0 520 4200 525
rect 0 475 4200 480
rect 0 445 85 475
rect 115 445 165 475
rect 195 445 245 475
rect 275 445 325 475
rect 355 445 405 475
rect 435 445 485 475
rect 515 445 565 475
rect 595 445 725 475
rect 755 445 805 475
rect 835 445 885 475
rect 915 445 965 475
rect 995 445 1045 475
rect 1075 445 1125 475
rect 1155 445 1205 475
rect 1235 445 1285 475
rect 1315 445 1365 475
rect 1395 445 1445 475
rect 1475 445 1525 475
rect 1555 445 1685 475
rect 1715 445 1765 475
rect 1795 445 1845 475
rect 1875 445 1925 475
rect 1955 445 2005 475
rect 2035 445 2085 475
rect 2115 445 2165 475
rect 2195 445 2245 475
rect 2275 445 2325 475
rect 2355 445 2405 475
rect 2435 445 2485 475
rect 2515 445 2645 475
rect 2675 445 2725 475
rect 2755 445 2805 475
rect 2835 445 2885 475
rect 2915 445 2965 475
rect 2995 445 3045 475
rect 3075 445 3125 475
rect 3155 445 3205 475
rect 3235 445 3285 475
rect 3315 445 3365 475
rect 3395 445 3445 475
rect 3475 445 3605 475
rect 3635 445 3685 475
rect 3715 445 3765 475
rect 3795 445 3845 475
rect 3875 445 3925 475
rect 3955 445 4085 475
rect 4115 445 4200 475
rect 0 440 4200 445
rect 0 395 4200 400
rect 0 365 4005 395
rect 4035 365 4200 395
rect 0 360 4200 365
rect 0 315 4200 320
rect 0 285 85 315
rect 115 285 165 315
rect 195 285 245 315
rect 275 285 325 315
rect 355 285 405 315
rect 435 285 485 315
rect 515 285 565 315
rect 595 285 725 315
rect 755 285 805 315
rect 835 285 885 315
rect 915 285 965 315
rect 995 285 1045 315
rect 1075 285 1125 315
rect 1155 285 1205 315
rect 1235 285 1285 315
rect 1315 285 1365 315
rect 1395 285 1445 315
rect 1475 285 1525 315
rect 1555 285 1685 315
rect 1715 285 1765 315
rect 1795 285 1845 315
rect 1875 285 1925 315
rect 1955 285 2005 315
rect 2035 285 2085 315
rect 2115 285 2165 315
rect 2195 285 2245 315
rect 2275 285 2325 315
rect 2355 285 2405 315
rect 2435 285 2485 315
rect 2515 285 2645 315
rect 2675 285 2725 315
rect 2755 285 2805 315
rect 2835 285 2885 315
rect 2915 285 2965 315
rect 2995 285 3045 315
rect 3075 285 3125 315
rect 3155 285 3205 315
rect 3235 285 3285 315
rect 3315 285 3365 315
rect 3395 285 3445 315
rect 3475 285 3605 315
rect 3635 285 3685 315
rect 3715 285 3765 315
rect 3795 285 3845 315
rect 3875 285 3925 315
rect 3955 285 4005 315
rect 4035 285 4085 315
rect 4115 285 4200 315
rect 0 280 4200 285
rect 160 170 200 180
rect 160 90 165 170
rect 195 90 200 170
rect 160 80 200 90
rect 0 -45 4200 -40
rect 0 -75 85 -45
rect 115 -75 165 -45
rect 195 -75 245 -45
rect 275 -75 325 -45
rect 355 -75 405 -45
rect 435 -75 485 -45
rect 515 -75 565 -45
rect 595 -75 725 -45
rect 755 -75 805 -45
rect 835 -75 885 -45
rect 915 -75 965 -45
rect 995 -75 1045 -45
rect 1075 -75 1125 -45
rect 1155 -75 1205 -45
rect 1235 -75 1285 -45
rect 1315 -75 1365 -45
rect 1395 -75 1445 -45
rect 1475 -75 1525 -45
rect 1555 -75 1685 -45
rect 1715 -75 1765 -45
rect 1795 -75 1845 -45
rect 1875 -75 1925 -45
rect 1955 -75 2005 -45
rect 2035 -75 2085 -45
rect 2115 -75 2165 -45
rect 2195 -75 2245 -45
rect 2275 -75 2325 -45
rect 2355 -75 2405 -45
rect 2435 -75 2485 -45
rect 2515 -75 2645 -45
rect 2675 -75 2725 -45
rect 2755 -75 2805 -45
rect 2835 -75 2885 -45
rect 2915 -75 2965 -45
rect 2995 -75 3045 -45
rect 3075 -75 3125 -45
rect 3155 -75 3205 -45
rect 3235 -75 3285 -45
rect 3315 -75 3365 -45
rect 3395 -75 3445 -45
rect 3475 -75 3605 -45
rect 3635 -75 3685 -45
rect 3715 -75 3765 -45
rect 3795 -75 3845 -45
rect 3875 -75 3925 -45
rect 3955 -75 4085 -45
rect 4115 -75 4200 -45
rect 0 -80 4200 -75
rect 0 -125 4200 -120
rect 0 -155 645 -125
rect 675 -155 1605 -125
rect 1635 -155 2565 -125
rect 2595 -155 3525 -125
rect 3555 -155 4005 -125
rect 4035 -155 4200 -125
rect 0 -160 4200 -155
rect 0 -205 4200 -200
rect 0 -235 85 -205
rect 115 -235 165 -205
rect 195 -235 245 -205
rect 275 -235 325 -205
rect 355 -235 405 -205
rect 435 -235 485 -205
rect 515 -235 565 -205
rect 595 -235 725 -205
rect 755 -235 805 -205
rect 835 -235 885 -205
rect 915 -235 965 -205
rect 995 -235 1045 -205
rect 1075 -235 1125 -205
rect 1155 -235 1205 -205
rect 1235 -235 1285 -205
rect 1315 -235 1365 -205
rect 1395 -235 1445 -205
rect 1475 -235 1525 -205
rect 1555 -235 1685 -205
rect 1715 -235 1765 -205
rect 1795 -235 1845 -205
rect 1875 -235 1925 -205
rect 1955 -235 2005 -205
rect 2035 -235 2085 -205
rect 2115 -235 2165 -205
rect 2195 -235 2245 -205
rect 2275 -235 2325 -205
rect 2355 -235 2405 -205
rect 2435 -235 2485 -205
rect 2515 -235 2645 -205
rect 2675 -235 2725 -205
rect 2755 -235 2805 -205
rect 2835 -235 2885 -205
rect 2915 -235 2965 -205
rect 2995 -235 3045 -205
rect 3075 -235 3125 -205
rect 3155 -235 3205 -205
rect 3235 -235 3285 -205
rect 3315 -235 3365 -205
rect 3395 -235 3445 -205
rect 3475 -235 3605 -205
rect 3635 -235 3685 -205
rect 3715 -235 3765 -205
rect 3795 -235 3845 -205
rect 3875 -235 3925 -205
rect 3955 -235 4085 -205
rect 4115 -235 4200 -205
rect 0 -240 4200 -235
rect 160 -350 200 -340
rect 160 -430 165 -350
rect 195 -430 200 -350
rect 160 -440 200 -430
<< via2 >>
rect 165 4690 195 4870
rect 85 4365 115 4395
rect 165 4365 195 4395
rect 245 4365 275 4395
rect 325 4365 355 4395
rect 405 4365 435 4395
rect 485 4365 515 4395
rect 565 4365 595 4395
rect 725 4365 755 4395
rect 805 4365 835 4395
rect 885 4365 915 4395
rect 965 4365 995 4395
rect 1045 4365 1075 4395
rect 1125 4365 1155 4395
rect 1205 4365 1235 4395
rect 1285 4365 1315 4395
rect 1365 4365 1395 4395
rect 1445 4365 1475 4395
rect 1525 4365 1555 4395
rect 1685 4365 1715 4395
rect 1765 4365 1795 4395
rect 1845 4365 1875 4395
rect 1925 4365 1955 4395
rect 2005 4365 2035 4395
rect 2085 4365 2115 4395
rect 2165 4365 2195 4395
rect 2245 4365 2275 4395
rect 2325 4365 2355 4395
rect 2405 4365 2435 4395
rect 2485 4365 2515 4395
rect 2645 4365 2675 4395
rect 2725 4365 2755 4395
rect 2805 4365 2835 4395
rect 2885 4365 2915 4395
rect 2965 4365 2995 4395
rect 3045 4365 3075 4395
rect 3125 4365 3155 4395
rect 3205 4365 3235 4395
rect 3285 4365 3315 4395
rect 3365 4365 3395 4395
rect 3445 4365 3475 4395
rect 3605 4365 3635 4395
rect 3685 4365 3715 4395
rect 3765 4365 3795 4395
rect 3845 4365 3875 4395
rect 3925 4365 3955 4395
rect 4005 4365 4035 4395
rect 4085 4365 4115 4395
rect 85 4205 115 4235
rect 165 4205 195 4235
rect 245 4205 275 4235
rect 325 4205 355 4235
rect 405 4205 435 4235
rect 485 4205 515 4235
rect 565 4205 595 4235
rect 725 4205 755 4235
rect 805 4205 835 4235
rect 885 4205 915 4235
rect 965 4205 995 4235
rect 1045 4205 1075 4235
rect 1125 4205 1155 4235
rect 1205 4205 1235 4235
rect 1285 4205 1315 4235
rect 1365 4205 1395 4235
rect 1445 4205 1475 4235
rect 1525 4205 1555 4235
rect 1685 4205 1715 4235
rect 1765 4205 1795 4235
rect 1845 4205 1875 4235
rect 1925 4205 1955 4235
rect 2005 4205 2035 4235
rect 2085 4205 2115 4235
rect 2165 4205 2195 4235
rect 2245 4205 2275 4235
rect 2325 4205 2355 4235
rect 2405 4205 2435 4235
rect 2485 4205 2515 4235
rect 2645 4205 2675 4235
rect 2725 4205 2755 4235
rect 2805 4205 2835 4235
rect 2885 4205 2915 4235
rect 2965 4205 2995 4235
rect 3045 4205 3075 4235
rect 3125 4205 3155 4235
rect 3205 4205 3235 4235
rect 3285 4205 3315 4235
rect 3365 4205 3395 4235
rect 3445 4205 3475 4235
rect 3605 4205 3635 4235
rect 3685 4205 3715 4235
rect 3765 4205 3795 4235
rect 3845 4205 3875 4235
rect 3925 4205 3955 4235
rect 4005 4205 4035 4235
rect 4085 4205 4115 4235
rect 85 4125 115 4155
rect 165 4125 195 4155
rect 245 4125 275 4155
rect 325 4125 355 4155
rect 405 4125 435 4155
rect 485 4125 515 4155
rect 565 4125 595 4155
rect 725 4125 755 4155
rect 805 4125 835 4155
rect 885 4125 915 4155
rect 965 4125 995 4155
rect 1045 4125 1075 4155
rect 1125 4125 1155 4155
rect 1205 4125 1235 4155
rect 1285 4125 1315 4155
rect 1365 4125 1395 4155
rect 1445 4125 1475 4155
rect 1525 4125 1555 4155
rect 1685 4125 1715 4155
rect 1765 4125 1795 4155
rect 1845 4125 1875 4155
rect 1925 4125 1955 4155
rect 2005 4125 2035 4155
rect 2085 4125 2115 4155
rect 2165 4125 2195 4155
rect 2245 4125 2275 4155
rect 2325 4125 2355 4155
rect 2405 4125 2435 4155
rect 2485 4125 2515 4155
rect 2645 4125 2675 4155
rect 2725 4125 2755 4155
rect 2805 4125 2835 4155
rect 2885 4125 2915 4155
rect 2965 4125 2995 4155
rect 3045 4125 3075 4155
rect 3125 4125 3155 4155
rect 3205 4125 3235 4155
rect 3285 4125 3315 4155
rect 3365 4125 3395 4155
rect 3445 4125 3475 4155
rect 3605 4125 3635 4155
rect 3685 4125 3715 4155
rect 3765 4125 3795 4155
rect 3845 4125 3875 4155
rect 3925 4125 3955 4155
rect 4005 4125 4035 4155
rect 4085 4125 4115 4155
rect 85 3965 115 3995
rect 165 3965 195 3995
rect 245 3965 275 3995
rect 325 3965 355 3995
rect 405 3965 435 3995
rect 485 3965 515 3995
rect 565 3965 595 3995
rect 725 3965 755 3995
rect 805 3965 835 3995
rect 885 3965 915 3995
rect 965 3965 995 3995
rect 1045 3965 1075 3995
rect 1125 3965 1155 3995
rect 1205 3965 1235 3995
rect 1285 3965 1315 3995
rect 1365 3965 1395 3995
rect 1445 3965 1475 3995
rect 1525 3965 1555 3995
rect 1685 3965 1715 3995
rect 1765 3965 1795 3995
rect 1845 3965 1875 3995
rect 1925 3965 1955 3995
rect 2005 3965 2035 3995
rect 2085 3965 2115 3995
rect 2165 3965 2195 3995
rect 2245 3965 2275 3995
rect 2325 3965 2355 3995
rect 2405 3965 2435 3995
rect 2485 3965 2515 3995
rect 2645 3965 2675 3995
rect 2725 3965 2755 3995
rect 2805 3965 2835 3995
rect 2885 3965 2915 3995
rect 2965 3965 2995 3995
rect 3045 3965 3075 3995
rect 3125 3965 3155 3995
rect 3205 3965 3235 3995
rect 3285 3965 3315 3995
rect 3365 3965 3395 3995
rect 3445 3965 3475 3995
rect 3605 3965 3635 3995
rect 3685 3965 3715 3995
rect 3765 3965 3795 3995
rect 3845 3965 3875 3995
rect 3925 3965 3955 3995
rect 4005 3965 4035 3995
rect 4085 3965 4115 3995
rect 165 3770 195 3850
rect 165 3470 195 3550
rect 85 3325 115 3355
rect 165 3325 195 3355
rect 245 3325 275 3355
rect 325 3325 355 3355
rect 405 3325 435 3355
rect 485 3325 515 3355
rect 565 3325 595 3355
rect 725 3325 755 3355
rect 805 3325 835 3355
rect 885 3325 915 3355
rect 965 3325 995 3355
rect 1045 3325 1075 3355
rect 1125 3325 1155 3355
rect 1205 3325 1235 3355
rect 1285 3325 1315 3355
rect 1365 3325 1395 3355
rect 1445 3325 1475 3355
rect 1525 3325 1555 3355
rect 1685 3325 1715 3355
rect 1765 3325 1795 3355
rect 1845 3325 1875 3355
rect 1925 3325 1955 3355
rect 2005 3325 2035 3355
rect 2085 3325 2115 3355
rect 2165 3325 2195 3355
rect 2245 3325 2275 3355
rect 2325 3325 2355 3355
rect 2405 3325 2435 3355
rect 2485 3325 2515 3355
rect 2645 3325 2675 3355
rect 2725 3325 2755 3355
rect 2805 3325 2835 3355
rect 2885 3325 2915 3355
rect 2965 3325 2995 3355
rect 3045 3325 3075 3355
rect 3125 3325 3155 3355
rect 3205 3325 3235 3355
rect 3285 3325 3315 3355
rect 3365 3325 3395 3355
rect 3445 3325 3475 3355
rect 3605 3325 3635 3355
rect 3685 3325 3715 3355
rect 3765 3325 3795 3355
rect 3845 3325 3875 3355
rect 3925 3325 3955 3355
rect 4085 3325 4115 3355
rect 85 3165 115 3195
rect 165 3165 195 3195
rect 245 3165 275 3195
rect 325 3165 355 3195
rect 405 3165 435 3195
rect 485 3165 515 3195
rect 565 3165 595 3195
rect 725 3165 755 3195
rect 805 3165 835 3195
rect 885 3165 915 3195
rect 965 3165 995 3195
rect 1045 3165 1075 3195
rect 1125 3165 1155 3195
rect 1205 3165 1235 3195
rect 1285 3165 1315 3195
rect 1365 3165 1395 3195
rect 1445 3165 1475 3195
rect 1525 3165 1555 3195
rect 1685 3165 1715 3195
rect 1765 3165 1795 3195
rect 1845 3165 1875 3195
rect 1925 3165 1955 3195
rect 2005 3165 2035 3195
rect 2085 3165 2115 3195
rect 2165 3165 2195 3195
rect 2245 3165 2275 3195
rect 2325 3165 2355 3195
rect 2405 3165 2435 3195
rect 2485 3165 2515 3195
rect 2645 3165 2675 3195
rect 2725 3165 2755 3195
rect 2805 3165 2835 3195
rect 2885 3165 2915 3195
rect 2965 3165 2995 3195
rect 3045 3165 3075 3195
rect 3125 3165 3155 3195
rect 3205 3165 3235 3195
rect 3285 3165 3315 3195
rect 3365 3165 3395 3195
rect 3445 3165 3475 3195
rect 3605 3165 3635 3195
rect 3685 3165 3715 3195
rect 3765 3165 3795 3195
rect 3845 3165 3875 3195
rect 3925 3165 3955 3195
rect 4085 3165 4115 3195
rect 85 3085 115 3115
rect 165 3085 195 3115
rect 245 3085 275 3115
rect 325 3085 355 3115
rect 405 3085 435 3115
rect 485 3085 515 3115
rect 565 3085 595 3115
rect 645 3085 675 3115
rect 725 3085 755 3115
rect 805 3085 835 3115
rect 885 3085 915 3115
rect 965 3085 995 3115
rect 1045 3085 1075 3115
rect 1125 3085 1155 3115
rect 1205 3085 1235 3115
rect 1285 3085 1315 3115
rect 1365 3085 1395 3115
rect 1445 3085 1475 3115
rect 1525 3085 1555 3115
rect 1605 3085 1635 3115
rect 1685 3085 1715 3115
rect 1765 3085 1795 3115
rect 1845 3085 1875 3115
rect 1925 3085 1955 3115
rect 2005 3085 2035 3115
rect 2085 3085 2115 3115
rect 2165 3085 2195 3115
rect 2245 3085 2275 3115
rect 2325 3085 2355 3115
rect 2405 3085 2435 3115
rect 2485 3085 2515 3115
rect 2565 3085 2595 3115
rect 2645 3085 2675 3115
rect 2725 3085 2755 3115
rect 2805 3085 2835 3115
rect 2885 3085 2915 3115
rect 2965 3085 2995 3115
rect 3045 3085 3075 3115
rect 3125 3085 3155 3115
rect 3205 3085 3235 3115
rect 3285 3085 3315 3115
rect 3365 3085 3395 3115
rect 3445 3085 3475 3115
rect 3525 3085 3555 3115
rect 3605 3085 3635 3115
rect 3685 3085 3715 3115
rect 3765 3085 3795 3115
rect 3845 3085 3875 3115
rect 3925 3085 3955 3115
rect 4085 3085 4115 3115
rect 85 2925 115 2955
rect 165 2925 195 2955
rect 245 2925 275 2955
rect 325 2925 355 2955
rect 405 2925 435 2955
rect 485 2925 515 2955
rect 565 2925 595 2955
rect 645 2925 675 2955
rect 725 2925 755 2955
rect 805 2925 835 2955
rect 885 2925 915 2955
rect 965 2925 995 2955
rect 1045 2925 1075 2955
rect 1125 2925 1155 2955
rect 1205 2925 1235 2955
rect 1285 2925 1315 2955
rect 1365 2925 1395 2955
rect 1445 2925 1475 2955
rect 1525 2925 1555 2955
rect 1605 2925 1635 2955
rect 1685 2925 1715 2955
rect 1765 2925 1795 2955
rect 1845 2925 1875 2955
rect 1925 2925 1955 2955
rect 2005 2925 2035 2955
rect 2085 2925 2115 2955
rect 2165 2925 2195 2955
rect 2245 2925 2275 2955
rect 2325 2925 2355 2955
rect 2405 2925 2435 2955
rect 2485 2925 2515 2955
rect 2565 2925 2595 2955
rect 2645 2925 2675 2955
rect 2725 2925 2755 2955
rect 2805 2925 2835 2955
rect 2885 2925 2915 2955
rect 2965 2925 2995 2955
rect 3045 2925 3075 2955
rect 3125 2925 3155 2955
rect 3205 2925 3235 2955
rect 3285 2925 3315 2955
rect 3365 2925 3395 2955
rect 3445 2925 3475 2955
rect 3525 2925 3555 2955
rect 3605 2925 3635 2955
rect 3685 2925 3715 2955
rect 3765 2925 3795 2955
rect 3845 2925 3875 2955
rect 3925 2925 3955 2955
rect 4085 2925 4115 2955
rect 85 2845 115 2875
rect 165 2845 195 2875
rect 245 2845 275 2875
rect 325 2845 355 2875
rect 405 2845 435 2875
rect 485 2845 515 2875
rect 565 2845 595 2875
rect 725 2845 755 2875
rect 805 2845 835 2875
rect 885 2845 915 2875
rect 965 2845 995 2875
rect 1045 2845 1075 2875
rect 1125 2845 1155 2875
rect 1205 2845 1235 2875
rect 1285 2845 1315 2875
rect 1365 2845 1395 2875
rect 1445 2845 1475 2875
rect 1525 2845 1555 2875
rect 1685 2845 1715 2875
rect 1765 2845 1795 2875
rect 1845 2845 1875 2875
rect 1925 2845 1955 2875
rect 2005 2845 2035 2875
rect 2085 2845 2115 2875
rect 2165 2845 2195 2875
rect 2245 2845 2275 2875
rect 2325 2845 2355 2875
rect 2405 2845 2435 2875
rect 2485 2845 2515 2875
rect 2645 2845 2675 2875
rect 2725 2845 2755 2875
rect 2805 2845 2835 2875
rect 2885 2845 2915 2875
rect 2965 2845 2995 2875
rect 3045 2845 3075 2875
rect 3125 2845 3155 2875
rect 3205 2845 3235 2875
rect 3285 2845 3315 2875
rect 3365 2845 3395 2875
rect 3445 2845 3475 2875
rect 3605 2845 3635 2875
rect 3685 2845 3715 2875
rect 3765 2845 3795 2875
rect 3845 2845 3875 2875
rect 3925 2845 3955 2875
rect 4085 2845 4115 2875
rect 85 2685 115 2715
rect 165 2685 195 2715
rect 245 2685 275 2715
rect 325 2685 355 2715
rect 405 2685 435 2715
rect 485 2685 515 2715
rect 565 2685 595 2715
rect 725 2685 755 2715
rect 805 2685 835 2715
rect 885 2685 915 2715
rect 965 2685 995 2715
rect 1045 2685 1075 2715
rect 1125 2685 1155 2715
rect 1205 2685 1235 2715
rect 1285 2685 1315 2715
rect 1365 2685 1395 2715
rect 1445 2685 1475 2715
rect 1525 2685 1555 2715
rect 1685 2685 1715 2715
rect 1765 2685 1795 2715
rect 1845 2685 1875 2715
rect 1925 2685 1955 2715
rect 2005 2685 2035 2715
rect 2085 2685 2115 2715
rect 2165 2685 2195 2715
rect 2245 2685 2275 2715
rect 2325 2685 2355 2715
rect 2405 2685 2435 2715
rect 2485 2685 2515 2715
rect 2645 2685 2675 2715
rect 2725 2685 2755 2715
rect 2805 2685 2835 2715
rect 2885 2685 2915 2715
rect 2965 2685 2995 2715
rect 3045 2685 3075 2715
rect 3125 2685 3155 2715
rect 3205 2685 3235 2715
rect 3285 2685 3315 2715
rect 3365 2685 3395 2715
rect 3445 2685 3475 2715
rect 3605 2685 3635 2715
rect 3685 2685 3715 2715
rect 3765 2685 3795 2715
rect 3845 2685 3875 2715
rect 3925 2685 3955 2715
rect 4085 2685 4115 2715
rect 165 2210 195 2390
rect 4005 1650 4035 1830
rect 5 1365 35 1395
rect 85 1365 115 1395
rect 165 1365 195 1395
rect 245 1365 275 1395
rect 325 1365 355 1395
rect 405 1365 435 1395
rect 485 1365 515 1395
rect 565 1365 595 1395
rect 725 1365 755 1395
rect 805 1365 835 1395
rect 885 1365 915 1395
rect 965 1365 995 1395
rect 1045 1365 1075 1395
rect 1125 1365 1155 1395
rect 1205 1365 1235 1395
rect 1285 1365 1315 1395
rect 1365 1365 1395 1395
rect 1445 1365 1475 1395
rect 1525 1365 1555 1395
rect 1685 1365 1715 1395
rect 1765 1365 1795 1395
rect 1845 1365 1875 1395
rect 1925 1365 1955 1395
rect 2005 1365 2035 1395
rect 2085 1365 2115 1395
rect 2165 1365 2195 1395
rect 2245 1365 2275 1395
rect 2325 1365 2355 1395
rect 2405 1365 2435 1395
rect 2485 1365 2515 1395
rect 2645 1365 2675 1395
rect 2725 1365 2755 1395
rect 2805 1365 2835 1395
rect 2885 1365 2915 1395
rect 2965 1365 2995 1395
rect 3045 1365 3075 1395
rect 3125 1365 3155 1395
rect 3205 1365 3235 1395
rect 3285 1365 3315 1395
rect 3365 1365 3395 1395
rect 3445 1365 3475 1395
rect 3605 1365 3635 1395
rect 3685 1365 3715 1395
rect 3765 1365 3795 1395
rect 3845 1365 3875 1395
rect 3925 1365 3955 1395
rect 4005 1365 4035 1395
rect 4085 1365 4115 1395
rect 4165 1365 4195 1395
rect 5 1205 35 1235
rect 85 1205 115 1235
rect 165 1205 195 1235
rect 245 1205 275 1235
rect 325 1205 355 1235
rect 405 1205 435 1235
rect 485 1205 515 1235
rect 565 1205 595 1235
rect 725 1205 755 1235
rect 805 1205 835 1235
rect 885 1205 915 1235
rect 965 1205 995 1235
rect 1045 1205 1075 1235
rect 1125 1205 1155 1235
rect 1205 1205 1235 1235
rect 1285 1205 1315 1235
rect 1365 1205 1395 1235
rect 1445 1205 1475 1235
rect 1525 1205 1555 1235
rect 1685 1205 1715 1235
rect 1765 1205 1795 1235
rect 1845 1205 1875 1235
rect 1925 1205 1955 1235
rect 2005 1205 2035 1235
rect 2085 1205 2115 1235
rect 2165 1205 2195 1235
rect 2245 1205 2275 1235
rect 2325 1205 2355 1235
rect 2405 1205 2435 1235
rect 2485 1205 2515 1235
rect 2645 1205 2675 1235
rect 2725 1205 2755 1235
rect 2805 1205 2835 1235
rect 2885 1205 2915 1235
rect 2965 1205 2995 1235
rect 3045 1205 3075 1235
rect 3125 1205 3155 1235
rect 3205 1205 3235 1235
rect 3285 1205 3315 1235
rect 3365 1205 3395 1235
rect 3445 1205 3475 1235
rect 3605 1205 3635 1235
rect 3685 1205 3715 1235
rect 3765 1205 3795 1235
rect 3845 1205 3875 1235
rect 3925 1205 3955 1235
rect 4005 1205 4035 1235
rect 4085 1205 4115 1235
rect 4165 1205 4195 1235
rect 85 605 115 635
rect 165 605 195 635
rect 245 605 275 635
rect 325 605 355 635
rect 405 605 435 635
rect 485 605 515 635
rect 565 605 595 635
rect 725 605 755 635
rect 805 605 835 635
rect 885 605 915 635
rect 965 605 995 635
rect 1045 605 1075 635
rect 1125 605 1155 635
rect 1205 605 1235 635
rect 1285 605 1315 635
rect 1365 605 1395 635
rect 1445 605 1475 635
rect 1525 605 1555 635
rect 1685 605 1715 635
rect 1765 605 1795 635
rect 1845 605 1875 635
rect 1925 605 1955 635
rect 2005 605 2035 635
rect 2085 605 2115 635
rect 2165 605 2195 635
rect 2245 605 2275 635
rect 2325 605 2355 635
rect 2405 605 2435 635
rect 2485 605 2515 635
rect 2645 605 2675 635
rect 2725 605 2755 635
rect 2805 605 2835 635
rect 2885 605 2915 635
rect 2965 605 2995 635
rect 3045 605 3075 635
rect 3125 605 3155 635
rect 3205 605 3235 635
rect 3285 605 3315 635
rect 3365 605 3395 635
rect 3445 605 3475 635
rect 3605 605 3635 635
rect 3685 605 3715 635
rect 3765 605 3795 635
rect 3845 605 3875 635
rect 3925 605 3955 635
rect 4005 605 4035 635
rect 4085 605 4115 635
rect 85 445 115 475
rect 165 445 195 475
rect 245 445 275 475
rect 325 445 355 475
rect 405 445 435 475
rect 485 445 515 475
rect 565 445 595 475
rect 725 445 755 475
rect 805 445 835 475
rect 885 445 915 475
rect 965 445 995 475
rect 1045 445 1075 475
rect 1125 445 1155 475
rect 1205 445 1235 475
rect 1285 445 1315 475
rect 1365 445 1395 475
rect 1445 445 1475 475
rect 1525 445 1555 475
rect 1685 445 1715 475
rect 1765 445 1795 475
rect 1845 445 1875 475
rect 1925 445 1955 475
rect 2005 445 2035 475
rect 2085 445 2115 475
rect 2165 445 2195 475
rect 2245 445 2275 475
rect 2325 445 2355 475
rect 2405 445 2435 475
rect 2485 445 2515 475
rect 2645 445 2675 475
rect 2725 445 2755 475
rect 2805 445 2835 475
rect 2885 445 2915 475
rect 2965 445 2995 475
rect 3045 445 3075 475
rect 3125 445 3155 475
rect 3205 445 3235 475
rect 3285 445 3315 475
rect 3365 445 3395 475
rect 3445 445 3475 475
rect 3605 445 3635 475
rect 3685 445 3715 475
rect 3765 445 3795 475
rect 3845 445 3875 475
rect 3925 445 3955 475
rect 4085 445 4115 475
rect 85 285 115 315
rect 165 285 195 315
rect 245 285 275 315
rect 325 285 355 315
rect 405 285 435 315
rect 485 285 515 315
rect 565 285 595 315
rect 725 285 755 315
rect 805 285 835 315
rect 885 285 915 315
rect 965 285 995 315
rect 1045 285 1075 315
rect 1125 285 1155 315
rect 1205 285 1235 315
rect 1285 285 1315 315
rect 1365 285 1395 315
rect 1445 285 1475 315
rect 1525 285 1555 315
rect 1685 285 1715 315
rect 1765 285 1795 315
rect 1845 285 1875 315
rect 1925 285 1955 315
rect 2005 285 2035 315
rect 2085 285 2115 315
rect 2165 285 2195 315
rect 2245 285 2275 315
rect 2325 285 2355 315
rect 2405 285 2435 315
rect 2485 285 2515 315
rect 2645 285 2675 315
rect 2725 285 2755 315
rect 2805 285 2835 315
rect 2885 285 2915 315
rect 2965 285 2995 315
rect 3045 285 3075 315
rect 3125 285 3155 315
rect 3205 285 3235 315
rect 3285 285 3315 315
rect 3365 285 3395 315
rect 3445 285 3475 315
rect 3605 285 3635 315
rect 3685 285 3715 315
rect 3765 285 3795 315
rect 3845 285 3875 315
rect 3925 285 3955 315
rect 4005 285 4035 315
rect 4085 285 4115 315
rect 165 90 195 170
rect 85 -75 115 -45
rect 165 -75 195 -45
rect 245 -75 275 -45
rect 325 -75 355 -45
rect 405 -75 435 -45
rect 485 -75 515 -45
rect 565 -75 595 -45
rect 725 -75 755 -45
rect 805 -75 835 -45
rect 885 -75 915 -45
rect 965 -75 995 -45
rect 1045 -75 1075 -45
rect 1125 -75 1155 -45
rect 1205 -75 1235 -45
rect 1285 -75 1315 -45
rect 1365 -75 1395 -45
rect 1445 -75 1475 -45
rect 1525 -75 1555 -45
rect 1685 -75 1715 -45
rect 1765 -75 1795 -45
rect 1845 -75 1875 -45
rect 1925 -75 1955 -45
rect 2005 -75 2035 -45
rect 2085 -75 2115 -45
rect 2165 -75 2195 -45
rect 2245 -75 2275 -45
rect 2325 -75 2355 -45
rect 2405 -75 2435 -45
rect 2485 -75 2515 -45
rect 2645 -75 2675 -45
rect 2725 -75 2755 -45
rect 2805 -75 2835 -45
rect 2885 -75 2915 -45
rect 2965 -75 2995 -45
rect 3045 -75 3075 -45
rect 3125 -75 3155 -45
rect 3205 -75 3235 -45
rect 3285 -75 3315 -45
rect 3365 -75 3395 -45
rect 3445 -75 3475 -45
rect 3605 -75 3635 -45
rect 3685 -75 3715 -45
rect 3765 -75 3795 -45
rect 3845 -75 3875 -45
rect 3925 -75 3955 -45
rect 4085 -75 4115 -45
rect 85 -235 115 -205
rect 165 -235 195 -205
rect 245 -235 275 -205
rect 325 -235 355 -205
rect 405 -235 435 -205
rect 485 -235 515 -205
rect 565 -235 595 -205
rect 725 -235 755 -205
rect 805 -235 835 -205
rect 885 -235 915 -205
rect 965 -235 995 -205
rect 1045 -235 1075 -205
rect 1125 -235 1155 -205
rect 1205 -235 1235 -205
rect 1285 -235 1315 -205
rect 1365 -235 1395 -205
rect 1445 -235 1475 -205
rect 1525 -235 1555 -205
rect 1685 -235 1715 -205
rect 1765 -235 1795 -205
rect 1845 -235 1875 -205
rect 1925 -235 1955 -205
rect 2005 -235 2035 -205
rect 2085 -235 2115 -205
rect 2165 -235 2195 -205
rect 2245 -235 2275 -205
rect 2325 -235 2355 -205
rect 2405 -235 2435 -205
rect 2485 -235 2515 -205
rect 2645 -235 2675 -205
rect 2725 -235 2755 -205
rect 2805 -235 2835 -205
rect 2885 -235 2915 -205
rect 2965 -235 2995 -205
rect 3045 -235 3075 -205
rect 3125 -235 3155 -205
rect 3205 -235 3235 -205
rect 3285 -235 3315 -205
rect 3365 -235 3395 -205
rect 3445 -235 3475 -205
rect 3605 -235 3635 -205
rect 3685 -235 3715 -205
rect 3765 -235 3795 -205
rect 3845 -235 3875 -205
rect 3925 -235 3955 -205
rect 4085 -235 4115 -205
rect 165 -430 195 -350
<< metal3 >>
rect 160 4871 200 4880
rect 160 4689 164 4871
rect 196 4689 200 4871
rect 160 4680 200 4689
rect 80 4396 120 4400
rect 80 4364 84 4396
rect 116 4364 120 4396
rect 80 4316 120 4364
rect 80 4284 84 4316
rect 116 4284 120 4316
rect 80 4236 120 4284
rect 80 4204 84 4236
rect 116 4204 120 4236
rect 80 4200 120 4204
rect 160 4396 200 4400
rect 160 4364 164 4396
rect 196 4364 200 4396
rect 160 4316 200 4364
rect 160 4284 164 4316
rect 196 4284 200 4316
rect 160 4236 200 4284
rect 160 4204 164 4236
rect 196 4204 200 4236
rect 160 4200 200 4204
rect 240 4396 280 4400
rect 240 4364 244 4396
rect 276 4364 280 4396
rect 240 4316 280 4364
rect 240 4284 244 4316
rect 276 4284 280 4316
rect 240 4236 280 4284
rect 240 4204 244 4236
rect 276 4204 280 4236
rect 240 4200 280 4204
rect 320 4396 360 4400
rect 320 4364 324 4396
rect 356 4364 360 4396
rect 320 4316 360 4364
rect 320 4284 324 4316
rect 356 4284 360 4316
rect 320 4236 360 4284
rect 320 4204 324 4236
rect 356 4204 360 4236
rect 320 4200 360 4204
rect 400 4396 440 4400
rect 400 4364 404 4396
rect 436 4364 440 4396
rect 400 4316 440 4364
rect 400 4284 404 4316
rect 436 4284 440 4316
rect 400 4236 440 4284
rect 400 4204 404 4236
rect 436 4204 440 4236
rect 400 4200 440 4204
rect 480 4396 520 4400
rect 480 4364 484 4396
rect 516 4364 520 4396
rect 480 4316 520 4364
rect 480 4284 484 4316
rect 516 4284 520 4316
rect 480 4236 520 4284
rect 480 4204 484 4236
rect 516 4204 520 4236
rect 480 4200 520 4204
rect 560 4396 600 4400
rect 560 4364 564 4396
rect 596 4364 600 4396
rect 560 4316 600 4364
rect 560 4284 564 4316
rect 596 4284 600 4316
rect 560 4236 600 4284
rect 560 4204 564 4236
rect 596 4204 600 4236
rect 560 4200 600 4204
rect 720 4396 760 4400
rect 720 4364 724 4396
rect 756 4364 760 4396
rect 720 4316 760 4364
rect 720 4284 724 4316
rect 756 4284 760 4316
rect 720 4236 760 4284
rect 720 4204 724 4236
rect 756 4204 760 4236
rect 720 4200 760 4204
rect 800 4396 840 4400
rect 800 4364 804 4396
rect 836 4364 840 4396
rect 800 4316 840 4364
rect 800 4284 804 4316
rect 836 4284 840 4316
rect 800 4236 840 4284
rect 800 4204 804 4236
rect 836 4204 840 4236
rect 800 4200 840 4204
rect 880 4396 920 4400
rect 880 4364 884 4396
rect 916 4364 920 4396
rect 880 4316 920 4364
rect 880 4284 884 4316
rect 916 4284 920 4316
rect 880 4236 920 4284
rect 880 4204 884 4236
rect 916 4204 920 4236
rect 880 4200 920 4204
rect 960 4396 1000 4400
rect 960 4364 964 4396
rect 996 4364 1000 4396
rect 960 4316 1000 4364
rect 960 4284 964 4316
rect 996 4284 1000 4316
rect 960 4236 1000 4284
rect 960 4204 964 4236
rect 996 4204 1000 4236
rect 960 4200 1000 4204
rect 1040 4396 1080 4400
rect 1040 4364 1044 4396
rect 1076 4364 1080 4396
rect 1040 4316 1080 4364
rect 1040 4284 1044 4316
rect 1076 4284 1080 4316
rect 1040 4236 1080 4284
rect 1040 4204 1044 4236
rect 1076 4204 1080 4236
rect 1040 4200 1080 4204
rect 1120 4396 1160 4400
rect 1120 4364 1124 4396
rect 1156 4364 1160 4396
rect 1120 4316 1160 4364
rect 1120 4284 1124 4316
rect 1156 4284 1160 4316
rect 1120 4236 1160 4284
rect 1120 4204 1124 4236
rect 1156 4204 1160 4236
rect 1120 4200 1160 4204
rect 1200 4396 1240 4400
rect 1200 4364 1204 4396
rect 1236 4364 1240 4396
rect 1200 4316 1240 4364
rect 1200 4284 1204 4316
rect 1236 4284 1240 4316
rect 1200 4236 1240 4284
rect 1200 4204 1204 4236
rect 1236 4204 1240 4236
rect 1200 4200 1240 4204
rect 1280 4396 1320 4400
rect 1280 4364 1284 4396
rect 1316 4364 1320 4396
rect 1280 4316 1320 4364
rect 1280 4284 1284 4316
rect 1316 4284 1320 4316
rect 1280 4236 1320 4284
rect 1280 4204 1284 4236
rect 1316 4204 1320 4236
rect 1280 4200 1320 4204
rect 1360 4396 1400 4400
rect 1360 4364 1364 4396
rect 1396 4364 1400 4396
rect 1360 4316 1400 4364
rect 1360 4284 1364 4316
rect 1396 4284 1400 4316
rect 1360 4236 1400 4284
rect 1360 4204 1364 4236
rect 1396 4204 1400 4236
rect 1360 4200 1400 4204
rect 1440 4396 1480 4400
rect 1440 4364 1444 4396
rect 1476 4364 1480 4396
rect 1440 4316 1480 4364
rect 1440 4284 1444 4316
rect 1476 4284 1480 4316
rect 1440 4236 1480 4284
rect 1440 4204 1444 4236
rect 1476 4204 1480 4236
rect 1440 4200 1480 4204
rect 1520 4396 1560 4400
rect 1520 4364 1524 4396
rect 1556 4364 1560 4396
rect 1520 4316 1560 4364
rect 1520 4284 1524 4316
rect 1556 4284 1560 4316
rect 1520 4236 1560 4284
rect 1520 4204 1524 4236
rect 1556 4204 1560 4236
rect 1520 4200 1560 4204
rect 1680 4396 1720 4400
rect 1680 4364 1684 4396
rect 1716 4364 1720 4396
rect 1680 4316 1720 4364
rect 1680 4284 1684 4316
rect 1716 4284 1720 4316
rect 1680 4236 1720 4284
rect 1680 4204 1684 4236
rect 1716 4204 1720 4236
rect 1680 4200 1720 4204
rect 1760 4396 1800 4400
rect 1760 4364 1764 4396
rect 1796 4364 1800 4396
rect 1760 4316 1800 4364
rect 1760 4284 1764 4316
rect 1796 4284 1800 4316
rect 1760 4236 1800 4284
rect 1760 4204 1764 4236
rect 1796 4204 1800 4236
rect 1760 4200 1800 4204
rect 1840 4396 1880 4400
rect 1840 4364 1844 4396
rect 1876 4364 1880 4396
rect 1840 4316 1880 4364
rect 1840 4284 1844 4316
rect 1876 4284 1880 4316
rect 1840 4236 1880 4284
rect 1840 4204 1844 4236
rect 1876 4204 1880 4236
rect 1840 4200 1880 4204
rect 1920 4396 1960 4400
rect 1920 4364 1924 4396
rect 1956 4364 1960 4396
rect 1920 4316 1960 4364
rect 1920 4284 1924 4316
rect 1956 4284 1960 4316
rect 1920 4236 1960 4284
rect 1920 4204 1924 4236
rect 1956 4204 1960 4236
rect 1920 4200 1960 4204
rect 2000 4396 2040 4400
rect 2000 4364 2004 4396
rect 2036 4364 2040 4396
rect 2000 4316 2040 4364
rect 2000 4284 2004 4316
rect 2036 4284 2040 4316
rect 2000 4236 2040 4284
rect 2000 4204 2004 4236
rect 2036 4204 2040 4236
rect 2000 4200 2040 4204
rect 2080 4396 2120 4400
rect 2080 4364 2084 4396
rect 2116 4364 2120 4396
rect 2080 4316 2120 4364
rect 2080 4284 2084 4316
rect 2116 4284 2120 4316
rect 2080 4236 2120 4284
rect 2080 4204 2084 4236
rect 2116 4204 2120 4236
rect 2080 4200 2120 4204
rect 2160 4396 2200 4400
rect 2160 4364 2164 4396
rect 2196 4364 2200 4396
rect 2160 4316 2200 4364
rect 2160 4284 2164 4316
rect 2196 4284 2200 4316
rect 2160 4236 2200 4284
rect 2160 4204 2164 4236
rect 2196 4204 2200 4236
rect 2160 4200 2200 4204
rect 2240 4396 2280 4400
rect 2240 4364 2244 4396
rect 2276 4364 2280 4396
rect 2240 4316 2280 4364
rect 2240 4284 2244 4316
rect 2276 4284 2280 4316
rect 2240 4236 2280 4284
rect 2240 4204 2244 4236
rect 2276 4204 2280 4236
rect 2240 4200 2280 4204
rect 2320 4396 2360 4400
rect 2320 4364 2324 4396
rect 2356 4364 2360 4396
rect 2320 4316 2360 4364
rect 2320 4284 2324 4316
rect 2356 4284 2360 4316
rect 2320 4236 2360 4284
rect 2320 4204 2324 4236
rect 2356 4204 2360 4236
rect 2320 4200 2360 4204
rect 2400 4396 2440 4400
rect 2400 4364 2404 4396
rect 2436 4364 2440 4396
rect 2400 4316 2440 4364
rect 2400 4284 2404 4316
rect 2436 4284 2440 4316
rect 2400 4236 2440 4284
rect 2400 4204 2404 4236
rect 2436 4204 2440 4236
rect 2400 4200 2440 4204
rect 2480 4396 2520 4400
rect 2480 4364 2484 4396
rect 2516 4364 2520 4396
rect 2480 4316 2520 4364
rect 2480 4284 2484 4316
rect 2516 4284 2520 4316
rect 2480 4236 2520 4284
rect 2480 4204 2484 4236
rect 2516 4204 2520 4236
rect 2480 4200 2520 4204
rect 2640 4396 2680 4400
rect 2640 4364 2644 4396
rect 2676 4364 2680 4396
rect 2640 4316 2680 4364
rect 2640 4284 2644 4316
rect 2676 4284 2680 4316
rect 2640 4236 2680 4284
rect 2640 4204 2644 4236
rect 2676 4204 2680 4236
rect 2640 4200 2680 4204
rect 2720 4396 2760 4400
rect 2720 4364 2724 4396
rect 2756 4364 2760 4396
rect 2720 4316 2760 4364
rect 2720 4284 2724 4316
rect 2756 4284 2760 4316
rect 2720 4236 2760 4284
rect 2720 4204 2724 4236
rect 2756 4204 2760 4236
rect 2720 4200 2760 4204
rect 2800 4396 2840 4400
rect 2800 4364 2804 4396
rect 2836 4364 2840 4396
rect 2800 4316 2840 4364
rect 2800 4284 2804 4316
rect 2836 4284 2840 4316
rect 2800 4236 2840 4284
rect 2800 4204 2804 4236
rect 2836 4204 2840 4236
rect 2800 4200 2840 4204
rect 2880 4396 2920 4400
rect 2880 4364 2884 4396
rect 2916 4364 2920 4396
rect 2880 4316 2920 4364
rect 2880 4284 2884 4316
rect 2916 4284 2920 4316
rect 2880 4236 2920 4284
rect 2880 4204 2884 4236
rect 2916 4204 2920 4236
rect 2880 4200 2920 4204
rect 2960 4396 3000 4400
rect 2960 4364 2964 4396
rect 2996 4364 3000 4396
rect 2960 4316 3000 4364
rect 2960 4284 2964 4316
rect 2996 4284 3000 4316
rect 2960 4236 3000 4284
rect 2960 4204 2964 4236
rect 2996 4204 3000 4236
rect 2960 4200 3000 4204
rect 3040 4396 3080 4400
rect 3040 4364 3044 4396
rect 3076 4364 3080 4396
rect 3040 4316 3080 4364
rect 3040 4284 3044 4316
rect 3076 4284 3080 4316
rect 3040 4236 3080 4284
rect 3040 4204 3044 4236
rect 3076 4204 3080 4236
rect 3040 4200 3080 4204
rect 3120 4396 3160 4400
rect 3120 4364 3124 4396
rect 3156 4364 3160 4396
rect 3120 4316 3160 4364
rect 3120 4284 3124 4316
rect 3156 4284 3160 4316
rect 3120 4236 3160 4284
rect 3120 4204 3124 4236
rect 3156 4204 3160 4236
rect 3120 4200 3160 4204
rect 3200 4396 3240 4400
rect 3200 4364 3204 4396
rect 3236 4364 3240 4396
rect 3200 4316 3240 4364
rect 3200 4284 3204 4316
rect 3236 4284 3240 4316
rect 3200 4236 3240 4284
rect 3200 4204 3204 4236
rect 3236 4204 3240 4236
rect 3200 4200 3240 4204
rect 3280 4396 3320 4400
rect 3280 4364 3284 4396
rect 3316 4364 3320 4396
rect 3280 4316 3320 4364
rect 3280 4284 3284 4316
rect 3316 4284 3320 4316
rect 3280 4236 3320 4284
rect 3280 4204 3284 4236
rect 3316 4204 3320 4236
rect 3280 4200 3320 4204
rect 3360 4396 3400 4400
rect 3360 4364 3364 4396
rect 3396 4364 3400 4396
rect 3360 4316 3400 4364
rect 3360 4284 3364 4316
rect 3396 4284 3400 4316
rect 3360 4236 3400 4284
rect 3360 4204 3364 4236
rect 3396 4204 3400 4236
rect 3360 4200 3400 4204
rect 3440 4396 3480 4400
rect 3440 4364 3444 4396
rect 3476 4364 3480 4396
rect 3440 4316 3480 4364
rect 3440 4284 3444 4316
rect 3476 4284 3480 4316
rect 3440 4236 3480 4284
rect 3440 4204 3444 4236
rect 3476 4204 3480 4236
rect 3440 4200 3480 4204
rect 3600 4396 3640 4400
rect 3600 4364 3604 4396
rect 3636 4364 3640 4396
rect 3600 4316 3640 4364
rect 3600 4284 3604 4316
rect 3636 4284 3640 4316
rect 3600 4236 3640 4284
rect 3600 4204 3604 4236
rect 3636 4204 3640 4236
rect 3600 4200 3640 4204
rect 3680 4396 3720 4400
rect 3680 4364 3684 4396
rect 3716 4364 3720 4396
rect 3680 4316 3720 4364
rect 3680 4284 3684 4316
rect 3716 4284 3720 4316
rect 3680 4236 3720 4284
rect 3680 4204 3684 4236
rect 3716 4204 3720 4236
rect 3680 4200 3720 4204
rect 3760 4396 3800 4400
rect 3760 4364 3764 4396
rect 3796 4364 3800 4396
rect 3760 4316 3800 4364
rect 3760 4284 3764 4316
rect 3796 4284 3800 4316
rect 3760 4236 3800 4284
rect 3760 4204 3764 4236
rect 3796 4204 3800 4236
rect 3760 4200 3800 4204
rect 3840 4396 3880 4400
rect 3840 4364 3844 4396
rect 3876 4364 3880 4396
rect 3840 4316 3880 4364
rect 3840 4284 3844 4316
rect 3876 4284 3880 4316
rect 3840 4236 3880 4284
rect 3840 4204 3844 4236
rect 3876 4204 3880 4236
rect 3840 4200 3880 4204
rect 3920 4396 3960 4400
rect 3920 4364 3924 4396
rect 3956 4364 3960 4396
rect 3920 4316 3960 4364
rect 3920 4284 3924 4316
rect 3956 4284 3960 4316
rect 3920 4236 3960 4284
rect 3920 4204 3924 4236
rect 3956 4204 3960 4236
rect 3920 4200 3960 4204
rect 4000 4396 4040 4400
rect 4000 4364 4004 4396
rect 4036 4364 4040 4396
rect 4000 4316 4040 4364
rect 4000 4284 4004 4316
rect 4036 4284 4040 4316
rect 4000 4236 4040 4284
rect 4000 4204 4004 4236
rect 4036 4204 4040 4236
rect 4000 4200 4040 4204
rect 4080 4396 4120 4400
rect 4080 4364 4084 4396
rect 4116 4364 4120 4396
rect 4080 4316 4120 4364
rect 4080 4284 4084 4316
rect 4116 4284 4120 4316
rect 4080 4236 4120 4284
rect 4080 4204 4084 4236
rect 4116 4204 4120 4236
rect 4080 4200 4120 4204
rect 80 4156 120 4160
rect 80 4124 84 4156
rect 116 4124 120 4156
rect 80 4076 120 4124
rect 80 4044 84 4076
rect 116 4044 120 4076
rect 80 3996 120 4044
rect 80 3964 84 3996
rect 116 3964 120 3996
rect 80 3960 120 3964
rect 160 4156 200 4160
rect 160 4124 164 4156
rect 196 4124 200 4156
rect 160 4076 200 4124
rect 160 4044 164 4076
rect 196 4044 200 4076
rect 160 3996 200 4044
rect 160 3964 164 3996
rect 196 3964 200 3996
rect 160 3960 200 3964
rect 240 4156 280 4160
rect 240 4124 244 4156
rect 276 4124 280 4156
rect 240 4076 280 4124
rect 240 4044 244 4076
rect 276 4044 280 4076
rect 240 3996 280 4044
rect 240 3964 244 3996
rect 276 3964 280 3996
rect 240 3960 280 3964
rect 320 4156 360 4160
rect 320 4124 324 4156
rect 356 4124 360 4156
rect 320 4076 360 4124
rect 320 4044 324 4076
rect 356 4044 360 4076
rect 320 3996 360 4044
rect 320 3964 324 3996
rect 356 3964 360 3996
rect 320 3960 360 3964
rect 400 4156 440 4160
rect 400 4124 404 4156
rect 436 4124 440 4156
rect 400 4076 440 4124
rect 400 4044 404 4076
rect 436 4044 440 4076
rect 400 3996 440 4044
rect 400 3964 404 3996
rect 436 3964 440 3996
rect 400 3960 440 3964
rect 480 4156 520 4160
rect 480 4124 484 4156
rect 516 4124 520 4156
rect 480 4076 520 4124
rect 480 4044 484 4076
rect 516 4044 520 4076
rect 480 3996 520 4044
rect 480 3964 484 3996
rect 516 3964 520 3996
rect 480 3960 520 3964
rect 560 4156 600 4160
rect 560 4124 564 4156
rect 596 4124 600 4156
rect 560 4076 600 4124
rect 560 4044 564 4076
rect 596 4044 600 4076
rect 560 3996 600 4044
rect 560 3964 564 3996
rect 596 3964 600 3996
rect 560 3960 600 3964
rect 720 4156 760 4160
rect 720 4124 724 4156
rect 756 4124 760 4156
rect 720 4076 760 4124
rect 720 4044 724 4076
rect 756 4044 760 4076
rect 720 3996 760 4044
rect 720 3964 724 3996
rect 756 3964 760 3996
rect 720 3960 760 3964
rect 800 4156 840 4160
rect 800 4124 804 4156
rect 836 4124 840 4156
rect 800 4076 840 4124
rect 800 4044 804 4076
rect 836 4044 840 4076
rect 800 3996 840 4044
rect 800 3964 804 3996
rect 836 3964 840 3996
rect 800 3960 840 3964
rect 880 4156 920 4160
rect 880 4124 884 4156
rect 916 4124 920 4156
rect 880 4076 920 4124
rect 880 4044 884 4076
rect 916 4044 920 4076
rect 880 3996 920 4044
rect 880 3964 884 3996
rect 916 3964 920 3996
rect 880 3960 920 3964
rect 960 4156 1000 4160
rect 960 4124 964 4156
rect 996 4124 1000 4156
rect 960 4076 1000 4124
rect 960 4044 964 4076
rect 996 4044 1000 4076
rect 960 3996 1000 4044
rect 960 3964 964 3996
rect 996 3964 1000 3996
rect 960 3960 1000 3964
rect 1040 4156 1080 4160
rect 1040 4124 1044 4156
rect 1076 4124 1080 4156
rect 1040 4076 1080 4124
rect 1040 4044 1044 4076
rect 1076 4044 1080 4076
rect 1040 3996 1080 4044
rect 1040 3964 1044 3996
rect 1076 3964 1080 3996
rect 1040 3960 1080 3964
rect 1120 4156 1160 4160
rect 1120 4124 1124 4156
rect 1156 4124 1160 4156
rect 1120 4076 1160 4124
rect 1120 4044 1124 4076
rect 1156 4044 1160 4076
rect 1120 3996 1160 4044
rect 1120 3964 1124 3996
rect 1156 3964 1160 3996
rect 1120 3960 1160 3964
rect 1200 4156 1240 4160
rect 1200 4124 1204 4156
rect 1236 4124 1240 4156
rect 1200 4076 1240 4124
rect 1200 4044 1204 4076
rect 1236 4044 1240 4076
rect 1200 3996 1240 4044
rect 1200 3964 1204 3996
rect 1236 3964 1240 3996
rect 1200 3960 1240 3964
rect 1280 4156 1320 4160
rect 1280 4124 1284 4156
rect 1316 4124 1320 4156
rect 1280 4076 1320 4124
rect 1280 4044 1284 4076
rect 1316 4044 1320 4076
rect 1280 3996 1320 4044
rect 1280 3964 1284 3996
rect 1316 3964 1320 3996
rect 1280 3960 1320 3964
rect 1360 4156 1400 4160
rect 1360 4124 1364 4156
rect 1396 4124 1400 4156
rect 1360 4076 1400 4124
rect 1360 4044 1364 4076
rect 1396 4044 1400 4076
rect 1360 3996 1400 4044
rect 1360 3964 1364 3996
rect 1396 3964 1400 3996
rect 1360 3960 1400 3964
rect 1440 4156 1480 4160
rect 1440 4124 1444 4156
rect 1476 4124 1480 4156
rect 1440 4076 1480 4124
rect 1440 4044 1444 4076
rect 1476 4044 1480 4076
rect 1440 3996 1480 4044
rect 1440 3964 1444 3996
rect 1476 3964 1480 3996
rect 1440 3960 1480 3964
rect 1520 4156 1560 4160
rect 1520 4124 1524 4156
rect 1556 4124 1560 4156
rect 1520 4076 1560 4124
rect 1520 4044 1524 4076
rect 1556 4044 1560 4076
rect 1520 3996 1560 4044
rect 1520 3964 1524 3996
rect 1556 3964 1560 3996
rect 1520 3960 1560 3964
rect 1680 4156 1720 4160
rect 1680 4124 1684 4156
rect 1716 4124 1720 4156
rect 1680 4076 1720 4124
rect 1680 4044 1684 4076
rect 1716 4044 1720 4076
rect 1680 3996 1720 4044
rect 1680 3964 1684 3996
rect 1716 3964 1720 3996
rect 1680 3960 1720 3964
rect 1760 4156 1800 4160
rect 1760 4124 1764 4156
rect 1796 4124 1800 4156
rect 1760 4076 1800 4124
rect 1760 4044 1764 4076
rect 1796 4044 1800 4076
rect 1760 3996 1800 4044
rect 1760 3964 1764 3996
rect 1796 3964 1800 3996
rect 1760 3960 1800 3964
rect 1840 4156 1880 4160
rect 1840 4124 1844 4156
rect 1876 4124 1880 4156
rect 1840 4076 1880 4124
rect 1840 4044 1844 4076
rect 1876 4044 1880 4076
rect 1840 3996 1880 4044
rect 1840 3964 1844 3996
rect 1876 3964 1880 3996
rect 1840 3960 1880 3964
rect 1920 4156 1960 4160
rect 1920 4124 1924 4156
rect 1956 4124 1960 4156
rect 1920 4076 1960 4124
rect 1920 4044 1924 4076
rect 1956 4044 1960 4076
rect 1920 3996 1960 4044
rect 1920 3964 1924 3996
rect 1956 3964 1960 3996
rect 1920 3960 1960 3964
rect 2000 4156 2040 4160
rect 2000 4124 2004 4156
rect 2036 4124 2040 4156
rect 2000 4076 2040 4124
rect 2000 4044 2004 4076
rect 2036 4044 2040 4076
rect 2000 3996 2040 4044
rect 2000 3964 2004 3996
rect 2036 3964 2040 3996
rect 2000 3960 2040 3964
rect 2080 4156 2120 4160
rect 2080 4124 2084 4156
rect 2116 4124 2120 4156
rect 2080 4076 2120 4124
rect 2080 4044 2084 4076
rect 2116 4044 2120 4076
rect 2080 3996 2120 4044
rect 2080 3964 2084 3996
rect 2116 3964 2120 3996
rect 2080 3960 2120 3964
rect 2160 4156 2200 4160
rect 2160 4124 2164 4156
rect 2196 4124 2200 4156
rect 2160 4076 2200 4124
rect 2160 4044 2164 4076
rect 2196 4044 2200 4076
rect 2160 3996 2200 4044
rect 2160 3964 2164 3996
rect 2196 3964 2200 3996
rect 2160 3960 2200 3964
rect 2240 4156 2280 4160
rect 2240 4124 2244 4156
rect 2276 4124 2280 4156
rect 2240 4076 2280 4124
rect 2240 4044 2244 4076
rect 2276 4044 2280 4076
rect 2240 3996 2280 4044
rect 2240 3964 2244 3996
rect 2276 3964 2280 3996
rect 2240 3960 2280 3964
rect 2320 4156 2360 4160
rect 2320 4124 2324 4156
rect 2356 4124 2360 4156
rect 2320 4076 2360 4124
rect 2320 4044 2324 4076
rect 2356 4044 2360 4076
rect 2320 3996 2360 4044
rect 2320 3964 2324 3996
rect 2356 3964 2360 3996
rect 2320 3960 2360 3964
rect 2400 4156 2440 4160
rect 2400 4124 2404 4156
rect 2436 4124 2440 4156
rect 2400 4076 2440 4124
rect 2400 4044 2404 4076
rect 2436 4044 2440 4076
rect 2400 3996 2440 4044
rect 2400 3964 2404 3996
rect 2436 3964 2440 3996
rect 2400 3960 2440 3964
rect 2480 4156 2520 4160
rect 2480 4124 2484 4156
rect 2516 4124 2520 4156
rect 2480 4076 2520 4124
rect 2480 4044 2484 4076
rect 2516 4044 2520 4076
rect 2480 3996 2520 4044
rect 2480 3964 2484 3996
rect 2516 3964 2520 3996
rect 2480 3960 2520 3964
rect 2640 4156 2680 4160
rect 2640 4124 2644 4156
rect 2676 4124 2680 4156
rect 2640 4076 2680 4124
rect 2640 4044 2644 4076
rect 2676 4044 2680 4076
rect 2640 3996 2680 4044
rect 2640 3964 2644 3996
rect 2676 3964 2680 3996
rect 2640 3960 2680 3964
rect 2720 4156 2760 4160
rect 2720 4124 2724 4156
rect 2756 4124 2760 4156
rect 2720 4076 2760 4124
rect 2720 4044 2724 4076
rect 2756 4044 2760 4076
rect 2720 3996 2760 4044
rect 2720 3964 2724 3996
rect 2756 3964 2760 3996
rect 2720 3960 2760 3964
rect 2800 4156 2840 4160
rect 2800 4124 2804 4156
rect 2836 4124 2840 4156
rect 2800 4076 2840 4124
rect 2800 4044 2804 4076
rect 2836 4044 2840 4076
rect 2800 3996 2840 4044
rect 2800 3964 2804 3996
rect 2836 3964 2840 3996
rect 2800 3960 2840 3964
rect 2880 4156 2920 4160
rect 2880 4124 2884 4156
rect 2916 4124 2920 4156
rect 2880 4076 2920 4124
rect 2880 4044 2884 4076
rect 2916 4044 2920 4076
rect 2880 3996 2920 4044
rect 2880 3964 2884 3996
rect 2916 3964 2920 3996
rect 2880 3960 2920 3964
rect 2960 4156 3000 4160
rect 2960 4124 2964 4156
rect 2996 4124 3000 4156
rect 2960 4076 3000 4124
rect 2960 4044 2964 4076
rect 2996 4044 3000 4076
rect 2960 3996 3000 4044
rect 2960 3964 2964 3996
rect 2996 3964 3000 3996
rect 2960 3960 3000 3964
rect 3040 4156 3080 4160
rect 3040 4124 3044 4156
rect 3076 4124 3080 4156
rect 3040 4076 3080 4124
rect 3040 4044 3044 4076
rect 3076 4044 3080 4076
rect 3040 3996 3080 4044
rect 3040 3964 3044 3996
rect 3076 3964 3080 3996
rect 3040 3960 3080 3964
rect 3120 4156 3160 4160
rect 3120 4124 3124 4156
rect 3156 4124 3160 4156
rect 3120 4076 3160 4124
rect 3120 4044 3124 4076
rect 3156 4044 3160 4076
rect 3120 3996 3160 4044
rect 3120 3964 3124 3996
rect 3156 3964 3160 3996
rect 3120 3960 3160 3964
rect 3200 4156 3240 4160
rect 3200 4124 3204 4156
rect 3236 4124 3240 4156
rect 3200 4076 3240 4124
rect 3200 4044 3204 4076
rect 3236 4044 3240 4076
rect 3200 3996 3240 4044
rect 3200 3964 3204 3996
rect 3236 3964 3240 3996
rect 3200 3960 3240 3964
rect 3280 4156 3320 4160
rect 3280 4124 3284 4156
rect 3316 4124 3320 4156
rect 3280 4076 3320 4124
rect 3280 4044 3284 4076
rect 3316 4044 3320 4076
rect 3280 3996 3320 4044
rect 3280 3964 3284 3996
rect 3316 3964 3320 3996
rect 3280 3960 3320 3964
rect 3360 4156 3400 4160
rect 3360 4124 3364 4156
rect 3396 4124 3400 4156
rect 3360 4076 3400 4124
rect 3360 4044 3364 4076
rect 3396 4044 3400 4076
rect 3360 3996 3400 4044
rect 3360 3964 3364 3996
rect 3396 3964 3400 3996
rect 3360 3960 3400 3964
rect 3440 4156 3480 4160
rect 3440 4124 3444 4156
rect 3476 4124 3480 4156
rect 3440 4076 3480 4124
rect 3440 4044 3444 4076
rect 3476 4044 3480 4076
rect 3440 3996 3480 4044
rect 3440 3964 3444 3996
rect 3476 3964 3480 3996
rect 3440 3960 3480 3964
rect 3600 4156 3640 4160
rect 3600 4124 3604 4156
rect 3636 4124 3640 4156
rect 3600 4076 3640 4124
rect 3600 4044 3604 4076
rect 3636 4044 3640 4076
rect 3600 3996 3640 4044
rect 3600 3964 3604 3996
rect 3636 3964 3640 3996
rect 3600 3960 3640 3964
rect 3680 4156 3720 4160
rect 3680 4124 3684 4156
rect 3716 4124 3720 4156
rect 3680 4076 3720 4124
rect 3680 4044 3684 4076
rect 3716 4044 3720 4076
rect 3680 3996 3720 4044
rect 3680 3964 3684 3996
rect 3716 3964 3720 3996
rect 3680 3960 3720 3964
rect 3760 4156 3800 4160
rect 3760 4124 3764 4156
rect 3796 4124 3800 4156
rect 3760 4076 3800 4124
rect 3760 4044 3764 4076
rect 3796 4044 3800 4076
rect 3760 3996 3800 4044
rect 3760 3964 3764 3996
rect 3796 3964 3800 3996
rect 3760 3960 3800 3964
rect 3840 4156 3880 4160
rect 3840 4124 3844 4156
rect 3876 4124 3880 4156
rect 3840 4076 3880 4124
rect 3840 4044 3844 4076
rect 3876 4044 3880 4076
rect 3840 3996 3880 4044
rect 3840 3964 3844 3996
rect 3876 3964 3880 3996
rect 3840 3960 3880 3964
rect 3920 4156 3960 4160
rect 3920 4124 3924 4156
rect 3956 4124 3960 4156
rect 3920 4076 3960 4124
rect 3920 4044 3924 4076
rect 3956 4044 3960 4076
rect 3920 3996 3960 4044
rect 3920 3964 3924 3996
rect 3956 3964 3960 3996
rect 3920 3960 3960 3964
rect 4000 4156 4040 4160
rect 4000 4124 4004 4156
rect 4036 4124 4040 4156
rect 4000 4076 4040 4124
rect 4000 4044 4004 4076
rect 4036 4044 4040 4076
rect 4000 3996 4040 4044
rect 4000 3964 4004 3996
rect 4036 3964 4040 3996
rect 4000 3960 4040 3964
rect 4080 4156 4120 4160
rect 4080 4124 4084 4156
rect 4116 4124 4120 4156
rect 4080 4076 4120 4124
rect 4080 4044 4084 4076
rect 4116 4044 4120 4076
rect 4080 3996 4120 4044
rect 4080 3964 4084 3996
rect 4116 3964 4120 3996
rect 4080 3960 4120 3964
rect 160 3851 200 3860
rect 160 3769 164 3851
rect 196 3769 200 3851
rect 160 3760 200 3769
rect 160 3551 200 3560
rect 160 3469 164 3551
rect 196 3469 200 3551
rect 160 3460 200 3469
rect 80 3356 120 3360
rect 80 3324 84 3356
rect 116 3324 120 3356
rect 80 3276 120 3324
rect 80 3244 84 3276
rect 116 3244 120 3276
rect 80 3196 120 3244
rect 80 3164 84 3196
rect 116 3164 120 3196
rect 80 3160 120 3164
rect 160 3356 200 3360
rect 160 3324 164 3356
rect 196 3324 200 3356
rect 160 3276 200 3324
rect 160 3244 164 3276
rect 196 3244 200 3276
rect 160 3196 200 3244
rect 160 3164 164 3196
rect 196 3164 200 3196
rect 160 3160 200 3164
rect 240 3356 280 3360
rect 240 3324 244 3356
rect 276 3324 280 3356
rect 240 3276 280 3324
rect 240 3244 244 3276
rect 276 3244 280 3276
rect 240 3196 280 3244
rect 240 3164 244 3196
rect 276 3164 280 3196
rect 240 3160 280 3164
rect 320 3356 360 3360
rect 320 3324 324 3356
rect 356 3324 360 3356
rect 320 3276 360 3324
rect 320 3244 324 3276
rect 356 3244 360 3276
rect 320 3196 360 3244
rect 320 3164 324 3196
rect 356 3164 360 3196
rect 320 3160 360 3164
rect 400 3356 440 3360
rect 400 3324 404 3356
rect 436 3324 440 3356
rect 400 3276 440 3324
rect 400 3244 404 3276
rect 436 3244 440 3276
rect 400 3196 440 3244
rect 400 3164 404 3196
rect 436 3164 440 3196
rect 400 3160 440 3164
rect 480 3356 520 3360
rect 480 3324 484 3356
rect 516 3324 520 3356
rect 480 3276 520 3324
rect 480 3244 484 3276
rect 516 3244 520 3276
rect 480 3196 520 3244
rect 480 3164 484 3196
rect 516 3164 520 3196
rect 480 3160 520 3164
rect 560 3356 600 3360
rect 560 3324 564 3356
rect 596 3324 600 3356
rect 560 3276 600 3324
rect 560 3244 564 3276
rect 596 3244 600 3276
rect 560 3196 600 3244
rect 560 3164 564 3196
rect 596 3164 600 3196
rect 560 3160 600 3164
rect 720 3356 760 3360
rect 720 3324 724 3356
rect 756 3324 760 3356
rect 720 3276 760 3324
rect 720 3244 724 3276
rect 756 3244 760 3276
rect 720 3196 760 3244
rect 720 3164 724 3196
rect 756 3164 760 3196
rect 720 3160 760 3164
rect 800 3356 840 3360
rect 800 3324 804 3356
rect 836 3324 840 3356
rect 800 3276 840 3324
rect 800 3244 804 3276
rect 836 3244 840 3276
rect 800 3196 840 3244
rect 800 3164 804 3196
rect 836 3164 840 3196
rect 800 3160 840 3164
rect 880 3356 920 3360
rect 880 3324 884 3356
rect 916 3324 920 3356
rect 880 3276 920 3324
rect 880 3244 884 3276
rect 916 3244 920 3276
rect 880 3196 920 3244
rect 880 3164 884 3196
rect 916 3164 920 3196
rect 880 3160 920 3164
rect 960 3356 1000 3360
rect 960 3324 964 3356
rect 996 3324 1000 3356
rect 960 3276 1000 3324
rect 960 3244 964 3276
rect 996 3244 1000 3276
rect 960 3196 1000 3244
rect 960 3164 964 3196
rect 996 3164 1000 3196
rect 960 3160 1000 3164
rect 1040 3356 1080 3360
rect 1040 3324 1044 3356
rect 1076 3324 1080 3356
rect 1040 3276 1080 3324
rect 1040 3244 1044 3276
rect 1076 3244 1080 3276
rect 1040 3196 1080 3244
rect 1040 3164 1044 3196
rect 1076 3164 1080 3196
rect 1040 3160 1080 3164
rect 1120 3356 1160 3360
rect 1120 3324 1124 3356
rect 1156 3324 1160 3356
rect 1120 3276 1160 3324
rect 1120 3244 1124 3276
rect 1156 3244 1160 3276
rect 1120 3196 1160 3244
rect 1120 3164 1124 3196
rect 1156 3164 1160 3196
rect 1120 3160 1160 3164
rect 1200 3356 1240 3360
rect 1200 3324 1204 3356
rect 1236 3324 1240 3356
rect 1200 3276 1240 3324
rect 1200 3244 1204 3276
rect 1236 3244 1240 3276
rect 1200 3196 1240 3244
rect 1200 3164 1204 3196
rect 1236 3164 1240 3196
rect 1200 3160 1240 3164
rect 1280 3356 1320 3360
rect 1280 3324 1284 3356
rect 1316 3324 1320 3356
rect 1280 3276 1320 3324
rect 1280 3244 1284 3276
rect 1316 3244 1320 3276
rect 1280 3196 1320 3244
rect 1280 3164 1284 3196
rect 1316 3164 1320 3196
rect 1280 3160 1320 3164
rect 1360 3356 1400 3360
rect 1360 3324 1364 3356
rect 1396 3324 1400 3356
rect 1360 3276 1400 3324
rect 1360 3244 1364 3276
rect 1396 3244 1400 3276
rect 1360 3196 1400 3244
rect 1360 3164 1364 3196
rect 1396 3164 1400 3196
rect 1360 3160 1400 3164
rect 1440 3356 1480 3360
rect 1440 3324 1444 3356
rect 1476 3324 1480 3356
rect 1440 3276 1480 3324
rect 1440 3244 1444 3276
rect 1476 3244 1480 3276
rect 1440 3196 1480 3244
rect 1440 3164 1444 3196
rect 1476 3164 1480 3196
rect 1440 3160 1480 3164
rect 1520 3356 1560 3360
rect 1520 3324 1524 3356
rect 1556 3324 1560 3356
rect 1520 3276 1560 3324
rect 1520 3244 1524 3276
rect 1556 3244 1560 3276
rect 1520 3196 1560 3244
rect 1520 3164 1524 3196
rect 1556 3164 1560 3196
rect 1520 3160 1560 3164
rect 1680 3356 1720 3360
rect 1680 3324 1684 3356
rect 1716 3324 1720 3356
rect 1680 3276 1720 3324
rect 1680 3244 1684 3276
rect 1716 3244 1720 3276
rect 1680 3196 1720 3244
rect 1680 3164 1684 3196
rect 1716 3164 1720 3196
rect 1680 3160 1720 3164
rect 1760 3356 1800 3360
rect 1760 3324 1764 3356
rect 1796 3324 1800 3356
rect 1760 3276 1800 3324
rect 1760 3244 1764 3276
rect 1796 3244 1800 3276
rect 1760 3196 1800 3244
rect 1760 3164 1764 3196
rect 1796 3164 1800 3196
rect 1760 3160 1800 3164
rect 1840 3356 1880 3360
rect 1840 3324 1844 3356
rect 1876 3324 1880 3356
rect 1840 3276 1880 3324
rect 1840 3244 1844 3276
rect 1876 3244 1880 3276
rect 1840 3196 1880 3244
rect 1840 3164 1844 3196
rect 1876 3164 1880 3196
rect 1840 3160 1880 3164
rect 1920 3356 1960 3360
rect 1920 3324 1924 3356
rect 1956 3324 1960 3356
rect 1920 3276 1960 3324
rect 1920 3244 1924 3276
rect 1956 3244 1960 3276
rect 1920 3196 1960 3244
rect 1920 3164 1924 3196
rect 1956 3164 1960 3196
rect 1920 3160 1960 3164
rect 2000 3356 2040 3360
rect 2000 3324 2004 3356
rect 2036 3324 2040 3356
rect 2000 3276 2040 3324
rect 2000 3244 2004 3276
rect 2036 3244 2040 3276
rect 2000 3196 2040 3244
rect 2000 3164 2004 3196
rect 2036 3164 2040 3196
rect 2000 3160 2040 3164
rect 2080 3356 2120 3360
rect 2080 3324 2084 3356
rect 2116 3324 2120 3356
rect 2080 3276 2120 3324
rect 2080 3244 2084 3276
rect 2116 3244 2120 3276
rect 2080 3196 2120 3244
rect 2080 3164 2084 3196
rect 2116 3164 2120 3196
rect 2080 3160 2120 3164
rect 2160 3356 2200 3360
rect 2160 3324 2164 3356
rect 2196 3324 2200 3356
rect 2160 3276 2200 3324
rect 2160 3244 2164 3276
rect 2196 3244 2200 3276
rect 2160 3196 2200 3244
rect 2160 3164 2164 3196
rect 2196 3164 2200 3196
rect 2160 3160 2200 3164
rect 2240 3356 2280 3360
rect 2240 3324 2244 3356
rect 2276 3324 2280 3356
rect 2240 3276 2280 3324
rect 2240 3244 2244 3276
rect 2276 3244 2280 3276
rect 2240 3196 2280 3244
rect 2240 3164 2244 3196
rect 2276 3164 2280 3196
rect 2240 3160 2280 3164
rect 2320 3356 2360 3360
rect 2320 3324 2324 3356
rect 2356 3324 2360 3356
rect 2320 3276 2360 3324
rect 2320 3244 2324 3276
rect 2356 3244 2360 3276
rect 2320 3196 2360 3244
rect 2320 3164 2324 3196
rect 2356 3164 2360 3196
rect 2320 3160 2360 3164
rect 2400 3356 2440 3360
rect 2400 3324 2404 3356
rect 2436 3324 2440 3356
rect 2400 3276 2440 3324
rect 2400 3244 2404 3276
rect 2436 3244 2440 3276
rect 2400 3196 2440 3244
rect 2400 3164 2404 3196
rect 2436 3164 2440 3196
rect 2400 3160 2440 3164
rect 2480 3356 2520 3360
rect 2480 3324 2484 3356
rect 2516 3324 2520 3356
rect 2480 3276 2520 3324
rect 2480 3244 2484 3276
rect 2516 3244 2520 3276
rect 2480 3196 2520 3244
rect 2480 3164 2484 3196
rect 2516 3164 2520 3196
rect 2480 3160 2520 3164
rect 2640 3356 2680 3360
rect 2640 3324 2644 3356
rect 2676 3324 2680 3356
rect 2640 3276 2680 3324
rect 2640 3244 2644 3276
rect 2676 3244 2680 3276
rect 2640 3196 2680 3244
rect 2640 3164 2644 3196
rect 2676 3164 2680 3196
rect 2640 3160 2680 3164
rect 2720 3356 2760 3360
rect 2720 3324 2724 3356
rect 2756 3324 2760 3356
rect 2720 3276 2760 3324
rect 2720 3244 2724 3276
rect 2756 3244 2760 3276
rect 2720 3196 2760 3244
rect 2720 3164 2724 3196
rect 2756 3164 2760 3196
rect 2720 3160 2760 3164
rect 2800 3356 2840 3360
rect 2800 3324 2804 3356
rect 2836 3324 2840 3356
rect 2800 3276 2840 3324
rect 2800 3244 2804 3276
rect 2836 3244 2840 3276
rect 2800 3196 2840 3244
rect 2800 3164 2804 3196
rect 2836 3164 2840 3196
rect 2800 3160 2840 3164
rect 2880 3356 2920 3360
rect 2880 3324 2884 3356
rect 2916 3324 2920 3356
rect 2880 3276 2920 3324
rect 2880 3244 2884 3276
rect 2916 3244 2920 3276
rect 2880 3196 2920 3244
rect 2880 3164 2884 3196
rect 2916 3164 2920 3196
rect 2880 3160 2920 3164
rect 2960 3356 3000 3360
rect 2960 3324 2964 3356
rect 2996 3324 3000 3356
rect 2960 3276 3000 3324
rect 2960 3244 2964 3276
rect 2996 3244 3000 3276
rect 2960 3196 3000 3244
rect 2960 3164 2964 3196
rect 2996 3164 3000 3196
rect 2960 3160 3000 3164
rect 3040 3356 3080 3360
rect 3040 3324 3044 3356
rect 3076 3324 3080 3356
rect 3040 3276 3080 3324
rect 3040 3244 3044 3276
rect 3076 3244 3080 3276
rect 3040 3196 3080 3244
rect 3040 3164 3044 3196
rect 3076 3164 3080 3196
rect 3040 3160 3080 3164
rect 3120 3356 3160 3360
rect 3120 3324 3124 3356
rect 3156 3324 3160 3356
rect 3120 3276 3160 3324
rect 3120 3244 3124 3276
rect 3156 3244 3160 3276
rect 3120 3196 3160 3244
rect 3120 3164 3124 3196
rect 3156 3164 3160 3196
rect 3120 3160 3160 3164
rect 3200 3356 3240 3360
rect 3200 3324 3204 3356
rect 3236 3324 3240 3356
rect 3200 3276 3240 3324
rect 3200 3244 3204 3276
rect 3236 3244 3240 3276
rect 3200 3196 3240 3244
rect 3200 3164 3204 3196
rect 3236 3164 3240 3196
rect 3200 3160 3240 3164
rect 3280 3356 3320 3360
rect 3280 3324 3284 3356
rect 3316 3324 3320 3356
rect 3280 3276 3320 3324
rect 3280 3244 3284 3276
rect 3316 3244 3320 3276
rect 3280 3196 3320 3244
rect 3280 3164 3284 3196
rect 3316 3164 3320 3196
rect 3280 3160 3320 3164
rect 3360 3356 3400 3360
rect 3360 3324 3364 3356
rect 3396 3324 3400 3356
rect 3360 3276 3400 3324
rect 3360 3244 3364 3276
rect 3396 3244 3400 3276
rect 3360 3196 3400 3244
rect 3360 3164 3364 3196
rect 3396 3164 3400 3196
rect 3360 3160 3400 3164
rect 3440 3356 3480 3360
rect 3440 3324 3444 3356
rect 3476 3324 3480 3356
rect 3440 3276 3480 3324
rect 3440 3244 3444 3276
rect 3476 3244 3480 3276
rect 3440 3196 3480 3244
rect 3440 3164 3444 3196
rect 3476 3164 3480 3196
rect 3440 3160 3480 3164
rect 3600 3356 3640 3360
rect 3600 3324 3604 3356
rect 3636 3324 3640 3356
rect 3600 3276 3640 3324
rect 3600 3244 3604 3276
rect 3636 3244 3640 3276
rect 3600 3196 3640 3244
rect 3600 3164 3604 3196
rect 3636 3164 3640 3196
rect 3600 3160 3640 3164
rect 3680 3356 3720 3360
rect 3680 3324 3684 3356
rect 3716 3324 3720 3356
rect 3680 3276 3720 3324
rect 3680 3244 3684 3276
rect 3716 3244 3720 3276
rect 3680 3196 3720 3244
rect 3680 3164 3684 3196
rect 3716 3164 3720 3196
rect 3680 3160 3720 3164
rect 3760 3356 3800 3360
rect 3760 3324 3764 3356
rect 3796 3324 3800 3356
rect 3760 3276 3800 3324
rect 3760 3244 3764 3276
rect 3796 3244 3800 3276
rect 3760 3196 3800 3244
rect 3760 3164 3764 3196
rect 3796 3164 3800 3196
rect 3760 3160 3800 3164
rect 3840 3356 3880 3360
rect 3840 3324 3844 3356
rect 3876 3324 3880 3356
rect 3840 3276 3880 3324
rect 3840 3244 3844 3276
rect 3876 3244 3880 3276
rect 3840 3196 3880 3244
rect 3840 3164 3844 3196
rect 3876 3164 3880 3196
rect 3840 3160 3880 3164
rect 3920 3356 3960 3360
rect 3920 3324 3924 3356
rect 3956 3324 3960 3356
rect 3920 3276 3960 3324
rect 3920 3244 3924 3276
rect 3956 3244 3960 3276
rect 3920 3196 3960 3244
rect 3920 3164 3924 3196
rect 3956 3164 3960 3196
rect 3920 3160 3960 3164
rect 4080 3356 4120 3360
rect 4080 3324 4084 3356
rect 4116 3324 4120 3356
rect 4080 3276 4120 3324
rect 4080 3244 4084 3276
rect 4116 3244 4120 3276
rect 4080 3196 4120 3244
rect 4080 3164 4084 3196
rect 4116 3164 4120 3196
rect 4080 3160 4120 3164
rect 80 3116 120 3120
rect 80 3084 84 3116
rect 116 3084 120 3116
rect 80 3036 120 3084
rect 80 3004 84 3036
rect 116 3004 120 3036
rect 80 2956 120 3004
rect 80 2924 84 2956
rect 116 2924 120 2956
rect 80 2920 120 2924
rect 160 3116 200 3120
rect 160 3084 164 3116
rect 196 3084 200 3116
rect 160 3036 200 3084
rect 160 3004 164 3036
rect 196 3004 200 3036
rect 160 2956 200 3004
rect 160 2924 164 2956
rect 196 2924 200 2956
rect 160 2920 200 2924
rect 240 3116 280 3120
rect 240 3084 244 3116
rect 276 3084 280 3116
rect 240 3036 280 3084
rect 240 3004 244 3036
rect 276 3004 280 3036
rect 240 2956 280 3004
rect 240 2924 244 2956
rect 276 2924 280 2956
rect 240 2920 280 2924
rect 320 3116 360 3120
rect 320 3084 324 3116
rect 356 3084 360 3116
rect 320 3036 360 3084
rect 320 3004 324 3036
rect 356 3004 360 3036
rect 320 2956 360 3004
rect 320 2924 324 2956
rect 356 2924 360 2956
rect 320 2920 360 2924
rect 400 3116 440 3120
rect 400 3084 404 3116
rect 436 3084 440 3116
rect 400 3036 440 3084
rect 400 3004 404 3036
rect 436 3004 440 3036
rect 400 2956 440 3004
rect 400 2924 404 2956
rect 436 2924 440 2956
rect 400 2920 440 2924
rect 480 3116 520 3120
rect 480 3084 484 3116
rect 516 3084 520 3116
rect 480 3036 520 3084
rect 480 3004 484 3036
rect 516 3004 520 3036
rect 480 2956 520 3004
rect 480 2924 484 2956
rect 516 2924 520 2956
rect 480 2920 520 2924
rect 560 3116 600 3120
rect 560 3084 564 3116
rect 596 3084 600 3116
rect 560 3036 600 3084
rect 560 3004 564 3036
rect 596 3004 600 3036
rect 560 2956 600 3004
rect 560 2924 564 2956
rect 596 2924 600 2956
rect 560 2920 600 2924
rect 640 3116 680 3120
rect 640 3084 644 3116
rect 676 3084 680 3116
rect 640 3036 680 3084
rect 640 3004 644 3036
rect 676 3004 680 3036
rect 640 2956 680 3004
rect 640 2924 644 2956
rect 676 2924 680 2956
rect 640 2920 680 2924
rect 720 3116 760 3120
rect 720 3084 724 3116
rect 756 3084 760 3116
rect 720 3036 760 3084
rect 720 3004 724 3036
rect 756 3004 760 3036
rect 720 2956 760 3004
rect 720 2924 724 2956
rect 756 2924 760 2956
rect 720 2920 760 2924
rect 800 3116 840 3120
rect 800 3084 804 3116
rect 836 3084 840 3116
rect 800 3036 840 3084
rect 800 3004 804 3036
rect 836 3004 840 3036
rect 800 2956 840 3004
rect 800 2924 804 2956
rect 836 2924 840 2956
rect 800 2920 840 2924
rect 880 3116 920 3120
rect 880 3084 884 3116
rect 916 3084 920 3116
rect 880 3036 920 3084
rect 880 3004 884 3036
rect 916 3004 920 3036
rect 880 2956 920 3004
rect 880 2924 884 2956
rect 916 2924 920 2956
rect 880 2920 920 2924
rect 960 3116 1000 3120
rect 960 3084 964 3116
rect 996 3084 1000 3116
rect 960 3036 1000 3084
rect 960 3004 964 3036
rect 996 3004 1000 3036
rect 960 2956 1000 3004
rect 960 2924 964 2956
rect 996 2924 1000 2956
rect 960 2920 1000 2924
rect 1040 3116 1080 3120
rect 1040 3084 1044 3116
rect 1076 3084 1080 3116
rect 1040 3036 1080 3084
rect 1040 3004 1044 3036
rect 1076 3004 1080 3036
rect 1040 2956 1080 3004
rect 1040 2924 1044 2956
rect 1076 2924 1080 2956
rect 1040 2920 1080 2924
rect 1120 3116 1160 3120
rect 1120 3084 1124 3116
rect 1156 3084 1160 3116
rect 1120 3036 1160 3084
rect 1120 3004 1124 3036
rect 1156 3004 1160 3036
rect 1120 2956 1160 3004
rect 1120 2924 1124 2956
rect 1156 2924 1160 2956
rect 1120 2920 1160 2924
rect 1200 3116 1240 3120
rect 1200 3084 1204 3116
rect 1236 3084 1240 3116
rect 1200 3036 1240 3084
rect 1200 3004 1204 3036
rect 1236 3004 1240 3036
rect 1200 2956 1240 3004
rect 1200 2924 1204 2956
rect 1236 2924 1240 2956
rect 1200 2920 1240 2924
rect 1280 3116 1320 3120
rect 1280 3084 1284 3116
rect 1316 3084 1320 3116
rect 1280 3036 1320 3084
rect 1280 3004 1284 3036
rect 1316 3004 1320 3036
rect 1280 2956 1320 3004
rect 1280 2924 1284 2956
rect 1316 2924 1320 2956
rect 1280 2920 1320 2924
rect 1360 3116 1400 3120
rect 1360 3084 1364 3116
rect 1396 3084 1400 3116
rect 1360 3036 1400 3084
rect 1360 3004 1364 3036
rect 1396 3004 1400 3036
rect 1360 2956 1400 3004
rect 1360 2924 1364 2956
rect 1396 2924 1400 2956
rect 1360 2920 1400 2924
rect 1440 3116 1480 3120
rect 1440 3084 1444 3116
rect 1476 3084 1480 3116
rect 1440 3036 1480 3084
rect 1440 3004 1444 3036
rect 1476 3004 1480 3036
rect 1440 2956 1480 3004
rect 1440 2924 1444 2956
rect 1476 2924 1480 2956
rect 1440 2920 1480 2924
rect 1520 3116 1560 3120
rect 1520 3084 1524 3116
rect 1556 3084 1560 3116
rect 1520 3036 1560 3084
rect 1520 3004 1524 3036
rect 1556 3004 1560 3036
rect 1520 2956 1560 3004
rect 1520 2924 1524 2956
rect 1556 2924 1560 2956
rect 1520 2920 1560 2924
rect 1600 3116 1640 3120
rect 1600 3084 1604 3116
rect 1636 3084 1640 3116
rect 1600 3036 1640 3084
rect 1600 3004 1604 3036
rect 1636 3004 1640 3036
rect 1600 2956 1640 3004
rect 1600 2924 1604 2956
rect 1636 2924 1640 2956
rect 1600 2920 1640 2924
rect 1680 3116 1720 3120
rect 1680 3084 1684 3116
rect 1716 3084 1720 3116
rect 1680 3036 1720 3084
rect 1680 3004 1684 3036
rect 1716 3004 1720 3036
rect 1680 2956 1720 3004
rect 1680 2924 1684 2956
rect 1716 2924 1720 2956
rect 1680 2920 1720 2924
rect 1760 3116 1800 3120
rect 1760 3084 1764 3116
rect 1796 3084 1800 3116
rect 1760 3036 1800 3084
rect 1760 3004 1764 3036
rect 1796 3004 1800 3036
rect 1760 2956 1800 3004
rect 1760 2924 1764 2956
rect 1796 2924 1800 2956
rect 1760 2920 1800 2924
rect 1840 3116 1880 3120
rect 1840 3084 1844 3116
rect 1876 3084 1880 3116
rect 1840 3036 1880 3084
rect 1840 3004 1844 3036
rect 1876 3004 1880 3036
rect 1840 2956 1880 3004
rect 1840 2924 1844 2956
rect 1876 2924 1880 2956
rect 1840 2920 1880 2924
rect 1920 3116 1960 3120
rect 1920 3084 1924 3116
rect 1956 3084 1960 3116
rect 1920 3036 1960 3084
rect 1920 3004 1924 3036
rect 1956 3004 1960 3036
rect 1920 2956 1960 3004
rect 1920 2924 1924 2956
rect 1956 2924 1960 2956
rect 1920 2920 1960 2924
rect 2000 3116 2040 3120
rect 2000 3084 2004 3116
rect 2036 3084 2040 3116
rect 2000 3036 2040 3084
rect 2000 3004 2004 3036
rect 2036 3004 2040 3036
rect 2000 2956 2040 3004
rect 2000 2924 2004 2956
rect 2036 2924 2040 2956
rect 2000 2920 2040 2924
rect 2080 3116 2120 3120
rect 2080 3084 2084 3116
rect 2116 3084 2120 3116
rect 2080 3036 2120 3084
rect 2080 3004 2084 3036
rect 2116 3004 2120 3036
rect 2080 2956 2120 3004
rect 2080 2924 2084 2956
rect 2116 2924 2120 2956
rect 2080 2920 2120 2924
rect 2160 3116 2200 3120
rect 2160 3084 2164 3116
rect 2196 3084 2200 3116
rect 2160 3036 2200 3084
rect 2160 3004 2164 3036
rect 2196 3004 2200 3036
rect 2160 2956 2200 3004
rect 2160 2924 2164 2956
rect 2196 2924 2200 2956
rect 2160 2920 2200 2924
rect 2240 3116 2280 3120
rect 2240 3084 2244 3116
rect 2276 3084 2280 3116
rect 2240 3036 2280 3084
rect 2240 3004 2244 3036
rect 2276 3004 2280 3036
rect 2240 2956 2280 3004
rect 2240 2924 2244 2956
rect 2276 2924 2280 2956
rect 2240 2920 2280 2924
rect 2320 3116 2360 3120
rect 2320 3084 2324 3116
rect 2356 3084 2360 3116
rect 2320 3036 2360 3084
rect 2320 3004 2324 3036
rect 2356 3004 2360 3036
rect 2320 2956 2360 3004
rect 2320 2924 2324 2956
rect 2356 2924 2360 2956
rect 2320 2920 2360 2924
rect 2400 3116 2440 3120
rect 2400 3084 2404 3116
rect 2436 3084 2440 3116
rect 2400 3036 2440 3084
rect 2400 3004 2404 3036
rect 2436 3004 2440 3036
rect 2400 2956 2440 3004
rect 2400 2924 2404 2956
rect 2436 2924 2440 2956
rect 2400 2920 2440 2924
rect 2480 3116 2520 3120
rect 2480 3084 2484 3116
rect 2516 3084 2520 3116
rect 2480 3036 2520 3084
rect 2480 3004 2484 3036
rect 2516 3004 2520 3036
rect 2480 2956 2520 3004
rect 2480 2924 2484 2956
rect 2516 2924 2520 2956
rect 2480 2920 2520 2924
rect 2560 3116 2600 3120
rect 2560 3084 2564 3116
rect 2596 3084 2600 3116
rect 2560 3036 2600 3084
rect 2560 3004 2564 3036
rect 2596 3004 2600 3036
rect 2560 2956 2600 3004
rect 2560 2924 2564 2956
rect 2596 2924 2600 2956
rect 2560 2920 2600 2924
rect 2640 3116 2680 3120
rect 2640 3084 2644 3116
rect 2676 3084 2680 3116
rect 2640 3036 2680 3084
rect 2640 3004 2644 3036
rect 2676 3004 2680 3036
rect 2640 2956 2680 3004
rect 2640 2924 2644 2956
rect 2676 2924 2680 2956
rect 2640 2920 2680 2924
rect 2720 3116 2760 3120
rect 2720 3084 2724 3116
rect 2756 3084 2760 3116
rect 2720 3036 2760 3084
rect 2720 3004 2724 3036
rect 2756 3004 2760 3036
rect 2720 2956 2760 3004
rect 2720 2924 2724 2956
rect 2756 2924 2760 2956
rect 2720 2920 2760 2924
rect 2800 3116 2840 3120
rect 2800 3084 2804 3116
rect 2836 3084 2840 3116
rect 2800 3036 2840 3084
rect 2800 3004 2804 3036
rect 2836 3004 2840 3036
rect 2800 2956 2840 3004
rect 2800 2924 2804 2956
rect 2836 2924 2840 2956
rect 2800 2920 2840 2924
rect 2880 3116 2920 3120
rect 2880 3084 2884 3116
rect 2916 3084 2920 3116
rect 2880 3036 2920 3084
rect 2880 3004 2884 3036
rect 2916 3004 2920 3036
rect 2880 2956 2920 3004
rect 2880 2924 2884 2956
rect 2916 2924 2920 2956
rect 2880 2920 2920 2924
rect 2960 3116 3000 3120
rect 2960 3084 2964 3116
rect 2996 3084 3000 3116
rect 2960 3036 3000 3084
rect 2960 3004 2964 3036
rect 2996 3004 3000 3036
rect 2960 2956 3000 3004
rect 2960 2924 2964 2956
rect 2996 2924 3000 2956
rect 2960 2920 3000 2924
rect 3040 3116 3080 3120
rect 3040 3084 3044 3116
rect 3076 3084 3080 3116
rect 3040 3036 3080 3084
rect 3040 3004 3044 3036
rect 3076 3004 3080 3036
rect 3040 2956 3080 3004
rect 3040 2924 3044 2956
rect 3076 2924 3080 2956
rect 3040 2920 3080 2924
rect 3120 3116 3160 3120
rect 3120 3084 3124 3116
rect 3156 3084 3160 3116
rect 3120 3036 3160 3084
rect 3120 3004 3124 3036
rect 3156 3004 3160 3036
rect 3120 2956 3160 3004
rect 3120 2924 3124 2956
rect 3156 2924 3160 2956
rect 3120 2920 3160 2924
rect 3200 3116 3240 3120
rect 3200 3084 3204 3116
rect 3236 3084 3240 3116
rect 3200 3036 3240 3084
rect 3200 3004 3204 3036
rect 3236 3004 3240 3036
rect 3200 2956 3240 3004
rect 3200 2924 3204 2956
rect 3236 2924 3240 2956
rect 3200 2920 3240 2924
rect 3280 3116 3320 3120
rect 3280 3084 3284 3116
rect 3316 3084 3320 3116
rect 3280 3036 3320 3084
rect 3280 3004 3284 3036
rect 3316 3004 3320 3036
rect 3280 2956 3320 3004
rect 3280 2924 3284 2956
rect 3316 2924 3320 2956
rect 3280 2920 3320 2924
rect 3360 3116 3400 3120
rect 3360 3084 3364 3116
rect 3396 3084 3400 3116
rect 3360 3036 3400 3084
rect 3360 3004 3364 3036
rect 3396 3004 3400 3036
rect 3360 2956 3400 3004
rect 3360 2924 3364 2956
rect 3396 2924 3400 2956
rect 3360 2920 3400 2924
rect 3440 3116 3480 3120
rect 3440 3084 3444 3116
rect 3476 3084 3480 3116
rect 3440 3036 3480 3084
rect 3440 3004 3444 3036
rect 3476 3004 3480 3036
rect 3440 2956 3480 3004
rect 3440 2924 3444 2956
rect 3476 2924 3480 2956
rect 3440 2920 3480 2924
rect 3520 3116 3560 3120
rect 3520 3084 3524 3116
rect 3556 3084 3560 3116
rect 3520 3036 3560 3084
rect 3520 3004 3524 3036
rect 3556 3004 3560 3036
rect 3520 2956 3560 3004
rect 3520 2924 3524 2956
rect 3556 2924 3560 2956
rect 3520 2920 3560 2924
rect 3600 3116 3640 3120
rect 3600 3084 3604 3116
rect 3636 3084 3640 3116
rect 3600 3036 3640 3084
rect 3600 3004 3604 3036
rect 3636 3004 3640 3036
rect 3600 2956 3640 3004
rect 3600 2924 3604 2956
rect 3636 2924 3640 2956
rect 3600 2920 3640 2924
rect 3680 3116 3720 3120
rect 3680 3084 3684 3116
rect 3716 3084 3720 3116
rect 3680 3036 3720 3084
rect 3680 3004 3684 3036
rect 3716 3004 3720 3036
rect 3680 2956 3720 3004
rect 3680 2924 3684 2956
rect 3716 2924 3720 2956
rect 3680 2920 3720 2924
rect 3760 3116 3800 3120
rect 3760 3084 3764 3116
rect 3796 3084 3800 3116
rect 3760 3036 3800 3084
rect 3760 3004 3764 3036
rect 3796 3004 3800 3036
rect 3760 2956 3800 3004
rect 3760 2924 3764 2956
rect 3796 2924 3800 2956
rect 3760 2920 3800 2924
rect 3840 3116 3880 3120
rect 3840 3084 3844 3116
rect 3876 3084 3880 3116
rect 3840 3036 3880 3084
rect 3840 3004 3844 3036
rect 3876 3004 3880 3036
rect 3840 2956 3880 3004
rect 3840 2924 3844 2956
rect 3876 2924 3880 2956
rect 3840 2920 3880 2924
rect 3920 3116 3960 3120
rect 3920 3084 3924 3116
rect 3956 3084 3960 3116
rect 3920 3036 3960 3084
rect 3920 3004 3924 3036
rect 3956 3004 3960 3036
rect 3920 2956 3960 3004
rect 3920 2924 3924 2956
rect 3956 2924 3960 2956
rect 3920 2920 3960 2924
rect 4080 3116 4120 3120
rect 4080 3084 4084 3116
rect 4116 3084 4120 3116
rect 4080 3036 4120 3084
rect 4080 3004 4084 3036
rect 4116 3004 4120 3036
rect 4080 2956 4120 3004
rect 4080 2924 4084 2956
rect 4116 2924 4120 2956
rect 4080 2920 4120 2924
rect 80 2876 120 2880
rect 80 2844 84 2876
rect 116 2844 120 2876
rect 80 2796 120 2844
rect 80 2764 84 2796
rect 116 2764 120 2796
rect 80 2716 120 2764
rect 80 2684 84 2716
rect 116 2684 120 2716
rect 80 2680 120 2684
rect 160 2876 200 2880
rect 160 2844 164 2876
rect 196 2844 200 2876
rect 160 2796 200 2844
rect 160 2764 164 2796
rect 196 2764 200 2796
rect 160 2716 200 2764
rect 160 2684 164 2716
rect 196 2684 200 2716
rect 160 2680 200 2684
rect 240 2876 280 2880
rect 240 2844 244 2876
rect 276 2844 280 2876
rect 240 2796 280 2844
rect 240 2764 244 2796
rect 276 2764 280 2796
rect 240 2716 280 2764
rect 240 2684 244 2716
rect 276 2684 280 2716
rect 240 2680 280 2684
rect 320 2876 360 2880
rect 320 2844 324 2876
rect 356 2844 360 2876
rect 320 2796 360 2844
rect 320 2764 324 2796
rect 356 2764 360 2796
rect 320 2716 360 2764
rect 320 2684 324 2716
rect 356 2684 360 2716
rect 320 2680 360 2684
rect 400 2876 440 2880
rect 400 2844 404 2876
rect 436 2844 440 2876
rect 400 2796 440 2844
rect 400 2764 404 2796
rect 436 2764 440 2796
rect 400 2716 440 2764
rect 400 2684 404 2716
rect 436 2684 440 2716
rect 400 2680 440 2684
rect 480 2876 520 2880
rect 480 2844 484 2876
rect 516 2844 520 2876
rect 480 2796 520 2844
rect 480 2764 484 2796
rect 516 2764 520 2796
rect 480 2716 520 2764
rect 480 2684 484 2716
rect 516 2684 520 2716
rect 480 2680 520 2684
rect 560 2876 600 2880
rect 560 2844 564 2876
rect 596 2844 600 2876
rect 560 2796 600 2844
rect 560 2764 564 2796
rect 596 2764 600 2796
rect 560 2716 600 2764
rect 560 2684 564 2716
rect 596 2684 600 2716
rect 560 2680 600 2684
rect 720 2876 760 2880
rect 720 2844 724 2876
rect 756 2844 760 2876
rect 720 2796 760 2844
rect 720 2764 724 2796
rect 756 2764 760 2796
rect 720 2716 760 2764
rect 720 2684 724 2716
rect 756 2684 760 2716
rect 720 2680 760 2684
rect 800 2876 840 2880
rect 800 2844 804 2876
rect 836 2844 840 2876
rect 800 2796 840 2844
rect 800 2764 804 2796
rect 836 2764 840 2796
rect 800 2716 840 2764
rect 800 2684 804 2716
rect 836 2684 840 2716
rect 800 2680 840 2684
rect 880 2876 920 2880
rect 880 2844 884 2876
rect 916 2844 920 2876
rect 880 2796 920 2844
rect 880 2764 884 2796
rect 916 2764 920 2796
rect 880 2716 920 2764
rect 880 2684 884 2716
rect 916 2684 920 2716
rect 880 2680 920 2684
rect 960 2876 1000 2880
rect 960 2844 964 2876
rect 996 2844 1000 2876
rect 960 2796 1000 2844
rect 960 2764 964 2796
rect 996 2764 1000 2796
rect 960 2716 1000 2764
rect 960 2684 964 2716
rect 996 2684 1000 2716
rect 960 2680 1000 2684
rect 1040 2876 1080 2880
rect 1040 2844 1044 2876
rect 1076 2844 1080 2876
rect 1040 2796 1080 2844
rect 1040 2764 1044 2796
rect 1076 2764 1080 2796
rect 1040 2716 1080 2764
rect 1040 2684 1044 2716
rect 1076 2684 1080 2716
rect 1040 2680 1080 2684
rect 1120 2876 1160 2880
rect 1120 2844 1124 2876
rect 1156 2844 1160 2876
rect 1120 2796 1160 2844
rect 1120 2764 1124 2796
rect 1156 2764 1160 2796
rect 1120 2716 1160 2764
rect 1120 2684 1124 2716
rect 1156 2684 1160 2716
rect 1120 2680 1160 2684
rect 1200 2876 1240 2880
rect 1200 2844 1204 2876
rect 1236 2844 1240 2876
rect 1200 2796 1240 2844
rect 1200 2764 1204 2796
rect 1236 2764 1240 2796
rect 1200 2716 1240 2764
rect 1200 2684 1204 2716
rect 1236 2684 1240 2716
rect 1200 2680 1240 2684
rect 1280 2876 1320 2880
rect 1280 2844 1284 2876
rect 1316 2844 1320 2876
rect 1280 2796 1320 2844
rect 1280 2764 1284 2796
rect 1316 2764 1320 2796
rect 1280 2716 1320 2764
rect 1280 2684 1284 2716
rect 1316 2684 1320 2716
rect 1280 2680 1320 2684
rect 1360 2876 1400 2880
rect 1360 2844 1364 2876
rect 1396 2844 1400 2876
rect 1360 2796 1400 2844
rect 1360 2764 1364 2796
rect 1396 2764 1400 2796
rect 1360 2716 1400 2764
rect 1360 2684 1364 2716
rect 1396 2684 1400 2716
rect 1360 2680 1400 2684
rect 1440 2876 1480 2880
rect 1440 2844 1444 2876
rect 1476 2844 1480 2876
rect 1440 2796 1480 2844
rect 1440 2764 1444 2796
rect 1476 2764 1480 2796
rect 1440 2716 1480 2764
rect 1440 2684 1444 2716
rect 1476 2684 1480 2716
rect 1440 2680 1480 2684
rect 1520 2876 1560 2880
rect 1520 2844 1524 2876
rect 1556 2844 1560 2876
rect 1520 2796 1560 2844
rect 1520 2764 1524 2796
rect 1556 2764 1560 2796
rect 1520 2716 1560 2764
rect 1520 2684 1524 2716
rect 1556 2684 1560 2716
rect 1520 2680 1560 2684
rect 1680 2876 1720 2880
rect 1680 2844 1684 2876
rect 1716 2844 1720 2876
rect 1680 2796 1720 2844
rect 1680 2764 1684 2796
rect 1716 2764 1720 2796
rect 1680 2716 1720 2764
rect 1680 2684 1684 2716
rect 1716 2684 1720 2716
rect 1680 2680 1720 2684
rect 1760 2876 1800 2880
rect 1760 2844 1764 2876
rect 1796 2844 1800 2876
rect 1760 2796 1800 2844
rect 1760 2764 1764 2796
rect 1796 2764 1800 2796
rect 1760 2716 1800 2764
rect 1760 2684 1764 2716
rect 1796 2684 1800 2716
rect 1760 2680 1800 2684
rect 1840 2876 1880 2880
rect 1840 2844 1844 2876
rect 1876 2844 1880 2876
rect 1840 2796 1880 2844
rect 1840 2764 1844 2796
rect 1876 2764 1880 2796
rect 1840 2716 1880 2764
rect 1840 2684 1844 2716
rect 1876 2684 1880 2716
rect 1840 2680 1880 2684
rect 1920 2876 1960 2880
rect 1920 2844 1924 2876
rect 1956 2844 1960 2876
rect 1920 2796 1960 2844
rect 1920 2764 1924 2796
rect 1956 2764 1960 2796
rect 1920 2716 1960 2764
rect 1920 2684 1924 2716
rect 1956 2684 1960 2716
rect 1920 2680 1960 2684
rect 2000 2876 2040 2880
rect 2000 2844 2004 2876
rect 2036 2844 2040 2876
rect 2000 2796 2040 2844
rect 2000 2764 2004 2796
rect 2036 2764 2040 2796
rect 2000 2716 2040 2764
rect 2000 2684 2004 2716
rect 2036 2684 2040 2716
rect 2000 2680 2040 2684
rect 2080 2876 2120 2880
rect 2080 2844 2084 2876
rect 2116 2844 2120 2876
rect 2080 2796 2120 2844
rect 2080 2764 2084 2796
rect 2116 2764 2120 2796
rect 2080 2716 2120 2764
rect 2080 2684 2084 2716
rect 2116 2684 2120 2716
rect 2080 2680 2120 2684
rect 2160 2876 2200 2880
rect 2160 2844 2164 2876
rect 2196 2844 2200 2876
rect 2160 2796 2200 2844
rect 2160 2764 2164 2796
rect 2196 2764 2200 2796
rect 2160 2716 2200 2764
rect 2160 2684 2164 2716
rect 2196 2684 2200 2716
rect 2160 2680 2200 2684
rect 2240 2876 2280 2880
rect 2240 2844 2244 2876
rect 2276 2844 2280 2876
rect 2240 2796 2280 2844
rect 2240 2764 2244 2796
rect 2276 2764 2280 2796
rect 2240 2716 2280 2764
rect 2240 2684 2244 2716
rect 2276 2684 2280 2716
rect 2240 2680 2280 2684
rect 2320 2876 2360 2880
rect 2320 2844 2324 2876
rect 2356 2844 2360 2876
rect 2320 2796 2360 2844
rect 2320 2764 2324 2796
rect 2356 2764 2360 2796
rect 2320 2716 2360 2764
rect 2320 2684 2324 2716
rect 2356 2684 2360 2716
rect 2320 2680 2360 2684
rect 2400 2876 2440 2880
rect 2400 2844 2404 2876
rect 2436 2844 2440 2876
rect 2400 2796 2440 2844
rect 2400 2764 2404 2796
rect 2436 2764 2440 2796
rect 2400 2716 2440 2764
rect 2400 2684 2404 2716
rect 2436 2684 2440 2716
rect 2400 2680 2440 2684
rect 2480 2876 2520 2880
rect 2480 2844 2484 2876
rect 2516 2844 2520 2876
rect 2480 2796 2520 2844
rect 2480 2764 2484 2796
rect 2516 2764 2520 2796
rect 2480 2716 2520 2764
rect 2480 2684 2484 2716
rect 2516 2684 2520 2716
rect 2480 2680 2520 2684
rect 2640 2876 2680 2880
rect 2640 2844 2644 2876
rect 2676 2844 2680 2876
rect 2640 2796 2680 2844
rect 2640 2764 2644 2796
rect 2676 2764 2680 2796
rect 2640 2716 2680 2764
rect 2640 2684 2644 2716
rect 2676 2684 2680 2716
rect 2640 2680 2680 2684
rect 2720 2876 2760 2880
rect 2720 2844 2724 2876
rect 2756 2844 2760 2876
rect 2720 2796 2760 2844
rect 2720 2764 2724 2796
rect 2756 2764 2760 2796
rect 2720 2716 2760 2764
rect 2720 2684 2724 2716
rect 2756 2684 2760 2716
rect 2720 2680 2760 2684
rect 2800 2876 2840 2880
rect 2800 2844 2804 2876
rect 2836 2844 2840 2876
rect 2800 2796 2840 2844
rect 2800 2764 2804 2796
rect 2836 2764 2840 2796
rect 2800 2716 2840 2764
rect 2800 2684 2804 2716
rect 2836 2684 2840 2716
rect 2800 2680 2840 2684
rect 2880 2876 2920 2880
rect 2880 2844 2884 2876
rect 2916 2844 2920 2876
rect 2880 2796 2920 2844
rect 2880 2764 2884 2796
rect 2916 2764 2920 2796
rect 2880 2716 2920 2764
rect 2880 2684 2884 2716
rect 2916 2684 2920 2716
rect 2880 2680 2920 2684
rect 2960 2876 3000 2880
rect 2960 2844 2964 2876
rect 2996 2844 3000 2876
rect 2960 2796 3000 2844
rect 2960 2764 2964 2796
rect 2996 2764 3000 2796
rect 2960 2716 3000 2764
rect 2960 2684 2964 2716
rect 2996 2684 3000 2716
rect 2960 2680 3000 2684
rect 3040 2876 3080 2880
rect 3040 2844 3044 2876
rect 3076 2844 3080 2876
rect 3040 2796 3080 2844
rect 3040 2764 3044 2796
rect 3076 2764 3080 2796
rect 3040 2716 3080 2764
rect 3040 2684 3044 2716
rect 3076 2684 3080 2716
rect 3040 2680 3080 2684
rect 3120 2876 3160 2880
rect 3120 2844 3124 2876
rect 3156 2844 3160 2876
rect 3120 2796 3160 2844
rect 3120 2764 3124 2796
rect 3156 2764 3160 2796
rect 3120 2716 3160 2764
rect 3120 2684 3124 2716
rect 3156 2684 3160 2716
rect 3120 2680 3160 2684
rect 3200 2876 3240 2880
rect 3200 2844 3204 2876
rect 3236 2844 3240 2876
rect 3200 2796 3240 2844
rect 3200 2764 3204 2796
rect 3236 2764 3240 2796
rect 3200 2716 3240 2764
rect 3200 2684 3204 2716
rect 3236 2684 3240 2716
rect 3200 2680 3240 2684
rect 3280 2876 3320 2880
rect 3280 2844 3284 2876
rect 3316 2844 3320 2876
rect 3280 2796 3320 2844
rect 3280 2764 3284 2796
rect 3316 2764 3320 2796
rect 3280 2716 3320 2764
rect 3280 2684 3284 2716
rect 3316 2684 3320 2716
rect 3280 2680 3320 2684
rect 3360 2876 3400 2880
rect 3360 2844 3364 2876
rect 3396 2844 3400 2876
rect 3360 2796 3400 2844
rect 3360 2764 3364 2796
rect 3396 2764 3400 2796
rect 3360 2716 3400 2764
rect 3360 2684 3364 2716
rect 3396 2684 3400 2716
rect 3360 2680 3400 2684
rect 3440 2876 3480 2880
rect 3440 2844 3444 2876
rect 3476 2844 3480 2876
rect 3440 2796 3480 2844
rect 3440 2764 3444 2796
rect 3476 2764 3480 2796
rect 3440 2716 3480 2764
rect 3440 2684 3444 2716
rect 3476 2684 3480 2716
rect 3440 2680 3480 2684
rect 3600 2876 3640 2880
rect 3600 2844 3604 2876
rect 3636 2844 3640 2876
rect 3600 2796 3640 2844
rect 3600 2764 3604 2796
rect 3636 2764 3640 2796
rect 3600 2716 3640 2764
rect 3600 2684 3604 2716
rect 3636 2684 3640 2716
rect 3600 2680 3640 2684
rect 3680 2876 3720 2880
rect 3680 2844 3684 2876
rect 3716 2844 3720 2876
rect 3680 2796 3720 2844
rect 3680 2764 3684 2796
rect 3716 2764 3720 2796
rect 3680 2716 3720 2764
rect 3680 2684 3684 2716
rect 3716 2684 3720 2716
rect 3680 2680 3720 2684
rect 3760 2876 3800 2880
rect 3760 2844 3764 2876
rect 3796 2844 3800 2876
rect 3760 2796 3800 2844
rect 3760 2764 3764 2796
rect 3796 2764 3800 2796
rect 3760 2716 3800 2764
rect 3760 2684 3764 2716
rect 3796 2684 3800 2716
rect 3760 2680 3800 2684
rect 3840 2876 3880 2880
rect 3840 2844 3844 2876
rect 3876 2844 3880 2876
rect 3840 2796 3880 2844
rect 3840 2764 3844 2796
rect 3876 2764 3880 2796
rect 3840 2716 3880 2764
rect 3840 2684 3844 2716
rect 3876 2684 3880 2716
rect 3840 2680 3880 2684
rect 3920 2876 3960 2880
rect 3920 2844 3924 2876
rect 3956 2844 3960 2876
rect 3920 2796 3960 2844
rect 3920 2764 3924 2796
rect 3956 2764 3960 2796
rect 3920 2716 3960 2764
rect 3920 2684 3924 2716
rect 3956 2684 3960 2716
rect 3920 2680 3960 2684
rect 4080 2876 4120 2880
rect 4080 2844 4084 2876
rect 4116 2844 4120 2876
rect 4080 2796 4120 2844
rect 4080 2764 4084 2796
rect 4116 2764 4120 2796
rect 4080 2716 4120 2764
rect 4080 2684 4084 2716
rect 4116 2684 4120 2716
rect 4080 2680 4120 2684
rect 160 2391 200 2400
rect 160 2209 164 2391
rect 196 2209 200 2391
rect 160 2200 200 2209
rect 4000 1831 4040 1840
rect 4000 1649 4004 1831
rect 4036 1649 4040 1831
rect 4000 1640 4040 1649
rect 0 1396 40 1400
rect 0 1364 4 1396
rect 36 1364 40 1396
rect 0 1236 40 1364
rect 0 1204 4 1236
rect 36 1204 40 1236
rect 0 1200 40 1204
rect 80 1396 120 1400
rect 80 1364 84 1396
rect 116 1364 120 1396
rect 80 1236 120 1364
rect 80 1204 84 1236
rect 116 1204 120 1236
rect 80 1200 120 1204
rect 160 1396 200 1400
rect 160 1364 164 1396
rect 196 1364 200 1396
rect 160 1236 200 1364
rect 160 1204 164 1236
rect 196 1204 200 1236
rect 160 1200 200 1204
rect 240 1396 280 1400
rect 240 1364 244 1396
rect 276 1364 280 1396
rect 240 1236 280 1364
rect 240 1204 244 1236
rect 276 1204 280 1236
rect 240 1200 280 1204
rect 320 1396 360 1400
rect 320 1364 324 1396
rect 356 1364 360 1396
rect 320 1236 360 1364
rect 320 1204 324 1236
rect 356 1204 360 1236
rect 320 1200 360 1204
rect 400 1396 440 1400
rect 400 1364 404 1396
rect 436 1364 440 1396
rect 400 1236 440 1364
rect 400 1204 404 1236
rect 436 1204 440 1236
rect 400 1200 440 1204
rect 480 1396 520 1400
rect 480 1364 484 1396
rect 516 1364 520 1396
rect 480 1236 520 1364
rect 480 1204 484 1236
rect 516 1204 520 1236
rect 480 1200 520 1204
rect 560 1396 600 1400
rect 560 1364 564 1396
rect 596 1364 600 1396
rect 560 1236 600 1364
rect 560 1204 564 1236
rect 596 1204 600 1236
rect 560 1200 600 1204
rect 720 1396 760 1400
rect 720 1364 724 1396
rect 756 1364 760 1396
rect 720 1236 760 1364
rect 720 1204 724 1236
rect 756 1204 760 1236
rect 720 1200 760 1204
rect 800 1396 840 1400
rect 800 1364 804 1396
rect 836 1364 840 1396
rect 800 1236 840 1364
rect 800 1204 804 1236
rect 836 1204 840 1236
rect 800 1200 840 1204
rect 880 1396 920 1400
rect 880 1364 884 1396
rect 916 1364 920 1396
rect 880 1236 920 1364
rect 880 1204 884 1236
rect 916 1204 920 1236
rect 880 1200 920 1204
rect 960 1396 1000 1400
rect 960 1364 964 1396
rect 996 1364 1000 1396
rect 960 1236 1000 1364
rect 960 1204 964 1236
rect 996 1204 1000 1236
rect 960 1200 1000 1204
rect 1040 1396 1080 1400
rect 1040 1364 1044 1396
rect 1076 1364 1080 1396
rect 1040 1236 1080 1364
rect 1040 1204 1044 1236
rect 1076 1204 1080 1236
rect 1040 1200 1080 1204
rect 1120 1396 1160 1400
rect 1120 1364 1124 1396
rect 1156 1364 1160 1396
rect 1120 1236 1160 1364
rect 1120 1204 1124 1236
rect 1156 1204 1160 1236
rect 1120 1200 1160 1204
rect 1200 1396 1240 1400
rect 1200 1364 1204 1396
rect 1236 1364 1240 1396
rect 1200 1236 1240 1364
rect 1200 1204 1204 1236
rect 1236 1204 1240 1236
rect 1200 1200 1240 1204
rect 1280 1396 1320 1400
rect 1280 1364 1284 1396
rect 1316 1364 1320 1396
rect 1280 1236 1320 1364
rect 1280 1204 1284 1236
rect 1316 1204 1320 1236
rect 1280 1200 1320 1204
rect 1360 1396 1400 1400
rect 1360 1364 1364 1396
rect 1396 1364 1400 1396
rect 1360 1236 1400 1364
rect 1360 1204 1364 1236
rect 1396 1204 1400 1236
rect 1360 1200 1400 1204
rect 1440 1396 1480 1400
rect 1440 1364 1444 1396
rect 1476 1364 1480 1396
rect 1440 1236 1480 1364
rect 1440 1204 1444 1236
rect 1476 1204 1480 1236
rect 1440 1200 1480 1204
rect 1520 1396 1560 1400
rect 1520 1364 1524 1396
rect 1556 1364 1560 1396
rect 1520 1236 1560 1364
rect 1520 1204 1524 1236
rect 1556 1204 1560 1236
rect 1520 1200 1560 1204
rect 1680 1396 1720 1400
rect 1680 1364 1684 1396
rect 1716 1364 1720 1396
rect 1680 1236 1720 1364
rect 1680 1204 1684 1236
rect 1716 1204 1720 1236
rect 1680 1200 1720 1204
rect 1760 1396 1800 1400
rect 1760 1364 1764 1396
rect 1796 1364 1800 1396
rect 1760 1236 1800 1364
rect 1760 1204 1764 1236
rect 1796 1204 1800 1236
rect 1760 1200 1800 1204
rect 1840 1396 1880 1400
rect 1840 1364 1844 1396
rect 1876 1364 1880 1396
rect 1840 1236 1880 1364
rect 1840 1204 1844 1236
rect 1876 1204 1880 1236
rect 1840 1200 1880 1204
rect 1920 1396 1960 1400
rect 1920 1364 1924 1396
rect 1956 1364 1960 1396
rect 1920 1236 1960 1364
rect 1920 1204 1924 1236
rect 1956 1204 1960 1236
rect 1920 1200 1960 1204
rect 2000 1396 2040 1400
rect 2000 1364 2004 1396
rect 2036 1364 2040 1396
rect 2000 1236 2040 1364
rect 2000 1204 2004 1236
rect 2036 1204 2040 1236
rect 2000 1200 2040 1204
rect 2080 1396 2120 1400
rect 2080 1364 2084 1396
rect 2116 1364 2120 1396
rect 2080 1236 2120 1364
rect 2080 1204 2084 1236
rect 2116 1204 2120 1236
rect 2080 1200 2120 1204
rect 2160 1396 2200 1400
rect 2160 1364 2164 1396
rect 2196 1364 2200 1396
rect 2160 1236 2200 1364
rect 2160 1204 2164 1236
rect 2196 1204 2200 1236
rect 2160 1200 2200 1204
rect 2240 1396 2280 1400
rect 2240 1364 2244 1396
rect 2276 1364 2280 1396
rect 2240 1236 2280 1364
rect 2240 1204 2244 1236
rect 2276 1204 2280 1236
rect 2240 1200 2280 1204
rect 2320 1396 2360 1400
rect 2320 1364 2324 1396
rect 2356 1364 2360 1396
rect 2320 1236 2360 1364
rect 2320 1204 2324 1236
rect 2356 1204 2360 1236
rect 2320 1200 2360 1204
rect 2400 1396 2440 1400
rect 2400 1364 2404 1396
rect 2436 1364 2440 1396
rect 2400 1236 2440 1364
rect 2400 1204 2404 1236
rect 2436 1204 2440 1236
rect 2400 1200 2440 1204
rect 2480 1396 2520 1400
rect 2480 1364 2484 1396
rect 2516 1364 2520 1396
rect 2480 1236 2520 1364
rect 2480 1204 2484 1236
rect 2516 1204 2520 1236
rect 2480 1200 2520 1204
rect 2640 1396 2680 1400
rect 2640 1364 2644 1396
rect 2676 1364 2680 1396
rect 2640 1236 2680 1364
rect 2640 1204 2644 1236
rect 2676 1204 2680 1236
rect 2640 1200 2680 1204
rect 2720 1396 2760 1400
rect 2720 1364 2724 1396
rect 2756 1364 2760 1396
rect 2720 1236 2760 1364
rect 2720 1204 2724 1236
rect 2756 1204 2760 1236
rect 2720 1200 2760 1204
rect 2800 1396 2840 1400
rect 2800 1364 2804 1396
rect 2836 1364 2840 1396
rect 2800 1236 2840 1364
rect 2800 1204 2804 1236
rect 2836 1204 2840 1236
rect 2800 1200 2840 1204
rect 2880 1396 2920 1400
rect 2880 1364 2884 1396
rect 2916 1364 2920 1396
rect 2880 1236 2920 1364
rect 2880 1204 2884 1236
rect 2916 1204 2920 1236
rect 2880 1200 2920 1204
rect 2960 1396 3000 1400
rect 2960 1364 2964 1396
rect 2996 1364 3000 1396
rect 2960 1236 3000 1364
rect 2960 1204 2964 1236
rect 2996 1204 3000 1236
rect 2960 1200 3000 1204
rect 3040 1396 3080 1400
rect 3040 1364 3044 1396
rect 3076 1364 3080 1396
rect 3040 1236 3080 1364
rect 3040 1204 3044 1236
rect 3076 1204 3080 1236
rect 3040 1200 3080 1204
rect 3120 1396 3160 1400
rect 3120 1364 3124 1396
rect 3156 1364 3160 1396
rect 3120 1236 3160 1364
rect 3120 1204 3124 1236
rect 3156 1204 3160 1236
rect 3120 1200 3160 1204
rect 3200 1396 3240 1400
rect 3200 1364 3204 1396
rect 3236 1364 3240 1396
rect 3200 1236 3240 1364
rect 3200 1204 3204 1236
rect 3236 1204 3240 1236
rect 3200 1200 3240 1204
rect 3280 1396 3320 1400
rect 3280 1364 3284 1396
rect 3316 1364 3320 1396
rect 3280 1236 3320 1364
rect 3280 1204 3284 1236
rect 3316 1204 3320 1236
rect 3280 1200 3320 1204
rect 3360 1396 3400 1400
rect 3360 1364 3364 1396
rect 3396 1364 3400 1396
rect 3360 1236 3400 1364
rect 3360 1204 3364 1236
rect 3396 1204 3400 1236
rect 3360 1200 3400 1204
rect 3440 1396 3480 1400
rect 3440 1364 3444 1396
rect 3476 1364 3480 1396
rect 3440 1236 3480 1364
rect 3440 1204 3444 1236
rect 3476 1204 3480 1236
rect 3440 1200 3480 1204
rect 3600 1396 3640 1400
rect 3600 1364 3604 1396
rect 3636 1364 3640 1396
rect 3600 1236 3640 1364
rect 3600 1204 3604 1236
rect 3636 1204 3640 1236
rect 3600 1200 3640 1204
rect 3680 1396 3720 1400
rect 3680 1364 3684 1396
rect 3716 1364 3720 1396
rect 3680 1236 3720 1364
rect 3680 1204 3684 1236
rect 3716 1204 3720 1236
rect 3680 1200 3720 1204
rect 3760 1396 3800 1400
rect 3760 1364 3764 1396
rect 3796 1364 3800 1396
rect 3760 1236 3800 1364
rect 3760 1204 3764 1236
rect 3796 1204 3800 1236
rect 3760 1200 3800 1204
rect 3840 1396 3880 1400
rect 3840 1364 3844 1396
rect 3876 1364 3880 1396
rect 3840 1236 3880 1364
rect 3840 1204 3844 1236
rect 3876 1204 3880 1236
rect 3840 1200 3880 1204
rect 3920 1396 3960 1400
rect 3920 1364 3924 1396
rect 3956 1364 3960 1396
rect 3920 1236 3960 1364
rect 3920 1204 3924 1236
rect 3956 1204 3960 1236
rect 3920 1200 3960 1204
rect 4000 1396 4040 1400
rect 4000 1364 4004 1396
rect 4036 1364 4040 1396
rect 4000 1236 4040 1364
rect 4000 1204 4004 1236
rect 4036 1204 4040 1236
rect 4000 1200 4040 1204
rect 4080 1396 4120 1400
rect 4080 1364 4084 1396
rect 4116 1364 4120 1396
rect 4080 1236 4120 1364
rect 4080 1204 4084 1236
rect 4116 1204 4120 1236
rect 4080 1200 4120 1204
rect 4160 1396 4200 1400
rect 4160 1364 4164 1396
rect 4196 1364 4200 1396
rect 4160 1236 4200 1364
rect 4160 1204 4164 1236
rect 4196 1204 4200 1236
rect 4160 1200 4200 1204
rect 80 635 120 640
rect 80 605 85 635
rect 115 605 120 635
rect 80 556 120 605
rect 80 524 84 556
rect 116 524 120 556
rect 80 476 120 524
rect 80 444 84 476
rect 116 444 120 476
rect 80 396 120 444
rect 80 364 84 396
rect 116 364 120 396
rect 80 315 120 364
rect 80 285 85 315
rect 115 285 120 315
rect 80 280 120 285
rect 160 635 200 640
rect 160 605 165 635
rect 195 605 200 635
rect 160 556 200 605
rect 160 524 164 556
rect 196 524 200 556
rect 160 476 200 524
rect 160 444 164 476
rect 196 444 200 476
rect 160 396 200 444
rect 160 364 164 396
rect 196 364 200 396
rect 160 315 200 364
rect 160 285 165 315
rect 195 285 200 315
rect 160 280 200 285
rect 240 635 280 640
rect 240 605 245 635
rect 275 605 280 635
rect 240 556 280 605
rect 240 524 244 556
rect 276 524 280 556
rect 240 476 280 524
rect 240 444 244 476
rect 276 444 280 476
rect 240 396 280 444
rect 240 364 244 396
rect 276 364 280 396
rect 240 315 280 364
rect 240 285 245 315
rect 275 285 280 315
rect 240 280 280 285
rect 320 635 360 640
rect 320 605 325 635
rect 355 605 360 635
rect 320 556 360 605
rect 320 524 324 556
rect 356 524 360 556
rect 320 476 360 524
rect 320 444 324 476
rect 356 444 360 476
rect 320 396 360 444
rect 320 364 324 396
rect 356 364 360 396
rect 320 315 360 364
rect 320 285 325 315
rect 355 285 360 315
rect 320 280 360 285
rect 400 635 440 640
rect 400 605 405 635
rect 435 605 440 635
rect 400 556 440 605
rect 400 524 404 556
rect 436 524 440 556
rect 400 476 440 524
rect 400 444 404 476
rect 436 444 440 476
rect 400 396 440 444
rect 400 364 404 396
rect 436 364 440 396
rect 400 315 440 364
rect 400 285 405 315
rect 435 285 440 315
rect 400 280 440 285
rect 480 635 520 640
rect 480 605 485 635
rect 515 605 520 635
rect 480 556 520 605
rect 480 524 484 556
rect 516 524 520 556
rect 480 476 520 524
rect 480 444 484 476
rect 516 444 520 476
rect 480 396 520 444
rect 480 364 484 396
rect 516 364 520 396
rect 480 315 520 364
rect 480 285 485 315
rect 515 285 520 315
rect 480 280 520 285
rect 560 635 600 640
rect 560 605 565 635
rect 595 605 600 635
rect 560 556 600 605
rect 560 524 564 556
rect 596 524 600 556
rect 560 476 600 524
rect 560 444 564 476
rect 596 444 600 476
rect 560 396 600 444
rect 560 364 564 396
rect 596 364 600 396
rect 560 315 600 364
rect 560 285 565 315
rect 595 285 600 315
rect 560 280 600 285
rect 720 635 760 640
rect 720 605 725 635
rect 755 605 760 635
rect 720 556 760 605
rect 720 524 724 556
rect 756 524 760 556
rect 720 476 760 524
rect 720 444 724 476
rect 756 444 760 476
rect 720 396 760 444
rect 720 364 724 396
rect 756 364 760 396
rect 720 315 760 364
rect 720 285 725 315
rect 755 285 760 315
rect 720 280 760 285
rect 800 635 840 640
rect 800 605 805 635
rect 835 605 840 635
rect 800 556 840 605
rect 800 524 804 556
rect 836 524 840 556
rect 800 476 840 524
rect 800 444 804 476
rect 836 444 840 476
rect 800 396 840 444
rect 800 364 804 396
rect 836 364 840 396
rect 800 315 840 364
rect 800 285 805 315
rect 835 285 840 315
rect 800 280 840 285
rect 880 635 920 640
rect 880 605 885 635
rect 915 605 920 635
rect 880 556 920 605
rect 880 524 884 556
rect 916 524 920 556
rect 880 476 920 524
rect 880 444 884 476
rect 916 444 920 476
rect 880 396 920 444
rect 880 364 884 396
rect 916 364 920 396
rect 880 315 920 364
rect 880 285 885 315
rect 915 285 920 315
rect 880 280 920 285
rect 960 635 1000 640
rect 960 605 965 635
rect 995 605 1000 635
rect 960 556 1000 605
rect 960 524 964 556
rect 996 524 1000 556
rect 960 476 1000 524
rect 960 444 964 476
rect 996 444 1000 476
rect 960 396 1000 444
rect 960 364 964 396
rect 996 364 1000 396
rect 960 315 1000 364
rect 960 285 965 315
rect 995 285 1000 315
rect 960 280 1000 285
rect 1040 635 1080 640
rect 1040 605 1045 635
rect 1075 605 1080 635
rect 1040 556 1080 605
rect 1040 524 1044 556
rect 1076 524 1080 556
rect 1040 476 1080 524
rect 1040 444 1044 476
rect 1076 444 1080 476
rect 1040 396 1080 444
rect 1040 364 1044 396
rect 1076 364 1080 396
rect 1040 315 1080 364
rect 1040 285 1045 315
rect 1075 285 1080 315
rect 1040 280 1080 285
rect 1120 635 1160 640
rect 1120 605 1125 635
rect 1155 605 1160 635
rect 1120 556 1160 605
rect 1120 524 1124 556
rect 1156 524 1160 556
rect 1120 476 1160 524
rect 1120 444 1124 476
rect 1156 444 1160 476
rect 1120 396 1160 444
rect 1120 364 1124 396
rect 1156 364 1160 396
rect 1120 315 1160 364
rect 1120 285 1125 315
rect 1155 285 1160 315
rect 1120 280 1160 285
rect 1200 635 1240 640
rect 1200 605 1205 635
rect 1235 605 1240 635
rect 1200 556 1240 605
rect 1200 524 1204 556
rect 1236 524 1240 556
rect 1200 476 1240 524
rect 1200 444 1204 476
rect 1236 444 1240 476
rect 1200 396 1240 444
rect 1200 364 1204 396
rect 1236 364 1240 396
rect 1200 315 1240 364
rect 1200 285 1205 315
rect 1235 285 1240 315
rect 1200 280 1240 285
rect 1280 635 1320 640
rect 1280 605 1285 635
rect 1315 605 1320 635
rect 1280 556 1320 605
rect 1280 524 1284 556
rect 1316 524 1320 556
rect 1280 476 1320 524
rect 1280 444 1284 476
rect 1316 444 1320 476
rect 1280 396 1320 444
rect 1280 364 1284 396
rect 1316 364 1320 396
rect 1280 315 1320 364
rect 1280 285 1285 315
rect 1315 285 1320 315
rect 1280 280 1320 285
rect 1360 635 1400 640
rect 1360 605 1365 635
rect 1395 605 1400 635
rect 1360 556 1400 605
rect 1360 524 1364 556
rect 1396 524 1400 556
rect 1360 476 1400 524
rect 1360 444 1364 476
rect 1396 444 1400 476
rect 1360 396 1400 444
rect 1360 364 1364 396
rect 1396 364 1400 396
rect 1360 315 1400 364
rect 1360 285 1365 315
rect 1395 285 1400 315
rect 1360 280 1400 285
rect 1440 635 1480 640
rect 1440 605 1445 635
rect 1475 605 1480 635
rect 1440 556 1480 605
rect 1440 524 1444 556
rect 1476 524 1480 556
rect 1440 476 1480 524
rect 1440 444 1444 476
rect 1476 444 1480 476
rect 1440 396 1480 444
rect 1440 364 1444 396
rect 1476 364 1480 396
rect 1440 315 1480 364
rect 1440 285 1445 315
rect 1475 285 1480 315
rect 1440 280 1480 285
rect 1520 635 1560 640
rect 1520 605 1525 635
rect 1555 605 1560 635
rect 1520 556 1560 605
rect 1520 524 1524 556
rect 1556 524 1560 556
rect 1520 476 1560 524
rect 1520 444 1524 476
rect 1556 444 1560 476
rect 1520 396 1560 444
rect 1520 364 1524 396
rect 1556 364 1560 396
rect 1520 315 1560 364
rect 1520 285 1525 315
rect 1555 285 1560 315
rect 1520 280 1560 285
rect 1680 635 1720 640
rect 1680 605 1685 635
rect 1715 605 1720 635
rect 1680 556 1720 605
rect 1680 524 1684 556
rect 1716 524 1720 556
rect 1680 476 1720 524
rect 1680 444 1684 476
rect 1716 444 1720 476
rect 1680 396 1720 444
rect 1680 364 1684 396
rect 1716 364 1720 396
rect 1680 315 1720 364
rect 1680 285 1685 315
rect 1715 285 1720 315
rect 1680 280 1720 285
rect 1760 635 1800 640
rect 1760 605 1765 635
rect 1795 605 1800 635
rect 1760 556 1800 605
rect 1760 524 1764 556
rect 1796 524 1800 556
rect 1760 476 1800 524
rect 1760 444 1764 476
rect 1796 444 1800 476
rect 1760 396 1800 444
rect 1760 364 1764 396
rect 1796 364 1800 396
rect 1760 315 1800 364
rect 1760 285 1765 315
rect 1795 285 1800 315
rect 1760 280 1800 285
rect 1840 635 1880 640
rect 1840 605 1845 635
rect 1875 605 1880 635
rect 1840 556 1880 605
rect 1840 524 1844 556
rect 1876 524 1880 556
rect 1840 476 1880 524
rect 1840 444 1844 476
rect 1876 444 1880 476
rect 1840 396 1880 444
rect 1840 364 1844 396
rect 1876 364 1880 396
rect 1840 315 1880 364
rect 1840 285 1845 315
rect 1875 285 1880 315
rect 1840 280 1880 285
rect 1920 635 1960 640
rect 1920 605 1925 635
rect 1955 605 1960 635
rect 1920 556 1960 605
rect 1920 524 1924 556
rect 1956 524 1960 556
rect 1920 476 1960 524
rect 1920 444 1924 476
rect 1956 444 1960 476
rect 1920 396 1960 444
rect 1920 364 1924 396
rect 1956 364 1960 396
rect 1920 315 1960 364
rect 1920 285 1925 315
rect 1955 285 1960 315
rect 1920 280 1960 285
rect 2000 635 2040 640
rect 2000 605 2005 635
rect 2035 605 2040 635
rect 2000 556 2040 605
rect 2000 524 2004 556
rect 2036 524 2040 556
rect 2000 476 2040 524
rect 2000 444 2004 476
rect 2036 444 2040 476
rect 2000 396 2040 444
rect 2000 364 2004 396
rect 2036 364 2040 396
rect 2000 315 2040 364
rect 2000 285 2005 315
rect 2035 285 2040 315
rect 2000 280 2040 285
rect 2080 635 2120 640
rect 2080 605 2085 635
rect 2115 605 2120 635
rect 2080 556 2120 605
rect 2080 524 2084 556
rect 2116 524 2120 556
rect 2080 476 2120 524
rect 2080 444 2084 476
rect 2116 444 2120 476
rect 2080 396 2120 444
rect 2080 364 2084 396
rect 2116 364 2120 396
rect 2080 315 2120 364
rect 2080 285 2085 315
rect 2115 285 2120 315
rect 2080 280 2120 285
rect 2160 635 2200 640
rect 2160 605 2165 635
rect 2195 605 2200 635
rect 2160 556 2200 605
rect 2160 524 2164 556
rect 2196 524 2200 556
rect 2160 476 2200 524
rect 2160 444 2164 476
rect 2196 444 2200 476
rect 2160 396 2200 444
rect 2160 364 2164 396
rect 2196 364 2200 396
rect 2160 315 2200 364
rect 2160 285 2165 315
rect 2195 285 2200 315
rect 2160 280 2200 285
rect 2240 635 2280 640
rect 2240 605 2245 635
rect 2275 605 2280 635
rect 2240 556 2280 605
rect 2240 524 2244 556
rect 2276 524 2280 556
rect 2240 476 2280 524
rect 2240 444 2244 476
rect 2276 444 2280 476
rect 2240 396 2280 444
rect 2240 364 2244 396
rect 2276 364 2280 396
rect 2240 315 2280 364
rect 2240 285 2245 315
rect 2275 285 2280 315
rect 2240 280 2280 285
rect 2320 635 2360 640
rect 2320 605 2325 635
rect 2355 605 2360 635
rect 2320 556 2360 605
rect 2320 524 2324 556
rect 2356 524 2360 556
rect 2320 476 2360 524
rect 2320 444 2324 476
rect 2356 444 2360 476
rect 2320 396 2360 444
rect 2320 364 2324 396
rect 2356 364 2360 396
rect 2320 315 2360 364
rect 2320 285 2325 315
rect 2355 285 2360 315
rect 2320 280 2360 285
rect 2400 635 2440 640
rect 2400 605 2405 635
rect 2435 605 2440 635
rect 2400 556 2440 605
rect 2400 524 2404 556
rect 2436 524 2440 556
rect 2400 476 2440 524
rect 2400 444 2404 476
rect 2436 444 2440 476
rect 2400 396 2440 444
rect 2400 364 2404 396
rect 2436 364 2440 396
rect 2400 315 2440 364
rect 2400 285 2405 315
rect 2435 285 2440 315
rect 2400 280 2440 285
rect 2480 635 2520 640
rect 2480 605 2485 635
rect 2515 605 2520 635
rect 2480 556 2520 605
rect 2480 524 2484 556
rect 2516 524 2520 556
rect 2480 476 2520 524
rect 2480 444 2484 476
rect 2516 444 2520 476
rect 2480 396 2520 444
rect 2480 364 2484 396
rect 2516 364 2520 396
rect 2480 315 2520 364
rect 2480 285 2485 315
rect 2515 285 2520 315
rect 2480 280 2520 285
rect 2640 635 2680 640
rect 2640 605 2645 635
rect 2675 605 2680 635
rect 2640 556 2680 605
rect 2640 524 2644 556
rect 2676 524 2680 556
rect 2640 476 2680 524
rect 2640 444 2644 476
rect 2676 444 2680 476
rect 2640 396 2680 444
rect 2640 364 2644 396
rect 2676 364 2680 396
rect 2640 315 2680 364
rect 2640 285 2645 315
rect 2675 285 2680 315
rect 2640 280 2680 285
rect 2720 635 2760 640
rect 2720 605 2725 635
rect 2755 605 2760 635
rect 2720 556 2760 605
rect 2720 524 2724 556
rect 2756 524 2760 556
rect 2720 476 2760 524
rect 2720 444 2724 476
rect 2756 444 2760 476
rect 2720 396 2760 444
rect 2720 364 2724 396
rect 2756 364 2760 396
rect 2720 315 2760 364
rect 2720 285 2725 315
rect 2755 285 2760 315
rect 2720 280 2760 285
rect 2800 635 2840 640
rect 2800 605 2805 635
rect 2835 605 2840 635
rect 2800 556 2840 605
rect 2800 524 2804 556
rect 2836 524 2840 556
rect 2800 476 2840 524
rect 2800 444 2804 476
rect 2836 444 2840 476
rect 2800 396 2840 444
rect 2800 364 2804 396
rect 2836 364 2840 396
rect 2800 315 2840 364
rect 2800 285 2805 315
rect 2835 285 2840 315
rect 2800 280 2840 285
rect 2880 635 2920 640
rect 2880 605 2885 635
rect 2915 605 2920 635
rect 2880 556 2920 605
rect 2880 524 2884 556
rect 2916 524 2920 556
rect 2880 476 2920 524
rect 2880 444 2884 476
rect 2916 444 2920 476
rect 2880 396 2920 444
rect 2880 364 2884 396
rect 2916 364 2920 396
rect 2880 315 2920 364
rect 2880 285 2885 315
rect 2915 285 2920 315
rect 2880 280 2920 285
rect 2960 635 3000 640
rect 2960 605 2965 635
rect 2995 605 3000 635
rect 2960 556 3000 605
rect 2960 524 2964 556
rect 2996 524 3000 556
rect 2960 476 3000 524
rect 2960 444 2964 476
rect 2996 444 3000 476
rect 2960 396 3000 444
rect 2960 364 2964 396
rect 2996 364 3000 396
rect 2960 315 3000 364
rect 2960 285 2965 315
rect 2995 285 3000 315
rect 2960 280 3000 285
rect 3040 635 3080 640
rect 3040 605 3045 635
rect 3075 605 3080 635
rect 3040 556 3080 605
rect 3040 524 3044 556
rect 3076 524 3080 556
rect 3040 476 3080 524
rect 3040 444 3044 476
rect 3076 444 3080 476
rect 3040 396 3080 444
rect 3040 364 3044 396
rect 3076 364 3080 396
rect 3040 315 3080 364
rect 3040 285 3045 315
rect 3075 285 3080 315
rect 3040 280 3080 285
rect 3120 635 3160 640
rect 3120 605 3125 635
rect 3155 605 3160 635
rect 3120 556 3160 605
rect 3120 524 3124 556
rect 3156 524 3160 556
rect 3120 476 3160 524
rect 3120 444 3124 476
rect 3156 444 3160 476
rect 3120 396 3160 444
rect 3120 364 3124 396
rect 3156 364 3160 396
rect 3120 315 3160 364
rect 3120 285 3125 315
rect 3155 285 3160 315
rect 3120 280 3160 285
rect 3200 635 3240 640
rect 3200 605 3205 635
rect 3235 605 3240 635
rect 3200 556 3240 605
rect 3200 524 3204 556
rect 3236 524 3240 556
rect 3200 476 3240 524
rect 3200 444 3204 476
rect 3236 444 3240 476
rect 3200 396 3240 444
rect 3200 364 3204 396
rect 3236 364 3240 396
rect 3200 315 3240 364
rect 3200 285 3205 315
rect 3235 285 3240 315
rect 3200 280 3240 285
rect 3280 635 3320 640
rect 3280 605 3285 635
rect 3315 605 3320 635
rect 3280 556 3320 605
rect 3280 524 3284 556
rect 3316 524 3320 556
rect 3280 476 3320 524
rect 3280 444 3284 476
rect 3316 444 3320 476
rect 3280 396 3320 444
rect 3280 364 3284 396
rect 3316 364 3320 396
rect 3280 315 3320 364
rect 3280 285 3285 315
rect 3315 285 3320 315
rect 3280 280 3320 285
rect 3360 635 3400 640
rect 3360 605 3365 635
rect 3395 605 3400 635
rect 3360 556 3400 605
rect 3360 524 3364 556
rect 3396 524 3400 556
rect 3360 476 3400 524
rect 3360 444 3364 476
rect 3396 444 3400 476
rect 3360 396 3400 444
rect 3360 364 3364 396
rect 3396 364 3400 396
rect 3360 315 3400 364
rect 3360 285 3365 315
rect 3395 285 3400 315
rect 3360 280 3400 285
rect 3440 635 3480 640
rect 3440 605 3445 635
rect 3475 605 3480 635
rect 3440 556 3480 605
rect 3440 524 3444 556
rect 3476 524 3480 556
rect 3440 476 3480 524
rect 3440 444 3444 476
rect 3476 444 3480 476
rect 3440 396 3480 444
rect 3440 364 3444 396
rect 3476 364 3480 396
rect 3440 315 3480 364
rect 3440 285 3445 315
rect 3475 285 3480 315
rect 3440 280 3480 285
rect 3600 635 3640 640
rect 3600 605 3605 635
rect 3635 605 3640 635
rect 3600 556 3640 605
rect 3600 524 3604 556
rect 3636 524 3640 556
rect 3600 476 3640 524
rect 3600 444 3604 476
rect 3636 444 3640 476
rect 3600 396 3640 444
rect 3600 364 3604 396
rect 3636 364 3640 396
rect 3600 315 3640 364
rect 3600 285 3605 315
rect 3635 285 3640 315
rect 3600 280 3640 285
rect 3680 635 3720 640
rect 3680 605 3685 635
rect 3715 605 3720 635
rect 3680 556 3720 605
rect 3680 524 3684 556
rect 3716 524 3720 556
rect 3680 476 3720 524
rect 3680 444 3684 476
rect 3716 444 3720 476
rect 3680 396 3720 444
rect 3680 364 3684 396
rect 3716 364 3720 396
rect 3680 315 3720 364
rect 3680 285 3685 315
rect 3715 285 3720 315
rect 3680 280 3720 285
rect 3760 635 3800 640
rect 3760 605 3765 635
rect 3795 605 3800 635
rect 3760 556 3800 605
rect 3760 524 3764 556
rect 3796 524 3800 556
rect 3760 476 3800 524
rect 3760 444 3764 476
rect 3796 444 3800 476
rect 3760 396 3800 444
rect 3760 364 3764 396
rect 3796 364 3800 396
rect 3760 315 3800 364
rect 3760 285 3765 315
rect 3795 285 3800 315
rect 3760 280 3800 285
rect 3840 635 3880 640
rect 3840 605 3845 635
rect 3875 605 3880 635
rect 3840 556 3880 605
rect 3840 524 3844 556
rect 3876 524 3880 556
rect 3840 476 3880 524
rect 3840 444 3844 476
rect 3876 444 3880 476
rect 3840 396 3880 444
rect 3840 364 3844 396
rect 3876 364 3880 396
rect 3840 315 3880 364
rect 3840 285 3845 315
rect 3875 285 3880 315
rect 3840 280 3880 285
rect 3920 635 3960 640
rect 3920 605 3925 635
rect 3955 605 3960 635
rect 3920 556 3960 605
rect 4000 635 4040 640
rect 4000 605 4005 635
rect 4035 605 4040 635
rect 4000 560 4040 605
rect 4080 635 4120 640
rect 4080 605 4085 635
rect 4115 605 4120 635
rect 3920 524 3924 556
rect 3956 524 3960 556
rect 3920 476 3960 524
rect 3920 444 3924 476
rect 3956 444 3960 476
rect 3920 396 3960 444
rect 3920 364 3924 396
rect 3956 364 3960 396
rect 3920 315 3960 364
rect 4080 556 4120 605
rect 4080 524 4084 556
rect 4116 524 4120 556
rect 4080 476 4120 524
rect 4080 444 4084 476
rect 4116 444 4120 476
rect 4080 396 4120 444
rect 4080 364 4084 396
rect 4116 364 4120 396
rect 3920 285 3925 315
rect 3955 285 3960 315
rect 3920 280 3960 285
rect 4000 315 4040 360
rect 4000 285 4005 315
rect 4035 285 4040 315
rect 4000 280 4040 285
rect 4080 315 4120 364
rect 4080 285 4085 315
rect 4115 285 4120 315
rect 4080 280 4120 285
rect 160 171 200 180
rect 160 89 164 171
rect 196 89 200 171
rect 160 80 200 89
rect 80 -44 120 -40
rect 80 -76 84 -44
rect 116 -76 120 -44
rect 80 -124 120 -76
rect 80 -156 84 -124
rect 116 -156 120 -124
rect 80 -204 120 -156
rect 80 -236 84 -204
rect 116 -236 120 -204
rect 80 -240 120 -236
rect 160 -44 200 -40
rect 160 -76 164 -44
rect 196 -76 200 -44
rect 160 -124 200 -76
rect 160 -156 164 -124
rect 196 -156 200 -124
rect 160 -204 200 -156
rect 160 -236 164 -204
rect 196 -236 200 -204
rect 160 -240 200 -236
rect 240 -44 280 -40
rect 240 -76 244 -44
rect 276 -76 280 -44
rect 240 -124 280 -76
rect 240 -156 244 -124
rect 276 -156 280 -124
rect 240 -204 280 -156
rect 240 -236 244 -204
rect 276 -236 280 -204
rect 240 -240 280 -236
rect 320 -44 360 -40
rect 320 -76 324 -44
rect 356 -76 360 -44
rect 320 -124 360 -76
rect 320 -156 324 -124
rect 356 -156 360 -124
rect 320 -204 360 -156
rect 320 -236 324 -204
rect 356 -236 360 -204
rect 320 -240 360 -236
rect 400 -44 440 -40
rect 400 -76 404 -44
rect 436 -76 440 -44
rect 400 -124 440 -76
rect 400 -156 404 -124
rect 436 -156 440 -124
rect 400 -204 440 -156
rect 400 -236 404 -204
rect 436 -236 440 -204
rect 400 -240 440 -236
rect 480 -44 520 -40
rect 480 -76 484 -44
rect 516 -76 520 -44
rect 480 -124 520 -76
rect 480 -156 484 -124
rect 516 -156 520 -124
rect 480 -204 520 -156
rect 480 -236 484 -204
rect 516 -236 520 -204
rect 480 -240 520 -236
rect 560 -44 600 -40
rect 560 -76 564 -44
rect 596 -76 600 -44
rect 560 -124 600 -76
rect 560 -156 564 -124
rect 596 -156 600 -124
rect 560 -204 600 -156
rect 560 -236 564 -204
rect 596 -236 600 -204
rect 560 -240 600 -236
rect 720 -44 760 -40
rect 720 -76 724 -44
rect 756 -76 760 -44
rect 720 -124 760 -76
rect 720 -156 724 -124
rect 756 -156 760 -124
rect 720 -204 760 -156
rect 720 -236 724 -204
rect 756 -236 760 -204
rect 720 -240 760 -236
rect 800 -44 840 -40
rect 800 -76 804 -44
rect 836 -76 840 -44
rect 800 -124 840 -76
rect 800 -156 804 -124
rect 836 -156 840 -124
rect 800 -204 840 -156
rect 800 -236 804 -204
rect 836 -236 840 -204
rect 800 -240 840 -236
rect 880 -44 920 -40
rect 880 -76 884 -44
rect 916 -76 920 -44
rect 880 -124 920 -76
rect 880 -156 884 -124
rect 916 -156 920 -124
rect 880 -204 920 -156
rect 880 -236 884 -204
rect 916 -236 920 -204
rect 880 -240 920 -236
rect 960 -44 1000 -40
rect 960 -76 964 -44
rect 996 -76 1000 -44
rect 960 -124 1000 -76
rect 960 -156 964 -124
rect 996 -156 1000 -124
rect 960 -204 1000 -156
rect 960 -236 964 -204
rect 996 -236 1000 -204
rect 960 -240 1000 -236
rect 1040 -44 1080 -40
rect 1040 -76 1044 -44
rect 1076 -76 1080 -44
rect 1040 -124 1080 -76
rect 1040 -156 1044 -124
rect 1076 -156 1080 -124
rect 1040 -204 1080 -156
rect 1040 -236 1044 -204
rect 1076 -236 1080 -204
rect 1040 -240 1080 -236
rect 1120 -44 1160 -40
rect 1120 -76 1124 -44
rect 1156 -76 1160 -44
rect 1120 -124 1160 -76
rect 1120 -156 1124 -124
rect 1156 -156 1160 -124
rect 1120 -204 1160 -156
rect 1120 -236 1124 -204
rect 1156 -236 1160 -204
rect 1120 -240 1160 -236
rect 1200 -44 1240 -40
rect 1200 -76 1204 -44
rect 1236 -76 1240 -44
rect 1200 -124 1240 -76
rect 1200 -156 1204 -124
rect 1236 -156 1240 -124
rect 1200 -204 1240 -156
rect 1200 -236 1204 -204
rect 1236 -236 1240 -204
rect 1200 -240 1240 -236
rect 1280 -44 1320 -40
rect 1280 -76 1284 -44
rect 1316 -76 1320 -44
rect 1280 -124 1320 -76
rect 1280 -156 1284 -124
rect 1316 -156 1320 -124
rect 1280 -204 1320 -156
rect 1280 -236 1284 -204
rect 1316 -236 1320 -204
rect 1280 -240 1320 -236
rect 1360 -44 1400 -40
rect 1360 -76 1364 -44
rect 1396 -76 1400 -44
rect 1360 -124 1400 -76
rect 1360 -156 1364 -124
rect 1396 -156 1400 -124
rect 1360 -204 1400 -156
rect 1360 -236 1364 -204
rect 1396 -236 1400 -204
rect 1360 -240 1400 -236
rect 1440 -44 1480 -40
rect 1440 -76 1444 -44
rect 1476 -76 1480 -44
rect 1440 -124 1480 -76
rect 1440 -156 1444 -124
rect 1476 -156 1480 -124
rect 1440 -204 1480 -156
rect 1440 -236 1444 -204
rect 1476 -236 1480 -204
rect 1440 -240 1480 -236
rect 1520 -44 1560 -40
rect 1520 -76 1524 -44
rect 1556 -76 1560 -44
rect 1520 -124 1560 -76
rect 1520 -156 1524 -124
rect 1556 -156 1560 -124
rect 1520 -204 1560 -156
rect 1520 -236 1524 -204
rect 1556 -236 1560 -204
rect 1520 -240 1560 -236
rect 1680 -44 1720 -40
rect 1680 -76 1684 -44
rect 1716 -76 1720 -44
rect 1680 -124 1720 -76
rect 1680 -156 1684 -124
rect 1716 -156 1720 -124
rect 1680 -204 1720 -156
rect 1680 -236 1684 -204
rect 1716 -236 1720 -204
rect 1680 -240 1720 -236
rect 1760 -44 1800 -40
rect 1760 -76 1764 -44
rect 1796 -76 1800 -44
rect 1760 -124 1800 -76
rect 1760 -156 1764 -124
rect 1796 -156 1800 -124
rect 1760 -204 1800 -156
rect 1760 -236 1764 -204
rect 1796 -236 1800 -204
rect 1760 -240 1800 -236
rect 1840 -44 1880 -40
rect 1840 -76 1844 -44
rect 1876 -76 1880 -44
rect 1840 -124 1880 -76
rect 1840 -156 1844 -124
rect 1876 -156 1880 -124
rect 1840 -204 1880 -156
rect 1840 -236 1844 -204
rect 1876 -236 1880 -204
rect 1840 -240 1880 -236
rect 1920 -44 1960 -40
rect 1920 -76 1924 -44
rect 1956 -76 1960 -44
rect 1920 -124 1960 -76
rect 1920 -156 1924 -124
rect 1956 -156 1960 -124
rect 1920 -204 1960 -156
rect 1920 -236 1924 -204
rect 1956 -236 1960 -204
rect 1920 -240 1960 -236
rect 2000 -44 2040 -40
rect 2000 -76 2004 -44
rect 2036 -76 2040 -44
rect 2000 -124 2040 -76
rect 2000 -156 2004 -124
rect 2036 -156 2040 -124
rect 2000 -204 2040 -156
rect 2000 -236 2004 -204
rect 2036 -236 2040 -204
rect 2000 -240 2040 -236
rect 2080 -44 2120 -40
rect 2080 -76 2084 -44
rect 2116 -76 2120 -44
rect 2080 -124 2120 -76
rect 2080 -156 2084 -124
rect 2116 -156 2120 -124
rect 2080 -204 2120 -156
rect 2080 -236 2084 -204
rect 2116 -236 2120 -204
rect 2080 -240 2120 -236
rect 2160 -44 2200 -40
rect 2160 -76 2164 -44
rect 2196 -76 2200 -44
rect 2160 -124 2200 -76
rect 2160 -156 2164 -124
rect 2196 -156 2200 -124
rect 2160 -204 2200 -156
rect 2160 -236 2164 -204
rect 2196 -236 2200 -204
rect 2160 -240 2200 -236
rect 2240 -44 2280 -40
rect 2240 -76 2244 -44
rect 2276 -76 2280 -44
rect 2240 -124 2280 -76
rect 2240 -156 2244 -124
rect 2276 -156 2280 -124
rect 2240 -204 2280 -156
rect 2240 -236 2244 -204
rect 2276 -236 2280 -204
rect 2240 -240 2280 -236
rect 2320 -44 2360 -40
rect 2320 -76 2324 -44
rect 2356 -76 2360 -44
rect 2320 -124 2360 -76
rect 2320 -156 2324 -124
rect 2356 -156 2360 -124
rect 2320 -204 2360 -156
rect 2320 -236 2324 -204
rect 2356 -236 2360 -204
rect 2320 -240 2360 -236
rect 2400 -44 2440 -40
rect 2400 -76 2404 -44
rect 2436 -76 2440 -44
rect 2400 -124 2440 -76
rect 2400 -156 2404 -124
rect 2436 -156 2440 -124
rect 2400 -204 2440 -156
rect 2400 -236 2404 -204
rect 2436 -236 2440 -204
rect 2400 -240 2440 -236
rect 2480 -44 2520 -40
rect 2480 -76 2484 -44
rect 2516 -76 2520 -44
rect 2480 -124 2520 -76
rect 2480 -156 2484 -124
rect 2516 -156 2520 -124
rect 2480 -204 2520 -156
rect 2480 -236 2484 -204
rect 2516 -236 2520 -204
rect 2480 -240 2520 -236
rect 2640 -44 2680 -40
rect 2640 -76 2644 -44
rect 2676 -76 2680 -44
rect 2640 -124 2680 -76
rect 2640 -156 2644 -124
rect 2676 -156 2680 -124
rect 2640 -204 2680 -156
rect 2640 -236 2644 -204
rect 2676 -236 2680 -204
rect 2640 -240 2680 -236
rect 2720 -44 2760 -40
rect 2720 -76 2724 -44
rect 2756 -76 2760 -44
rect 2720 -124 2760 -76
rect 2720 -156 2724 -124
rect 2756 -156 2760 -124
rect 2720 -204 2760 -156
rect 2720 -236 2724 -204
rect 2756 -236 2760 -204
rect 2720 -240 2760 -236
rect 2800 -44 2840 -40
rect 2800 -76 2804 -44
rect 2836 -76 2840 -44
rect 2800 -124 2840 -76
rect 2800 -156 2804 -124
rect 2836 -156 2840 -124
rect 2800 -204 2840 -156
rect 2800 -236 2804 -204
rect 2836 -236 2840 -204
rect 2800 -240 2840 -236
rect 2880 -44 2920 -40
rect 2880 -76 2884 -44
rect 2916 -76 2920 -44
rect 2880 -124 2920 -76
rect 2880 -156 2884 -124
rect 2916 -156 2920 -124
rect 2880 -204 2920 -156
rect 2880 -236 2884 -204
rect 2916 -236 2920 -204
rect 2880 -240 2920 -236
rect 2960 -44 3000 -40
rect 2960 -76 2964 -44
rect 2996 -76 3000 -44
rect 2960 -124 3000 -76
rect 2960 -156 2964 -124
rect 2996 -156 3000 -124
rect 2960 -204 3000 -156
rect 2960 -236 2964 -204
rect 2996 -236 3000 -204
rect 2960 -240 3000 -236
rect 3040 -44 3080 -40
rect 3040 -76 3044 -44
rect 3076 -76 3080 -44
rect 3040 -124 3080 -76
rect 3040 -156 3044 -124
rect 3076 -156 3080 -124
rect 3040 -204 3080 -156
rect 3040 -236 3044 -204
rect 3076 -236 3080 -204
rect 3040 -240 3080 -236
rect 3120 -44 3160 -40
rect 3120 -76 3124 -44
rect 3156 -76 3160 -44
rect 3120 -124 3160 -76
rect 3120 -156 3124 -124
rect 3156 -156 3160 -124
rect 3120 -204 3160 -156
rect 3120 -236 3124 -204
rect 3156 -236 3160 -204
rect 3120 -240 3160 -236
rect 3200 -44 3240 -40
rect 3200 -76 3204 -44
rect 3236 -76 3240 -44
rect 3200 -124 3240 -76
rect 3200 -156 3204 -124
rect 3236 -156 3240 -124
rect 3200 -204 3240 -156
rect 3200 -236 3204 -204
rect 3236 -236 3240 -204
rect 3200 -240 3240 -236
rect 3280 -44 3320 -40
rect 3280 -76 3284 -44
rect 3316 -76 3320 -44
rect 3280 -124 3320 -76
rect 3280 -156 3284 -124
rect 3316 -156 3320 -124
rect 3280 -204 3320 -156
rect 3280 -236 3284 -204
rect 3316 -236 3320 -204
rect 3280 -240 3320 -236
rect 3360 -44 3400 -40
rect 3360 -76 3364 -44
rect 3396 -76 3400 -44
rect 3360 -124 3400 -76
rect 3360 -156 3364 -124
rect 3396 -156 3400 -124
rect 3360 -204 3400 -156
rect 3360 -236 3364 -204
rect 3396 -236 3400 -204
rect 3360 -240 3400 -236
rect 3440 -44 3480 -40
rect 3440 -76 3444 -44
rect 3476 -76 3480 -44
rect 3440 -124 3480 -76
rect 3440 -156 3444 -124
rect 3476 -156 3480 -124
rect 3440 -204 3480 -156
rect 3440 -236 3444 -204
rect 3476 -236 3480 -204
rect 3440 -240 3480 -236
rect 3600 -44 3640 -40
rect 3600 -76 3604 -44
rect 3636 -76 3640 -44
rect 3600 -124 3640 -76
rect 3600 -156 3604 -124
rect 3636 -156 3640 -124
rect 3600 -204 3640 -156
rect 3600 -236 3604 -204
rect 3636 -236 3640 -204
rect 3600 -240 3640 -236
rect 3680 -44 3720 -40
rect 3680 -76 3684 -44
rect 3716 -76 3720 -44
rect 3680 -124 3720 -76
rect 3680 -156 3684 -124
rect 3716 -156 3720 -124
rect 3680 -204 3720 -156
rect 3680 -236 3684 -204
rect 3716 -236 3720 -204
rect 3680 -240 3720 -236
rect 3760 -44 3800 -40
rect 3760 -76 3764 -44
rect 3796 -76 3800 -44
rect 3760 -124 3800 -76
rect 3760 -156 3764 -124
rect 3796 -156 3800 -124
rect 3760 -204 3800 -156
rect 3760 -236 3764 -204
rect 3796 -236 3800 -204
rect 3760 -240 3800 -236
rect 3840 -44 3880 -40
rect 3840 -76 3844 -44
rect 3876 -76 3880 -44
rect 3840 -124 3880 -76
rect 3840 -156 3844 -124
rect 3876 -156 3880 -124
rect 3840 -204 3880 -156
rect 3840 -236 3844 -204
rect 3876 -236 3880 -204
rect 3840 -240 3880 -236
rect 3920 -44 3960 -40
rect 3920 -76 3924 -44
rect 3956 -76 3960 -44
rect 3920 -124 3960 -76
rect 3920 -156 3924 -124
rect 3956 -156 3960 -124
rect 3920 -204 3960 -156
rect 3920 -236 3924 -204
rect 3956 -236 3960 -204
rect 3920 -240 3960 -236
rect 4080 -44 4120 -40
rect 4080 -76 4084 -44
rect 4116 -76 4120 -44
rect 4080 -124 4120 -76
rect 4080 -156 4084 -124
rect 4116 -156 4120 -124
rect 4080 -204 4120 -156
rect 4080 -236 4084 -204
rect 4116 -236 4120 -204
rect 4080 -240 4120 -236
rect 160 -349 200 -340
rect 160 -431 164 -349
rect 196 -431 200 -349
rect 160 -440 200 -431
<< via3 >>
rect 164 4870 196 4871
rect 164 4690 165 4870
rect 165 4690 195 4870
rect 195 4690 196 4870
rect 164 4689 196 4690
rect 84 4395 116 4396
rect 84 4365 85 4395
rect 85 4365 115 4395
rect 115 4365 116 4395
rect 84 4364 116 4365
rect 84 4284 116 4316
rect 84 4235 116 4236
rect 84 4205 85 4235
rect 85 4205 115 4235
rect 115 4205 116 4235
rect 84 4204 116 4205
rect 164 4395 196 4396
rect 164 4365 165 4395
rect 165 4365 195 4395
rect 195 4365 196 4395
rect 164 4364 196 4365
rect 164 4284 196 4316
rect 164 4235 196 4236
rect 164 4205 165 4235
rect 165 4205 195 4235
rect 195 4205 196 4235
rect 164 4204 196 4205
rect 244 4395 276 4396
rect 244 4365 245 4395
rect 245 4365 275 4395
rect 275 4365 276 4395
rect 244 4364 276 4365
rect 244 4284 276 4316
rect 244 4235 276 4236
rect 244 4205 245 4235
rect 245 4205 275 4235
rect 275 4205 276 4235
rect 244 4204 276 4205
rect 324 4395 356 4396
rect 324 4365 325 4395
rect 325 4365 355 4395
rect 355 4365 356 4395
rect 324 4364 356 4365
rect 324 4284 356 4316
rect 324 4235 356 4236
rect 324 4205 325 4235
rect 325 4205 355 4235
rect 355 4205 356 4235
rect 324 4204 356 4205
rect 404 4395 436 4396
rect 404 4365 405 4395
rect 405 4365 435 4395
rect 435 4365 436 4395
rect 404 4364 436 4365
rect 404 4284 436 4316
rect 404 4235 436 4236
rect 404 4205 405 4235
rect 405 4205 435 4235
rect 435 4205 436 4235
rect 404 4204 436 4205
rect 484 4395 516 4396
rect 484 4365 485 4395
rect 485 4365 515 4395
rect 515 4365 516 4395
rect 484 4364 516 4365
rect 484 4284 516 4316
rect 484 4235 516 4236
rect 484 4205 485 4235
rect 485 4205 515 4235
rect 515 4205 516 4235
rect 484 4204 516 4205
rect 564 4395 596 4396
rect 564 4365 565 4395
rect 565 4365 595 4395
rect 595 4365 596 4395
rect 564 4364 596 4365
rect 564 4284 596 4316
rect 564 4235 596 4236
rect 564 4205 565 4235
rect 565 4205 595 4235
rect 595 4205 596 4235
rect 564 4204 596 4205
rect 724 4395 756 4396
rect 724 4365 725 4395
rect 725 4365 755 4395
rect 755 4365 756 4395
rect 724 4364 756 4365
rect 724 4284 756 4316
rect 724 4235 756 4236
rect 724 4205 725 4235
rect 725 4205 755 4235
rect 755 4205 756 4235
rect 724 4204 756 4205
rect 804 4395 836 4396
rect 804 4365 805 4395
rect 805 4365 835 4395
rect 835 4365 836 4395
rect 804 4364 836 4365
rect 804 4284 836 4316
rect 804 4235 836 4236
rect 804 4205 805 4235
rect 805 4205 835 4235
rect 835 4205 836 4235
rect 804 4204 836 4205
rect 884 4395 916 4396
rect 884 4365 885 4395
rect 885 4365 915 4395
rect 915 4365 916 4395
rect 884 4364 916 4365
rect 884 4284 916 4316
rect 884 4235 916 4236
rect 884 4205 885 4235
rect 885 4205 915 4235
rect 915 4205 916 4235
rect 884 4204 916 4205
rect 964 4395 996 4396
rect 964 4365 965 4395
rect 965 4365 995 4395
rect 995 4365 996 4395
rect 964 4364 996 4365
rect 964 4284 996 4316
rect 964 4235 996 4236
rect 964 4205 965 4235
rect 965 4205 995 4235
rect 995 4205 996 4235
rect 964 4204 996 4205
rect 1044 4395 1076 4396
rect 1044 4365 1045 4395
rect 1045 4365 1075 4395
rect 1075 4365 1076 4395
rect 1044 4364 1076 4365
rect 1044 4284 1076 4316
rect 1044 4235 1076 4236
rect 1044 4205 1045 4235
rect 1045 4205 1075 4235
rect 1075 4205 1076 4235
rect 1044 4204 1076 4205
rect 1124 4395 1156 4396
rect 1124 4365 1125 4395
rect 1125 4365 1155 4395
rect 1155 4365 1156 4395
rect 1124 4364 1156 4365
rect 1124 4284 1156 4316
rect 1124 4235 1156 4236
rect 1124 4205 1125 4235
rect 1125 4205 1155 4235
rect 1155 4205 1156 4235
rect 1124 4204 1156 4205
rect 1204 4395 1236 4396
rect 1204 4365 1205 4395
rect 1205 4365 1235 4395
rect 1235 4365 1236 4395
rect 1204 4364 1236 4365
rect 1204 4284 1236 4316
rect 1204 4235 1236 4236
rect 1204 4205 1205 4235
rect 1205 4205 1235 4235
rect 1235 4205 1236 4235
rect 1204 4204 1236 4205
rect 1284 4395 1316 4396
rect 1284 4365 1285 4395
rect 1285 4365 1315 4395
rect 1315 4365 1316 4395
rect 1284 4364 1316 4365
rect 1284 4284 1316 4316
rect 1284 4235 1316 4236
rect 1284 4205 1285 4235
rect 1285 4205 1315 4235
rect 1315 4205 1316 4235
rect 1284 4204 1316 4205
rect 1364 4395 1396 4396
rect 1364 4365 1365 4395
rect 1365 4365 1395 4395
rect 1395 4365 1396 4395
rect 1364 4364 1396 4365
rect 1364 4284 1396 4316
rect 1364 4235 1396 4236
rect 1364 4205 1365 4235
rect 1365 4205 1395 4235
rect 1395 4205 1396 4235
rect 1364 4204 1396 4205
rect 1444 4395 1476 4396
rect 1444 4365 1445 4395
rect 1445 4365 1475 4395
rect 1475 4365 1476 4395
rect 1444 4364 1476 4365
rect 1444 4284 1476 4316
rect 1444 4235 1476 4236
rect 1444 4205 1445 4235
rect 1445 4205 1475 4235
rect 1475 4205 1476 4235
rect 1444 4204 1476 4205
rect 1524 4395 1556 4396
rect 1524 4365 1525 4395
rect 1525 4365 1555 4395
rect 1555 4365 1556 4395
rect 1524 4364 1556 4365
rect 1524 4284 1556 4316
rect 1524 4235 1556 4236
rect 1524 4205 1525 4235
rect 1525 4205 1555 4235
rect 1555 4205 1556 4235
rect 1524 4204 1556 4205
rect 1684 4395 1716 4396
rect 1684 4365 1685 4395
rect 1685 4365 1715 4395
rect 1715 4365 1716 4395
rect 1684 4364 1716 4365
rect 1684 4284 1716 4316
rect 1684 4235 1716 4236
rect 1684 4205 1685 4235
rect 1685 4205 1715 4235
rect 1715 4205 1716 4235
rect 1684 4204 1716 4205
rect 1764 4395 1796 4396
rect 1764 4365 1765 4395
rect 1765 4365 1795 4395
rect 1795 4365 1796 4395
rect 1764 4364 1796 4365
rect 1764 4284 1796 4316
rect 1764 4235 1796 4236
rect 1764 4205 1765 4235
rect 1765 4205 1795 4235
rect 1795 4205 1796 4235
rect 1764 4204 1796 4205
rect 1844 4395 1876 4396
rect 1844 4365 1845 4395
rect 1845 4365 1875 4395
rect 1875 4365 1876 4395
rect 1844 4364 1876 4365
rect 1844 4284 1876 4316
rect 1844 4235 1876 4236
rect 1844 4205 1845 4235
rect 1845 4205 1875 4235
rect 1875 4205 1876 4235
rect 1844 4204 1876 4205
rect 1924 4395 1956 4396
rect 1924 4365 1925 4395
rect 1925 4365 1955 4395
rect 1955 4365 1956 4395
rect 1924 4364 1956 4365
rect 1924 4284 1956 4316
rect 1924 4235 1956 4236
rect 1924 4205 1925 4235
rect 1925 4205 1955 4235
rect 1955 4205 1956 4235
rect 1924 4204 1956 4205
rect 2004 4395 2036 4396
rect 2004 4365 2005 4395
rect 2005 4365 2035 4395
rect 2035 4365 2036 4395
rect 2004 4364 2036 4365
rect 2004 4284 2036 4316
rect 2004 4235 2036 4236
rect 2004 4205 2005 4235
rect 2005 4205 2035 4235
rect 2035 4205 2036 4235
rect 2004 4204 2036 4205
rect 2084 4395 2116 4396
rect 2084 4365 2085 4395
rect 2085 4365 2115 4395
rect 2115 4365 2116 4395
rect 2084 4364 2116 4365
rect 2084 4284 2116 4316
rect 2084 4235 2116 4236
rect 2084 4205 2085 4235
rect 2085 4205 2115 4235
rect 2115 4205 2116 4235
rect 2084 4204 2116 4205
rect 2164 4395 2196 4396
rect 2164 4365 2165 4395
rect 2165 4365 2195 4395
rect 2195 4365 2196 4395
rect 2164 4364 2196 4365
rect 2164 4284 2196 4316
rect 2164 4235 2196 4236
rect 2164 4205 2165 4235
rect 2165 4205 2195 4235
rect 2195 4205 2196 4235
rect 2164 4204 2196 4205
rect 2244 4395 2276 4396
rect 2244 4365 2245 4395
rect 2245 4365 2275 4395
rect 2275 4365 2276 4395
rect 2244 4364 2276 4365
rect 2244 4284 2276 4316
rect 2244 4235 2276 4236
rect 2244 4205 2245 4235
rect 2245 4205 2275 4235
rect 2275 4205 2276 4235
rect 2244 4204 2276 4205
rect 2324 4395 2356 4396
rect 2324 4365 2325 4395
rect 2325 4365 2355 4395
rect 2355 4365 2356 4395
rect 2324 4364 2356 4365
rect 2324 4284 2356 4316
rect 2324 4235 2356 4236
rect 2324 4205 2325 4235
rect 2325 4205 2355 4235
rect 2355 4205 2356 4235
rect 2324 4204 2356 4205
rect 2404 4395 2436 4396
rect 2404 4365 2405 4395
rect 2405 4365 2435 4395
rect 2435 4365 2436 4395
rect 2404 4364 2436 4365
rect 2404 4284 2436 4316
rect 2404 4235 2436 4236
rect 2404 4205 2405 4235
rect 2405 4205 2435 4235
rect 2435 4205 2436 4235
rect 2404 4204 2436 4205
rect 2484 4395 2516 4396
rect 2484 4365 2485 4395
rect 2485 4365 2515 4395
rect 2515 4365 2516 4395
rect 2484 4364 2516 4365
rect 2484 4284 2516 4316
rect 2484 4235 2516 4236
rect 2484 4205 2485 4235
rect 2485 4205 2515 4235
rect 2515 4205 2516 4235
rect 2484 4204 2516 4205
rect 2644 4395 2676 4396
rect 2644 4365 2645 4395
rect 2645 4365 2675 4395
rect 2675 4365 2676 4395
rect 2644 4364 2676 4365
rect 2644 4284 2676 4316
rect 2644 4235 2676 4236
rect 2644 4205 2645 4235
rect 2645 4205 2675 4235
rect 2675 4205 2676 4235
rect 2644 4204 2676 4205
rect 2724 4395 2756 4396
rect 2724 4365 2725 4395
rect 2725 4365 2755 4395
rect 2755 4365 2756 4395
rect 2724 4364 2756 4365
rect 2724 4284 2756 4316
rect 2724 4235 2756 4236
rect 2724 4205 2725 4235
rect 2725 4205 2755 4235
rect 2755 4205 2756 4235
rect 2724 4204 2756 4205
rect 2804 4395 2836 4396
rect 2804 4365 2805 4395
rect 2805 4365 2835 4395
rect 2835 4365 2836 4395
rect 2804 4364 2836 4365
rect 2804 4284 2836 4316
rect 2804 4235 2836 4236
rect 2804 4205 2805 4235
rect 2805 4205 2835 4235
rect 2835 4205 2836 4235
rect 2804 4204 2836 4205
rect 2884 4395 2916 4396
rect 2884 4365 2885 4395
rect 2885 4365 2915 4395
rect 2915 4365 2916 4395
rect 2884 4364 2916 4365
rect 2884 4284 2916 4316
rect 2884 4235 2916 4236
rect 2884 4205 2885 4235
rect 2885 4205 2915 4235
rect 2915 4205 2916 4235
rect 2884 4204 2916 4205
rect 2964 4395 2996 4396
rect 2964 4365 2965 4395
rect 2965 4365 2995 4395
rect 2995 4365 2996 4395
rect 2964 4364 2996 4365
rect 2964 4284 2996 4316
rect 2964 4235 2996 4236
rect 2964 4205 2965 4235
rect 2965 4205 2995 4235
rect 2995 4205 2996 4235
rect 2964 4204 2996 4205
rect 3044 4395 3076 4396
rect 3044 4365 3045 4395
rect 3045 4365 3075 4395
rect 3075 4365 3076 4395
rect 3044 4364 3076 4365
rect 3044 4284 3076 4316
rect 3044 4235 3076 4236
rect 3044 4205 3045 4235
rect 3045 4205 3075 4235
rect 3075 4205 3076 4235
rect 3044 4204 3076 4205
rect 3124 4395 3156 4396
rect 3124 4365 3125 4395
rect 3125 4365 3155 4395
rect 3155 4365 3156 4395
rect 3124 4364 3156 4365
rect 3124 4284 3156 4316
rect 3124 4235 3156 4236
rect 3124 4205 3125 4235
rect 3125 4205 3155 4235
rect 3155 4205 3156 4235
rect 3124 4204 3156 4205
rect 3204 4395 3236 4396
rect 3204 4365 3205 4395
rect 3205 4365 3235 4395
rect 3235 4365 3236 4395
rect 3204 4364 3236 4365
rect 3204 4284 3236 4316
rect 3204 4235 3236 4236
rect 3204 4205 3205 4235
rect 3205 4205 3235 4235
rect 3235 4205 3236 4235
rect 3204 4204 3236 4205
rect 3284 4395 3316 4396
rect 3284 4365 3285 4395
rect 3285 4365 3315 4395
rect 3315 4365 3316 4395
rect 3284 4364 3316 4365
rect 3284 4284 3316 4316
rect 3284 4235 3316 4236
rect 3284 4205 3285 4235
rect 3285 4205 3315 4235
rect 3315 4205 3316 4235
rect 3284 4204 3316 4205
rect 3364 4395 3396 4396
rect 3364 4365 3365 4395
rect 3365 4365 3395 4395
rect 3395 4365 3396 4395
rect 3364 4364 3396 4365
rect 3364 4284 3396 4316
rect 3364 4235 3396 4236
rect 3364 4205 3365 4235
rect 3365 4205 3395 4235
rect 3395 4205 3396 4235
rect 3364 4204 3396 4205
rect 3444 4395 3476 4396
rect 3444 4365 3445 4395
rect 3445 4365 3475 4395
rect 3475 4365 3476 4395
rect 3444 4364 3476 4365
rect 3444 4284 3476 4316
rect 3444 4235 3476 4236
rect 3444 4205 3445 4235
rect 3445 4205 3475 4235
rect 3475 4205 3476 4235
rect 3444 4204 3476 4205
rect 3604 4395 3636 4396
rect 3604 4365 3605 4395
rect 3605 4365 3635 4395
rect 3635 4365 3636 4395
rect 3604 4364 3636 4365
rect 3604 4284 3636 4316
rect 3604 4235 3636 4236
rect 3604 4205 3605 4235
rect 3605 4205 3635 4235
rect 3635 4205 3636 4235
rect 3604 4204 3636 4205
rect 3684 4395 3716 4396
rect 3684 4365 3685 4395
rect 3685 4365 3715 4395
rect 3715 4365 3716 4395
rect 3684 4364 3716 4365
rect 3684 4284 3716 4316
rect 3684 4235 3716 4236
rect 3684 4205 3685 4235
rect 3685 4205 3715 4235
rect 3715 4205 3716 4235
rect 3684 4204 3716 4205
rect 3764 4395 3796 4396
rect 3764 4365 3765 4395
rect 3765 4365 3795 4395
rect 3795 4365 3796 4395
rect 3764 4364 3796 4365
rect 3764 4284 3796 4316
rect 3764 4235 3796 4236
rect 3764 4205 3765 4235
rect 3765 4205 3795 4235
rect 3795 4205 3796 4235
rect 3764 4204 3796 4205
rect 3844 4395 3876 4396
rect 3844 4365 3845 4395
rect 3845 4365 3875 4395
rect 3875 4365 3876 4395
rect 3844 4364 3876 4365
rect 3844 4284 3876 4316
rect 3844 4235 3876 4236
rect 3844 4205 3845 4235
rect 3845 4205 3875 4235
rect 3875 4205 3876 4235
rect 3844 4204 3876 4205
rect 3924 4395 3956 4396
rect 3924 4365 3925 4395
rect 3925 4365 3955 4395
rect 3955 4365 3956 4395
rect 3924 4364 3956 4365
rect 3924 4284 3956 4316
rect 3924 4235 3956 4236
rect 3924 4205 3925 4235
rect 3925 4205 3955 4235
rect 3955 4205 3956 4235
rect 3924 4204 3956 4205
rect 4004 4395 4036 4396
rect 4004 4365 4005 4395
rect 4005 4365 4035 4395
rect 4035 4365 4036 4395
rect 4004 4364 4036 4365
rect 4004 4284 4036 4316
rect 4004 4235 4036 4236
rect 4004 4205 4005 4235
rect 4005 4205 4035 4235
rect 4035 4205 4036 4235
rect 4004 4204 4036 4205
rect 4084 4395 4116 4396
rect 4084 4365 4085 4395
rect 4085 4365 4115 4395
rect 4115 4365 4116 4395
rect 4084 4364 4116 4365
rect 4084 4284 4116 4316
rect 4084 4235 4116 4236
rect 4084 4205 4085 4235
rect 4085 4205 4115 4235
rect 4115 4205 4116 4235
rect 4084 4204 4116 4205
rect 84 4155 116 4156
rect 84 4125 85 4155
rect 85 4125 115 4155
rect 115 4125 116 4155
rect 84 4124 116 4125
rect 84 4044 116 4076
rect 84 3995 116 3996
rect 84 3965 85 3995
rect 85 3965 115 3995
rect 115 3965 116 3995
rect 84 3964 116 3965
rect 164 4155 196 4156
rect 164 4125 165 4155
rect 165 4125 195 4155
rect 195 4125 196 4155
rect 164 4124 196 4125
rect 164 4044 196 4076
rect 164 3995 196 3996
rect 164 3965 165 3995
rect 165 3965 195 3995
rect 195 3965 196 3995
rect 164 3964 196 3965
rect 244 4155 276 4156
rect 244 4125 245 4155
rect 245 4125 275 4155
rect 275 4125 276 4155
rect 244 4124 276 4125
rect 244 4044 276 4076
rect 244 3995 276 3996
rect 244 3965 245 3995
rect 245 3965 275 3995
rect 275 3965 276 3995
rect 244 3964 276 3965
rect 324 4155 356 4156
rect 324 4125 325 4155
rect 325 4125 355 4155
rect 355 4125 356 4155
rect 324 4124 356 4125
rect 324 4044 356 4076
rect 324 3995 356 3996
rect 324 3965 325 3995
rect 325 3965 355 3995
rect 355 3965 356 3995
rect 324 3964 356 3965
rect 404 4155 436 4156
rect 404 4125 405 4155
rect 405 4125 435 4155
rect 435 4125 436 4155
rect 404 4124 436 4125
rect 404 4044 436 4076
rect 404 3995 436 3996
rect 404 3965 405 3995
rect 405 3965 435 3995
rect 435 3965 436 3995
rect 404 3964 436 3965
rect 484 4155 516 4156
rect 484 4125 485 4155
rect 485 4125 515 4155
rect 515 4125 516 4155
rect 484 4124 516 4125
rect 484 4044 516 4076
rect 484 3995 516 3996
rect 484 3965 485 3995
rect 485 3965 515 3995
rect 515 3965 516 3995
rect 484 3964 516 3965
rect 564 4155 596 4156
rect 564 4125 565 4155
rect 565 4125 595 4155
rect 595 4125 596 4155
rect 564 4124 596 4125
rect 564 4044 596 4076
rect 564 3995 596 3996
rect 564 3965 565 3995
rect 565 3965 595 3995
rect 595 3965 596 3995
rect 564 3964 596 3965
rect 724 4155 756 4156
rect 724 4125 725 4155
rect 725 4125 755 4155
rect 755 4125 756 4155
rect 724 4124 756 4125
rect 724 4044 756 4076
rect 724 3995 756 3996
rect 724 3965 725 3995
rect 725 3965 755 3995
rect 755 3965 756 3995
rect 724 3964 756 3965
rect 804 4155 836 4156
rect 804 4125 805 4155
rect 805 4125 835 4155
rect 835 4125 836 4155
rect 804 4124 836 4125
rect 804 4044 836 4076
rect 804 3995 836 3996
rect 804 3965 805 3995
rect 805 3965 835 3995
rect 835 3965 836 3995
rect 804 3964 836 3965
rect 884 4155 916 4156
rect 884 4125 885 4155
rect 885 4125 915 4155
rect 915 4125 916 4155
rect 884 4124 916 4125
rect 884 4044 916 4076
rect 884 3995 916 3996
rect 884 3965 885 3995
rect 885 3965 915 3995
rect 915 3965 916 3995
rect 884 3964 916 3965
rect 964 4155 996 4156
rect 964 4125 965 4155
rect 965 4125 995 4155
rect 995 4125 996 4155
rect 964 4124 996 4125
rect 964 4044 996 4076
rect 964 3995 996 3996
rect 964 3965 965 3995
rect 965 3965 995 3995
rect 995 3965 996 3995
rect 964 3964 996 3965
rect 1044 4155 1076 4156
rect 1044 4125 1045 4155
rect 1045 4125 1075 4155
rect 1075 4125 1076 4155
rect 1044 4124 1076 4125
rect 1044 4044 1076 4076
rect 1044 3995 1076 3996
rect 1044 3965 1045 3995
rect 1045 3965 1075 3995
rect 1075 3965 1076 3995
rect 1044 3964 1076 3965
rect 1124 4155 1156 4156
rect 1124 4125 1125 4155
rect 1125 4125 1155 4155
rect 1155 4125 1156 4155
rect 1124 4124 1156 4125
rect 1124 4044 1156 4076
rect 1124 3995 1156 3996
rect 1124 3965 1125 3995
rect 1125 3965 1155 3995
rect 1155 3965 1156 3995
rect 1124 3964 1156 3965
rect 1204 4155 1236 4156
rect 1204 4125 1205 4155
rect 1205 4125 1235 4155
rect 1235 4125 1236 4155
rect 1204 4124 1236 4125
rect 1204 4044 1236 4076
rect 1204 3995 1236 3996
rect 1204 3965 1205 3995
rect 1205 3965 1235 3995
rect 1235 3965 1236 3995
rect 1204 3964 1236 3965
rect 1284 4155 1316 4156
rect 1284 4125 1285 4155
rect 1285 4125 1315 4155
rect 1315 4125 1316 4155
rect 1284 4124 1316 4125
rect 1284 4044 1316 4076
rect 1284 3995 1316 3996
rect 1284 3965 1285 3995
rect 1285 3965 1315 3995
rect 1315 3965 1316 3995
rect 1284 3964 1316 3965
rect 1364 4155 1396 4156
rect 1364 4125 1365 4155
rect 1365 4125 1395 4155
rect 1395 4125 1396 4155
rect 1364 4124 1396 4125
rect 1364 4044 1396 4076
rect 1364 3995 1396 3996
rect 1364 3965 1365 3995
rect 1365 3965 1395 3995
rect 1395 3965 1396 3995
rect 1364 3964 1396 3965
rect 1444 4155 1476 4156
rect 1444 4125 1445 4155
rect 1445 4125 1475 4155
rect 1475 4125 1476 4155
rect 1444 4124 1476 4125
rect 1444 4044 1476 4076
rect 1444 3995 1476 3996
rect 1444 3965 1445 3995
rect 1445 3965 1475 3995
rect 1475 3965 1476 3995
rect 1444 3964 1476 3965
rect 1524 4155 1556 4156
rect 1524 4125 1525 4155
rect 1525 4125 1555 4155
rect 1555 4125 1556 4155
rect 1524 4124 1556 4125
rect 1524 4044 1556 4076
rect 1524 3995 1556 3996
rect 1524 3965 1525 3995
rect 1525 3965 1555 3995
rect 1555 3965 1556 3995
rect 1524 3964 1556 3965
rect 1684 4155 1716 4156
rect 1684 4125 1685 4155
rect 1685 4125 1715 4155
rect 1715 4125 1716 4155
rect 1684 4124 1716 4125
rect 1684 4044 1716 4076
rect 1684 3995 1716 3996
rect 1684 3965 1685 3995
rect 1685 3965 1715 3995
rect 1715 3965 1716 3995
rect 1684 3964 1716 3965
rect 1764 4155 1796 4156
rect 1764 4125 1765 4155
rect 1765 4125 1795 4155
rect 1795 4125 1796 4155
rect 1764 4124 1796 4125
rect 1764 4044 1796 4076
rect 1764 3995 1796 3996
rect 1764 3965 1765 3995
rect 1765 3965 1795 3995
rect 1795 3965 1796 3995
rect 1764 3964 1796 3965
rect 1844 4155 1876 4156
rect 1844 4125 1845 4155
rect 1845 4125 1875 4155
rect 1875 4125 1876 4155
rect 1844 4124 1876 4125
rect 1844 4044 1876 4076
rect 1844 3995 1876 3996
rect 1844 3965 1845 3995
rect 1845 3965 1875 3995
rect 1875 3965 1876 3995
rect 1844 3964 1876 3965
rect 1924 4155 1956 4156
rect 1924 4125 1925 4155
rect 1925 4125 1955 4155
rect 1955 4125 1956 4155
rect 1924 4124 1956 4125
rect 1924 4044 1956 4076
rect 1924 3995 1956 3996
rect 1924 3965 1925 3995
rect 1925 3965 1955 3995
rect 1955 3965 1956 3995
rect 1924 3964 1956 3965
rect 2004 4155 2036 4156
rect 2004 4125 2005 4155
rect 2005 4125 2035 4155
rect 2035 4125 2036 4155
rect 2004 4124 2036 4125
rect 2004 4044 2036 4076
rect 2004 3995 2036 3996
rect 2004 3965 2005 3995
rect 2005 3965 2035 3995
rect 2035 3965 2036 3995
rect 2004 3964 2036 3965
rect 2084 4155 2116 4156
rect 2084 4125 2085 4155
rect 2085 4125 2115 4155
rect 2115 4125 2116 4155
rect 2084 4124 2116 4125
rect 2084 4044 2116 4076
rect 2084 3995 2116 3996
rect 2084 3965 2085 3995
rect 2085 3965 2115 3995
rect 2115 3965 2116 3995
rect 2084 3964 2116 3965
rect 2164 4155 2196 4156
rect 2164 4125 2165 4155
rect 2165 4125 2195 4155
rect 2195 4125 2196 4155
rect 2164 4124 2196 4125
rect 2164 4044 2196 4076
rect 2164 3995 2196 3996
rect 2164 3965 2165 3995
rect 2165 3965 2195 3995
rect 2195 3965 2196 3995
rect 2164 3964 2196 3965
rect 2244 4155 2276 4156
rect 2244 4125 2245 4155
rect 2245 4125 2275 4155
rect 2275 4125 2276 4155
rect 2244 4124 2276 4125
rect 2244 4044 2276 4076
rect 2244 3995 2276 3996
rect 2244 3965 2245 3995
rect 2245 3965 2275 3995
rect 2275 3965 2276 3995
rect 2244 3964 2276 3965
rect 2324 4155 2356 4156
rect 2324 4125 2325 4155
rect 2325 4125 2355 4155
rect 2355 4125 2356 4155
rect 2324 4124 2356 4125
rect 2324 4044 2356 4076
rect 2324 3995 2356 3996
rect 2324 3965 2325 3995
rect 2325 3965 2355 3995
rect 2355 3965 2356 3995
rect 2324 3964 2356 3965
rect 2404 4155 2436 4156
rect 2404 4125 2405 4155
rect 2405 4125 2435 4155
rect 2435 4125 2436 4155
rect 2404 4124 2436 4125
rect 2404 4044 2436 4076
rect 2404 3995 2436 3996
rect 2404 3965 2405 3995
rect 2405 3965 2435 3995
rect 2435 3965 2436 3995
rect 2404 3964 2436 3965
rect 2484 4155 2516 4156
rect 2484 4125 2485 4155
rect 2485 4125 2515 4155
rect 2515 4125 2516 4155
rect 2484 4124 2516 4125
rect 2484 4044 2516 4076
rect 2484 3995 2516 3996
rect 2484 3965 2485 3995
rect 2485 3965 2515 3995
rect 2515 3965 2516 3995
rect 2484 3964 2516 3965
rect 2644 4155 2676 4156
rect 2644 4125 2645 4155
rect 2645 4125 2675 4155
rect 2675 4125 2676 4155
rect 2644 4124 2676 4125
rect 2644 4044 2676 4076
rect 2644 3995 2676 3996
rect 2644 3965 2645 3995
rect 2645 3965 2675 3995
rect 2675 3965 2676 3995
rect 2644 3964 2676 3965
rect 2724 4155 2756 4156
rect 2724 4125 2725 4155
rect 2725 4125 2755 4155
rect 2755 4125 2756 4155
rect 2724 4124 2756 4125
rect 2724 4044 2756 4076
rect 2724 3995 2756 3996
rect 2724 3965 2725 3995
rect 2725 3965 2755 3995
rect 2755 3965 2756 3995
rect 2724 3964 2756 3965
rect 2804 4155 2836 4156
rect 2804 4125 2805 4155
rect 2805 4125 2835 4155
rect 2835 4125 2836 4155
rect 2804 4124 2836 4125
rect 2804 4044 2836 4076
rect 2804 3995 2836 3996
rect 2804 3965 2805 3995
rect 2805 3965 2835 3995
rect 2835 3965 2836 3995
rect 2804 3964 2836 3965
rect 2884 4155 2916 4156
rect 2884 4125 2885 4155
rect 2885 4125 2915 4155
rect 2915 4125 2916 4155
rect 2884 4124 2916 4125
rect 2884 4044 2916 4076
rect 2884 3995 2916 3996
rect 2884 3965 2885 3995
rect 2885 3965 2915 3995
rect 2915 3965 2916 3995
rect 2884 3964 2916 3965
rect 2964 4155 2996 4156
rect 2964 4125 2965 4155
rect 2965 4125 2995 4155
rect 2995 4125 2996 4155
rect 2964 4124 2996 4125
rect 2964 4044 2996 4076
rect 2964 3995 2996 3996
rect 2964 3965 2965 3995
rect 2965 3965 2995 3995
rect 2995 3965 2996 3995
rect 2964 3964 2996 3965
rect 3044 4155 3076 4156
rect 3044 4125 3045 4155
rect 3045 4125 3075 4155
rect 3075 4125 3076 4155
rect 3044 4124 3076 4125
rect 3044 4044 3076 4076
rect 3044 3995 3076 3996
rect 3044 3965 3045 3995
rect 3045 3965 3075 3995
rect 3075 3965 3076 3995
rect 3044 3964 3076 3965
rect 3124 4155 3156 4156
rect 3124 4125 3125 4155
rect 3125 4125 3155 4155
rect 3155 4125 3156 4155
rect 3124 4124 3156 4125
rect 3124 4044 3156 4076
rect 3124 3995 3156 3996
rect 3124 3965 3125 3995
rect 3125 3965 3155 3995
rect 3155 3965 3156 3995
rect 3124 3964 3156 3965
rect 3204 4155 3236 4156
rect 3204 4125 3205 4155
rect 3205 4125 3235 4155
rect 3235 4125 3236 4155
rect 3204 4124 3236 4125
rect 3204 4044 3236 4076
rect 3204 3995 3236 3996
rect 3204 3965 3205 3995
rect 3205 3965 3235 3995
rect 3235 3965 3236 3995
rect 3204 3964 3236 3965
rect 3284 4155 3316 4156
rect 3284 4125 3285 4155
rect 3285 4125 3315 4155
rect 3315 4125 3316 4155
rect 3284 4124 3316 4125
rect 3284 4044 3316 4076
rect 3284 3995 3316 3996
rect 3284 3965 3285 3995
rect 3285 3965 3315 3995
rect 3315 3965 3316 3995
rect 3284 3964 3316 3965
rect 3364 4155 3396 4156
rect 3364 4125 3365 4155
rect 3365 4125 3395 4155
rect 3395 4125 3396 4155
rect 3364 4124 3396 4125
rect 3364 4044 3396 4076
rect 3364 3995 3396 3996
rect 3364 3965 3365 3995
rect 3365 3965 3395 3995
rect 3395 3965 3396 3995
rect 3364 3964 3396 3965
rect 3444 4155 3476 4156
rect 3444 4125 3445 4155
rect 3445 4125 3475 4155
rect 3475 4125 3476 4155
rect 3444 4124 3476 4125
rect 3444 4044 3476 4076
rect 3444 3995 3476 3996
rect 3444 3965 3445 3995
rect 3445 3965 3475 3995
rect 3475 3965 3476 3995
rect 3444 3964 3476 3965
rect 3604 4155 3636 4156
rect 3604 4125 3605 4155
rect 3605 4125 3635 4155
rect 3635 4125 3636 4155
rect 3604 4124 3636 4125
rect 3604 4044 3636 4076
rect 3604 3995 3636 3996
rect 3604 3965 3605 3995
rect 3605 3965 3635 3995
rect 3635 3965 3636 3995
rect 3604 3964 3636 3965
rect 3684 4155 3716 4156
rect 3684 4125 3685 4155
rect 3685 4125 3715 4155
rect 3715 4125 3716 4155
rect 3684 4124 3716 4125
rect 3684 4044 3716 4076
rect 3684 3995 3716 3996
rect 3684 3965 3685 3995
rect 3685 3965 3715 3995
rect 3715 3965 3716 3995
rect 3684 3964 3716 3965
rect 3764 4155 3796 4156
rect 3764 4125 3765 4155
rect 3765 4125 3795 4155
rect 3795 4125 3796 4155
rect 3764 4124 3796 4125
rect 3764 4044 3796 4076
rect 3764 3995 3796 3996
rect 3764 3965 3765 3995
rect 3765 3965 3795 3995
rect 3795 3965 3796 3995
rect 3764 3964 3796 3965
rect 3844 4155 3876 4156
rect 3844 4125 3845 4155
rect 3845 4125 3875 4155
rect 3875 4125 3876 4155
rect 3844 4124 3876 4125
rect 3844 4044 3876 4076
rect 3844 3995 3876 3996
rect 3844 3965 3845 3995
rect 3845 3965 3875 3995
rect 3875 3965 3876 3995
rect 3844 3964 3876 3965
rect 3924 4155 3956 4156
rect 3924 4125 3925 4155
rect 3925 4125 3955 4155
rect 3955 4125 3956 4155
rect 3924 4124 3956 4125
rect 3924 4044 3956 4076
rect 3924 3995 3956 3996
rect 3924 3965 3925 3995
rect 3925 3965 3955 3995
rect 3955 3965 3956 3995
rect 3924 3964 3956 3965
rect 4004 4155 4036 4156
rect 4004 4125 4005 4155
rect 4005 4125 4035 4155
rect 4035 4125 4036 4155
rect 4004 4124 4036 4125
rect 4004 4044 4036 4076
rect 4004 3995 4036 3996
rect 4004 3965 4005 3995
rect 4005 3965 4035 3995
rect 4035 3965 4036 3995
rect 4004 3964 4036 3965
rect 4084 4155 4116 4156
rect 4084 4125 4085 4155
rect 4085 4125 4115 4155
rect 4115 4125 4116 4155
rect 4084 4124 4116 4125
rect 4084 4044 4116 4076
rect 4084 3995 4116 3996
rect 4084 3965 4085 3995
rect 4085 3965 4115 3995
rect 4115 3965 4116 3995
rect 4084 3964 4116 3965
rect 164 3850 196 3851
rect 164 3770 165 3850
rect 165 3770 195 3850
rect 195 3770 196 3850
rect 164 3769 196 3770
rect 164 3550 196 3551
rect 164 3470 165 3550
rect 165 3470 195 3550
rect 195 3470 196 3550
rect 164 3469 196 3470
rect 84 3355 116 3356
rect 84 3325 85 3355
rect 85 3325 115 3355
rect 115 3325 116 3355
rect 84 3324 116 3325
rect 84 3244 116 3276
rect 84 3195 116 3196
rect 84 3165 85 3195
rect 85 3165 115 3195
rect 115 3165 116 3195
rect 84 3164 116 3165
rect 164 3355 196 3356
rect 164 3325 165 3355
rect 165 3325 195 3355
rect 195 3325 196 3355
rect 164 3324 196 3325
rect 164 3244 196 3276
rect 164 3195 196 3196
rect 164 3165 165 3195
rect 165 3165 195 3195
rect 195 3165 196 3195
rect 164 3164 196 3165
rect 244 3355 276 3356
rect 244 3325 245 3355
rect 245 3325 275 3355
rect 275 3325 276 3355
rect 244 3324 276 3325
rect 244 3244 276 3276
rect 244 3195 276 3196
rect 244 3165 245 3195
rect 245 3165 275 3195
rect 275 3165 276 3195
rect 244 3164 276 3165
rect 324 3355 356 3356
rect 324 3325 325 3355
rect 325 3325 355 3355
rect 355 3325 356 3355
rect 324 3324 356 3325
rect 324 3244 356 3276
rect 324 3195 356 3196
rect 324 3165 325 3195
rect 325 3165 355 3195
rect 355 3165 356 3195
rect 324 3164 356 3165
rect 404 3355 436 3356
rect 404 3325 405 3355
rect 405 3325 435 3355
rect 435 3325 436 3355
rect 404 3324 436 3325
rect 404 3244 436 3276
rect 404 3195 436 3196
rect 404 3165 405 3195
rect 405 3165 435 3195
rect 435 3165 436 3195
rect 404 3164 436 3165
rect 484 3355 516 3356
rect 484 3325 485 3355
rect 485 3325 515 3355
rect 515 3325 516 3355
rect 484 3324 516 3325
rect 484 3244 516 3276
rect 484 3195 516 3196
rect 484 3165 485 3195
rect 485 3165 515 3195
rect 515 3165 516 3195
rect 484 3164 516 3165
rect 564 3355 596 3356
rect 564 3325 565 3355
rect 565 3325 595 3355
rect 595 3325 596 3355
rect 564 3324 596 3325
rect 564 3244 596 3276
rect 564 3195 596 3196
rect 564 3165 565 3195
rect 565 3165 595 3195
rect 595 3165 596 3195
rect 564 3164 596 3165
rect 724 3355 756 3356
rect 724 3325 725 3355
rect 725 3325 755 3355
rect 755 3325 756 3355
rect 724 3324 756 3325
rect 724 3244 756 3276
rect 724 3195 756 3196
rect 724 3165 725 3195
rect 725 3165 755 3195
rect 755 3165 756 3195
rect 724 3164 756 3165
rect 804 3355 836 3356
rect 804 3325 805 3355
rect 805 3325 835 3355
rect 835 3325 836 3355
rect 804 3324 836 3325
rect 804 3244 836 3276
rect 804 3195 836 3196
rect 804 3165 805 3195
rect 805 3165 835 3195
rect 835 3165 836 3195
rect 804 3164 836 3165
rect 884 3355 916 3356
rect 884 3325 885 3355
rect 885 3325 915 3355
rect 915 3325 916 3355
rect 884 3324 916 3325
rect 884 3244 916 3276
rect 884 3195 916 3196
rect 884 3165 885 3195
rect 885 3165 915 3195
rect 915 3165 916 3195
rect 884 3164 916 3165
rect 964 3355 996 3356
rect 964 3325 965 3355
rect 965 3325 995 3355
rect 995 3325 996 3355
rect 964 3324 996 3325
rect 964 3244 996 3276
rect 964 3195 996 3196
rect 964 3165 965 3195
rect 965 3165 995 3195
rect 995 3165 996 3195
rect 964 3164 996 3165
rect 1044 3355 1076 3356
rect 1044 3325 1045 3355
rect 1045 3325 1075 3355
rect 1075 3325 1076 3355
rect 1044 3324 1076 3325
rect 1044 3244 1076 3276
rect 1044 3195 1076 3196
rect 1044 3165 1045 3195
rect 1045 3165 1075 3195
rect 1075 3165 1076 3195
rect 1044 3164 1076 3165
rect 1124 3355 1156 3356
rect 1124 3325 1125 3355
rect 1125 3325 1155 3355
rect 1155 3325 1156 3355
rect 1124 3324 1156 3325
rect 1124 3244 1156 3276
rect 1124 3195 1156 3196
rect 1124 3165 1125 3195
rect 1125 3165 1155 3195
rect 1155 3165 1156 3195
rect 1124 3164 1156 3165
rect 1204 3355 1236 3356
rect 1204 3325 1205 3355
rect 1205 3325 1235 3355
rect 1235 3325 1236 3355
rect 1204 3324 1236 3325
rect 1204 3244 1236 3276
rect 1204 3195 1236 3196
rect 1204 3165 1205 3195
rect 1205 3165 1235 3195
rect 1235 3165 1236 3195
rect 1204 3164 1236 3165
rect 1284 3355 1316 3356
rect 1284 3325 1285 3355
rect 1285 3325 1315 3355
rect 1315 3325 1316 3355
rect 1284 3324 1316 3325
rect 1284 3244 1316 3276
rect 1284 3195 1316 3196
rect 1284 3165 1285 3195
rect 1285 3165 1315 3195
rect 1315 3165 1316 3195
rect 1284 3164 1316 3165
rect 1364 3355 1396 3356
rect 1364 3325 1365 3355
rect 1365 3325 1395 3355
rect 1395 3325 1396 3355
rect 1364 3324 1396 3325
rect 1364 3244 1396 3276
rect 1364 3195 1396 3196
rect 1364 3165 1365 3195
rect 1365 3165 1395 3195
rect 1395 3165 1396 3195
rect 1364 3164 1396 3165
rect 1444 3355 1476 3356
rect 1444 3325 1445 3355
rect 1445 3325 1475 3355
rect 1475 3325 1476 3355
rect 1444 3324 1476 3325
rect 1444 3244 1476 3276
rect 1444 3195 1476 3196
rect 1444 3165 1445 3195
rect 1445 3165 1475 3195
rect 1475 3165 1476 3195
rect 1444 3164 1476 3165
rect 1524 3355 1556 3356
rect 1524 3325 1525 3355
rect 1525 3325 1555 3355
rect 1555 3325 1556 3355
rect 1524 3324 1556 3325
rect 1524 3244 1556 3276
rect 1524 3195 1556 3196
rect 1524 3165 1525 3195
rect 1525 3165 1555 3195
rect 1555 3165 1556 3195
rect 1524 3164 1556 3165
rect 1684 3355 1716 3356
rect 1684 3325 1685 3355
rect 1685 3325 1715 3355
rect 1715 3325 1716 3355
rect 1684 3324 1716 3325
rect 1684 3244 1716 3276
rect 1684 3195 1716 3196
rect 1684 3165 1685 3195
rect 1685 3165 1715 3195
rect 1715 3165 1716 3195
rect 1684 3164 1716 3165
rect 1764 3355 1796 3356
rect 1764 3325 1765 3355
rect 1765 3325 1795 3355
rect 1795 3325 1796 3355
rect 1764 3324 1796 3325
rect 1764 3244 1796 3276
rect 1764 3195 1796 3196
rect 1764 3165 1765 3195
rect 1765 3165 1795 3195
rect 1795 3165 1796 3195
rect 1764 3164 1796 3165
rect 1844 3355 1876 3356
rect 1844 3325 1845 3355
rect 1845 3325 1875 3355
rect 1875 3325 1876 3355
rect 1844 3324 1876 3325
rect 1844 3244 1876 3276
rect 1844 3195 1876 3196
rect 1844 3165 1845 3195
rect 1845 3165 1875 3195
rect 1875 3165 1876 3195
rect 1844 3164 1876 3165
rect 1924 3355 1956 3356
rect 1924 3325 1925 3355
rect 1925 3325 1955 3355
rect 1955 3325 1956 3355
rect 1924 3324 1956 3325
rect 1924 3244 1956 3276
rect 1924 3195 1956 3196
rect 1924 3165 1925 3195
rect 1925 3165 1955 3195
rect 1955 3165 1956 3195
rect 1924 3164 1956 3165
rect 2004 3355 2036 3356
rect 2004 3325 2005 3355
rect 2005 3325 2035 3355
rect 2035 3325 2036 3355
rect 2004 3324 2036 3325
rect 2004 3244 2036 3276
rect 2004 3195 2036 3196
rect 2004 3165 2005 3195
rect 2005 3165 2035 3195
rect 2035 3165 2036 3195
rect 2004 3164 2036 3165
rect 2084 3355 2116 3356
rect 2084 3325 2085 3355
rect 2085 3325 2115 3355
rect 2115 3325 2116 3355
rect 2084 3324 2116 3325
rect 2084 3244 2116 3276
rect 2084 3195 2116 3196
rect 2084 3165 2085 3195
rect 2085 3165 2115 3195
rect 2115 3165 2116 3195
rect 2084 3164 2116 3165
rect 2164 3355 2196 3356
rect 2164 3325 2165 3355
rect 2165 3325 2195 3355
rect 2195 3325 2196 3355
rect 2164 3324 2196 3325
rect 2164 3244 2196 3276
rect 2164 3195 2196 3196
rect 2164 3165 2165 3195
rect 2165 3165 2195 3195
rect 2195 3165 2196 3195
rect 2164 3164 2196 3165
rect 2244 3355 2276 3356
rect 2244 3325 2245 3355
rect 2245 3325 2275 3355
rect 2275 3325 2276 3355
rect 2244 3324 2276 3325
rect 2244 3244 2276 3276
rect 2244 3195 2276 3196
rect 2244 3165 2245 3195
rect 2245 3165 2275 3195
rect 2275 3165 2276 3195
rect 2244 3164 2276 3165
rect 2324 3355 2356 3356
rect 2324 3325 2325 3355
rect 2325 3325 2355 3355
rect 2355 3325 2356 3355
rect 2324 3324 2356 3325
rect 2324 3244 2356 3276
rect 2324 3195 2356 3196
rect 2324 3165 2325 3195
rect 2325 3165 2355 3195
rect 2355 3165 2356 3195
rect 2324 3164 2356 3165
rect 2404 3355 2436 3356
rect 2404 3325 2405 3355
rect 2405 3325 2435 3355
rect 2435 3325 2436 3355
rect 2404 3324 2436 3325
rect 2404 3244 2436 3276
rect 2404 3195 2436 3196
rect 2404 3165 2405 3195
rect 2405 3165 2435 3195
rect 2435 3165 2436 3195
rect 2404 3164 2436 3165
rect 2484 3355 2516 3356
rect 2484 3325 2485 3355
rect 2485 3325 2515 3355
rect 2515 3325 2516 3355
rect 2484 3324 2516 3325
rect 2484 3244 2516 3276
rect 2484 3195 2516 3196
rect 2484 3165 2485 3195
rect 2485 3165 2515 3195
rect 2515 3165 2516 3195
rect 2484 3164 2516 3165
rect 2644 3355 2676 3356
rect 2644 3325 2645 3355
rect 2645 3325 2675 3355
rect 2675 3325 2676 3355
rect 2644 3324 2676 3325
rect 2644 3244 2676 3276
rect 2644 3195 2676 3196
rect 2644 3165 2645 3195
rect 2645 3165 2675 3195
rect 2675 3165 2676 3195
rect 2644 3164 2676 3165
rect 2724 3355 2756 3356
rect 2724 3325 2725 3355
rect 2725 3325 2755 3355
rect 2755 3325 2756 3355
rect 2724 3324 2756 3325
rect 2724 3244 2756 3276
rect 2724 3195 2756 3196
rect 2724 3165 2725 3195
rect 2725 3165 2755 3195
rect 2755 3165 2756 3195
rect 2724 3164 2756 3165
rect 2804 3355 2836 3356
rect 2804 3325 2805 3355
rect 2805 3325 2835 3355
rect 2835 3325 2836 3355
rect 2804 3324 2836 3325
rect 2804 3244 2836 3276
rect 2804 3195 2836 3196
rect 2804 3165 2805 3195
rect 2805 3165 2835 3195
rect 2835 3165 2836 3195
rect 2804 3164 2836 3165
rect 2884 3355 2916 3356
rect 2884 3325 2885 3355
rect 2885 3325 2915 3355
rect 2915 3325 2916 3355
rect 2884 3324 2916 3325
rect 2884 3244 2916 3276
rect 2884 3195 2916 3196
rect 2884 3165 2885 3195
rect 2885 3165 2915 3195
rect 2915 3165 2916 3195
rect 2884 3164 2916 3165
rect 2964 3355 2996 3356
rect 2964 3325 2965 3355
rect 2965 3325 2995 3355
rect 2995 3325 2996 3355
rect 2964 3324 2996 3325
rect 2964 3244 2996 3276
rect 2964 3195 2996 3196
rect 2964 3165 2965 3195
rect 2965 3165 2995 3195
rect 2995 3165 2996 3195
rect 2964 3164 2996 3165
rect 3044 3355 3076 3356
rect 3044 3325 3045 3355
rect 3045 3325 3075 3355
rect 3075 3325 3076 3355
rect 3044 3324 3076 3325
rect 3044 3244 3076 3276
rect 3044 3195 3076 3196
rect 3044 3165 3045 3195
rect 3045 3165 3075 3195
rect 3075 3165 3076 3195
rect 3044 3164 3076 3165
rect 3124 3355 3156 3356
rect 3124 3325 3125 3355
rect 3125 3325 3155 3355
rect 3155 3325 3156 3355
rect 3124 3324 3156 3325
rect 3124 3244 3156 3276
rect 3124 3195 3156 3196
rect 3124 3165 3125 3195
rect 3125 3165 3155 3195
rect 3155 3165 3156 3195
rect 3124 3164 3156 3165
rect 3204 3355 3236 3356
rect 3204 3325 3205 3355
rect 3205 3325 3235 3355
rect 3235 3325 3236 3355
rect 3204 3324 3236 3325
rect 3204 3244 3236 3276
rect 3204 3195 3236 3196
rect 3204 3165 3205 3195
rect 3205 3165 3235 3195
rect 3235 3165 3236 3195
rect 3204 3164 3236 3165
rect 3284 3355 3316 3356
rect 3284 3325 3285 3355
rect 3285 3325 3315 3355
rect 3315 3325 3316 3355
rect 3284 3324 3316 3325
rect 3284 3244 3316 3276
rect 3284 3195 3316 3196
rect 3284 3165 3285 3195
rect 3285 3165 3315 3195
rect 3315 3165 3316 3195
rect 3284 3164 3316 3165
rect 3364 3355 3396 3356
rect 3364 3325 3365 3355
rect 3365 3325 3395 3355
rect 3395 3325 3396 3355
rect 3364 3324 3396 3325
rect 3364 3244 3396 3276
rect 3364 3195 3396 3196
rect 3364 3165 3365 3195
rect 3365 3165 3395 3195
rect 3395 3165 3396 3195
rect 3364 3164 3396 3165
rect 3444 3355 3476 3356
rect 3444 3325 3445 3355
rect 3445 3325 3475 3355
rect 3475 3325 3476 3355
rect 3444 3324 3476 3325
rect 3444 3244 3476 3276
rect 3444 3195 3476 3196
rect 3444 3165 3445 3195
rect 3445 3165 3475 3195
rect 3475 3165 3476 3195
rect 3444 3164 3476 3165
rect 3604 3355 3636 3356
rect 3604 3325 3605 3355
rect 3605 3325 3635 3355
rect 3635 3325 3636 3355
rect 3604 3324 3636 3325
rect 3604 3244 3636 3276
rect 3604 3195 3636 3196
rect 3604 3165 3605 3195
rect 3605 3165 3635 3195
rect 3635 3165 3636 3195
rect 3604 3164 3636 3165
rect 3684 3355 3716 3356
rect 3684 3325 3685 3355
rect 3685 3325 3715 3355
rect 3715 3325 3716 3355
rect 3684 3324 3716 3325
rect 3684 3244 3716 3276
rect 3684 3195 3716 3196
rect 3684 3165 3685 3195
rect 3685 3165 3715 3195
rect 3715 3165 3716 3195
rect 3684 3164 3716 3165
rect 3764 3355 3796 3356
rect 3764 3325 3765 3355
rect 3765 3325 3795 3355
rect 3795 3325 3796 3355
rect 3764 3324 3796 3325
rect 3764 3244 3796 3276
rect 3764 3195 3796 3196
rect 3764 3165 3765 3195
rect 3765 3165 3795 3195
rect 3795 3165 3796 3195
rect 3764 3164 3796 3165
rect 3844 3355 3876 3356
rect 3844 3325 3845 3355
rect 3845 3325 3875 3355
rect 3875 3325 3876 3355
rect 3844 3324 3876 3325
rect 3844 3244 3876 3276
rect 3844 3195 3876 3196
rect 3844 3165 3845 3195
rect 3845 3165 3875 3195
rect 3875 3165 3876 3195
rect 3844 3164 3876 3165
rect 3924 3355 3956 3356
rect 3924 3325 3925 3355
rect 3925 3325 3955 3355
rect 3955 3325 3956 3355
rect 3924 3324 3956 3325
rect 3924 3244 3956 3276
rect 3924 3195 3956 3196
rect 3924 3165 3925 3195
rect 3925 3165 3955 3195
rect 3955 3165 3956 3195
rect 3924 3164 3956 3165
rect 4084 3355 4116 3356
rect 4084 3325 4085 3355
rect 4085 3325 4115 3355
rect 4115 3325 4116 3355
rect 4084 3324 4116 3325
rect 4084 3244 4116 3276
rect 4084 3195 4116 3196
rect 4084 3165 4085 3195
rect 4085 3165 4115 3195
rect 4115 3165 4116 3195
rect 4084 3164 4116 3165
rect 84 3115 116 3116
rect 84 3085 85 3115
rect 85 3085 115 3115
rect 115 3085 116 3115
rect 84 3084 116 3085
rect 84 3004 116 3036
rect 84 2955 116 2956
rect 84 2925 85 2955
rect 85 2925 115 2955
rect 115 2925 116 2955
rect 84 2924 116 2925
rect 164 3115 196 3116
rect 164 3085 165 3115
rect 165 3085 195 3115
rect 195 3085 196 3115
rect 164 3084 196 3085
rect 164 3004 196 3036
rect 164 2955 196 2956
rect 164 2925 165 2955
rect 165 2925 195 2955
rect 195 2925 196 2955
rect 164 2924 196 2925
rect 244 3115 276 3116
rect 244 3085 245 3115
rect 245 3085 275 3115
rect 275 3085 276 3115
rect 244 3084 276 3085
rect 244 3004 276 3036
rect 244 2955 276 2956
rect 244 2925 245 2955
rect 245 2925 275 2955
rect 275 2925 276 2955
rect 244 2924 276 2925
rect 324 3115 356 3116
rect 324 3085 325 3115
rect 325 3085 355 3115
rect 355 3085 356 3115
rect 324 3084 356 3085
rect 324 3004 356 3036
rect 324 2955 356 2956
rect 324 2925 325 2955
rect 325 2925 355 2955
rect 355 2925 356 2955
rect 324 2924 356 2925
rect 404 3115 436 3116
rect 404 3085 405 3115
rect 405 3085 435 3115
rect 435 3085 436 3115
rect 404 3084 436 3085
rect 404 3004 436 3036
rect 404 2955 436 2956
rect 404 2925 405 2955
rect 405 2925 435 2955
rect 435 2925 436 2955
rect 404 2924 436 2925
rect 484 3115 516 3116
rect 484 3085 485 3115
rect 485 3085 515 3115
rect 515 3085 516 3115
rect 484 3084 516 3085
rect 484 3004 516 3036
rect 484 2955 516 2956
rect 484 2925 485 2955
rect 485 2925 515 2955
rect 515 2925 516 2955
rect 484 2924 516 2925
rect 564 3115 596 3116
rect 564 3085 565 3115
rect 565 3085 595 3115
rect 595 3085 596 3115
rect 564 3084 596 3085
rect 564 3004 596 3036
rect 564 2955 596 2956
rect 564 2925 565 2955
rect 565 2925 595 2955
rect 595 2925 596 2955
rect 564 2924 596 2925
rect 644 3115 676 3116
rect 644 3085 645 3115
rect 645 3085 675 3115
rect 675 3085 676 3115
rect 644 3084 676 3085
rect 644 3004 676 3036
rect 644 2955 676 2956
rect 644 2925 645 2955
rect 645 2925 675 2955
rect 675 2925 676 2955
rect 644 2924 676 2925
rect 724 3115 756 3116
rect 724 3085 725 3115
rect 725 3085 755 3115
rect 755 3085 756 3115
rect 724 3084 756 3085
rect 724 3004 756 3036
rect 724 2955 756 2956
rect 724 2925 725 2955
rect 725 2925 755 2955
rect 755 2925 756 2955
rect 724 2924 756 2925
rect 804 3115 836 3116
rect 804 3085 805 3115
rect 805 3085 835 3115
rect 835 3085 836 3115
rect 804 3084 836 3085
rect 804 3004 836 3036
rect 804 2955 836 2956
rect 804 2925 805 2955
rect 805 2925 835 2955
rect 835 2925 836 2955
rect 804 2924 836 2925
rect 884 3115 916 3116
rect 884 3085 885 3115
rect 885 3085 915 3115
rect 915 3085 916 3115
rect 884 3084 916 3085
rect 884 3004 916 3036
rect 884 2955 916 2956
rect 884 2925 885 2955
rect 885 2925 915 2955
rect 915 2925 916 2955
rect 884 2924 916 2925
rect 964 3115 996 3116
rect 964 3085 965 3115
rect 965 3085 995 3115
rect 995 3085 996 3115
rect 964 3084 996 3085
rect 964 3004 996 3036
rect 964 2955 996 2956
rect 964 2925 965 2955
rect 965 2925 995 2955
rect 995 2925 996 2955
rect 964 2924 996 2925
rect 1044 3115 1076 3116
rect 1044 3085 1045 3115
rect 1045 3085 1075 3115
rect 1075 3085 1076 3115
rect 1044 3084 1076 3085
rect 1044 3004 1076 3036
rect 1044 2955 1076 2956
rect 1044 2925 1045 2955
rect 1045 2925 1075 2955
rect 1075 2925 1076 2955
rect 1044 2924 1076 2925
rect 1124 3115 1156 3116
rect 1124 3085 1125 3115
rect 1125 3085 1155 3115
rect 1155 3085 1156 3115
rect 1124 3084 1156 3085
rect 1124 3004 1156 3036
rect 1124 2955 1156 2956
rect 1124 2925 1125 2955
rect 1125 2925 1155 2955
rect 1155 2925 1156 2955
rect 1124 2924 1156 2925
rect 1204 3115 1236 3116
rect 1204 3085 1205 3115
rect 1205 3085 1235 3115
rect 1235 3085 1236 3115
rect 1204 3084 1236 3085
rect 1204 3004 1236 3036
rect 1204 2955 1236 2956
rect 1204 2925 1205 2955
rect 1205 2925 1235 2955
rect 1235 2925 1236 2955
rect 1204 2924 1236 2925
rect 1284 3115 1316 3116
rect 1284 3085 1285 3115
rect 1285 3085 1315 3115
rect 1315 3085 1316 3115
rect 1284 3084 1316 3085
rect 1284 3004 1316 3036
rect 1284 2955 1316 2956
rect 1284 2925 1285 2955
rect 1285 2925 1315 2955
rect 1315 2925 1316 2955
rect 1284 2924 1316 2925
rect 1364 3115 1396 3116
rect 1364 3085 1365 3115
rect 1365 3085 1395 3115
rect 1395 3085 1396 3115
rect 1364 3084 1396 3085
rect 1364 3004 1396 3036
rect 1364 2955 1396 2956
rect 1364 2925 1365 2955
rect 1365 2925 1395 2955
rect 1395 2925 1396 2955
rect 1364 2924 1396 2925
rect 1444 3115 1476 3116
rect 1444 3085 1445 3115
rect 1445 3085 1475 3115
rect 1475 3085 1476 3115
rect 1444 3084 1476 3085
rect 1444 3004 1476 3036
rect 1444 2955 1476 2956
rect 1444 2925 1445 2955
rect 1445 2925 1475 2955
rect 1475 2925 1476 2955
rect 1444 2924 1476 2925
rect 1524 3115 1556 3116
rect 1524 3085 1525 3115
rect 1525 3085 1555 3115
rect 1555 3085 1556 3115
rect 1524 3084 1556 3085
rect 1524 3004 1556 3036
rect 1524 2955 1556 2956
rect 1524 2925 1525 2955
rect 1525 2925 1555 2955
rect 1555 2925 1556 2955
rect 1524 2924 1556 2925
rect 1604 3115 1636 3116
rect 1604 3085 1605 3115
rect 1605 3085 1635 3115
rect 1635 3085 1636 3115
rect 1604 3084 1636 3085
rect 1604 3004 1636 3036
rect 1604 2955 1636 2956
rect 1604 2925 1605 2955
rect 1605 2925 1635 2955
rect 1635 2925 1636 2955
rect 1604 2924 1636 2925
rect 1684 3115 1716 3116
rect 1684 3085 1685 3115
rect 1685 3085 1715 3115
rect 1715 3085 1716 3115
rect 1684 3084 1716 3085
rect 1684 3004 1716 3036
rect 1684 2955 1716 2956
rect 1684 2925 1685 2955
rect 1685 2925 1715 2955
rect 1715 2925 1716 2955
rect 1684 2924 1716 2925
rect 1764 3115 1796 3116
rect 1764 3085 1765 3115
rect 1765 3085 1795 3115
rect 1795 3085 1796 3115
rect 1764 3084 1796 3085
rect 1764 3004 1796 3036
rect 1764 2955 1796 2956
rect 1764 2925 1765 2955
rect 1765 2925 1795 2955
rect 1795 2925 1796 2955
rect 1764 2924 1796 2925
rect 1844 3115 1876 3116
rect 1844 3085 1845 3115
rect 1845 3085 1875 3115
rect 1875 3085 1876 3115
rect 1844 3084 1876 3085
rect 1844 3004 1876 3036
rect 1844 2955 1876 2956
rect 1844 2925 1845 2955
rect 1845 2925 1875 2955
rect 1875 2925 1876 2955
rect 1844 2924 1876 2925
rect 1924 3115 1956 3116
rect 1924 3085 1925 3115
rect 1925 3085 1955 3115
rect 1955 3085 1956 3115
rect 1924 3084 1956 3085
rect 1924 3004 1956 3036
rect 1924 2955 1956 2956
rect 1924 2925 1925 2955
rect 1925 2925 1955 2955
rect 1955 2925 1956 2955
rect 1924 2924 1956 2925
rect 2004 3115 2036 3116
rect 2004 3085 2005 3115
rect 2005 3085 2035 3115
rect 2035 3085 2036 3115
rect 2004 3084 2036 3085
rect 2004 3004 2036 3036
rect 2004 2955 2036 2956
rect 2004 2925 2005 2955
rect 2005 2925 2035 2955
rect 2035 2925 2036 2955
rect 2004 2924 2036 2925
rect 2084 3115 2116 3116
rect 2084 3085 2085 3115
rect 2085 3085 2115 3115
rect 2115 3085 2116 3115
rect 2084 3084 2116 3085
rect 2084 3004 2116 3036
rect 2084 2955 2116 2956
rect 2084 2925 2085 2955
rect 2085 2925 2115 2955
rect 2115 2925 2116 2955
rect 2084 2924 2116 2925
rect 2164 3115 2196 3116
rect 2164 3085 2165 3115
rect 2165 3085 2195 3115
rect 2195 3085 2196 3115
rect 2164 3084 2196 3085
rect 2164 3004 2196 3036
rect 2164 2955 2196 2956
rect 2164 2925 2165 2955
rect 2165 2925 2195 2955
rect 2195 2925 2196 2955
rect 2164 2924 2196 2925
rect 2244 3115 2276 3116
rect 2244 3085 2245 3115
rect 2245 3085 2275 3115
rect 2275 3085 2276 3115
rect 2244 3084 2276 3085
rect 2244 3004 2276 3036
rect 2244 2955 2276 2956
rect 2244 2925 2245 2955
rect 2245 2925 2275 2955
rect 2275 2925 2276 2955
rect 2244 2924 2276 2925
rect 2324 3115 2356 3116
rect 2324 3085 2325 3115
rect 2325 3085 2355 3115
rect 2355 3085 2356 3115
rect 2324 3084 2356 3085
rect 2324 3004 2356 3036
rect 2324 2955 2356 2956
rect 2324 2925 2325 2955
rect 2325 2925 2355 2955
rect 2355 2925 2356 2955
rect 2324 2924 2356 2925
rect 2404 3115 2436 3116
rect 2404 3085 2405 3115
rect 2405 3085 2435 3115
rect 2435 3085 2436 3115
rect 2404 3084 2436 3085
rect 2404 3004 2436 3036
rect 2404 2955 2436 2956
rect 2404 2925 2405 2955
rect 2405 2925 2435 2955
rect 2435 2925 2436 2955
rect 2404 2924 2436 2925
rect 2484 3115 2516 3116
rect 2484 3085 2485 3115
rect 2485 3085 2515 3115
rect 2515 3085 2516 3115
rect 2484 3084 2516 3085
rect 2484 3004 2516 3036
rect 2484 2955 2516 2956
rect 2484 2925 2485 2955
rect 2485 2925 2515 2955
rect 2515 2925 2516 2955
rect 2484 2924 2516 2925
rect 2564 3115 2596 3116
rect 2564 3085 2565 3115
rect 2565 3085 2595 3115
rect 2595 3085 2596 3115
rect 2564 3084 2596 3085
rect 2564 3004 2596 3036
rect 2564 2955 2596 2956
rect 2564 2925 2565 2955
rect 2565 2925 2595 2955
rect 2595 2925 2596 2955
rect 2564 2924 2596 2925
rect 2644 3115 2676 3116
rect 2644 3085 2645 3115
rect 2645 3085 2675 3115
rect 2675 3085 2676 3115
rect 2644 3084 2676 3085
rect 2644 3004 2676 3036
rect 2644 2955 2676 2956
rect 2644 2925 2645 2955
rect 2645 2925 2675 2955
rect 2675 2925 2676 2955
rect 2644 2924 2676 2925
rect 2724 3115 2756 3116
rect 2724 3085 2725 3115
rect 2725 3085 2755 3115
rect 2755 3085 2756 3115
rect 2724 3084 2756 3085
rect 2724 3004 2756 3036
rect 2724 2955 2756 2956
rect 2724 2925 2725 2955
rect 2725 2925 2755 2955
rect 2755 2925 2756 2955
rect 2724 2924 2756 2925
rect 2804 3115 2836 3116
rect 2804 3085 2805 3115
rect 2805 3085 2835 3115
rect 2835 3085 2836 3115
rect 2804 3084 2836 3085
rect 2804 3004 2836 3036
rect 2804 2955 2836 2956
rect 2804 2925 2805 2955
rect 2805 2925 2835 2955
rect 2835 2925 2836 2955
rect 2804 2924 2836 2925
rect 2884 3115 2916 3116
rect 2884 3085 2885 3115
rect 2885 3085 2915 3115
rect 2915 3085 2916 3115
rect 2884 3084 2916 3085
rect 2884 3004 2916 3036
rect 2884 2955 2916 2956
rect 2884 2925 2885 2955
rect 2885 2925 2915 2955
rect 2915 2925 2916 2955
rect 2884 2924 2916 2925
rect 2964 3115 2996 3116
rect 2964 3085 2965 3115
rect 2965 3085 2995 3115
rect 2995 3085 2996 3115
rect 2964 3084 2996 3085
rect 2964 3004 2996 3036
rect 2964 2955 2996 2956
rect 2964 2925 2965 2955
rect 2965 2925 2995 2955
rect 2995 2925 2996 2955
rect 2964 2924 2996 2925
rect 3044 3115 3076 3116
rect 3044 3085 3045 3115
rect 3045 3085 3075 3115
rect 3075 3085 3076 3115
rect 3044 3084 3076 3085
rect 3044 3004 3076 3036
rect 3044 2955 3076 2956
rect 3044 2925 3045 2955
rect 3045 2925 3075 2955
rect 3075 2925 3076 2955
rect 3044 2924 3076 2925
rect 3124 3115 3156 3116
rect 3124 3085 3125 3115
rect 3125 3085 3155 3115
rect 3155 3085 3156 3115
rect 3124 3084 3156 3085
rect 3124 3004 3156 3036
rect 3124 2955 3156 2956
rect 3124 2925 3125 2955
rect 3125 2925 3155 2955
rect 3155 2925 3156 2955
rect 3124 2924 3156 2925
rect 3204 3115 3236 3116
rect 3204 3085 3205 3115
rect 3205 3085 3235 3115
rect 3235 3085 3236 3115
rect 3204 3084 3236 3085
rect 3204 3004 3236 3036
rect 3204 2955 3236 2956
rect 3204 2925 3205 2955
rect 3205 2925 3235 2955
rect 3235 2925 3236 2955
rect 3204 2924 3236 2925
rect 3284 3115 3316 3116
rect 3284 3085 3285 3115
rect 3285 3085 3315 3115
rect 3315 3085 3316 3115
rect 3284 3084 3316 3085
rect 3284 3004 3316 3036
rect 3284 2955 3316 2956
rect 3284 2925 3285 2955
rect 3285 2925 3315 2955
rect 3315 2925 3316 2955
rect 3284 2924 3316 2925
rect 3364 3115 3396 3116
rect 3364 3085 3365 3115
rect 3365 3085 3395 3115
rect 3395 3085 3396 3115
rect 3364 3084 3396 3085
rect 3364 3004 3396 3036
rect 3364 2955 3396 2956
rect 3364 2925 3365 2955
rect 3365 2925 3395 2955
rect 3395 2925 3396 2955
rect 3364 2924 3396 2925
rect 3444 3115 3476 3116
rect 3444 3085 3445 3115
rect 3445 3085 3475 3115
rect 3475 3085 3476 3115
rect 3444 3084 3476 3085
rect 3444 3004 3476 3036
rect 3444 2955 3476 2956
rect 3444 2925 3445 2955
rect 3445 2925 3475 2955
rect 3475 2925 3476 2955
rect 3444 2924 3476 2925
rect 3524 3115 3556 3116
rect 3524 3085 3525 3115
rect 3525 3085 3555 3115
rect 3555 3085 3556 3115
rect 3524 3084 3556 3085
rect 3524 3004 3556 3036
rect 3524 2955 3556 2956
rect 3524 2925 3525 2955
rect 3525 2925 3555 2955
rect 3555 2925 3556 2955
rect 3524 2924 3556 2925
rect 3604 3115 3636 3116
rect 3604 3085 3605 3115
rect 3605 3085 3635 3115
rect 3635 3085 3636 3115
rect 3604 3084 3636 3085
rect 3604 3004 3636 3036
rect 3604 2955 3636 2956
rect 3604 2925 3605 2955
rect 3605 2925 3635 2955
rect 3635 2925 3636 2955
rect 3604 2924 3636 2925
rect 3684 3115 3716 3116
rect 3684 3085 3685 3115
rect 3685 3085 3715 3115
rect 3715 3085 3716 3115
rect 3684 3084 3716 3085
rect 3684 3004 3716 3036
rect 3684 2955 3716 2956
rect 3684 2925 3685 2955
rect 3685 2925 3715 2955
rect 3715 2925 3716 2955
rect 3684 2924 3716 2925
rect 3764 3115 3796 3116
rect 3764 3085 3765 3115
rect 3765 3085 3795 3115
rect 3795 3085 3796 3115
rect 3764 3084 3796 3085
rect 3764 3004 3796 3036
rect 3764 2955 3796 2956
rect 3764 2925 3765 2955
rect 3765 2925 3795 2955
rect 3795 2925 3796 2955
rect 3764 2924 3796 2925
rect 3844 3115 3876 3116
rect 3844 3085 3845 3115
rect 3845 3085 3875 3115
rect 3875 3085 3876 3115
rect 3844 3084 3876 3085
rect 3844 3004 3876 3036
rect 3844 2955 3876 2956
rect 3844 2925 3845 2955
rect 3845 2925 3875 2955
rect 3875 2925 3876 2955
rect 3844 2924 3876 2925
rect 3924 3115 3956 3116
rect 3924 3085 3925 3115
rect 3925 3085 3955 3115
rect 3955 3085 3956 3115
rect 3924 3084 3956 3085
rect 3924 3004 3956 3036
rect 3924 2955 3956 2956
rect 3924 2925 3925 2955
rect 3925 2925 3955 2955
rect 3955 2925 3956 2955
rect 3924 2924 3956 2925
rect 4084 3115 4116 3116
rect 4084 3085 4085 3115
rect 4085 3085 4115 3115
rect 4115 3085 4116 3115
rect 4084 3084 4116 3085
rect 4084 3004 4116 3036
rect 4084 2955 4116 2956
rect 4084 2925 4085 2955
rect 4085 2925 4115 2955
rect 4115 2925 4116 2955
rect 4084 2924 4116 2925
rect 84 2875 116 2876
rect 84 2845 85 2875
rect 85 2845 115 2875
rect 115 2845 116 2875
rect 84 2844 116 2845
rect 84 2764 116 2796
rect 84 2715 116 2716
rect 84 2685 85 2715
rect 85 2685 115 2715
rect 115 2685 116 2715
rect 84 2684 116 2685
rect 164 2875 196 2876
rect 164 2845 165 2875
rect 165 2845 195 2875
rect 195 2845 196 2875
rect 164 2844 196 2845
rect 164 2764 196 2796
rect 164 2715 196 2716
rect 164 2685 165 2715
rect 165 2685 195 2715
rect 195 2685 196 2715
rect 164 2684 196 2685
rect 244 2875 276 2876
rect 244 2845 245 2875
rect 245 2845 275 2875
rect 275 2845 276 2875
rect 244 2844 276 2845
rect 244 2764 276 2796
rect 244 2715 276 2716
rect 244 2685 245 2715
rect 245 2685 275 2715
rect 275 2685 276 2715
rect 244 2684 276 2685
rect 324 2875 356 2876
rect 324 2845 325 2875
rect 325 2845 355 2875
rect 355 2845 356 2875
rect 324 2844 356 2845
rect 324 2764 356 2796
rect 324 2715 356 2716
rect 324 2685 325 2715
rect 325 2685 355 2715
rect 355 2685 356 2715
rect 324 2684 356 2685
rect 404 2875 436 2876
rect 404 2845 405 2875
rect 405 2845 435 2875
rect 435 2845 436 2875
rect 404 2844 436 2845
rect 404 2764 436 2796
rect 404 2715 436 2716
rect 404 2685 405 2715
rect 405 2685 435 2715
rect 435 2685 436 2715
rect 404 2684 436 2685
rect 484 2875 516 2876
rect 484 2845 485 2875
rect 485 2845 515 2875
rect 515 2845 516 2875
rect 484 2844 516 2845
rect 484 2764 516 2796
rect 484 2715 516 2716
rect 484 2685 485 2715
rect 485 2685 515 2715
rect 515 2685 516 2715
rect 484 2684 516 2685
rect 564 2875 596 2876
rect 564 2845 565 2875
rect 565 2845 595 2875
rect 595 2845 596 2875
rect 564 2844 596 2845
rect 564 2764 596 2796
rect 564 2715 596 2716
rect 564 2685 565 2715
rect 565 2685 595 2715
rect 595 2685 596 2715
rect 564 2684 596 2685
rect 724 2875 756 2876
rect 724 2845 725 2875
rect 725 2845 755 2875
rect 755 2845 756 2875
rect 724 2844 756 2845
rect 724 2764 756 2796
rect 724 2715 756 2716
rect 724 2685 725 2715
rect 725 2685 755 2715
rect 755 2685 756 2715
rect 724 2684 756 2685
rect 804 2875 836 2876
rect 804 2845 805 2875
rect 805 2845 835 2875
rect 835 2845 836 2875
rect 804 2844 836 2845
rect 804 2764 836 2796
rect 804 2715 836 2716
rect 804 2685 805 2715
rect 805 2685 835 2715
rect 835 2685 836 2715
rect 804 2684 836 2685
rect 884 2875 916 2876
rect 884 2845 885 2875
rect 885 2845 915 2875
rect 915 2845 916 2875
rect 884 2844 916 2845
rect 884 2764 916 2796
rect 884 2715 916 2716
rect 884 2685 885 2715
rect 885 2685 915 2715
rect 915 2685 916 2715
rect 884 2684 916 2685
rect 964 2875 996 2876
rect 964 2845 965 2875
rect 965 2845 995 2875
rect 995 2845 996 2875
rect 964 2844 996 2845
rect 964 2764 996 2796
rect 964 2715 996 2716
rect 964 2685 965 2715
rect 965 2685 995 2715
rect 995 2685 996 2715
rect 964 2684 996 2685
rect 1044 2875 1076 2876
rect 1044 2845 1045 2875
rect 1045 2845 1075 2875
rect 1075 2845 1076 2875
rect 1044 2844 1076 2845
rect 1044 2764 1076 2796
rect 1044 2715 1076 2716
rect 1044 2685 1045 2715
rect 1045 2685 1075 2715
rect 1075 2685 1076 2715
rect 1044 2684 1076 2685
rect 1124 2875 1156 2876
rect 1124 2845 1125 2875
rect 1125 2845 1155 2875
rect 1155 2845 1156 2875
rect 1124 2844 1156 2845
rect 1124 2764 1156 2796
rect 1124 2715 1156 2716
rect 1124 2685 1125 2715
rect 1125 2685 1155 2715
rect 1155 2685 1156 2715
rect 1124 2684 1156 2685
rect 1204 2875 1236 2876
rect 1204 2845 1205 2875
rect 1205 2845 1235 2875
rect 1235 2845 1236 2875
rect 1204 2844 1236 2845
rect 1204 2764 1236 2796
rect 1204 2715 1236 2716
rect 1204 2685 1205 2715
rect 1205 2685 1235 2715
rect 1235 2685 1236 2715
rect 1204 2684 1236 2685
rect 1284 2875 1316 2876
rect 1284 2845 1285 2875
rect 1285 2845 1315 2875
rect 1315 2845 1316 2875
rect 1284 2844 1316 2845
rect 1284 2764 1316 2796
rect 1284 2715 1316 2716
rect 1284 2685 1285 2715
rect 1285 2685 1315 2715
rect 1315 2685 1316 2715
rect 1284 2684 1316 2685
rect 1364 2875 1396 2876
rect 1364 2845 1365 2875
rect 1365 2845 1395 2875
rect 1395 2845 1396 2875
rect 1364 2844 1396 2845
rect 1364 2764 1396 2796
rect 1364 2715 1396 2716
rect 1364 2685 1365 2715
rect 1365 2685 1395 2715
rect 1395 2685 1396 2715
rect 1364 2684 1396 2685
rect 1444 2875 1476 2876
rect 1444 2845 1445 2875
rect 1445 2845 1475 2875
rect 1475 2845 1476 2875
rect 1444 2844 1476 2845
rect 1444 2764 1476 2796
rect 1444 2715 1476 2716
rect 1444 2685 1445 2715
rect 1445 2685 1475 2715
rect 1475 2685 1476 2715
rect 1444 2684 1476 2685
rect 1524 2875 1556 2876
rect 1524 2845 1525 2875
rect 1525 2845 1555 2875
rect 1555 2845 1556 2875
rect 1524 2844 1556 2845
rect 1524 2764 1556 2796
rect 1524 2715 1556 2716
rect 1524 2685 1525 2715
rect 1525 2685 1555 2715
rect 1555 2685 1556 2715
rect 1524 2684 1556 2685
rect 1684 2875 1716 2876
rect 1684 2845 1685 2875
rect 1685 2845 1715 2875
rect 1715 2845 1716 2875
rect 1684 2844 1716 2845
rect 1684 2764 1716 2796
rect 1684 2715 1716 2716
rect 1684 2685 1685 2715
rect 1685 2685 1715 2715
rect 1715 2685 1716 2715
rect 1684 2684 1716 2685
rect 1764 2875 1796 2876
rect 1764 2845 1765 2875
rect 1765 2845 1795 2875
rect 1795 2845 1796 2875
rect 1764 2844 1796 2845
rect 1764 2764 1796 2796
rect 1764 2715 1796 2716
rect 1764 2685 1765 2715
rect 1765 2685 1795 2715
rect 1795 2685 1796 2715
rect 1764 2684 1796 2685
rect 1844 2875 1876 2876
rect 1844 2845 1845 2875
rect 1845 2845 1875 2875
rect 1875 2845 1876 2875
rect 1844 2844 1876 2845
rect 1844 2764 1876 2796
rect 1844 2715 1876 2716
rect 1844 2685 1845 2715
rect 1845 2685 1875 2715
rect 1875 2685 1876 2715
rect 1844 2684 1876 2685
rect 1924 2875 1956 2876
rect 1924 2845 1925 2875
rect 1925 2845 1955 2875
rect 1955 2845 1956 2875
rect 1924 2844 1956 2845
rect 1924 2764 1956 2796
rect 1924 2715 1956 2716
rect 1924 2685 1925 2715
rect 1925 2685 1955 2715
rect 1955 2685 1956 2715
rect 1924 2684 1956 2685
rect 2004 2875 2036 2876
rect 2004 2845 2005 2875
rect 2005 2845 2035 2875
rect 2035 2845 2036 2875
rect 2004 2844 2036 2845
rect 2004 2764 2036 2796
rect 2004 2715 2036 2716
rect 2004 2685 2005 2715
rect 2005 2685 2035 2715
rect 2035 2685 2036 2715
rect 2004 2684 2036 2685
rect 2084 2875 2116 2876
rect 2084 2845 2085 2875
rect 2085 2845 2115 2875
rect 2115 2845 2116 2875
rect 2084 2844 2116 2845
rect 2084 2764 2116 2796
rect 2084 2715 2116 2716
rect 2084 2685 2085 2715
rect 2085 2685 2115 2715
rect 2115 2685 2116 2715
rect 2084 2684 2116 2685
rect 2164 2875 2196 2876
rect 2164 2845 2165 2875
rect 2165 2845 2195 2875
rect 2195 2845 2196 2875
rect 2164 2844 2196 2845
rect 2164 2764 2196 2796
rect 2164 2715 2196 2716
rect 2164 2685 2165 2715
rect 2165 2685 2195 2715
rect 2195 2685 2196 2715
rect 2164 2684 2196 2685
rect 2244 2875 2276 2876
rect 2244 2845 2245 2875
rect 2245 2845 2275 2875
rect 2275 2845 2276 2875
rect 2244 2844 2276 2845
rect 2244 2764 2276 2796
rect 2244 2715 2276 2716
rect 2244 2685 2245 2715
rect 2245 2685 2275 2715
rect 2275 2685 2276 2715
rect 2244 2684 2276 2685
rect 2324 2875 2356 2876
rect 2324 2845 2325 2875
rect 2325 2845 2355 2875
rect 2355 2845 2356 2875
rect 2324 2844 2356 2845
rect 2324 2764 2356 2796
rect 2324 2715 2356 2716
rect 2324 2685 2325 2715
rect 2325 2685 2355 2715
rect 2355 2685 2356 2715
rect 2324 2684 2356 2685
rect 2404 2875 2436 2876
rect 2404 2845 2405 2875
rect 2405 2845 2435 2875
rect 2435 2845 2436 2875
rect 2404 2844 2436 2845
rect 2404 2764 2436 2796
rect 2404 2715 2436 2716
rect 2404 2685 2405 2715
rect 2405 2685 2435 2715
rect 2435 2685 2436 2715
rect 2404 2684 2436 2685
rect 2484 2875 2516 2876
rect 2484 2845 2485 2875
rect 2485 2845 2515 2875
rect 2515 2845 2516 2875
rect 2484 2844 2516 2845
rect 2484 2764 2516 2796
rect 2484 2715 2516 2716
rect 2484 2685 2485 2715
rect 2485 2685 2515 2715
rect 2515 2685 2516 2715
rect 2484 2684 2516 2685
rect 2644 2875 2676 2876
rect 2644 2845 2645 2875
rect 2645 2845 2675 2875
rect 2675 2845 2676 2875
rect 2644 2844 2676 2845
rect 2644 2764 2676 2796
rect 2644 2715 2676 2716
rect 2644 2685 2645 2715
rect 2645 2685 2675 2715
rect 2675 2685 2676 2715
rect 2644 2684 2676 2685
rect 2724 2875 2756 2876
rect 2724 2845 2725 2875
rect 2725 2845 2755 2875
rect 2755 2845 2756 2875
rect 2724 2844 2756 2845
rect 2724 2764 2756 2796
rect 2724 2715 2756 2716
rect 2724 2685 2725 2715
rect 2725 2685 2755 2715
rect 2755 2685 2756 2715
rect 2724 2684 2756 2685
rect 2804 2875 2836 2876
rect 2804 2845 2805 2875
rect 2805 2845 2835 2875
rect 2835 2845 2836 2875
rect 2804 2844 2836 2845
rect 2804 2764 2836 2796
rect 2804 2715 2836 2716
rect 2804 2685 2805 2715
rect 2805 2685 2835 2715
rect 2835 2685 2836 2715
rect 2804 2684 2836 2685
rect 2884 2875 2916 2876
rect 2884 2845 2885 2875
rect 2885 2845 2915 2875
rect 2915 2845 2916 2875
rect 2884 2844 2916 2845
rect 2884 2764 2916 2796
rect 2884 2715 2916 2716
rect 2884 2685 2885 2715
rect 2885 2685 2915 2715
rect 2915 2685 2916 2715
rect 2884 2684 2916 2685
rect 2964 2875 2996 2876
rect 2964 2845 2965 2875
rect 2965 2845 2995 2875
rect 2995 2845 2996 2875
rect 2964 2844 2996 2845
rect 2964 2764 2996 2796
rect 2964 2715 2996 2716
rect 2964 2685 2965 2715
rect 2965 2685 2995 2715
rect 2995 2685 2996 2715
rect 2964 2684 2996 2685
rect 3044 2875 3076 2876
rect 3044 2845 3045 2875
rect 3045 2845 3075 2875
rect 3075 2845 3076 2875
rect 3044 2844 3076 2845
rect 3044 2764 3076 2796
rect 3044 2715 3076 2716
rect 3044 2685 3045 2715
rect 3045 2685 3075 2715
rect 3075 2685 3076 2715
rect 3044 2684 3076 2685
rect 3124 2875 3156 2876
rect 3124 2845 3125 2875
rect 3125 2845 3155 2875
rect 3155 2845 3156 2875
rect 3124 2844 3156 2845
rect 3124 2764 3156 2796
rect 3124 2715 3156 2716
rect 3124 2685 3125 2715
rect 3125 2685 3155 2715
rect 3155 2685 3156 2715
rect 3124 2684 3156 2685
rect 3204 2875 3236 2876
rect 3204 2845 3205 2875
rect 3205 2845 3235 2875
rect 3235 2845 3236 2875
rect 3204 2844 3236 2845
rect 3204 2764 3236 2796
rect 3204 2715 3236 2716
rect 3204 2685 3205 2715
rect 3205 2685 3235 2715
rect 3235 2685 3236 2715
rect 3204 2684 3236 2685
rect 3284 2875 3316 2876
rect 3284 2845 3285 2875
rect 3285 2845 3315 2875
rect 3315 2845 3316 2875
rect 3284 2844 3316 2845
rect 3284 2764 3316 2796
rect 3284 2715 3316 2716
rect 3284 2685 3285 2715
rect 3285 2685 3315 2715
rect 3315 2685 3316 2715
rect 3284 2684 3316 2685
rect 3364 2875 3396 2876
rect 3364 2845 3365 2875
rect 3365 2845 3395 2875
rect 3395 2845 3396 2875
rect 3364 2844 3396 2845
rect 3364 2764 3396 2796
rect 3364 2715 3396 2716
rect 3364 2685 3365 2715
rect 3365 2685 3395 2715
rect 3395 2685 3396 2715
rect 3364 2684 3396 2685
rect 3444 2875 3476 2876
rect 3444 2845 3445 2875
rect 3445 2845 3475 2875
rect 3475 2845 3476 2875
rect 3444 2844 3476 2845
rect 3444 2764 3476 2796
rect 3444 2715 3476 2716
rect 3444 2685 3445 2715
rect 3445 2685 3475 2715
rect 3475 2685 3476 2715
rect 3444 2684 3476 2685
rect 3604 2875 3636 2876
rect 3604 2845 3605 2875
rect 3605 2845 3635 2875
rect 3635 2845 3636 2875
rect 3604 2844 3636 2845
rect 3604 2764 3636 2796
rect 3604 2715 3636 2716
rect 3604 2685 3605 2715
rect 3605 2685 3635 2715
rect 3635 2685 3636 2715
rect 3604 2684 3636 2685
rect 3684 2875 3716 2876
rect 3684 2845 3685 2875
rect 3685 2845 3715 2875
rect 3715 2845 3716 2875
rect 3684 2844 3716 2845
rect 3684 2764 3716 2796
rect 3684 2715 3716 2716
rect 3684 2685 3685 2715
rect 3685 2685 3715 2715
rect 3715 2685 3716 2715
rect 3684 2684 3716 2685
rect 3764 2875 3796 2876
rect 3764 2845 3765 2875
rect 3765 2845 3795 2875
rect 3795 2845 3796 2875
rect 3764 2844 3796 2845
rect 3764 2764 3796 2796
rect 3764 2715 3796 2716
rect 3764 2685 3765 2715
rect 3765 2685 3795 2715
rect 3795 2685 3796 2715
rect 3764 2684 3796 2685
rect 3844 2875 3876 2876
rect 3844 2845 3845 2875
rect 3845 2845 3875 2875
rect 3875 2845 3876 2875
rect 3844 2844 3876 2845
rect 3844 2764 3876 2796
rect 3844 2715 3876 2716
rect 3844 2685 3845 2715
rect 3845 2685 3875 2715
rect 3875 2685 3876 2715
rect 3844 2684 3876 2685
rect 3924 2875 3956 2876
rect 3924 2845 3925 2875
rect 3925 2845 3955 2875
rect 3955 2845 3956 2875
rect 3924 2844 3956 2845
rect 3924 2764 3956 2796
rect 3924 2715 3956 2716
rect 3924 2685 3925 2715
rect 3925 2685 3955 2715
rect 3955 2685 3956 2715
rect 3924 2684 3956 2685
rect 4084 2875 4116 2876
rect 4084 2845 4085 2875
rect 4085 2845 4115 2875
rect 4115 2845 4116 2875
rect 4084 2844 4116 2845
rect 4084 2764 4116 2796
rect 4084 2715 4116 2716
rect 4084 2685 4085 2715
rect 4085 2685 4115 2715
rect 4115 2685 4116 2715
rect 4084 2684 4116 2685
rect 164 2390 196 2391
rect 164 2210 165 2390
rect 165 2210 195 2390
rect 195 2210 196 2390
rect 164 2209 196 2210
rect 4004 1830 4036 1831
rect 4004 1650 4005 1830
rect 4005 1650 4035 1830
rect 4035 1650 4036 1830
rect 4004 1649 4036 1650
rect 4 1395 36 1396
rect 4 1365 5 1395
rect 5 1365 35 1395
rect 35 1365 36 1395
rect 4 1364 36 1365
rect 4 1235 36 1236
rect 4 1205 5 1235
rect 5 1205 35 1235
rect 35 1205 36 1235
rect 4 1204 36 1205
rect 84 1395 116 1396
rect 84 1365 85 1395
rect 85 1365 115 1395
rect 115 1365 116 1395
rect 84 1364 116 1365
rect 84 1235 116 1236
rect 84 1205 85 1235
rect 85 1205 115 1235
rect 115 1205 116 1235
rect 84 1204 116 1205
rect 164 1395 196 1396
rect 164 1365 165 1395
rect 165 1365 195 1395
rect 195 1365 196 1395
rect 164 1364 196 1365
rect 164 1235 196 1236
rect 164 1205 165 1235
rect 165 1205 195 1235
rect 195 1205 196 1235
rect 164 1204 196 1205
rect 244 1395 276 1396
rect 244 1365 245 1395
rect 245 1365 275 1395
rect 275 1365 276 1395
rect 244 1364 276 1365
rect 244 1235 276 1236
rect 244 1205 245 1235
rect 245 1205 275 1235
rect 275 1205 276 1235
rect 244 1204 276 1205
rect 324 1395 356 1396
rect 324 1365 325 1395
rect 325 1365 355 1395
rect 355 1365 356 1395
rect 324 1364 356 1365
rect 324 1235 356 1236
rect 324 1205 325 1235
rect 325 1205 355 1235
rect 355 1205 356 1235
rect 324 1204 356 1205
rect 404 1395 436 1396
rect 404 1365 405 1395
rect 405 1365 435 1395
rect 435 1365 436 1395
rect 404 1364 436 1365
rect 404 1235 436 1236
rect 404 1205 405 1235
rect 405 1205 435 1235
rect 435 1205 436 1235
rect 404 1204 436 1205
rect 484 1395 516 1396
rect 484 1365 485 1395
rect 485 1365 515 1395
rect 515 1365 516 1395
rect 484 1364 516 1365
rect 484 1235 516 1236
rect 484 1205 485 1235
rect 485 1205 515 1235
rect 515 1205 516 1235
rect 484 1204 516 1205
rect 564 1395 596 1396
rect 564 1365 565 1395
rect 565 1365 595 1395
rect 595 1365 596 1395
rect 564 1364 596 1365
rect 564 1235 596 1236
rect 564 1205 565 1235
rect 565 1205 595 1235
rect 595 1205 596 1235
rect 564 1204 596 1205
rect 724 1395 756 1396
rect 724 1365 725 1395
rect 725 1365 755 1395
rect 755 1365 756 1395
rect 724 1364 756 1365
rect 724 1235 756 1236
rect 724 1205 725 1235
rect 725 1205 755 1235
rect 755 1205 756 1235
rect 724 1204 756 1205
rect 804 1395 836 1396
rect 804 1365 805 1395
rect 805 1365 835 1395
rect 835 1365 836 1395
rect 804 1364 836 1365
rect 804 1235 836 1236
rect 804 1205 805 1235
rect 805 1205 835 1235
rect 835 1205 836 1235
rect 804 1204 836 1205
rect 884 1395 916 1396
rect 884 1365 885 1395
rect 885 1365 915 1395
rect 915 1365 916 1395
rect 884 1364 916 1365
rect 884 1235 916 1236
rect 884 1205 885 1235
rect 885 1205 915 1235
rect 915 1205 916 1235
rect 884 1204 916 1205
rect 964 1395 996 1396
rect 964 1365 965 1395
rect 965 1365 995 1395
rect 995 1365 996 1395
rect 964 1364 996 1365
rect 964 1235 996 1236
rect 964 1205 965 1235
rect 965 1205 995 1235
rect 995 1205 996 1235
rect 964 1204 996 1205
rect 1044 1395 1076 1396
rect 1044 1365 1045 1395
rect 1045 1365 1075 1395
rect 1075 1365 1076 1395
rect 1044 1364 1076 1365
rect 1044 1235 1076 1236
rect 1044 1205 1045 1235
rect 1045 1205 1075 1235
rect 1075 1205 1076 1235
rect 1044 1204 1076 1205
rect 1124 1395 1156 1396
rect 1124 1365 1125 1395
rect 1125 1365 1155 1395
rect 1155 1365 1156 1395
rect 1124 1364 1156 1365
rect 1124 1235 1156 1236
rect 1124 1205 1125 1235
rect 1125 1205 1155 1235
rect 1155 1205 1156 1235
rect 1124 1204 1156 1205
rect 1204 1395 1236 1396
rect 1204 1365 1205 1395
rect 1205 1365 1235 1395
rect 1235 1365 1236 1395
rect 1204 1364 1236 1365
rect 1204 1235 1236 1236
rect 1204 1205 1205 1235
rect 1205 1205 1235 1235
rect 1235 1205 1236 1235
rect 1204 1204 1236 1205
rect 1284 1395 1316 1396
rect 1284 1365 1285 1395
rect 1285 1365 1315 1395
rect 1315 1365 1316 1395
rect 1284 1364 1316 1365
rect 1284 1235 1316 1236
rect 1284 1205 1285 1235
rect 1285 1205 1315 1235
rect 1315 1205 1316 1235
rect 1284 1204 1316 1205
rect 1364 1395 1396 1396
rect 1364 1365 1365 1395
rect 1365 1365 1395 1395
rect 1395 1365 1396 1395
rect 1364 1364 1396 1365
rect 1364 1235 1396 1236
rect 1364 1205 1365 1235
rect 1365 1205 1395 1235
rect 1395 1205 1396 1235
rect 1364 1204 1396 1205
rect 1444 1395 1476 1396
rect 1444 1365 1445 1395
rect 1445 1365 1475 1395
rect 1475 1365 1476 1395
rect 1444 1364 1476 1365
rect 1444 1235 1476 1236
rect 1444 1205 1445 1235
rect 1445 1205 1475 1235
rect 1475 1205 1476 1235
rect 1444 1204 1476 1205
rect 1524 1395 1556 1396
rect 1524 1365 1525 1395
rect 1525 1365 1555 1395
rect 1555 1365 1556 1395
rect 1524 1364 1556 1365
rect 1524 1235 1556 1236
rect 1524 1205 1525 1235
rect 1525 1205 1555 1235
rect 1555 1205 1556 1235
rect 1524 1204 1556 1205
rect 1684 1395 1716 1396
rect 1684 1365 1685 1395
rect 1685 1365 1715 1395
rect 1715 1365 1716 1395
rect 1684 1364 1716 1365
rect 1684 1235 1716 1236
rect 1684 1205 1685 1235
rect 1685 1205 1715 1235
rect 1715 1205 1716 1235
rect 1684 1204 1716 1205
rect 1764 1395 1796 1396
rect 1764 1365 1765 1395
rect 1765 1365 1795 1395
rect 1795 1365 1796 1395
rect 1764 1364 1796 1365
rect 1764 1235 1796 1236
rect 1764 1205 1765 1235
rect 1765 1205 1795 1235
rect 1795 1205 1796 1235
rect 1764 1204 1796 1205
rect 1844 1395 1876 1396
rect 1844 1365 1845 1395
rect 1845 1365 1875 1395
rect 1875 1365 1876 1395
rect 1844 1364 1876 1365
rect 1844 1235 1876 1236
rect 1844 1205 1845 1235
rect 1845 1205 1875 1235
rect 1875 1205 1876 1235
rect 1844 1204 1876 1205
rect 1924 1395 1956 1396
rect 1924 1365 1925 1395
rect 1925 1365 1955 1395
rect 1955 1365 1956 1395
rect 1924 1364 1956 1365
rect 1924 1235 1956 1236
rect 1924 1205 1925 1235
rect 1925 1205 1955 1235
rect 1955 1205 1956 1235
rect 1924 1204 1956 1205
rect 2004 1395 2036 1396
rect 2004 1365 2005 1395
rect 2005 1365 2035 1395
rect 2035 1365 2036 1395
rect 2004 1364 2036 1365
rect 2004 1235 2036 1236
rect 2004 1205 2005 1235
rect 2005 1205 2035 1235
rect 2035 1205 2036 1235
rect 2004 1204 2036 1205
rect 2084 1395 2116 1396
rect 2084 1365 2085 1395
rect 2085 1365 2115 1395
rect 2115 1365 2116 1395
rect 2084 1364 2116 1365
rect 2084 1235 2116 1236
rect 2084 1205 2085 1235
rect 2085 1205 2115 1235
rect 2115 1205 2116 1235
rect 2084 1204 2116 1205
rect 2164 1395 2196 1396
rect 2164 1365 2165 1395
rect 2165 1365 2195 1395
rect 2195 1365 2196 1395
rect 2164 1364 2196 1365
rect 2164 1235 2196 1236
rect 2164 1205 2165 1235
rect 2165 1205 2195 1235
rect 2195 1205 2196 1235
rect 2164 1204 2196 1205
rect 2244 1395 2276 1396
rect 2244 1365 2245 1395
rect 2245 1365 2275 1395
rect 2275 1365 2276 1395
rect 2244 1364 2276 1365
rect 2244 1235 2276 1236
rect 2244 1205 2245 1235
rect 2245 1205 2275 1235
rect 2275 1205 2276 1235
rect 2244 1204 2276 1205
rect 2324 1395 2356 1396
rect 2324 1365 2325 1395
rect 2325 1365 2355 1395
rect 2355 1365 2356 1395
rect 2324 1364 2356 1365
rect 2324 1235 2356 1236
rect 2324 1205 2325 1235
rect 2325 1205 2355 1235
rect 2355 1205 2356 1235
rect 2324 1204 2356 1205
rect 2404 1395 2436 1396
rect 2404 1365 2405 1395
rect 2405 1365 2435 1395
rect 2435 1365 2436 1395
rect 2404 1364 2436 1365
rect 2404 1235 2436 1236
rect 2404 1205 2405 1235
rect 2405 1205 2435 1235
rect 2435 1205 2436 1235
rect 2404 1204 2436 1205
rect 2484 1395 2516 1396
rect 2484 1365 2485 1395
rect 2485 1365 2515 1395
rect 2515 1365 2516 1395
rect 2484 1364 2516 1365
rect 2484 1235 2516 1236
rect 2484 1205 2485 1235
rect 2485 1205 2515 1235
rect 2515 1205 2516 1235
rect 2484 1204 2516 1205
rect 2644 1395 2676 1396
rect 2644 1365 2645 1395
rect 2645 1365 2675 1395
rect 2675 1365 2676 1395
rect 2644 1364 2676 1365
rect 2644 1235 2676 1236
rect 2644 1205 2645 1235
rect 2645 1205 2675 1235
rect 2675 1205 2676 1235
rect 2644 1204 2676 1205
rect 2724 1395 2756 1396
rect 2724 1365 2725 1395
rect 2725 1365 2755 1395
rect 2755 1365 2756 1395
rect 2724 1364 2756 1365
rect 2724 1235 2756 1236
rect 2724 1205 2725 1235
rect 2725 1205 2755 1235
rect 2755 1205 2756 1235
rect 2724 1204 2756 1205
rect 2804 1395 2836 1396
rect 2804 1365 2805 1395
rect 2805 1365 2835 1395
rect 2835 1365 2836 1395
rect 2804 1364 2836 1365
rect 2804 1235 2836 1236
rect 2804 1205 2805 1235
rect 2805 1205 2835 1235
rect 2835 1205 2836 1235
rect 2804 1204 2836 1205
rect 2884 1395 2916 1396
rect 2884 1365 2885 1395
rect 2885 1365 2915 1395
rect 2915 1365 2916 1395
rect 2884 1364 2916 1365
rect 2884 1235 2916 1236
rect 2884 1205 2885 1235
rect 2885 1205 2915 1235
rect 2915 1205 2916 1235
rect 2884 1204 2916 1205
rect 2964 1395 2996 1396
rect 2964 1365 2965 1395
rect 2965 1365 2995 1395
rect 2995 1365 2996 1395
rect 2964 1364 2996 1365
rect 2964 1235 2996 1236
rect 2964 1205 2965 1235
rect 2965 1205 2995 1235
rect 2995 1205 2996 1235
rect 2964 1204 2996 1205
rect 3044 1395 3076 1396
rect 3044 1365 3045 1395
rect 3045 1365 3075 1395
rect 3075 1365 3076 1395
rect 3044 1364 3076 1365
rect 3044 1235 3076 1236
rect 3044 1205 3045 1235
rect 3045 1205 3075 1235
rect 3075 1205 3076 1235
rect 3044 1204 3076 1205
rect 3124 1395 3156 1396
rect 3124 1365 3125 1395
rect 3125 1365 3155 1395
rect 3155 1365 3156 1395
rect 3124 1364 3156 1365
rect 3124 1235 3156 1236
rect 3124 1205 3125 1235
rect 3125 1205 3155 1235
rect 3155 1205 3156 1235
rect 3124 1204 3156 1205
rect 3204 1395 3236 1396
rect 3204 1365 3205 1395
rect 3205 1365 3235 1395
rect 3235 1365 3236 1395
rect 3204 1364 3236 1365
rect 3204 1235 3236 1236
rect 3204 1205 3205 1235
rect 3205 1205 3235 1235
rect 3235 1205 3236 1235
rect 3204 1204 3236 1205
rect 3284 1395 3316 1396
rect 3284 1365 3285 1395
rect 3285 1365 3315 1395
rect 3315 1365 3316 1395
rect 3284 1364 3316 1365
rect 3284 1235 3316 1236
rect 3284 1205 3285 1235
rect 3285 1205 3315 1235
rect 3315 1205 3316 1235
rect 3284 1204 3316 1205
rect 3364 1395 3396 1396
rect 3364 1365 3365 1395
rect 3365 1365 3395 1395
rect 3395 1365 3396 1395
rect 3364 1364 3396 1365
rect 3364 1235 3396 1236
rect 3364 1205 3365 1235
rect 3365 1205 3395 1235
rect 3395 1205 3396 1235
rect 3364 1204 3396 1205
rect 3444 1395 3476 1396
rect 3444 1365 3445 1395
rect 3445 1365 3475 1395
rect 3475 1365 3476 1395
rect 3444 1364 3476 1365
rect 3444 1235 3476 1236
rect 3444 1205 3445 1235
rect 3445 1205 3475 1235
rect 3475 1205 3476 1235
rect 3444 1204 3476 1205
rect 3604 1395 3636 1396
rect 3604 1365 3605 1395
rect 3605 1365 3635 1395
rect 3635 1365 3636 1395
rect 3604 1364 3636 1365
rect 3604 1235 3636 1236
rect 3604 1205 3605 1235
rect 3605 1205 3635 1235
rect 3635 1205 3636 1235
rect 3604 1204 3636 1205
rect 3684 1395 3716 1396
rect 3684 1365 3685 1395
rect 3685 1365 3715 1395
rect 3715 1365 3716 1395
rect 3684 1364 3716 1365
rect 3684 1235 3716 1236
rect 3684 1205 3685 1235
rect 3685 1205 3715 1235
rect 3715 1205 3716 1235
rect 3684 1204 3716 1205
rect 3764 1395 3796 1396
rect 3764 1365 3765 1395
rect 3765 1365 3795 1395
rect 3795 1365 3796 1395
rect 3764 1364 3796 1365
rect 3764 1235 3796 1236
rect 3764 1205 3765 1235
rect 3765 1205 3795 1235
rect 3795 1205 3796 1235
rect 3764 1204 3796 1205
rect 3844 1395 3876 1396
rect 3844 1365 3845 1395
rect 3845 1365 3875 1395
rect 3875 1365 3876 1395
rect 3844 1364 3876 1365
rect 3844 1235 3876 1236
rect 3844 1205 3845 1235
rect 3845 1205 3875 1235
rect 3875 1205 3876 1235
rect 3844 1204 3876 1205
rect 3924 1395 3956 1396
rect 3924 1365 3925 1395
rect 3925 1365 3955 1395
rect 3955 1365 3956 1395
rect 3924 1364 3956 1365
rect 3924 1235 3956 1236
rect 3924 1205 3925 1235
rect 3925 1205 3955 1235
rect 3955 1205 3956 1235
rect 3924 1204 3956 1205
rect 4004 1395 4036 1396
rect 4004 1365 4005 1395
rect 4005 1365 4035 1395
rect 4035 1365 4036 1395
rect 4004 1364 4036 1365
rect 4004 1235 4036 1236
rect 4004 1205 4005 1235
rect 4005 1205 4035 1235
rect 4035 1205 4036 1235
rect 4004 1204 4036 1205
rect 4084 1395 4116 1396
rect 4084 1365 4085 1395
rect 4085 1365 4115 1395
rect 4115 1365 4116 1395
rect 4084 1364 4116 1365
rect 4084 1235 4116 1236
rect 4084 1205 4085 1235
rect 4085 1205 4115 1235
rect 4115 1205 4116 1235
rect 4084 1204 4116 1205
rect 4164 1395 4196 1396
rect 4164 1365 4165 1395
rect 4165 1365 4195 1395
rect 4195 1365 4196 1395
rect 4164 1364 4196 1365
rect 4164 1235 4196 1236
rect 4164 1205 4165 1235
rect 4165 1205 4195 1235
rect 4195 1205 4196 1235
rect 4164 1204 4196 1205
rect 84 524 116 556
rect 84 475 116 476
rect 84 445 85 475
rect 85 445 115 475
rect 115 445 116 475
rect 84 444 116 445
rect 84 364 116 396
rect 164 524 196 556
rect 164 475 196 476
rect 164 445 165 475
rect 165 445 195 475
rect 195 445 196 475
rect 164 444 196 445
rect 164 364 196 396
rect 244 524 276 556
rect 244 475 276 476
rect 244 445 245 475
rect 245 445 275 475
rect 275 445 276 475
rect 244 444 276 445
rect 244 364 276 396
rect 324 524 356 556
rect 324 475 356 476
rect 324 445 325 475
rect 325 445 355 475
rect 355 445 356 475
rect 324 444 356 445
rect 324 364 356 396
rect 404 524 436 556
rect 404 475 436 476
rect 404 445 405 475
rect 405 445 435 475
rect 435 445 436 475
rect 404 444 436 445
rect 404 364 436 396
rect 484 524 516 556
rect 484 475 516 476
rect 484 445 485 475
rect 485 445 515 475
rect 515 445 516 475
rect 484 444 516 445
rect 484 364 516 396
rect 564 524 596 556
rect 564 475 596 476
rect 564 445 565 475
rect 565 445 595 475
rect 595 445 596 475
rect 564 444 596 445
rect 564 364 596 396
rect 724 524 756 556
rect 724 475 756 476
rect 724 445 725 475
rect 725 445 755 475
rect 755 445 756 475
rect 724 444 756 445
rect 724 364 756 396
rect 804 524 836 556
rect 804 475 836 476
rect 804 445 805 475
rect 805 445 835 475
rect 835 445 836 475
rect 804 444 836 445
rect 804 364 836 396
rect 884 524 916 556
rect 884 475 916 476
rect 884 445 885 475
rect 885 445 915 475
rect 915 445 916 475
rect 884 444 916 445
rect 884 364 916 396
rect 964 524 996 556
rect 964 475 996 476
rect 964 445 965 475
rect 965 445 995 475
rect 995 445 996 475
rect 964 444 996 445
rect 964 364 996 396
rect 1044 524 1076 556
rect 1044 475 1076 476
rect 1044 445 1045 475
rect 1045 445 1075 475
rect 1075 445 1076 475
rect 1044 444 1076 445
rect 1044 364 1076 396
rect 1124 524 1156 556
rect 1124 475 1156 476
rect 1124 445 1125 475
rect 1125 445 1155 475
rect 1155 445 1156 475
rect 1124 444 1156 445
rect 1124 364 1156 396
rect 1204 524 1236 556
rect 1204 475 1236 476
rect 1204 445 1205 475
rect 1205 445 1235 475
rect 1235 445 1236 475
rect 1204 444 1236 445
rect 1204 364 1236 396
rect 1284 524 1316 556
rect 1284 475 1316 476
rect 1284 445 1285 475
rect 1285 445 1315 475
rect 1315 445 1316 475
rect 1284 444 1316 445
rect 1284 364 1316 396
rect 1364 524 1396 556
rect 1364 475 1396 476
rect 1364 445 1365 475
rect 1365 445 1395 475
rect 1395 445 1396 475
rect 1364 444 1396 445
rect 1364 364 1396 396
rect 1444 524 1476 556
rect 1444 475 1476 476
rect 1444 445 1445 475
rect 1445 445 1475 475
rect 1475 445 1476 475
rect 1444 444 1476 445
rect 1444 364 1476 396
rect 1524 524 1556 556
rect 1524 475 1556 476
rect 1524 445 1525 475
rect 1525 445 1555 475
rect 1555 445 1556 475
rect 1524 444 1556 445
rect 1524 364 1556 396
rect 1684 524 1716 556
rect 1684 475 1716 476
rect 1684 445 1685 475
rect 1685 445 1715 475
rect 1715 445 1716 475
rect 1684 444 1716 445
rect 1684 364 1716 396
rect 1764 524 1796 556
rect 1764 475 1796 476
rect 1764 445 1765 475
rect 1765 445 1795 475
rect 1795 445 1796 475
rect 1764 444 1796 445
rect 1764 364 1796 396
rect 1844 524 1876 556
rect 1844 475 1876 476
rect 1844 445 1845 475
rect 1845 445 1875 475
rect 1875 445 1876 475
rect 1844 444 1876 445
rect 1844 364 1876 396
rect 1924 524 1956 556
rect 1924 475 1956 476
rect 1924 445 1925 475
rect 1925 445 1955 475
rect 1955 445 1956 475
rect 1924 444 1956 445
rect 1924 364 1956 396
rect 2004 524 2036 556
rect 2004 475 2036 476
rect 2004 445 2005 475
rect 2005 445 2035 475
rect 2035 445 2036 475
rect 2004 444 2036 445
rect 2004 364 2036 396
rect 2084 524 2116 556
rect 2084 475 2116 476
rect 2084 445 2085 475
rect 2085 445 2115 475
rect 2115 445 2116 475
rect 2084 444 2116 445
rect 2084 364 2116 396
rect 2164 524 2196 556
rect 2164 475 2196 476
rect 2164 445 2165 475
rect 2165 445 2195 475
rect 2195 445 2196 475
rect 2164 444 2196 445
rect 2164 364 2196 396
rect 2244 524 2276 556
rect 2244 475 2276 476
rect 2244 445 2245 475
rect 2245 445 2275 475
rect 2275 445 2276 475
rect 2244 444 2276 445
rect 2244 364 2276 396
rect 2324 524 2356 556
rect 2324 475 2356 476
rect 2324 445 2325 475
rect 2325 445 2355 475
rect 2355 445 2356 475
rect 2324 444 2356 445
rect 2324 364 2356 396
rect 2404 524 2436 556
rect 2404 475 2436 476
rect 2404 445 2405 475
rect 2405 445 2435 475
rect 2435 445 2436 475
rect 2404 444 2436 445
rect 2404 364 2436 396
rect 2484 524 2516 556
rect 2484 475 2516 476
rect 2484 445 2485 475
rect 2485 445 2515 475
rect 2515 445 2516 475
rect 2484 444 2516 445
rect 2484 364 2516 396
rect 2644 524 2676 556
rect 2644 475 2676 476
rect 2644 445 2645 475
rect 2645 445 2675 475
rect 2675 445 2676 475
rect 2644 444 2676 445
rect 2644 364 2676 396
rect 2724 524 2756 556
rect 2724 475 2756 476
rect 2724 445 2725 475
rect 2725 445 2755 475
rect 2755 445 2756 475
rect 2724 444 2756 445
rect 2724 364 2756 396
rect 2804 524 2836 556
rect 2804 475 2836 476
rect 2804 445 2805 475
rect 2805 445 2835 475
rect 2835 445 2836 475
rect 2804 444 2836 445
rect 2804 364 2836 396
rect 2884 524 2916 556
rect 2884 475 2916 476
rect 2884 445 2885 475
rect 2885 445 2915 475
rect 2915 445 2916 475
rect 2884 444 2916 445
rect 2884 364 2916 396
rect 2964 524 2996 556
rect 2964 475 2996 476
rect 2964 445 2965 475
rect 2965 445 2995 475
rect 2995 445 2996 475
rect 2964 444 2996 445
rect 2964 364 2996 396
rect 3044 524 3076 556
rect 3044 475 3076 476
rect 3044 445 3045 475
rect 3045 445 3075 475
rect 3075 445 3076 475
rect 3044 444 3076 445
rect 3044 364 3076 396
rect 3124 524 3156 556
rect 3124 475 3156 476
rect 3124 445 3125 475
rect 3125 445 3155 475
rect 3155 445 3156 475
rect 3124 444 3156 445
rect 3124 364 3156 396
rect 3204 524 3236 556
rect 3204 475 3236 476
rect 3204 445 3205 475
rect 3205 445 3235 475
rect 3235 445 3236 475
rect 3204 444 3236 445
rect 3204 364 3236 396
rect 3284 524 3316 556
rect 3284 475 3316 476
rect 3284 445 3285 475
rect 3285 445 3315 475
rect 3315 445 3316 475
rect 3284 444 3316 445
rect 3284 364 3316 396
rect 3364 524 3396 556
rect 3364 475 3396 476
rect 3364 445 3365 475
rect 3365 445 3395 475
rect 3395 445 3396 475
rect 3364 444 3396 445
rect 3364 364 3396 396
rect 3444 524 3476 556
rect 3444 475 3476 476
rect 3444 445 3445 475
rect 3445 445 3475 475
rect 3475 445 3476 475
rect 3444 444 3476 445
rect 3444 364 3476 396
rect 3604 524 3636 556
rect 3604 475 3636 476
rect 3604 445 3605 475
rect 3605 445 3635 475
rect 3635 445 3636 475
rect 3604 444 3636 445
rect 3604 364 3636 396
rect 3684 524 3716 556
rect 3684 475 3716 476
rect 3684 445 3685 475
rect 3685 445 3715 475
rect 3715 445 3716 475
rect 3684 444 3716 445
rect 3684 364 3716 396
rect 3764 524 3796 556
rect 3764 475 3796 476
rect 3764 445 3765 475
rect 3765 445 3795 475
rect 3795 445 3796 475
rect 3764 444 3796 445
rect 3764 364 3796 396
rect 3844 524 3876 556
rect 3844 475 3876 476
rect 3844 445 3845 475
rect 3845 445 3875 475
rect 3875 445 3876 475
rect 3844 444 3876 445
rect 3844 364 3876 396
rect 3924 524 3956 556
rect 3924 475 3956 476
rect 3924 445 3925 475
rect 3925 445 3955 475
rect 3955 445 3956 475
rect 3924 444 3956 445
rect 3924 364 3956 396
rect 4084 524 4116 556
rect 4084 475 4116 476
rect 4084 445 4085 475
rect 4085 445 4115 475
rect 4115 445 4116 475
rect 4084 444 4116 445
rect 4084 364 4116 396
rect 164 170 196 171
rect 164 90 165 170
rect 165 90 195 170
rect 195 90 196 170
rect 164 89 196 90
rect 84 -45 116 -44
rect 84 -75 85 -45
rect 85 -75 115 -45
rect 115 -75 116 -45
rect 84 -76 116 -75
rect 84 -156 116 -124
rect 84 -205 116 -204
rect 84 -235 85 -205
rect 85 -235 115 -205
rect 115 -235 116 -205
rect 84 -236 116 -235
rect 164 -45 196 -44
rect 164 -75 165 -45
rect 165 -75 195 -45
rect 195 -75 196 -45
rect 164 -76 196 -75
rect 164 -156 196 -124
rect 164 -205 196 -204
rect 164 -235 165 -205
rect 165 -235 195 -205
rect 195 -235 196 -205
rect 164 -236 196 -235
rect 244 -45 276 -44
rect 244 -75 245 -45
rect 245 -75 275 -45
rect 275 -75 276 -45
rect 244 -76 276 -75
rect 244 -156 276 -124
rect 244 -205 276 -204
rect 244 -235 245 -205
rect 245 -235 275 -205
rect 275 -235 276 -205
rect 244 -236 276 -235
rect 324 -45 356 -44
rect 324 -75 325 -45
rect 325 -75 355 -45
rect 355 -75 356 -45
rect 324 -76 356 -75
rect 324 -156 356 -124
rect 324 -205 356 -204
rect 324 -235 325 -205
rect 325 -235 355 -205
rect 355 -235 356 -205
rect 324 -236 356 -235
rect 404 -45 436 -44
rect 404 -75 405 -45
rect 405 -75 435 -45
rect 435 -75 436 -45
rect 404 -76 436 -75
rect 404 -156 436 -124
rect 404 -205 436 -204
rect 404 -235 405 -205
rect 405 -235 435 -205
rect 435 -235 436 -205
rect 404 -236 436 -235
rect 484 -45 516 -44
rect 484 -75 485 -45
rect 485 -75 515 -45
rect 515 -75 516 -45
rect 484 -76 516 -75
rect 484 -156 516 -124
rect 484 -205 516 -204
rect 484 -235 485 -205
rect 485 -235 515 -205
rect 515 -235 516 -205
rect 484 -236 516 -235
rect 564 -45 596 -44
rect 564 -75 565 -45
rect 565 -75 595 -45
rect 595 -75 596 -45
rect 564 -76 596 -75
rect 564 -156 596 -124
rect 564 -205 596 -204
rect 564 -235 565 -205
rect 565 -235 595 -205
rect 595 -235 596 -205
rect 564 -236 596 -235
rect 724 -45 756 -44
rect 724 -75 725 -45
rect 725 -75 755 -45
rect 755 -75 756 -45
rect 724 -76 756 -75
rect 724 -156 756 -124
rect 724 -205 756 -204
rect 724 -235 725 -205
rect 725 -235 755 -205
rect 755 -235 756 -205
rect 724 -236 756 -235
rect 804 -45 836 -44
rect 804 -75 805 -45
rect 805 -75 835 -45
rect 835 -75 836 -45
rect 804 -76 836 -75
rect 804 -156 836 -124
rect 804 -205 836 -204
rect 804 -235 805 -205
rect 805 -235 835 -205
rect 835 -235 836 -205
rect 804 -236 836 -235
rect 884 -45 916 -44
rect 884 -75 885 -45
rect 885 -75 915 -45
rect 915 -75 916 -45
rect 884 -76 916 -75
rect 884 -156 916 -124
rect 884 -205 916 -204
rect 884 -235 885 -205
rect 885 -235 915 -205
rect 915 -235 916 -205
rect 884 -236 916 -235
rect 964 -45 996 -44
rect 964 -75 965 -45
rect 965 -75 995 -45
rect 995 -75 996 -45
rect 964 -76 996 -75
rect 964 -156 996 -124
rect 964 -205 996 -204
rect 964 -235 965 -205
rect 965 -235 995 -205
rect 995 -235 996 -205
rect 964 -236 996 -235
rect 1044 -45 1076 -44
rect 1044 -75 1045 -45
rect 1045 -75 1075 -45
rect 1075 -75 1076 -45
rect 1044 -76 1076 -75
rect 1044 -156 1076 -124
rect 1044 -205 1076 -204
rect 1044 -235 1045 -205
rect 1045 -235 1075 -205
rect 1075 -235 1076 -205
rect 1044 -236 1076 -235
rect 1124 -45 1156 -44
rect 1124 -75 1125 -45
rect 1125 -75 1155 -45
rect 1155 -75 1156 -45
rect 1124 -76 1156 -75
rect 1124 -156 1156 -124
rect 1124 -205 1156 -204
rect 1124 -235 1125 -205
rect 1125 -235 1155 -205
rect 1155 -235 1156 -205
rect 1124 -236 1156 -235
rect 1204 -45 1236 -44
rect 1204 -75 1205 -45
rect 1205 -75 1235 -45
rect 1235 -75 1236 -45
rect 1204 -76 1236 -75
rect 1204 -156 1236 -124
rect 1204 -205 1236 -204
rect 1204 -235 1205 -205
rect 1205 -235 1235 -205
rect 1235 -235 1236 -205
rect 1204 -236 1236 -235
rect 1284 -45 1316 -44
rect 1284 -75 1285 -45
rect 1285 -75 1315 -45
rect 1315 -75 1316 -45
rect 1284 -76 1316 -75
rect 1284 -156 1316 -124
rect 1284 -205 1316 -204
rect 1284 -235 1285 -205
rect 1285 -235 1315 -205
rect 1315 -235 1316 -205
rect 1284 -236 1316 -235
rect 1364 -45 1396 -44
rect 1364 -75 1365 -45
rect 1365 -75 1395 -45
rect 1395 -75 1396 -45
rect 1364 -76 1396 -75
rect 1364 -156 1396 -124
rect 1364 -205 1396 -204
rect 1364 -235 1365 -205
rect 1365 -235 1395 -205
rect 1395 -235 1396 -205
rect 1364 -236 1396 -235
rect 1444 -45 1476 -44
rect 1444 -75 1445 -45
rect 1445 -75 1475 -45
rect 1475 -75 1476 -45
rect 1444 -76 1476 -75
rect 1444 -156 1476 -124
rect 1444 -205 1476 -204
rect 1444 -235 1445 -205
rect 1445 -235 1475 -205
rect 1475 -235 1476 -205
rect 1444 -236 1476 -235
rect 1524 -45 1556 -44
rect 1524 -75 1525 -45
rect 1525 -75 1555 -45
rect 1555 -75 1556 -45
rect 1524 -76 1556 -75
rect 1524 -156 1556 -124
rect 1524 -205 1556 -204
rect 1524 -235 1525 -205
rect 1525 -235 1555 -205
rect 1555 -235 1556 -205
rect 1524 -236 1556 -235
rect 1684 -45 1716 -44
rect 1684 -75 1685 -45
rect 1685 -75 1715 -45
rect 1715 -75 1716 -45
rect 1684 -76 1716 -75
rect 1684 -156 1716 -124
rect 1684 -205 1716 -204
rect 1684 -235 1685 -205
rect 1685 -235 1715 -205
rect 1715 -235 1716 -205
rect 1684 -236 1716 -235
rect 1764 -45 1796 -44
rect 1764 -75 1765 -45
rect 1765 -75 1795 -45
rect 1795 -75 1796 -45
rect 1764 -76 1796 -75
rect 1764 -156 1796 -124
rect 1764 -205 1796 -204
rect 1764 -235 1765 -205
rect 1765 -235 1795 -205
rect 1795 -235 1796 -205
rect 1764 -236 1796 -235
rect 1844 -45 1876 -44
rect 1844 -75 1845 -45
rect 1845 -75 1875 -45
rect 1875 -75 1876 -45
rect 1844 -76 1876 -75
rect 1844 -156 1876 -124
rect 1844 -205 1876 -204
rect 1844 -235 1845 -205
rect 1845 -235 1875 -205
rect 1875 -235 1876 -205
rect 1844 -236 1876 -235
rect 1924 -45 1956 -44
rect 1924 -75 1925 -45
rect 1925 -75 1955 -45
rect 1955 -75 1956 -45
rect 1924 -76 1956 -75
rect 1924 -156 1956 -124
rect 1924 -205 1956 -204
rect 1924 -235 1925 -205
rect 1925 -235 1955 -205
rect 1955 -235 1956 -205
rect 1924 -236 1956 -235
rect 2004 -45 2036 -44
rect 2004 -75 2005 -45
rect 2005 -75 2035 -45
rect 2035 -75 2036 -45
rect 2004 -76 2036 -75
rect 2004 -156 2036 -124
rect 2004 -205 2036 -204
rect 2004 -235 2005 -205
rect 2005 -235 2035 -205
rect 2035 -235 2036 -205
rect 2004 -236 2036 -235
rect 2084 -45 2116 -44
rect 2084 -75 2085 -45
rect 2085 -75 2115 -45
rect 2115 -75 2116 -45
rect 2084 -76 2116 -75
rect 2084 -156 2116 -124
rect 2084 -205 2116 -204
rect 2084 -235 2085 -205
rect 2085 -235 2115 -205
rect 2115 -235 2116 -205
rect 2084 -236 2116 -235
rect 2164 -45 2196 -44
rect 2164 -75 2165 -45
rect 2165 -75 2195 -45
rect 2195 -75 2196 -45
rect 2164 -76 2196 -75
rect 2164 -156 2196 -124
rect 2164 -205 2196 -204
rect 2164 -235 2165 -205
rect 2165 -235 2195 -205
rect 2195 -235 2196 -205
rect 2164 -236 2196 -235
rect 2244 -45 2276 -44
rect 2244 -75 2245 -45
rect 2245 -75 2275 -45
rect 2275 -75 2276 -45
rect 2244 -76 2276 -75
rect 2244 -156 2276 -124
rect 2244 -205 2276 -204
rect 2244 -235 2245 -205
rect 2245 -235 2275 -205
rect 2275 -235 2276 -205
rect 2244 -236 2276 -235
rect 2324 -45 2356 -44
rect 2324 -75 2325 -45
rect 2325 -75 2355 -45
rect 2355 -75 2356 -45
rect 2324 -76 2356 -75
rect 2324 -156 2356 -124
rect 2324 -205 2356 -204
rect 2324 -235 2325 -205
rect 2325 -235 2355 -205
rect 2355 -235 2356 -205
rect 2324 -236 2356 -235
rect 2404 -45 2436 -44
rect 2404 -75 2405 -45
rect 2405 -75 2435 -45
rect 2435 -75 2436 -45
rect 2404 -76 2436 -75
rect 2404 -156 2436 -124
rect 2404 -205 2436 -204
rect 2404 -235 2405 -205
rect 2405 -235 2435 -205
rect 2435 -235 2436 -205
rect 2404 -236 2436 -235
rect 2484 -45 2516 -44
rect 2484 -75 2485 -45
rect 2485 -75 2515 -45
rect 2515 -75 2516 -45
rect 2484 -76 2516 -75
rect 2484 -156 2516 -124
rect 2484 -205 2516 -204
rect 2484 -235 2485 -205
rect 2485 -235 2515 -205
rect 2515 -235 2516 -205
rect 2484 -236 2516 -235
rect 2644 -45 2676 -44
rect 2644 -75 2645 -45
rect 2645 -75 2675 -45
rect 2675 -75 2676 -45
rect 2644 -76 2676 -75
rect 2644 -156 2676 -124
rect 2644 -205 2676 -204
rect 2644 -235 2645 -205
rect 2645 -235 2675 -205
rect 2675 -235 2676 -205
rect 2644 -236 2676 -235
rect 2724 -45 2756 -44
rect 2724 -75 2725 -45
rect 2725 -75 2755 -45
rect 2755 -75 2756 -45
rect 2724 -76 2756 -75
rect 2724 -156 2756 -124
rect 2724 -205 2756 -204
rect 2724 -235 2725 -205
rect 2725 -235 2755 -205
rect 2755 -235 2756 -205
rect 2724 -236 2756 -235
rect 2804 -45 2836 -44
rect 2804 -75 2805 -45
rect 2805 -75 2835 -45
rect 2835 -75 2836 -45
rect 2804 -76 2836 -75
rect 2804 -156 2836 -124
rect 2804 -205 2836 -204
rect 2804 -235 2805 -205
rect 2805 -235 2835 -205
rect 2835 -235 2836 -205
rect 2804 -236 2836 -235
rect 2884 -45 2916 -44
rect 2884 -75 2885 -45
rect 2885 -75 2915 -45
rect 2915 -75 2916 -45
rect 2884 -76 2916 -75
rect 2884 -156 2916 -124
rect 2884 -205 2916 -204
rect 2884 -235 2885 -205
rect 2885 -235 2915 -205
rect 2915 -235 2916 -205
rect 2884 -236 2916 -235
rect 2964 -45 2996 -44
rect 2964 -75 2965 -45
rect 2965 -75 2995 -45
rect 2995 -75 2996 -45
rect 2964 -76 2996 -75
rect 2964 -156 2996 -124
rect 2964 -205 2996 -204
rect 2964 -235 2965 -205
rect 2965 -235 2995 -205
rect 2995 -235 2996 -205
rect 2964 -236 2996 -235
rect 3044 -45 3076 -44
rect 3044 -75 3045 -45
rect 3045 -75 3075 -45
rect 3075 -75 3076 -45
rect 3044 -76 3076 -75
rect 3044 -156 3076 -124
rect 3044 -205 3076 -204
rect 3044 -235 3045 -205
rect 3045 -235 3075 -205
rect 3075 -235 3076 -205
rect 3044 -236 3076 -235
rect 3124 -45 3156 -44
rect 3124 -75 3125 -45
rect 3125 -75 3155 -45
rect 3155 -75 3156 -45
rect 3124 -76 3156 -75
rect 3124 -156 3156 -124
rect 3124 -205 3156 -204
rect 3124 -235 3125 -205
rect 3125 -235 3155 -205
rect 3155 -235 3156 -205
rect 3124 -236 3156 -235
rect 3204 -45 3236 -44
rect 3204 -75 3205 -45
rect 3205 -75 3235 -45
rect 3235 -75 3236 -45
rect 3204 -76 3236 -75
rect 3204 -156 3236 -124
rect 3204 -205 3236 -204
rect 3204 -235 3205 -205
rect 3205 -235 3235 -205
rect 3235 -235 3236 -205
rect 3204 -236 3236 -235
rect 3284 -45 3316 -44
rect 3284 -75 3285 -45
rect 3285 -75 3315 -45
rect 3315 -75 3316 -45
rect 3284 -76 3316 -75
rect 3284 -156 3316 -124
rect 3284 -205 3316 -204
rect 3284 -235 3285 -205
rect 3285 -235 3315 -205
rect 3315 -235 3316 -205
rect 3284 -236 3316 -235
rect 3364 -45 3396 -44
rect 3364 -75 3365 -45
rect 3365 -75 3395 -45
rect 3395 -75 3396 -45
rect 3364 -76 3396 -75
rect 3364 -156 3396 -124
rect 3364 -205 3396 -204
rect 3364 -235 3365 -205
rect 3365 -235 3395 -205
rect 3395 -235 3396 -205
rect 3364 -236 3396 -235
rect 3444 -45 3476 -44
rect 3444 -75 3445 -45
rect 3445 -75 3475 -45
rect 3475 -75 3476 -45
rect 3444 -76 3476 -75
rect 3444 -156 3476 -124
rect 3444 -205 3476 -204
rect 3444 -235 3445 -205
rect 3445 -235 3475 -205
rect 3475 -235 3476 -205
rect 3444 -236 3476 -235
rect 3604 -45 3636 -44
rect 3604 -75 3605 -45
rect 3605 -75 3635 -45
rect 3635 -75 3636 -45
rect 3604 -76 3636 -75
rect 3604 -156 3636 -124
rect 3604 -205 3636 -204
rect 3604 -235 3605 -205
rect 3605 -235 3635 -205
rect 3635 -235 3636 -205
rect 3604 -236 3636 -235
rect 3684 -45 3716 -44
rect 3684 -75 3685 -45
rect 3685 -75 3715 -45
rect 3715 -75 3716 -45
rect 3684 -76 3716 -75
rect 3684 -156 3716 -124
rect 3684 -205 3716 -204
rect 3684 -235 3685 -205
rect 3685 -235 3715 -205
rect 3715 -235 3716 -205
rect 3684 -236 3716 -235
rect 3764 -45 3796 -44
rect 3764 -75 3765 -45
rect 3765 -75 3795 -45
rect 3795 -75 3796 -45
rect 3764 -76 3796 -75
rect 3764 -156 3796 -124
rect 3764 -205 3796 -204
rect 3764 -235 3765 -205
rect 3765 -235 3795 -205
rect 3795 -235 3796 -205
rect 3764 -236 3796 -235
rect 3844 -45 3876 -44
rect 3844 -75 3845 -45
rect 3845 -75 3875 -45
rect 3875 -75 3876 -45
rect 3844 -76 3876 -75
rect 3844 -156 3876 -124
rect 3844 -205 3876 -204
rect 3844 -235 3845 -205
rect 3845 -235 3875 -205
rect 3875 -235 3876 -205
rect 3844 -236 3876 -235
rect 3924 -45 3956 -44
rect 3924 -75 3925 -45
rect 3925 -75 3955 -45
rect 3955 -75 3956 -45
rect 3924 -76 3956 -75
rect 3924 -156 3956 -124
rect 3924 -205 3956 -204
rect 3924 -235 3925 -205
rect 3925 -235 3955 -205
rect 3955 -235 3956 -205
rect 3924 -236 3956 -235
rect 4084 -45 4116 -44
rect 4084 -75 4085 -45
rect 4085 -75 4115 -45
rect 4115 -75 4116 -45
rect 4084 -76 4116 -75
rect 4084 -156 4116 -124
rect 4084 -205 4116 -204
rect 4084 -235 4085 -205
rect 4085 -235 4115 -205
rect 4115 -235 4116 -205
rect 4084 -236 4116 -235
rect 164 -350 196 -349
rect 164 -430 165 -350
rect 165 -430 195 -350
rect 195 -430 196 -350
rect 164 -431 196 -430
<< metal4 >>
rect 0 4871 4200 4880
rect 0 4840 164 4871
rect 196 4840 4200 4871
rect 0 4720 120 4840
rect 240 4720 3960 4840
rect 4080 4720 4200 4840
rect 0 4689 164 4720
rect 196 4689 4200 4720
rect 0 4680 4200 4689
rect 0 4396 4200 4400
rect 0 4364 84 4396
rect 116 4364 164 4396
rect 196 4364 244 4396
rect 276 4364 324 4396
rect 356 4364 404 4396
rect 436 4364 484 4396
rect 516 4364 564 4396
rect 596 4364 724 4396
rect 756 4364 804 4396
rect 836 4364 884 4396
rect 916 4364 964 4396
rect 996 4364 1044 4396
rect 1076 4364 1124 4396
rect 1156 4364 1204 4396
rect 1236 4364 1284 4396
rect 1316 4364 1364 4396
rect 1396 4364 1444 4396
rect 1476 4364 1524 4396
rect 1556 4364 1684 4396
rect 1716 4364 1764 4396
rect 1796 4364 1844 4396
rect 1876 4364 1924 4396
rect 1956 4364 2004 4396
rect 2036 4364 2084 4396
rect 2116 4364 2164 4396
rect 2196 4364 2244 4396
rect 2276 4364 2324 4396
rect 2356 4364 2404 4396
rect 2436 4364 2484 4396
rect 2516 4364 2644 4396
rect 2676 4364 2724 4396
rect 2756 4364 2804 4396
rect 2836 4364 2884 4396
rect 2916 4364 2964 4396
rect 2996 4364 3044 4396
rect 3076 4364 3124 4396
rect 3156 4364 3204 4396
rect 3236 4364 3284 4396
rect 3316 4364 3364 4396
rect 3396 4364 3444 4396
rect 3476 4364 3604 4396
rect 3636 4364 3684 4396
rect 3716 4364 3764 4396
rect 3796 4364 3844 4396
rect 3876 4364 3924 4396
rect 3956 4364 4004 4396
rect 4036 4364 4084 4396
rect 4116 4364 4200 4396
rect 0 4360 4200 4364
rect 0 4316 120 4360
rect 240 4316 3960 4360
rect 4080 4316 4200 4360
rect 0 4284 84 4316
rect 116 4284 120 4316
rect 240 4284 244 4316
rect 276 4284 324 4316
rect 356 4284 404 4316
rect 436 4284 484 4316
rect 516 4284 564 4316
rect 596 4284 724 4316
rect 756 4284 804 4316
rect 836 4284 884 4316
rect 916 4284 964 4316
rect 996 4284 1044 4316
rect 1076 4284 1124 4316
rect 1156 4284 1204 4316
rect 1236 4284 1284 4316
rect 1316 4284 1364 4316
rect 1396 4284 1444 4316
rect 1476 4284 1524 4316
rect 1556 4284 1684 4316
rect 1716 4284 1764 4316
rect 1796 4284 1844 4316
rect 1876 4284 1924 4316
rect 1956 4284 2004 4316
rect 2036 4284 2084 4316
rect 2116 4284 2164 4316
rect 2196 4284 2244 4316
rect 2276 4284 2324 4316
rect 2356 4284 2404 4316
rect 2436 4284 2484 4316
rect 2516 4284 2644 4316
rect 2676 4284 2724 4316
rect 2756 4284 2804 4316
rect 2836 4284 2884 4316
rect 2916 4284 2964 4316
rect 2996 4284 3044 4316
rect 3076 4284 3124 4316
rect 3156 4284 3204 4316
rect 3236 4284 3284 4316
rect 3316 4284 3364 4316
rect 3396 4284 3444 4316
rect 3476 4284 3604 4316
rect 3636 4284 3684 4316
rect 3716 4284 3764 4316
rect 3796 4284 3844 4316
rect 3876 4284 3924 4316
rect 3956 4284 3960 4316
rect 4080 4284 4084 4316
rect 4116 4284 4200 4316
rect 0 4240 120 4284
rect 240 4240 3960 4284
rect 4080 4240 4200 4284
rect 0 4236 4200 4240
rect 0 4204 84 4236
rect 116 4204 164 4236
rect 196 4204 244 4236
rect 276 4204 324 4236
rect 356 4204 404 4236
rect 436 4204 484 4236
rect 516 4204 564 4236
rect 596 4204 724 4236
rect 756 4204 804 4236
rect 836 4204 884 4236
rect 916 4204 964 4236
rect 996 4204 1044 4236
rect 1076 4204 1124 4236
rect 1156 4204 1204 4236
rect 1236 4204 1284 4236
rect 1316 4204 1364 4236
rect 1396 4204 1444 4236
rect 1476 4204 1524 4236
rect 1556 4204 1684 4236
rect 1716 4204 1764 4236
rect 1796 4204 1844 4236
rect 1876 4204 1924 4236
rect 1956 4204 2004 4236
rect 2036 4204 2084 4236
rect 2116 4204 2164 4236
rect 2196 4204 2244 4236
rect 2276 4204 2324 4236
rect 2356 4204 2404 4236
rect 2436 4204 2484 4236
rect 2516 4204 2644 4236
rect 2676 4204 2724 4236
rect 2756 4204 2804 4236
rect 2836 4204 2884 4236
rect 2916 4204 2964 4236
rect 2996 4204 3044 4236
rect 3076 4204 3124 4236
rect 3156 4204 3204 4236
rect 3236 4204 3284 4236
rect 3316 4204 3364 4236
rect 3396 4204 3444 4236
rect 3476 4204 3604 4236
rect 3636 4204 3684 4236
rect 3716 4204 3764 4236
rect 3796 4204 3844 4236
rect 3876 4204 3924 4236
rect 3956 4204 4004 4236
rect 4036 4204 4084 4236
rect 4116 4204 4200 4236
rect 0 4200 4200 4204
rect 0 4156 4200 4160
rect 0 4124 84 4156
rect 116 4124 164 4156
rect 196 4124 244 4156
rect 276 4124 324 4156
rect 356 4124 404 4156
rect 436 4124 484 4156
rect 516 4124 564 4156
rect 596 4124 724 4156
rect 756 4124 804 4156
rect 836 4124 884 4156
rect 916 4124 964 4156
rect 996 4124 1044 4156
rect 1076 4124 1124 4156
rect 1156 4124 1204 4156
rect 1236 4124 1284 4156
rect 1316 4124 1364 4156
rect 1396 4124 1444 4156
rect 1476 4124 1524 4156
rect 1556 4124 1684 4156
rect 1716 4124 1764 4156
rect 1796 4124 1844 4156
rect 1876 4124 1924 4156
rect 1956 4124 2004 4156
rect 2036 4124 2084 4156
rect 2116 4124 2164 4156
rect 2196 4124 2244 4156
rect 2276 4124 2324 4156
rect 2356 4124 2404 4156
rect 2436 4124 2484 4156
rect 2516 4124 2644 4156
rect 2676 4124 2724 4156
rect 2756 4124 2804 4156
rect 2836 4124 2884 4156
rect 2916 4124 2964 4156
rect 2996 4124 3044 4156
rect 3076 4124 3124 4156
rect 3156 4124 3204 4156
rect 3236 4124 3284 4156
rect 3316 4124 3364 4156
rect 3396 4124 3444 4156
rect 3476 4124 3604 4156
rect 3636 4124 3684 4156
rect 3716 4124 3764 4156
rect 3796 4124 3844 4156
rect 3876 4124 3924 4156
rect 3956 4124 4004 4156
rect 4036 4124 4084 4156
rect 4116 4124 4200 4156
rect 0 4120 4200 4124
rect 0 4076 1560 4120
rect 0 4044 84 4076
rect 116 4044 164 4076
rect 196 4044 244 4076
rect 276 4044 324 4076
rect 356 4044 404 4076
rect 436 4044 484 4076
rect 516 4044 564 4076
rect 596 4044 724 4076
rect 756 4044 804 4076
rect 836 4044 884 4076
rect 916 4044 964 4076
rect 996 4044 1044 4076
rect 1076 4044 1124 4076
rect 1156 4044 1204 4076
rect 1236 4044 1284 4076
rect 1316 4044 1364 4076
rect 1396 4044 1444 4076
rect 1476 4044 1524 4076
rect 1556 4044 1560 4076
rect 0 4000 1560 4044
rect 1680 4076 2520 4120
rect 1680 4044 1684 4076
rect 1716 4044 1764 4076
rect 1796 4044 1844 4076
rect 1876 4044 1924 4076
rect 1956 4044 2004 4076
rect 2036 4044 2084 4076
rect 2116 4044 2164 4076
rect 2196 4044 2244 4076
rect 2276 4044 2324 4076
rect 2356 4044 2404 4076
rect 2436 4044 2484 4076
rect 2516 4044 2520 4076
rect 1680 4000 2520 4044
rect 2640 4076 4200 4120
rect 2640 4044 2644 4076
rect 2676 4044 2724 4076
rect 2756 4044 2804 4076
rect 2836 4044 2884 4076
rect 2916 4044 2964 4076
rect 2996 4044 3044 4076
rect 3076 4044 3124 4076
rect 3156 4044 3204 4076
rect 3236 4044 3284 4076
rect 3316 4044 3364 4076
rect 3396 4044 3444 4076
rect 3476 4044 3604 4076
rect 3636 4044 3684 4076
rect 3716 4044 3764 4076
rect 3796 4044 3844 4076
rect 3876 4044 3924 4076
rect 3956 4044 4004 4076
rect 4036 4044 4084 4076
rect 4116 4044 4200 4076
rect 2640 4000 4200 4044
rect 0 3996 4200 4000
rect 0 3964 84 3996
rect 116 3964 164 3996
rect 196 3964 244 3996
rect 276 3964 324 3996
rect 356 3964 404 3996
rect 436 3964 484 3996
rect 516 3964 564 3996
rect 596 3964 724 3996
rect 756 3964 804 3996
rect 836 3964 884 3996
rect 916 3964 964 3996
rect 996 3964 1044 3996
rect 1076 3964 1124 3996
rect 1156 3964 1204 3996
rect 1236 3964 1284 3996
rect 1316 3964 1364 3996
rect 1396 3964 1444 3996
rect 1476 3964 1524 3996
rect 1556 3964 1684 3996
rect 1716 3964 1764 3996
rect 1796 3964 1844 3996
rect 1876 3964 1924 3996
rect 1956 3964 2004 3996
rect 2036 3964 2084 3996
rect 2116 3964 2164 3996
rect 2196 3964 2244 3996
rect 2276 3964 2324 3996
rect 2356 3964 2404 3996
rect 2436 3964 2484 3996
rect 2516 3964 2644 3996
rect 2676 3964 2724 3996
rect 2756 3964 2804 3996
rect 2836 3964 2884 3996
rect 2916 3964 2964 3996
rect 2996 3964 3044 3996
rect 3076 3964 3124 3996
rect 3156 3964 3204 3996
rect 3236 3964 3284 3996
rect 3316 3964 3364 3996
rect 3396 3964 3444 3996
rect 3476 3964 3604 3996
rect 3636 3964 3684 3996
rect 3716 3964 3764 3996
rect 3796 3964 3844 3996
rect 3876 3964 3924 3996
rect 3956 3964 4004 3996
rect 4036 3964 4084 3996
rect 4116 3964 4200 3996
rect 0 3960 4200 3964
rect 0 3851 4200 3880
rect 0 3769 164 3851
rect 196 3840 4200 3851
rect 196 3769 1560 3840
rect 0 3720 1560 3769
rect 1680 3720 2520 3840
rect 2640 3720 4200 3840
rect 0 3680 4200 3720
rect 0 3600 4200 3640
rect 0 3551 1560 3600
rect 0 3469 164 3551
rect 196 3480 1560 3551
rect 1680 3480 2520 3600
rect 2640 3480 4200 3600
rect 196 3469 4200 3480
rect 0 3440 4200 3469
rect 0 3356 4200 3360
rect 0 3324 84 3356
rect 116 3324 164 3356
rect 196 3324 244 3356
rect 276 3324 324 3356
rect 356 3324 404 3356
rect 436 3324 484 3356
rect 516 3324 564 3356
rect 596 3324 724 3356
rect 756 3324 804 3356
rect 836 3324 884 3356
rect 916 3324 964 3356
rect 996 3324 1044 3356
rect 1076 3324 1124 3356
rect 1156 3324 1204 3356
rect 1236 3324 1284 3356
rect 1316 3324 1364 3356
rect 1396 3324 1444 3356
rect 1476 3324 1524 3356
rect 1556 3324 1684 3356
rect 1716 3324 1764 3356
rect 1796 3324 1844 3356
rect 1876 3324 1924 3356
rect 1956 3324 2004 3356
rect 2036 3324 2084 3356
rect 2116 3324 2164 3356
rect 2196 3324 2244 3356
rect 2276 3324 2324 3356
rect 2356 3324 2404 3356
rect 2436 3324 2484 3356
rect 2516 3324 2644 3356
rect 2676 3324 2724 3356
rect 2756 3324 2804 3356
rect 2836 3324 2884 3356
rect 2916 3324 2964 3356
rect 2996 3324 3044 3356
rect 3076 3324 3124 3356
rect 3156 3324 3204 3356
rect 3236 3324 3284 3356
rect 3316 3324 3364 3356
rect 3396 3324 3444 3356
rect 3476 3324 3604 3356
rect 3636 3324 3684 3356
rect 3716 3324 3764 3356
rect 3796 3324 3844 3356
rect 3876 3324 3924 3356
rect 3956 3324 4084 3356
rect 4116 3324 4200 3356
rect 0 3320 4200 3324
rect 0 3276 1560 3320
rect 0 3244 84 3276
rect 116 3244 164 3276
rect 196 3244 244 3276
rect 276 3244 324 3276
rect 356 3244 404 3276
rect 436 3244 484 3276
rect 516 3244 564 3276
rect 596 3244 724 3276
rect 756 3244 804 3276
rect 836 3244 884 3276
rect 916 3244 964 3276
rect 996 3244 1044 3276
rect 1076 3244 1124 3276
rect 1156 3244 1204 3276
rect 1236 3244 1284 3276
rect 1316 3244 1364 3276
rect 1396 3244 1444 3276
rect 1476 3244 1524 3276
rect 1556 3244 1560 3276
rect 0 3200 1560 3244
rect 1680 3276 2520 3320
rect 1680 3244 1684 3276
rect 1716 3244 1764 3276
rect 1796 3244 1844 3276
rect 1876 3244 1924 3276
rect 1956 3244 2004 3276
rect 2036 3244 2084 3276
rect 2116 3244 2164 3276
rect 2196 3244 2244 3276
rect 2276 3244 2324 3276
rect 2356 3244 2404 3276
rect 2436 3244 2484 3276
rect 2516 3244 2520 3276
rect 1680 3200 2520 3244
rect 2640 3276 4200 3320
rect 2640 3244 2644 3276
rect 2676 3244 2724 3276
rect 2756 3244 2804 3276
rect 2836 3244 2884 3276
rect 2916 3244 2964 3276
rect 2996 3244 3044 3276
rect 3076 3244 3124 3276
rect 3156 3244 3204 3276
rect 3236 3244 3284 3276
rect 3316 3244 3364 3276
rect 3396 3244 3444 3276
rect 3476 3244 3604 3276
rect 3636 3244 3684 3276
rect 3716 3244 3764 3276
rect 3796 3244 3844 3276
rect 3876 3244 3924 3276
rect 3956 3244 4084 3276
rect 4116 3244 4200 3276
rect 2640 3200 4200 3244
rect 0 3196 4200 3200
rect 0 3164 84 3196
rect 116 3164 164 3196
rect 196 3164 244 3196
rect 276 3164 324 3196
rect 356 3164 404 3196
rect 436 3164 484 3196
rect 516 3164 564 3196
rect 596 3164 724 3196
rect 756 3164 804 3196
rect 836 3164 884 3196
rect 916 3164 964 3196
rect 996 3164 1044 3196
rect 1076 3164 1124 3196
rect 1156 3164 1204 3196
rect 1236 3164 1284 3196
rect 1316 3164 1364 3196
rect 1396 3164 1444 3196
rect 1476 3164 1524 3196
rect 1556 3164 1684 3196
rect 1716 3164 1764 3196
rect 1796 3164 1844 3196
rect 1876 3164 1924 3196
rect 1956 3164 2004 3196
rect 2036 3164 2084 3196
rect 2116 3164 2164 3196
rect 2196 3164 2244 3196
rect 2276 3164 2324 3196
rect 2356 3164 2404 3196
rect 2436 3164 2484 3196
rect 2516 3164 2644 3196
rect 2676 3164 2724 3196
rect 2756 3164 2804 3196
rect 2836 3164 2884 3196
rect 2916 3164 2964 3196
rect 2996 3164 3044 3196
rect 3076 3164 3124 3196
rect 3156 3164 3204 3196
rect 3236 3164 3284 3196
rect 3316 3164 3364 3196
rect 3396 3164 3444 3196
rect 3476 3164 3604 3196
rect 3636 3164 3684 3196
rect 3716 3164 3764 3196
rect 3796 3164 3844 3196
rect 3876 3164 3924 3196
rect 3956 3164 4084 3196
rect 4116 3164 4200 3196
rect 0 3160 4200 3164
rect 0 3116 4200 3120
rect 0 3084 84 3116
rect 116 3084 164 3116
rect 196 3084 244 3116
rect 276 3084 324 3116
rect 356 3084 404 3116
rect 436 3084 484 3116
rect 516 3084 564 3116
rect 596 3084 644 3116
rect 676 3084 724 3116
rect 756 3084 804 3116
rect 836 3084 884 3116
rect 916 3084 964 3116
rect 996 3084 1044 3116
rect 1076 3084 1124 3116
rect 1156 3084 1204 3116
rect 1236 3084 1284 3116
rect 1316 3084 1364 3116
rect 1396 3084 1444 3116
rect 1476 3084 1524 3116
rect 1556 3084 1604 3116
rect 1636 3084 1684 3116
rect 1716 3084 1764 3116
rect 1796 3084 1844 3116
rect 1876 3084 1924 3116
rect 1956 3084 2004 3116
rect 2036 3084 2084 3116
rect 2116 3084 2164 3116
rect 2196 3084 2244 3116
rect 2276 3084 2324 3116
rect 2356 3084 2404 3116
rect 2436 3084 2484 3116
rect 2516 3084 2564 3116
rect 2596 3084 2644 3116
rect 2676 3084 2724 3116
rect 2756 3084 2804 3116
rect 2836 3084 2884 3116
rect 2916 3084 2964 3116
rect 2996 3084 3044 3116
rect 3076 3084 3124 3116
rect 3156 3084 3204 3116
rect 3236 3084 3284 3116
rect 3316 3084 3364 3116
rect 3396 3084 3444 3116
rect 3476 3084 3524 3116
rect 3556 3084 3604 3116
rect 3636 3084 3684 3116
rect 3716 3084 3764 3116
rect 3796 3084 3844 3116
rect 3876 3084 3924 3116
rect 3956 3084 4084 3116
rect 4116 3084 4200 3116
rect 0 3080 4200 3084
rect 0 3036 600 3080
rect 720 3036 3480 3080
rect 3600 3036 4200 3080
rect 0 3004 84 3036
rect 116 3004 164 3036
rect 196 3004 244 3036
rect 276 3004 324 3036
rect 356 3004 404 3036
rect 436 3004 484 3036
rect 516 3004 564 3036
rect 596 3004 600 3036
rect 720 3004 724 3036
rect 756 3004 804 3036
rect 836 3004 884 3036
rect 916 3004 964 3036
rect 996 3004 1044 3036
rect 1076 3004 1124 3036
rect 1156 3004 1204 3036
rect 1236 3004 1284 3036
rect 1316 3004 1364 3036
rect 1396 3004 1444 3036
rect 1476 3004 1524 3036
rect 1556 3004 1604 3036
rect 1636 3004 1684 3036
rect 1716 3004 1764 3036
rect 1796 3004 1844 3036
rect 1876 3004 1924 3036
rect 1956 3004 2004 3036
rect 2036 3004 2084 3036
rect 2116 3004 2164 3036
rect 2196 3004 2244 3036
rect 2276 3004 2324 3036
rect 2356 3004 2404 3036
rect 2436 3004 2484 3036
rect 2516 3004 2564 3036
rect 2596 3004 2644 3036
rect 2676 3004 2724 3036
rect 2756 3004 2804 3036
rect 2836 3004 2884 3036
rect 2916 3004 2964 3036
rect 2996 3004 3044 3036
rect 3076 3004 3124 3036
rect 3156 3004 3204 3036
rect 3236 3004 3284 3036
rect 3316 3004 3364 3036
rect 3396 3004 3444 3036
rect 3476 3004 3480 3036
rect 3600 3004 3604 3036
rect 3636 3004 3684 3036
rect 3716 3004 3764 3036
rect 3796 3004 3844 3036
rect 3876 3004 3924 3036
rect 3956 3004 4084 3036
rect 4116 3004 4200 3036
rect 0 2960 600 3004
rect 720 2960 3480 3004
rect 3600 2960 4200 3004
rect 0 2956 4200 2960
rect 0 2924 84 2956
rect 116 2924 164 2956
rect 196 2924 244 2956
rect 276 2924 324 2956
rect 356 2924 404 2956
rect 436 2924 484 2956
rect 516 2924 564 2956
rect 596 2924 644 2956
rect 676 2924 724 2956
rect 756 2924 804 2956
rect 836 2924 884 2956
rect 916 2924 964 2956
rect 996 2924 1044 2956
rect 1076 2924 1124 2956
rect 1156 2924 1204 2956
rect 1236 2924 1284 2956
rect 1316 2924 1364 2956
rect 1396 2924 1444 2956
rect 1476 2924 1524 2956
rect 1556 2924 1604 2956
rect 1636 2924 1684 2956
rect 1716 2924 1764 2956
rect 1796 2924 1844 2956
rect 1876 2924 1924 2956
rect 1956 2924 2004 2956
rect 2036 2924 2084 2956
rect 2116 2924 2164 2956
rect 2196 2924 2244 2956
rect 2276 2924 2324 2956
rect 2356 2924 2404 2956
rect 2436 2924 2484 2956
rect 2516 2924 2564 2956
rect 2596 2924 2644 2956
rect 2676 2924 2724 2956
rect 2756 2924 2804 2956
rect 2836 2924 2884 2956
rect 2916 2924 2964 2956
rect 2996 2924 3044 2956
rect 3076 2924 3124 2956
rect 3156 2924 3204 2956
rect 3236 2924 3284 2956
rect 3316 2924 3364 2956
rect 3396 2924 3444 2956
rect 3476 2924 3524 2956
rect 3556 2924 3604 2956
rect 3636 2924 3684 2956
rect 3716 2924 3764 2956
rect 3796 2924 3844 2956
rect 3876 2924 3924 2956
rect 3956 2924 4084 2956
rect 4116 2924 4200 2956
rect 0 2920 4200 2924
rect 0 2876 4200 2880
rect 0 2844 84 2876
rect 116 2844 164 2876
rect 196 2844 244 2876
rect 276 2844 324 2876
rect 356 2844 404 2876
rect 436 2844 484 2876
rect 516 2844 564 2876
rect 596 2844 724 2876
rect 756 2844 804 2876
rect 836 2844 884 2876
rect 916 2844 964 2876
rect 996 2844 1044 2876
rect 1076 2844 1124 2876
rect 1156 2844 1204 2876
rect 1236 2844 1284 2876
rect 1316 2844 1364 2876
rect 1396 2844 1444 2876
rect 1476 2844 1524 2876
rect 1556 2844 1684 2876
rect 1716 2844 1764 2876
rect 1796 2844 1844 2876
rect 1876 2844 1924 2876
rect 1956 2844 2004 2876
rect 2036 2844 2084 2876
rect 2116 2844 2164 2876
rect 2196 2844 2244 2876
rect 2276 2844 2324 2876
rect 2356 2844 2404 2876
rect 2436 2844 2484 2876
rect 2516 2844 2644 2876
rect 2676 2844 2724 2876
rect 2756 2844 2804 2876
rect 2836 2844 2884 2876
rect 2916 2844 2964 2876
rect 2996 2844 3044 2876
rect 3076 2844 3124 2876
rect 3156 2844 3204 2876
rect 3236 2844 3284 2876
rect 3316 2844 3364 2876
rect 3396 2844 3444 2876
rect 3476 2844 3604 2876
rect 3636 2844 3684 2876
rect 3716 2844 3764 2876
rect 3796 2844 3844 2876
rect 3876 2844 3924 2876
rect 3956 2844 4084 2876
rect 4116 2844 4200 2876
rect 0 2840 4200 2844
rect 0 2796 120 2840
rect 240 2796 3960 2840
rect 0 2764 84 2796
rect 116 2764 120 2796
rect 240 2764 244 2796
rect 276 2764 324 2796
rect 356 2764 404 2796
rect 436 2764 484 2796
rect 516 2764 564 2796
rect 596 2764 724 2796
rect 756 2764 804 2796
rect 836 2764 884 2796
rect 916 2764 964 2796
rect 996 2764 1044 2796
rect 1076 2764 1124 2796
rect 1156 2764 1204 2796
rect 1236 2764 1284 2796
rect 1316 2764 1364 2796
rect 1396 2764 1444 2796
rect 1476 2764 1524 2796
rect 1556 2764 1684 2796
rect 1716 2764 1764 2796
rect 1796 2764 1844 2796
rect 1876 2764 1924 2796
rect 1956 2764 2004 2796
rect 2036 2764 2084 2796
rect 2116 2764 2164 2796
rect 2196 2764 2244 2796
rect 2276 2764 2324 2796
rect 2356 2764 2404 2796
rect 2436 2764 2484 2796
rect 2516 2764 2644 2796
rect 2676 2764 2724 2796
rect 2756 2764 2804 2796
rect 2836 2764 2884 2796
rect 2916 2764 2964 2796
rect 2996 2764 3044 2796
rect 3076 2764 3124 2796
rect 3156 2764 3204 2796
rect 3236 2764 3284 2796
rect 3316 2764 3364 2796
rect 3396 2764 3444 2796
rect 3476 2764 3604 2796
rect 3636 2764 3684 2796
rect 3716 2764 3764 2796
rect 3796 2764 3844 2796
rect 3876 2764 3924 2796
rect 3956 2764 3960 2796
rect 0 2720 120 2764
rect 240 2720 3960 2764
rect 4080 2796 4200 2840
rect 4080 2764 4084 2796
rect 4116 2764 4200 2796
rect 4080 2720 4200 2764
rect 0 2716 4200 2720
rect 0 2684 84 2716
rect 116 2684 164 2716
rect 196 2684 244 2716
rect 276 2684 324 2716
rect 356 2684 404 2716
rect 436 2684 484 2716
rect 516 2684 564 2716
rect 596 2684 724 2716
rect 756 2684 804 2716
rect 836 2684 884 2716
rect 916 2684 964 2716
rect 996 2684 1044 2716
rect 1076 2684 1124 2716
rect 1156 2684 1204 2716
rect 1236 2684 1284 2716
rect 1316 2684 1364 2716
rect 1396 2684 1444 2716
rect 1476 2684 1524 2716
rect 1556 2684 1684 2716
rect 1716 2684 1764 2716
rect 1796 2684 1844 2716
rect 1876 2684 1924 2716
rect 1956 2684 2004 2716
rect 2036 2684 2084 2716
rect 2116 2684 2164 2716
rect 2196 2684 2244 2716
rect 2276 2684 2324 2716
rect 2356 2684 2404 2716
rect 2436 2684 2484 2716
rect 2516 2684 2644 2716
rect 2676 2684 2724 2716
rect 2756 2684 2804 2716
rect 2836 2684 2884 2716
rect 2916 2684 2964 2716
rect 2996 2684 3044 2716
rect 3076 2684 3124 2716
rect 3156 2684 3204 2716
rect 3236 2684 3284 2716
rect 3316 2684 3364 2716
rect 3396 2684 3444 2716
rect 3476 2684 3604 2716
rect 3636 2684 3684 2716
rect 3716 2684 3764 2716
rect 3796 2684 3844 2716
rect 3876 2684 3924 2716
rect 3956 2684 4084 2716
rect 4116 2684 4200 2716
rect 0 2680 4200 2684
rect 0 2391 4200 2400
rect 0 2360 164 2391
rect 196 2360 4200 2391
rect 0 2240 120 2360
rect 240 2240 3960 2360
rect 4080 2240 4200 2360
rect 0 2209 164 2240
rect 196 2209 4200 2240
rect 0 2200 4200 2209
rect 0 1831 4200 1840
rect 0 1800 4004 1831
rect 4036 1800 4200 1831
rect 0 1680 120 1800
rect 240 1680 3960 1800
rect 4080 1680 4200 1800
rect 0 1649 4004 1680
rect 4036 1649 4200 1680
rect 0 1640 4200 1649
rect 0 1396 4200 1400
rect 0 1364 4 1396
rect 36 1364 84 1396
rect 116 1364 164 1396
rect 196 1364 244 1396
rect 276 1364 324 1396
rect 356 1364 404 1396
rect 436 1364 484 1396
rect 516 1364 564 1396
rect 596 1364 724 1396
rect 756 1364 804 1396
rect 836 1364 884 1396
rect 916 1364 964 1396
rect 996 1364 1044 1396
rect 1076 1364 1124 1396
rect 1156 1364 1204 1396
rect 1236 1364 1284 1396
rect 1316 1364 1364 1396
rect 1396 1364 1444 1396
rect 1476 1364 1524 1396
rect 1556 1364 1684 1396
rect 1716 1364 1764 1396
rect 1796 1364 1844 1396
rect 1876 1364 1924 1396
rect 1956 1364 2004 1396
rect 2036 1364 2084 1396
rect 2116 1364 2164 1396
rect 2196 1364 2244 1396
rect 2276 1364 2324 1396
rect 2356 1364 2404 1396
rect 2436 1364 2484 1396
rect 2516 1364 2644 1396
rect 2676 1364 2724 1396
rect 2756 1364 2804 1396
rect 2836 1364 2884 1396
rect 2916 1364 2964 1396
rect 2996 1364 3044 1396
rect 3076 1364 3124 1396
rect 3156 1364 3204 1396
rect 3236 1364 3284 1396
rect 3316 1364 3364 1396
rect 3396 1364 3444 1396
rect 3476 1364 3604 1396
rect 3636 1364 3684 1396
rect 3716 1364 3764 1396
rect 3796 1364 3844 1396
rect 3876 1364 3924 1396
rect 3956 1364 4004 1396
rect 4036 1364 4084 1396
rect 4116 1364 4164 1396
rect 4196 1364 4200 1396
rect 0 1360 4200 1364
rect 0 1240 600 1360
rect 720 1240 3480 1360
rect 3600 1240 4200 1360
rect 0 1236 4200 1240
rect 0 1204 4 1236
rect 36 1204 84 1236
rect 116 1204 164 1236
rect 196 1204 244 1236
rect 276 1204 324 1236
rect 356 1204 404 1236
rect 436 1204 484 1236
rect 516 1204 564 1236
rect 596 1204 724 1236
rect 756 1204 804 1236
rect 836 1204 884 1236
rect 916 1204 964 1236
rect 996 1204 1044 1236
rect 1076 1204 1124 1236
rect 1156 1204 1204 1236
rect 1236 1204 1284 1236
rect 1316 1204 1364 1236
rect 1396 1204 1444 1236
rect 1476 1204 1524 1236
rect 1556 1204 1684 1236
rect 1716 1204 1764 1236
rect 1796 1204 1844 1236
rect 1876 1204 1924 1236
rect 1956 1204 2004 1236
rect 2036 1204 2084 1236
rect 2116 1204 2164 1236
rect 2196 1204 2244 1236
rect 2276 1204 2324 1236
rect 2356 1204 2404 1236
rect 2436 1204 2484 1236
rect 2516 1204 2644 1236
rect 2676 1204 2724 1236
rect 2756 1204 2804 1236
rect 2836 1204 2884 1236
rect 2916 1204 2964 1236
rect 2996 1204 3044 1236
rect 3076 1204 3124 1236
rect 3156 1204 3204 1236
rect 3236 1204 3284 1236
rect 3316 1204 3364 1236
rect 3396 1204 3444 1236
rect 3476 1204 3604 1236
rect 3636 1204 3684 1236
rect 3716 1204 3764 1236
rect 3796 1204 3844 1236
rect 3876 1204 3924 1236
rect 3956 1204 4004 1236
rect 4036 1204 4084 1236
rect 4116 1204 4164 1236
rect 4196 1204 4200 1236
rect 0 1200 4200 1204
rect 0 556 4200 560
rect 0 524 84 556
rect 116 524 164 556
rect 196 524 244 556
rect 276 524 324 556
rect 356 524 404 556
rect 436 524 484 556
rect 516 524 564 556
rect 596 524 724 556
rect 756 524 804 556
rect 836 524 884 556
rect 916 524 964 556
rect 996 524 1044 556
rect 1076 524 1124 556
rect 1156 524 1204 556
rect 1236 524 1284 556
rect 1316 524 1364 556
rect 1396 524 1444 556
rect 1476 524 1524 556
rect 1556 524 1684 556
rect 1716 524 1764 556
rect 1796 524 1844 556
rect 1876 524 1924 556
rect 1956 524 2004 556
rect 2036 524 2084 556
rect 2116 524 2164 556
rect 2196 524 2244 556
rect 2276 524 2324 556
rect 2356 524 2404 556
rect 2436 524 2484 556
rect 2516 524 2644 556
rect 2676 524 2724 556
rect 2756 524 2804 556
rect 2836 524 2884 556
rect 2916 524 2964 556
rect 2996 524 3044 556
rect 3076 524 3124 556
rect 3156 524 3204 556
rect 3236 524 3284 556
rect 3316 524 3364 556
rect 3396 524 3444 556
rect 3476 524 3604 556
rect 3636 524 3684 556
rect 3716 524 3764 556
rect 3796 524 3844 556
rect 3876 524 3924 556
rect 3956 524 4084 556
rect 4116 524 4200 556
rect 0 520 4200 524
rect 0 476 1080 520
rect 1200 476 2040 520
rect 2160 476 3000 520
rect 3120 476 4200 520
rect 0 444 84 476
rect 116 444 164 476
rect 196 444 244 476
rect 276 444 324 476
rect 356 444 404 476
rect 436 444 484 476
rect 516 444 564 476
rect 596 444 724 476
rect 756 444 804 476
rect 836 444 884 476
rect 916 444 964 476
rect 996 444 1044 476
rect 1076 444 1080 476
rect 1200 444 1204 476
rect 1236 444 1284 476
rect 1316 444 1364 476
rect 1396 444 1444 476
rect 1476 444 1524 476
rect 1556 444 1684 476
rect 1716 444 1764 476
rect 1796 444 1844 476
rect 1876 444 1924 476
rect 1956 444 2004 476
rect 2036 444 2040 476
rect 2160 444 2164 476
rect 2196 444 2244 476
rect 2276 444 2324 476
rect 2356 444 2404 476
rect 2436 444 2484 476
rect 2516 444 2644 476
rect 2676 444 2724 476
rect 2756 444 2804 476
rect 2836 444 2884 476
rect 2916 444 2964 476
rect 2996 444 3000 476
rect 3120 444 3124 476
rect 3156 444 3204 476
rect 3236 444 3284 476
rect 3316 444 3364 476
rect 3396 444 3444 476
rect 3476 444 3604 476
rect 3636 444 3684 476
rect 3716 444 3764 476
rect 3796 444 3844 476
rect 3876 444 3924 476
rect 3956 444 4084 476
rect 4116 444 4200 476
rect 0 400 1080 444
rect 1200 400 2040 444
rect 2160 400 3000 444
rect 3120 400 4200 444
rect 0 396 4200 400
rect 0 364 84 396
rect 116 364 164 396
rect 196 364 244 396
rect 276 364 324 396
rect 356 364 404 396
rect 436 364 484 396
rect 516 364 564 396
rect 596 364 724 396
rect 756 364 804 396
rect 836 364 884 396
rect 916 364 964 396
rect 996 364 1044 396
rect 1076 364 1124 396
rect 1156 364 1204 396
rect 1236 364 1284 396
rect 1316 364 1364 396
rect 1396 364 1444 396
rect 1476 364 1524 396
rect 1556 364 1684 396
rect 1716 364 1764 396
rect 1796 364 1844 396
rect 1876 364 1924 396
rect 1956 364 2004 396
rect 2036 364 2084 396
rect 2116 364 2164 396
rect 2196 364 2244 396
rect 2276 364 2324 396
rect 2356 364 2404 396
rect 2436 364 2484 396
rect 2516 364 2644 396
rect 2676 364 2724 396
rect 2756 364 2804 396
rect 2836 364 2884 396
rect 2916 364 2964 396
rect 2996 364 3044 396
rect 3076 364 3124 396
rect 3156 364 3204 396
rect 3236 364 3284 396
rect 3316 364 3364 396
rect 3396 364 3444 396
rect 3476 364 3604 396
rect 3636 364 3684 396
rect 3716 364 3764 396
rect 3796 364 3844 396
rect 3876 364 3924 396
rect 3956 364 4084 396
rect 4116 364 4200 396
rect 0 360 4200 364
rect 0 171 4200 200
rect 0 89 164 171
rect 196 160 4200 171
rect 196 89 1560 160
rect 0 40 1560 89
rect 1680 40 2520 160
rect 2640 40 4200 160
rect 0 0 4200 40
rect 0 -44 4200 -40
rect 0 -76 84 -44
rect 116 -76 164 -44
rect 196 -76 244 -44
rect 276 -76 324 -44
rect 356 -76 404 -44
rect 436 -76 484 -44
rect 516 -76 564 -44
rect 596 -76 724 -44
rect 756 -76 804 -44
rect 836 -76 884 -44
rect 916 -76 964 -44
rect 996 -76 1044 -44
rect 1076 -76 1124 -44
rect 1156 -76 1204 -44
rect 1236 -76 1284 -44
rect 1316 -76 1364 -44
rect 1396 -76 1444 -44
rect 1476 -76 1524 -44
rect 1556 -76 1684 -44
rect 1716 -76 1764 -44
rect 1796 -76 1844 -44
rect 1876 -76 1924 -44
rect 1956 -76 2004 -44
rect 2036 -76 2084 -44
rect 2116 -76 2164 -44
rect 2196 -76 2244 -44
rect 2276 -76 2324 -44
rect 2356 -76 2404 -44
rect 2436 -76 2484 -44
rect 2516 -76 2644 -44
rect 2676 -76 2724 -44
rect 2756 -76 2804 -44
rect 2836 -76 2884 -44
rect 2916 -76 2964 -44
rect 2996 -76 3044 -44
rect 3076 -76 3124 -44
rect 3156 -76 3204 -44
rect 3236 -76 3284 -44
rect 3316 -76 3364 -44
rect 3396 -76 3444 -44
rect 3476 -76 3604 -44
rect 3636 -76 3684 -44
rect 3716 -76 3764 -44
rect 3796 -76 3844 -44
rect 3876 -76 3924 -44
rect 3956 -76 4084 -44
rect 4116 -76 4200 -44
rect 0 -80 4200 -76
rect 0 -124 1560 -80
rect 0 -156 84 -124
rect 116 -156 164 -124
rect 196 -156 244 -124
rect 276 -156 324 -124
rect 356 -156 404 -124
rect 436 -156 484 -124
rect 516 -156 564 -124
rect 596 -156 724 -124
rect 756 -156 804 -124
rect 836 -156 884 -124
rect 916 -156 964 -124
rect 996 -156 1044 -124
rect 1076 -156 1124 -124
rect 1156 -156 1204 -124
rect 1236 -156 1284 -124
rect 1316 -156 1364 -124
rect 1396 -156 1444 -124
rect 1476 -156 1524 -124
rect 1556 -156 1560 -124
rect 0 -200 1560 -156
rect 1680 -124 2520 -80
rect 1680 -156 1684 -124
rect 1716 -156 1764 -124
rect 1796 -156 1844 -124
rect 1876 -156 1924 -124
rect 1956 -156 2004 -124
rect 2036 -156 2084 -124
rect 2116 -156 2164 -124
rect 2196 -156 2244 -124
rect 2276 -156 2324 -124
rect 2356 -156 2404 -124
rect 2436 -156 2484 -124
rect 2516 -156 2520 -124
rect 1680 -200 2520 -156
rect 2640 -124 4200 -80
rect 2640 -156 2644 -124
rect 2676 -156 2724 -124
rect 2756 -156 2804 -124
rect 2836 -156 2884 -124
rect 2916 -156 2964 -124
rect 2996 -156 3044 -124
rect 3076 -156 3124 -124
rect 3156 -156 3204 -124
rect 3236 -156 3284 -124
rect 3316 -156 3364 -124
rect 3396 -156 3444 -124
rect 3476 -156 3604 -124
rect 3636 -156 3684 -124
rect 3716 -156 3764 -124
rect 3796 -156 3844 -124
rect 3876 -156 3924 -124
rect 3956 -156 4084 -124
rect 4116 -156 4200 -124
rect 2640 -200 4200 -156
rect 0 -204 4200 -200
rect 0 -236 84 -204
rect 116 -236 164 -204
rect 196 -236 244 -204
rect 276 -236 324 -204
rect 356 -236 404 -204
rect 436 -236 484 -204
rect 516 -236 564 -204
rect 596 -236 724 -204
rect 756 -236 804 -204
rect 836 -236 884 -204
rect 916 -236 964 -204
rect 996 -236 1044 -204
rect 1076 -236 1124 -204
rect 1156 -236 1204 -204
rect 1236 -236 1284 -204
rect 1316 -236 1364 -204
rect 1396 -236 1444 -204
rect 1476 -236 1524 -204
rect 1556 -236 1684 -204
rect 1716 -236 1764 -204
rect 1796 -236 1844 -204
rect 1876 -236 1924 -204
rect 1956 -236 2004 -204
rect 2036 -236 2084 -204
rect 2116 -236 2164 -204
rect 2196 -236 2244 -204
rect 2276 -236 2324 -204
rect 2356 -236 2404 -204
rect 2436 -236 2484 -204
rect 2516 -236 2644 -204
rect 2676 -236 2724 -204
rect 2756 -236 2804 -204
rect 2836 -236 2884 -204
rect 2916 -236 2964 -204
rect 2996 -236 3044 -204
rect 3076 -236 3124 -204
rect 3156 -236 3204 -204
rect 3236 -236 3284 -204
rect 3316 -236 3364 -204
rect 3396 -236 3444 -204
rect 3476 -236 3604 -204
rect 3636 -236 3684 -204
rect 3716 -236 3764 -204
rect 3796 -236 3844 -204
rect 3876 -236 3924 -204
rect 3956 -236 4084 -204
rect 4116 -236 4200 -204
rect 0 -240 4200 -236
rect 0 -349 4200 -320
rect 0 -431 164 -349
rect 196 -360 4200 -349
rect 196 -431 1560 -360
rect 0 -480 1560 -431
rect 1680 -480 2520 -360
rect 2640 -480 4200 -360
rect 0 -520 4200 -480
<< via4 >>
rect 120 4720 164 4840
rect 164 4720 196 4840
rect 196 4720 240 4840
rect 3960 4720 4080 4840
rect 120 4316 240 4360
rect 3960 4316 4080 4360
rect 120 4284 164 4316
rect 164 4284 196 4316
rect 196 4284 240 4316
rect 3960 4284 4004 4316
rect 4004 4284 4036 4316
rect 4036 4284 4080 4316
rect 120 4240 240 4284
rect 3960 4240 4080 4284
rect 1560 4000 1680 4120
rect 2520 4000 2640 4120
rect 1560 3720 1680 3840
rect 2520 3720 2640 3840
rect 1560 3480 1680 3600
rect 2520 3480 2640 3600
rect 1560 3200 1680 3320
rect 2520 3200 2640 3320
rect 600 3036 720 3080
rect 3480 3036 3600 3080
rect 600 3004 644 3036
rect 644 3004 676 3036
rect 676 3004 720 3036
rect 3480 3004 3524 3036
rect 3524 3004 3556 3036
rect 3556 3004 3600 3036
rect 600 2960 720 3004
rect 3480 2960 3600 3004
rect 120 2796 240 2840
rect 120 2764 164 2796
rect 164 2764 196 2796
rect 196 2764 240 2796
rect 120 2720 240 2764
rect 3960 2720 4080 2840
rect 120 2240 164 2360
rect 164 2240 196 2360
rect 196 2240 240 2360
rect 3960 2240 4080 2360
rect 120 1680 240 1800
rect 3960 1680 4004 1800
rect 4004 1680 4036 1800
rect 4036 1680 4080 1800
rect 600 1240 720 1360
rect 3480 1240 3600 1360
rect 1080 476 1200 520
rect 2040 476 2160 520
rect 3000 476 3120 520
rect 1080 444 1124 476
rect 1124 444 1156 476
rect 1156 444 1200 476
rect 2040 444 2084 476
rect 2084 444 2116 476
rect 2116 444 2160 476
rect 3000 444 3044 476
rect 3044 444 3076 476
rect 3076 444 3120 476
rect 1080 400 1200 444
rect 2040 400 2160 444
rect 3000 400 3120 444
rect 1560 40 1680 160
rect 2520 40 2640 160
rect 1560 -200 1680 -80
rect 2520 -200 2640 -80
rect 1560 -480 1680 -360
rect 2520 -480 2640 -360
<< metal5 >>
rect 80 4840 280 5040
rect 80 4720 120 4840
rect 240 4720 280 4840
rect 80 4360 280 4720
rect 80 4240 120 4360
rect 240 4240 280 4360
rect 80 2840 280 4240
rect 80 2720 120 2840
rect 240 2720 280 2840
rect 80 2360 280 2720
rect 80 2240 120 2360
rect 240 2240 280 2360
rect 80 1800 280 2240
rect 80 1680 120 1800
rect 240 1680 280 1800
rect 80 -520 280 1680
rect 560 3080 760 5040
rect 560 2960 600 3080
rect 720 2960 760 3080
rect 560 1360 760 2960
rect 560 1240 600 1360
rect 720 1240 760 1360
rect 560 -520 760 1240
rect 1040 520 1240 5040
rect 1040 400 1080 520
rect 1200 400 1240 520
rect 1040 -520 1240 400
rect 1520 4120 1720 5040
rect 1520 4000 1560 4120
rect 1680 4000 1720 4120
rect 1520 3840 1720 4000
rect 1520 3720 1560 3840
rect 1680 3720 1720 3840
rect 1520 3600 1720 3720
rect 1520 3480 1560 3600
rect 1680 3480 1720 3600
rect 1520 3320 1720 3480
rect 1520 3200 1560 3320
rect 1680 3200 1720 3320
rect 1520 160 1720 3200
rect 1520 40 1560 160
rect 1680 40 1720 160
rect 1520 -80 1720 40
rect 1520 -200 1560 -80
rect 1680 -200 1720 -80
rect 1520 -360 1720 -200
rect 1520 -480 1560 -360
rect 1680 -480 1720 -360
rect 1520 -520 1720 -480
rect 2000 520 2200 5040
rect 2000 400 2040 520
rect 2160 400 2200 520
rect 2000 -520 2200 400
rect 2480 4120 2680 5040
rect 2480 4000 2520 4120
rect 2640 4000 2680 4120
rect 2480 3840 2680 4000
rect 2480 3720 2520 3840
rect 2640 3720 2680 3840
rect 2480 3600 2680 3720
rect 2480 3480 2520 3600
rect 2640 3480 2680 3600
rect 2480 3320 2680 3480
rect 2480 3200 2520 3320
rect 2640 3200 2680 3320
rect 2480 160 2680 3200
rect 2480 40 2520 160
rect 2640 40 2680 160
rect 2480 -80 2680 40
rect 2480 -200 2520 -80
rect 2640 -200 2680 -80
rect 2480 -360 2680 -200
rect 2480 -480 2520 -360
rect 2640 -480 2680 -360
rect 2480 -520 2680 -480
rect 2960 520 3160 5040
rect 2960 400 3000 520
rect 3120 400 3160 520
rect 2960 -520 3160 400
rect 3440 3080 3640 5040
rect 3440 2960 3480 3080
rect 3600 2960 3640 3080
rect 3440 1360 3640 2960
rect 3440 1240 3480 1360
rect 3600 1240 3640 1360
rect 3440 -520 3640 1240
rect 3920 4840 4120 5040
rect 3920 4720 3960 4840
rect 4080 4720 4120 4840
rect 3920 4360 4120 4720
rect 3920 4240 3960 4360
rect 4080 4240 4120 4360
rect 3920 2840 4120 4240
rect 3920 2720 3960 2840
rect 4080 2720 4120 2840
rect 3920 2360 4120 2720
rect 3920 2240 3960 2360
rect 4080 2240 4120 2360
rect 3920 1800 4120 2240
rect 3920 1680 3960 1800
rect 4080 1680 4120 1800
rect 3920 -520 4120 1680
<< labels >>
rlabel metal2 0 -160 4200 -120 0 na
port 3 nsew
rlabel metal2 0 360 4200 400 0 qa
port 5 nsew
rlabel metal2 0 1280 4200 1320 0 bpa
port 0 nsew
rlabel metal2 0 2760 4200 2800 0 xa
port 10 nsew
rlabel metal2 0 3000 4200 3040 0 bpb
port 1 nsew
rlabel metal2 0 3240 4200 3280 0 nb
port 4 nsew
rlabel metal5 80 -520 280 5040 0 vdda
port 7 nsew
rlabel metal5 560 -520 760 5040 0 vddx
port 8 nsew
rlabel metal5 1040 -520 1240 5040 0 gnda
port 2 nsew
rlabel metal5 1520 -520 1720 5040 0 vssa
port 9 nsew
rlabel metal1 1120 -440 1160 -340 0 na1
rlabel metal1 2080 -440 2120 -340 0 na2
rlabel metal1 3040 -440 3080 -340 0 na3
rlabel metal1 1120 80 1160 180 0 qa1
rlabel metal1 2080 80 2120 180 0 qa2
rlabel metal1 3040 80 3080 180 0 qa3
rlabel metal1 3040 820 3080 1120 0 qa4
rlabel metal1 2080 820 2120 1120 0 qa5
rlabel metal1 1120 820 1160 1120 0 qa6
rlabel metal1 3040 1540 3080 1840 0 bpa1
rlabel metal1 2080 1540 2120 1840 0 bpa2
rlabel metal1 1120 1540 1160 1840 0 bpa3
rlabel metal1 1120 2200 1160 2500 0 xa1
rlabel metal1 2080 2200 2120 2500 0 xa2
rlabel metal1 3040 2200 3080 2500 0 xa3
rlabel metal1 1120 3460 1160 3560 0 nb1
rlabel metal1 2080 3460 2120 3560 0 nb2
rlabel metal1 3040 3460 3080 3560 0 nb3
rlabel metal1 1120 3760 1160 3860 0 qb1
rlabel metal1 2080 3760 2120 3860 0 qb2
rlabel metal1 3040 3760 3080 3860 0 qb3
rlabel metal1 1120 4580 1160 4880 0 xb1
rlabel metal1 2080 4580 2120 4880 0 xb2
rlabel metal1 3040 4580 3080 4880 0 xb3
rlabel metal2 0 4280 4200 4320 0 xb
port 11 nsew
rlabel metal2 0 4040 4200 4080 0 qb
port 6 nsew
<< end >>
