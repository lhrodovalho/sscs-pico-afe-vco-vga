magic
tech sky130A
magscale 1 2
timestamp 1634821592
<< error_p >>
rect -607 -638 -549 -632
rect -607 -672 -595 -638
rect -607 -678 -549 -672
<< pwell >>
rect -631 -526 631 526
<< nmos >>
rect -543 -500 -513 500
rect -447 -500 -417 500
rect -351 -500 -321 500
rect -255 -500 -225 500
rect -159 -500 -129 500
rect -63 -500 -33 500
rect 33 -500 63 500
rect 129 -500 159 500
rect 225 -500 255 500
rect 321 -500 351 500
rect 417 -500 447 500
rect 513 -500 543 500
<< ndiff >>
rect -605 459 -543 500
rect -605 425 -593 459
rect -559 425 -543 459
rect -605 391 -543 425
rect -605 357 -593 391
rect -559 357 -543 391
rect -605 323 -543 357
rect -605 289 -593 323
rect -559 289 -543 323
rect -605 255 -543 289
rect -605 221 -593 255
rect -559 221 -543 255
rect -605 187 -543 221
rect -605 153 -593 187
rect -559 153 -543 187
rect -605 119 -543 153
rect -605 85 -593 119
rect -559 85 -543 119
rect -605 51 -543 85
rect -605 17 -593 51
rect -559 17 -543 51
rect -605 -17 -543 17
rect -605 -51 -593 -17
rect -559 -51 -543 -17
rect -605 -85 -543 -51
rect -605 -119 -593 -85
rect -559 -119 -543 -85
rect -605 -153 -543 -119
rect -605 -187 -593 -153
rect -559 -187 -543 -153
rect -605 -221 -543 -187
rect -605 -255 -593 -221
rect -559 -255 -543 -221
rect -605 -289 -543 -255
rect -605 -323 -593 -289
rect -559 -323 -543 -289
rect -605 -357 -543 -323
rect -605 -391 -593 -357
rect -559 -391 -543 -357
rect -605 -425 -543 -391
rect -605 -459 -593 -425
rect -559 -459 -543 -425
rect -605 -500 -543 -459
rect -513 459 -447 500
rect -513 425 -497 459
rect -463 425 -447 459
rect -513 391 -447 425
rect -513 357 -497 391
rect -463 357 -447 391
rect -513 323 -447 357
rect -513 289 -497 323
rect -463 289 -447 323
rect -513 255 -447 289
rect -513 221 -497 255
rect -463 221 -447 255
rect -513 187 -447 221
rect -513 153 -497 187
rect -463 153 -447 187
rect -513 119 -447 153
rect -513 85 -497 119
rect -463 85 -447 119
rect -513 51 -447 85
rect -513 17 -497 51
rect -463 17 -447 51
rect -513 -17 -447 17
rect -513 -51 -497 -17
rect -463 -51 -447 -17
rect -513 -85 -447 -51
rect -513 -119 -497 -85
rect -463 -119 -447 -85
rect -513 -153 -447 -119
rect -513 -187 -497 -153
rect -463 -187 -447 -153
rect -513 -221 -447 -187
rect -513 -255 -497 -221
rect -463 -255 -447 -221
rect -513 -289 -447 -255
rect -513 -323 -497 -289
rect -463 -323 -447 -289
rect -513 -357 -447 -323
rect -513 -391 -497 -357
rect -463 -391 -447 -357
rect -513 -425 -447 -391
rect -513 -459 -497 -425
rect -463 -459 -447 -425
rect -513 -500 -447 -459
rect -417 459 -351 500
rect -417 425 -401 459
rect -367 425 -351 459
rect -417 391 -351 425
rect -417 357 -401 391
rect -367 357 -351 391
rect -417 323 -351 357
rect -417 289 -401 323
rect -367 289 -351 323
rect -417 255 -351 289
rect -417 221 -401 255
rect -367 221 -351 255
rect -417 187 -351 221
rect -417 153 -401 187
rect -367 153 -351 187
rect -417 119 -351 153
rect -417 85 -401 119
rect -367 85 -351 119
rect -417 51 -351 85
rect -417 17 -401 51
rect -367 17 -351 51
rect -417 -17 -351 17
rect -417 -51 -401 -17
rect -367 -51 -351 -17
rect -417 -85 -351 -51
rect -417 -119 -401 -85
rect -367 -119 -351 -85
rect -417 -153 -351 -119
rect -417 -187 -401 -153
rect -367 -187 -351 -153
rect -417 -221 -351 -187
rect -417 -255 -401 -221
rect -367 -255 -351 -221
rect -417 -289 -351 -255
rect -417 -323 -401 -289
rect -367 -323 -351 -289
rect -417 -357 -351 -323
rect -417 -391 -401 -357
rect -367 -391 -351 -357
rect -417 -425 -351 -391
rect -417 -459 -401 -425
rect -367 -459 -351 -425
rect -417 -500 -351 -459
rect -321 459 -255 500
rect -321 425 -305 459
rect -271 425 -255 459
rect -321 391 -255 425
rect -321 357 -305 391
rect -271 357 -255 391
rect -321 323 -255 357
rect -321 289 -305 323
rect -271 289 -255 323
rect -321 255 -255 289
rect -321 221 -305 255
rect -271 221 -255 255
rect -321 187 -255 221
rect -321 153 -305 187
rect -271 153 -255 187
rect -321 119 -255 153
rect -321 85 -305 119
rect -271 85 -255 119
rect -321 51 -255 85
rect -321 17 -305 51
rect -271 17 -255 51
rect -321 -17 -255 17
rect -321 -51 -305 -17
rect -271 -51 -255 -17
rect -321 -85 -255 -51
rect -321 -119 -305 -85
rect -271 -119 -255 -85
rect -321 -153 -255 -119
rect -321 -187 -305 -153
rect -271 -187 -255 -153
rect -321 -221 -255 -187
rect -321 -255 -305 -221
rect -271 -255 -255 -221
rect -321 -289 -255 -255
rect -321 -323 -305 -289
rect -271 -323 -255 -289
rect -321 -357 -255 -323
rect -321 -391 -305 -357
rect -271 -391 -255 -357
rect -321 -425 -255 -391
rect -321 -459 -305 -425
rect -271 -459 -255 -425
rect -321 -500 -255 -459
rect -225 459 -159 500
rect -225 425 -209 459
rect -175 425 -159 459
rect -225 391 -159 425
rect -225 357 -209 391
rect -175 357 -159 391
rect -225 323 -159 357
rect -225 289 -209 323
rect -175 289 -159 323
rect -225 255 -159 289
rect -225 221 -209 255
rect -175 221 -159 255
rect -225 187 -159 221
rect -225 153 -209 187
rect -175 153 -159 187
rect -225 119 -159 153
rect -225 85 -209 119
rect -175 85 -159 119
rect -225 51 -159 85
rect -225 17 -209 51
rect -175 17 -159 51
rect -225 -17 -159 17
rect -225 -51 -209 -17
rect -175 -51 -159 -17
rect -225 -85 -159 -51
rect -225 -119 -209 -85
rect -175 -119 -159 -85
rect -225 -153 -159 -119
rect -225 -187 -209 -153
rect -175 -187 -159 -153
rect -225 -221 -159 -187
rect -225 -255 -209 -221
rect -175 -255 -159 -221
rect -225 -289 -159 -255
rect -225 -323 -209 -289
rect -175 -323 -159 -289
rect -225 -357 -159 -323
rect -225 -391 -209 -357
rect -175 -391 -159 -357
rect -225 -425 -159 -391
rect -225 -459 -209 -425
rect -175 -459 -159 -425
rect -225 -500 -159 -459
rect -129 459 -63 500
rect -129 425 -113 459
rect -79 425 -63 459
rect -129 391 -63 425
rect -129 357 -113 391
rect -79 357 -63 391
rect -129 323 -63 357
rect -129 289 -113 323
rect -79 289 -63 323
rect -129 255 -63 289
rect -129 221 -113 255
rect -79 221 -63 255
rect -129 187 -63 221
rect -129 153 -113 187
rect -79 153 -63 187
rect -129 119 -63 153
rect -129 85 -113 119
rect -79 85 -63 119
rect -129 51 -63 85
rect -129 17 -113 51
rect -79 17 -63 51
rect -129 -17 -63 17
rect -129 -51 -113 -17
rect -79 -51 -63 -17
rect -129 -85 -63 -51
rect -129 -119 -113 -85
rect -79 -119 -63 -85
rect -129 -153 -63 -119
rect -129 -187 -113 -153
rect -79 -187 -63 -153
rect -129 -221 -63 -187
rect -129 -255 -113 -221
rect -79 -255 -63 -221
rect -129 -289 -63 -255
rect -129 -323 -113 -289
rect -79 -323 -63 -289
rect -129 -357 -63 -323
rect -129 -391 -113 -357
rect -79 -391 -63 -357
rect -129 -425 -63 -391
rect -129 -459 -113 -425
rect -79 -459 -63 -425
rect -129 -500 -63 -459
rect -33 459 33 500
rect -33 425 -17 459
rect 17 425 33 459
rect -33 391 33 425
rect -33 357 -17 391
rect 17 357 33 391
rect -33 323 33 357
rect -33 289 -17 323
rect 17 289 33 323
rect -33 255 33 289
rect -33 221 -17 255
rect 17 221 33 255
rect -33 187 33 221
rect -33 153 -17 187
rect 17 153 33 187
rect -33 119 33 153
rect -33 85 -17 119
rect 17 85 33 119
rect -33 51 33 85
rect -33 17 -17 51
rect 17 17 33 51
rect -33 -17 33 17
rect -33 -51 -17 -17
rect 17 -51 33 -17
rect -33 -85 33 -51
rect -33 -119 -17 -85
rect 17 -119 33 -85
rect -33 -153 33 -119
rect -33 -187 -17 -153
rect 17 -187 33 -153
rect -33 -221 33 -187
rect -33 -255 -17 -221
rect 17 -255 33 -221
rect -33 -289 33 -255
rect -33 -323 -17 -289
rect 17 -323 33 -289
rect -33 -357 33 -323
rect -33 -391 -17 -357
rect 17 -391 33 -357
rect -33 -425 33 -391
rect -33 -459 -17 -425
rect 17 -459 33 -425
rect -33 -500 33 -459
rect 63 459 129 500
rect 63 425 79 459
rect 113 425 129 459
rect 63 391 129 425
rect 63 357 79 391
rect 113 357 129 391
rect 63 323 129 357
rect 63 289 79 323
rect 113 289 129 323
rect 63 255 129 289
rect 63 221 79 255
rect 113 221 129 255
rect 63 187 129 221
rect 63 153 79 187
rect 113 153 129 187
rect 63 119 129 153
rect 63 85 79 119
rect 113 85 129 119
rect 63 51 129 85
rect 63 17 79 51
rect 113 17 129 51
rect 63 -17 129 17
rect 63 -51 79 -17
rect 113 -51 129 -17
rect 63 -85 129 -51
rect 63 -119 79 -85
rect 113 -119 129 -85
rect 63 -153 129 -119
rect 63 -187 79 -153
rect 113 -187 129 -153
rect 63 -221 129 -187
rect 63 -255 79 -221
rect 113 -255 129 -221
rect 63 -289 129 -255
rect 63 -323 79 -289
rect 113 -323 129 -289
rect 63 -357 129 -323
rect 63 -391 79 -357
rect 113 -391 129 -357
rect 63 -425 129 -391
rect 63 -459 79 -425
rect 113 -459 129 -425
rect 63 -500 129 -459
rect 159 459 225 500
rect 159 425 175 459
rect 209 425 225 459
rect 159 391 225 425
rect 159 357 175 391
rect 209 357 225 391
rect 159 323 225 357
rect 159 289 175 323
rect 209 289 225 323
rect 159 255 225 289
rect 159 221 175 255
rect 209 221 225 255
rect 159 187 225 221
rect 159 153 175 187
rect 209 153 225 187
rect 159 119 225 153
rect 159 85 175 119
rect 209 85 225 119
rect 159 51 225 85
rect 159 17 175 51
rect 209 17 225 51
rect 159 -17 225 17
rect 159 -51 175 -17
rect 209 -51 225 -17
rect 159 -85 225 -51
rect 159 -119 175 -85
rect 209 -119 225 -85
rect 159 -153 225 -119
rect 159 -187 175 -153
rect 209 -187 225 -153
rect 159 -221 225 -187
rect 159 -255 175 -221
rect 209 -255 225 -221
rect 159 -289 225 -255
rect 159 -323 175 -289
rect 209 -323 225 -289
rect 159 -357 225 -323
rect 159 -391 175 -357
rect 209 -391 225 -357
rect 159 -425 225 -391
rect 159 -459 175 -425
rect 209 -459 225 -425
rect 159 -500 225 -459
rect 255 459 321 500
rect 255 425 271 459
rect 305 425 321 459
rect 255 391 321 425
rect 255 357 271 391
rect 305 357 321 391
rect 255 323 321 357
rect 255 289 271 323
rect 305 289 321 323
rect 255 255 321 289
rect 255 221 271 255
rect 305 221 321 255
rect 255 187 321 221
rect 255 153 271 187
rect 305 153 321 187
rect 255 119 321 153
rect 255 85 271 119
rect 305 85 321 119
rect 255 51 321 85
rect 255 17 271 51
rect 305 17 321 51
rect 255 -17 321 17
rect 255 -51 271 -17
rect 305 -51 321 -17
rect 255 -85 321 -51
rect 255 -119 271 -85
rect 305 -119 321 -85
rect 255 -153 321 -119
rect 255 -187 271 -153
rect 305 -187 321 -153
rect 255 -221 321 -187
rect 255 -255 271 -221
rect 305 -255 321 -221
rect 255 -289 321 -255
rect 255 -323 271 -289
rect 305 -323 321 -289
rect 255 -357 321 -323
rect 255 -391 271 -357
rect 305 -391 321 -357
rect 255 -425 321 -391
rect 255 -459 271 -425
rect 305 -459 321 -425
rect 255 -500 321 -459
rect 351 459 417 500
rect 351 425 367 459
rect 401 425 417 459
rect 351 391 417 425
rect 351 357 367 391
rect 401 357 417 391
rect 351 323 417 357
rect 351 289 367 323
rect 401 289 417 323
rect 351 255 417 289
rect 351 221 367 255
rect 401 221 417 255
rect 351 187 417 221
rect 351 153 367 187
rect 401 153 417 187
rect 351 119 417 153
rect 351 85 367 119
rect 401 85 417 119
rect 351 51 417 85
rect 351 17 367 51
rect 401 17 417 51
rect 351 -17 417 17
rect 351 -51 367 -17
rect 401 -51 417 -17
rect 351 -85 417 -51
rect 351 -119 367 -85
rect 401 -119 417 -85
rect 351 -153 417 -119
rect 351 -187 367 -153
rect 401 -187 417 -153
rect 351 -221 417 -187
rect 351 -255 367 -221
rect 401 -255 417 -221
rect 351 -289 417 -255
rect 351 -323 367 -289
rect 401 -323 417 -289
rect 351 -357 417 -323
rect 351 -391 367 -357
rect 401 -391 417 -357
rect 351 -425 417 -391
rect 351 -459 367 -425
rect 401 -459 417 -425
rect 351 -500 417 -459
rect 447 459 513 500
rect 447 425 463 459
rect 497 425 513 459
rect 447 391 513 425
rect 447 357 463 391
rect 497 357 513 391
rect 447 323 513 357
rect 447 289 463 323
rect 497 289 513 323
rect 447 255 513 289
rect 447 221 463 255
rect 497 221 513 255
rect 447 187 513 221
rect 447 153 463 187
rect 497 153 513 187
rect 447 119 513 153
rect 447 85 463 119
rect 497 85 513 119
rect 447 51 513 85
rect 447 17 463 51
rect 497 17 513 51
rect 447 -17 513 17
rect 447 -51 463 -17
rect 497 -51 513 -17
rect 447 -85 513 -51
rect 447 -119 463 -85
rect 497 -119 513 -85
rect 447 -153 513 -119
rect 447 -187 463 -153
rect 497 -187 513 -153
rect 447 -221 513 -187
rect 447 -255 463 -221
rect 497 -255 513 -221
rect 447 -289 513 -255
rect 447 -323 463 -289
rect 497 -323 513 -289
rect 447 -357 513 -323
rect 447 -391 463 -357
rect 497 -391 513 -357
rect 447 -425 513 -391
rect 447 -459 463 -425
rect 497 -459 513 -425
rect 447 -500 513 -459
rect 543 459 605 500
rect 543 425 559 459
rect 593 425 605 459
rect 543 391 605 425
rect 543 357 559 391
rect 593 357 605 391
rect 543 323 605 357
rect 543 289 559 323
rect 593 289 605 323
rect 543 255 605 289
rect 543 221 559 255
rect 593 221 605 255
rect 543 187 605 221
rect 543 153 559 187
rect 593 153 605 187
rect 543 119 605 153
rect 543 85 559 119
rect 593 85 605 119
rect 543 51 605 85
rect 543 17 559 51
rect 593 17 605 51
rect 543 -17 605 17
rect 543 -51 559 -17
rect 593 -51 605 -17
rect 543 -85 605 -51
rect 543 -119 559 -85
rect 593 -119 605 -85
rect 543 -153 605 -119
rect 543 -187 559 -153
rect 593 -187 605 -153
rect 543 -221 605 -187
rect 543 -255 559 -221
rect 593 -255 605 -221
rect 543 -289 605 -255
rect 543 -323 559 -289
rect 593 -323 605 -289
rect 543 -357 605 -323
rect 543 -391 559 -357
rect 593 -391 605 -357
rect 543 -425 605 -391
rect 543 -459 559 -425
rect 593 -459 605 -425
rect 543 -500 605 -459
<< ndiffc >>
rect -593 425 -559 459
rect -593 357 -559 391
rect -593 289 -559 323
rect -593 221 -559 255
rect -593 153 -559 187
rect -593 85 -559 119
rect -593 17 -559 51
rect -593 -51 -559 -17
rect -593 -119 -559 -85
rect -593 -187 -559 -153
rect -593 -255 -559 -221
rect -593 -323 -559 -289
rect -593 -391 -559 -357
rect -593 -459 -559 -425
rect -497 425 -463 459
rect -497 357 -463 391
rect -497 289 -463 323
rect -497 221 -463 255
rect -497 153 -463 187
rect -497 85 -463 119
rect -497 17 -463 51
rect -497 -51 -463 -17
rect -497 -119 -463 -85
rect -497 -187 -463 -153
rect -497 -255 -463 -221
rect -497 -323 -463 -289
rect -497 -391 -463 -357
rect -497 -459 -463 -425
rect -401 425 -367 459
rect -401 357 -367 391
rect -401 289 -367 323
rect -401 221 -367 255
rect -401 153 -367 187
rect -401 85 -367 119
rect -401 17 -367 51
rect -401 -51 -367 -17
rect -401 -119 -367 -85
rect -401 -187 -367 -153
rect -401 -255 -367 -221
rect -401 -323 -367 -289
rect -401 -391 -367 -357
rect -401 -459 -367 -425
rect -305 425 -271 459
rect -305 357 -271 391
rect -305 289 -271 323
rect -305 221 -271 255
rect -305 153 -271 187
rect -305 85 -271 119
rect -305 17 -271 51
rect -305 -51 -271 -17
rect -305 -119 -271 -85
rect -305 -187 -271 -153
rect -305 -255 -271 -221
rect -305 -323 -271 -289
rect -305 -391 -271 -357
rect -305 -459 -271 -425
rect -209 425 -175 459
rect -209 357 -175 391
rect -209 289 -175 323
rect -209 221 -175 255
rect -209 153 -175 187
rect -209 85 -175 119
rect -209 17 -175 51
rect -209 -51 -175 -17
rect -209 -119 -175 -85
rect -209 -187 -175 -153
rect -209 -255 -175 -221
rect -209 -323 -175 -289
rect -209 -391 -175 -357
rect -209 -459 -175 -425
rect -113 425 -79 459
rect -113 357 -79 391
rect -113 289 -79 323
rect -113 221 -79 255
rect -113 153 -79 187
rect -113 85 -79 119
rect -113 17 -79 51
rect -113 -51 -79 -17
rect -113 -119 -79 -85
rect -113 -187 -79 -153
rect -113 -255 -79 -221
rect -113 -323 -79 -289
rect -113 -391 -79 -357
rect -113 -459 -79 -425
rect -17 425 17 459
rect -17 357 17 391
rect -17 289 17 323
rect -17 221 17 255
rect -17 153 17 187
rect -17 85 17 119
rect -17 17 17 51
rect -17 -51 17 -17
rect -17 -119 17 -85
rect -17 -187 17 -153
rect -17 -255 17 -221
rect -17 -323 17 -289
rect -17 -391 17 -357
rect -17 -459 17 -425
rect 79 425 113 459
rect 79 357 113 391
rect 79 289 113 323
rect 79 221 113 255
rect 79 153 113 187
rect 79 85 113 119
rect 79 17 113 51
rect 79 -51 113 -17
rect 79 -119 113 -85
rect 79 -187 113 -153
rect 79 -255 113 -221
rect 79 -323 113 -289
rect 79 -391 113 -357
rect 79 -459 113 -425
rect 175 425 209 459
rect 175 357 209 391
rect 175 289 209 323
rect 175 221 209 255
rect 175 153 209 187
rect 175 85 209 119
rect 175 17 209 51
rect 175 -51 209 -17
rect 175 -119 209 -85
rect 175 -187 209 -153
rect 175 -255 209 -221
rect 175 -323 209 -289
rect 175 -391 209 -357
rect 175 -459 209 -425
rect 271 425 305 459
rect 271 357 305 391
rect 271 289 305 323
rect 271 221 305 255
rect 271 153 305 187
rect 271 85 305 119
rect 271 17 305 51
rect 271 -51 305 -17
rect 271 -119 305 -85
rect 271 -187 305 -153
rect 271 -255 305 -221
rect 271 -323 305 -289
rect 271 -391 305 -357
rect 271 -459 305 -425
rect 367 425 401 459
rect 367 357 401 391
rect 367 289 401 323
rect 367 221 401 255
rect 367 153 401 187
rect 367 85 401 119
rect 367 17 401 51
rect 367 -51 401 -17
rect 367 -119 401 -85
rect 367 -187 401 -153
rect 367 -255 401 -221
rect 367 -323 401 -289
rect 367 -391 401 -357
rect 367 -459 401 -425
rect 463 425 497 459
rect 463 357 497 391
rect 463 289 497 323
rect 463 221 497 255
rect 463 153 497 187
rect 463 85 497 119
rect 463 17 497 51
rect 463 -51 497 -17
rect 463 -119 497 -85
rect 463 -187 497 -153
rect 463 -255 497 -221
rect 463 -323 497 -289
rect 463 -391 497 -357
rect 463 -459 497 -425
rect 559 425 593 459
rect 559 357 593 391
rect 559 289 593 323
rect 559 221 593 255
rect 559 153 593 187
rect 559 85 593 119
rect 559 17 593 51
rect 559 -51 593 -17
rect 559 -119 593 -85
rect 559 -187 593 -153
rect 559 -255 593 -221
rect 559 -323 593 -289
rect 559 -391 593 -357
rect 559 -459 593 -425
<< poly >>
rect -543 538 543 568
rect -543 500 -513 538
rect -447 500 -417 538
rect -351 500 -321 538
rect -255 500 -225 538
rect -159 500 -129 538
rect -63 500 -33 538
rect 33 500 63 538
rect 129 500 159 538
rect 225 500 255 538
rect 321 500 351 538
rect 417 500 447 538
rect 513 500 543 538
rect -543 -554 -513 -500
rect -447 -526 -417 -500
rect -351 -526 -321 -500
rect -255 -526 -225 -500
rect -159 -526 -129 -500
rect -63 -526 -33 -500
rect 33 -526 63 -500
rect 129 -526 159 -500
rect 225 -526 255 -500
rect 321 -526 351 -500
rect 417 -526 447 -500
rect 513 -526 543 -500
rect -575 -584 -513 -554
rect -575 -622 -545 -584
rect -611 -638 -545 -622
rect -611 -672 -595 -638
rect -561 -672 -545 -638
rect -611 -688 -545 -672
<< polycont >>
rect -595 -672 -561 -638
<< locali >>
rect -499 544 497 578
rect -593 485 -559 504
rect -593 413 -559 425
rect -593 341 -559 357
rect -593 269 -559 289
rect -593 197 -559 221
rect -593 125 -559 153
rect -593 53 -559 85
rect -593 -17 -559 17
rect -593 -85 -559 -53
rect -593 -153 -559 -125
rect -593 -221 -559 -197
rect -593 -289 -559 -269
rect -593 -357 -559 -341
rect -593 -425 -559 -413
rect -593 -554 -559 -485
rect -497 485 -463 544
rect -497 413 -463 425
rect -497 341 -463 357
rect -497 269 -463 289
rect -497 197 -463 221
rect -497 125 -463 153
rect -497 53 -463 85
rect -497 -17 -463 17
rect -497 -85 -463 -53
rect -497 -153 -463 -125
rect -497 -221 -463 -197
rect -497 -289 -463 -269
rect -497 -357 -463 -341
rect -497 -425 -463 -413
rect -497 -504 -463 -485
rect -401 485 -367 502
rect -401 413 -367 425
rect -401 341 -367 357
rect -401 269 -367 289
rect -401 197 -367 221
rect -401 125 -367 153
rect -401 53 -367 85
rect -401 -17 -367 17
rect -401 -85 -367 -53
rect -401 -153 -367 -125
rect -401 -221 -367 -197
rect -401 -289 -367 -269
rect -401 -357 -367 -341
rect -401 -425 -367 -413
rect -401 -554 -367 -485
rect -305 485 -271 544
rect -305 413 -271 425
rect -305 341 -271 357
rect -305 269 -271 289
rect -305 197 -271 221
rect -305 125 -271 153
rect -305 53 -271 85
rect -305 -17 -271 17
rect -305 -85 -271 -53
rect -305 -153 -271 -125
rect -305 -221 -271 -197
rect -305 -289 -271 -269
rect -305 -357 -271 -341
rect -305 -425 -271 -413
rect -305 -504 -271 -485
rect -209 485 -175 502
rect -209 413 -175 425
rect -209 341 -175 357
rect -209 269 -175 289
rect -209 197 -175 221
rect -209 125 -175 153
rect -209 53 -175 85
rect -209 -17 -175 17
rect -209 -85 -175 -53
rect -209 -153 -175 -125
rect -209 -221 -175 -197
rect -209 -289 -175 -269
rect -209 -357 -175 -341
rect -209 -425 -175 -413
rect -209 -554 -175 -485
rect -113 485 -79 544
rect -113 413 -79 425
rect -113 341 -79 357
rect -113 269 -79 289
rect -113 197 -79 221
rect -113 125 -79 153
rect -113 53 -79 85
rect -113 -17 -79 17
rect -113 -85 -79 -53
rect -113 -153 -79 -125
rect -113 -221 -79 -197
rect -113 -289 -79 -269
rect -113 -357 -79 -341
rect -113 -425 -79 -413
rect -113 -504 -79 -485
rect -17 485 17 502
rect -17 413 17 425
rect -17 341 17 357
rect -17 269 17 289
rect -17 197 17 221
rect -17 125 17 153
rect -17 53 17 85
rect -17 -17 17 17
rect -17 -85 17 -53
rect -17 -153 17 -125
rect -17 -221 17 -197
rect -17 -289 17 -269
rect -17 -357 17 -341
rect -17 -425 17 -413
rect -17 -554 17 -485
rect 79 485 113 544
rect 79 413 113 425
rect 79 341 113 357
rect 79 269 113 289
rect 79 197 113 221
rect 79 125 113 153
rect 79 53 113 85
rect 79 -17 113 17
rect 79 -85 113 -53
rect 79 -153 113 -125
rect 79 -221 113 -197
rect 79 -289 113 -269
rect 79 -357 113 -341
rect 79 -425 113 -413
rect 79 -504 113 -485
rect 175 485 209 502
rect 175 413 209 425
rect 175 341 209 357
rect 175 269 209 289
rect 175 197 209 221
rect 175 125 209 153
rect 175 53 209 85
rect 175 -17 209 17
rect 175 -85 209 -53
rect 175 -153 209 -125
rect 175 -221 209 -197
rect 175 -289 209 -269
rect 175 -357 209 -341
rect 175 -425 209 -413
rect 175 -554 209 -485
rect 271 485 305 544
rect 271 413 305 425
rect 271 341 305 357
rect 271 269 305 289
rect 271 197 305 221
rect 271 125 305 153
rect 271 53 305 85
rect 271 -17 305 17
rect 271 -85 305 -53
rect 271 -153 305 -125
rect 271 -221 305 -197
rect 271 -289 305 -269
rect 271 -357 305 -341
rect 271 -425 305 -413
rect 271 -504 305 -485
rect 367 485 401 502
rect 367 413 401 425
rect 367 341 401 357
rect 367 269 401 289
rect 367 197 401 221
rect 367 125 401 153
rect 367 53 401 85
rect 367 -17 401 17
rect 367 -85 401 -53
rect 367 -153 401 -125
rect 367 -221 401 -197
rect 367 -289 401 -269
rect 367 -357 401 -341
rect 367 -425 401 -413
rect 367 -554 401 -485
rect 463 485 497 544
rect 463 413 497 425
rect 463 341 497 357
rect 463 269 497 289
rect 463 197 497 221
rect 463 125 497 153
rect 463 53 497 85
rect 463 -17 497 17
rect 463 -85 497 -53
rect 463 -153 497 -125
rect 463 -221 497 -197
rect 463 -289 497 -269
rect 463 -357 497 -341
rect 463 -425 497 -413
rect 463 -502 497 -485
rect 559 485 593 502
rect 559 413 593 425
rect 559 341 593 357
rect 559 269 593 289
rect 559 197 593 221
rect 559 125 593 153
rect 559 53 593 85
rect 559 -17 593 17
rect 559 -85 593 -53
rect 559 -153 593 -125
rect 559 -221 593 -197
rect 559 -289 593 -269
rect 559 -357 593 -341
rect 559 -425 593 -413
rect 559 -554 593 -485
rect -593 -588 593 -554
rect -611 -672 -595 -638
rect -561 -672 -545 -638
<< viali >>
rect -593 459 -559 485
rect -593 451 -559 459
rect -593 391 -559 413
rect -593 379 -559 391
rect -593 323 -559 341
rect -593 307 -559 323
rect -593 255 -559 269
rect -593 235 -559 255
rect -593 187 -559 197
rect -593 163 -559 187
rect -593 119 -559 125
rect -593 91 -559 119
rect -593 51 -559 53
rect -593 19 -559 51
rect -593 -51 -559 -19
rect -593 -53 -559 -51
rect -593 -119 -559 -91
rect -593 -125 -559 -119
rect -593 -187 -559 -163
rect -593 -197 -559 -187
rect -593 -255 -559 -235
rect -593 -269 -559 -255
rect -593 -323 -559 -307
rect -593 -341 -559 -323
rect -593 -391 -559 -379
rect -593 -413 -559 -391
rect -593 -459 -559 -451
rect -593 -485 -559 -459
rect -497 459 -463 485
rect -497 451 -463 459
rect -497 391 -463 413
rect -497 379 -463 391
rect -497 323 -463 341
rect -497 307 -463 323
rect -497 255 -463 269
rect -497 235 -463 255
rect -497 187 -463 197
rect -497 163 -463 187
rect -497 119 -463 125
rect -497 91 -463 119
rect -497 51 -463 53
rect -497 19 -463 51
rect -497 -51 -463 -19
rect -497 -53 -463 -51
rect -497 -119 -463 -91
rect -497 -125 -463 -119
rect -497 -187 -463 -163
rect -497 -197 -463 -187
rect -497 -255 -463 -235
rect -497 -269 -463 -255
rect -497 -323 -463 -307
rect -497 -341 -463 -323
rect -497 -391 -463 -379
rect -497 -413 -463 -391
rect -497 -459 -463 -451
rect -497 -485 -463 -459
rect -401 459 -367 485
rect -401 451 -367 459
rect -401 391 -367 413
rect -401 379 -367 391
rect -401 323 -367 341
rect -401 307 -367 323
rect -401 255 -367 269
rect -401 235 -367 255
rect -401 187 -367 197
rect -401 163 -367 187
rect -401 119 -367 125
rect -401 91 -367 119
rect -401 51 -367 53
rect -401 19 -367 51
rect -401 -51 -367 -19
rect -401 -53 -367 -51
rect -401 -119 -367 -91
rect -401 -125 -367 -119
rect -401 -187 -367 -163
rect -401 -197 -367 -187
rect -401 -255 -367 -235
rect -401 -269 -367 -255
rect -401 -323 -367 -307
rect -401 -341 -367 -323
rect -401 -391 -367 -379
rect -401 -413 -367 -391
rect -401 -459 -367 -451
rect -401 -485 -367 -459
rect -305 459 -271 485
rect -305 451 -271 459
rect -305 391 -271 413
rect -305 379 -271 391
rect -305 323 -271 341
rect -305 307 -271 323
rect -305 255 -271 269
rect -305 235 -271 255
rect -305 187 -271 197
rect -305 163 -271 187
rect -305 119 -271 125
rect -305 91 -271 119
rect -305 51 -271 53
rect -305 19 -271 51
rect -305 -51 -271 -19
rect -305 -53 -271 -51
rect -305 -119 -271 -91
rect -305 -125 -271 -119
rect -305 -187 -271 -163
rect -305 -197 -271 -187
rect -305 -255 -271 -235
rect -305 -269 -271 -255
rect -305 -323 -271 -307
rect -305 -341 -271 -323
rect -305 -391 -271 -379
rect -305 -413 -271 -391
rect -305 -459 -271 -451
rect -305 -485 -271 -459
rect -209 459 -175 485
rect -209 451 -175 459
rect -209 391 -175 413
rect -209 379 -175 391
rect -209 323 -175 341
rect -209 307 -175 323
rect -209 255 -175 269
rect -209 235 -175 255
rect -209 187 -175 197
rect -209 163 -175 187
rect -209 119 -175 125
rect -209 91 -175 119
rect -209 51 -175 53
rect -209 19 -175 51
rect -209 -51 -175 -19
rect -209 -53 -175 -51
rect -209 -119 -175 -91
rect -209 -125 -175 -119
rect -209 -187 -175 -163
rect -209 -197 -175 -187
rect -209 -255 -175 -235
rect -209 -269 -175 -255
rect -209 -323 -175 -307
rect -209 -341 -175 -323
rect -209 -391 -175 -379
rect -209 -413 -175 -391
rect -209 -459 -175 -451
rect -209 -485 -175 -459
rect -113 459 -79 485
rect -113 451 -79 459
rect -113 391 -79 413
rect -113 379 -79 391
rect -113 323 -79 341
rect -113 307 -79 323
rect -113 255 -79 269
rect -113 235 -79 255
rect -113 187 -79 197
rect -113 163 -79 187
rect -113 119 -79 125
rect -113 91 -79 119
rect -113 51 -79 53
rect -113 19 -79 51
rect -113 -51 -79 -19
rect -113 -53 -79 -51
rect -113 -119 -79 -91
rect -113 -125 -79 -119
rect -113 -187 -79 -163
rect -113 -197 -79 -187
rect -113 -255 -79 -235
rect -113 -269 -79 -255
rect -113 -323 -79 -307
rect -113 -341 -79 -323
rect -113 -391 -79 -379
rect -113 -413 -79 -391
rect -113 -459 -79 -451
rect -113 -485 -79 -459
rect -17 459 17 485
rect -17 451 17 459
rect -17 391 17 413
rect -17 379 17 391
rect -17 323 17 341
rect -17 307 17 323
rect -17 255 17 269
rect -17 235 17 255
rect -17 187 17 197
rect -17 163 17 187
rect -17 119 17 125
rect -17 91 17 119
rect -17 51 17 53
rect -17 19 17 51
rect -17 -51 17 -19
rect -17 -53 17 -51
rect -17 -119 17 -91
rect -17 -125 17 -119
rect -17 -187 17 -163
rect -17 -197 17 -187
rect -17 -255 17 -235
rect -17 -269 17 -255
rect -17 -323 17 -307
rect -17 -341 17 -323
rect -17 -391 17 -379
rect -17 -413 17 -391
rect -17 -459 17 -451
rect -17 -485 17 -459
rect 79 459 113 485
rect 79 451 113 459
rect 79 391 113 413
rect 79 379 113 391
rect 79 323 113 341
rect 79 307 113 323
rect 79 255 113 269
rect 79 235 113 255
rect 79 187 113 197
rect 79 163 113 187
rect 79 119 113 125
rect 79 91 113 119
rect 79 51 113 53
rect 79 19 113 51
rect 79 -51 113 -19
rect 79 -53 113 -51
rect 79 -119 113 -91
rect 79 -125 113 -119
rect 79 -187 113 -163
rect 79 -197 113 -187
rect 79 -255 113 -235
rect 79 -269 113 -255
rect 79 -323 113 -307
rect 79 -341 113 -323
rect 79 -391 113 -379
rect 79 -413 113 -391
rect 79 -459 113 -451
rect 79 -485 113 -459
rect 175 459 209 485
rect 175 451 209 459
rect 175 391 209 413
rect 175 379 209 391
rect 175 323 209 341
rect 175 307 209 323
rect 175 255 209 269
rect 175 235 209 255
rect 175 187 209 197
rect 175 163 209 187
rect 175 119 209 125
rect 175 91 209 119
rect 175 51 209 53
rect 175 19 209 51
rect 175 -51 209 -19
rect 175 -53 209 -51
rect 175 -119 209 -91
rect 175 -125 209 -119
rect 175 -187 209 -163
rect 175 -197 209 -187
rect 175 -255 209 -235
rect 175 -269 209 -255
rect 175 -323 209 -307
rect 175 -341 209 -323
rect 175 -391 209 -379
rect 175 -413 209 -391
rect 175 -459 209 -451
rect 175 -485 209 -459
rect 271 459 305 485
rect 271 451 305 459
rect 271 391 305 413
rect 271 379 305 391
rect 271 323 305 341
rect 271 307 305 323
rect 271 255 305 269
rect 271 235 305 255
rect 271 187 305 197
rect 271 163 305 187
rect 271 119 305 125
rect 271 91 305 119
rect 271 51 305 53
rect 271 19 305 51
rect 271 -51 305 -19
rect 271 -53 305 -51
rect 271 -119 305 -91
rect 271 -125 305 -119
rect 271 -187 305 -163
rect 271 -197 305 -187
rect 271 -255 305 -235
rect 271 -269 305 -255
rect 271 -323 305 -307
rect 271 -341 305 -323
rect 271 -391 305 -379
rect 271 -413 305 -391
rect 271 -459 305 -451
rect 271 -485 305 -459
rect 367 459 401 485
rect 367 451 401 459
rect 367 391 401 413
rect 367 379 401 391
rect 367 323 401 341
rect 367 307 401 323
rect 367 255 401 269
rect 367 235 401 255
rect 367 187 401 197
rect 367 163 401 187
rect 367 119 401 125
rect 367 91 401 119
rect 367 51 401 53
rect 367 19 401 51
rect 367 -51 401 -19
rect 367 -53 401 -51
rect 367 -119 401 -91
rect 367 -125 401 -119
rect 367 -187 401 -163
rect 367 -197 401 -187
rect 367 -255 401 -235
rect 367 -269 401 -255
rect 367 -323 401 -307
rect 367 -341 401 -323
rect 367 -391 401 -379
rect 367 -413 401 -391
rect 367 -459 401 -451
rect 367 -485 401 -459
rect 463 459 497 485
rect 463 451 497 459
rect 463 391 497 413
rect 463 379 497 391
rect 463 323 497 341
rect 463 307 497 323
rect 463 255 497 269
rect 463 235 497 255
rect 463 187 497 197
rect 463 163 497 187
rect 463 119 497 125
rect 463 91 497 119
rect 463 51 497 53
rect 463 19 497 51
rect 463 -51 497 -19
rect 463 -53 497 -51
rect 463 -119 497 -91
rect 463 -125 497 -119
rect 463 -187 497 -163
rect 463 -197 497 -187
rect 463 -255 497 -235
rect 463 -269 497 -255
rect 463 -323 497 -307
rect 463 -341 497 -323
rect 463 -391 497 -379
rect 463 -413 497 -391
rect 463 -459 497 -451
rect 463 -485 497 -459
rect 559 459 593 485
rect 559 451 593 459
rect 559 391 593 413
rect 559 379 593 391
rect 559 323 593 341
rect 559 307 593 323
rect 559 255 593 269
rect 559 235 593 255
rect 559 187 593 197
rect 559 163 593 187
rect 559 119 593 125
rect 559 91 593 119
rect 559 51 593 53
rect 559 19 593 51
rect 559 -51 593 -19
rect 559 -53 593 -51
rect 559 -119 593 -91
rect 559 -125 593 -119
rect 559 -187 593 -163
rect 559 -197 593 -187
rect 559 -255 593 -235
rect 559 -269 593 -255
rect 559 -323 593 -307
rect 559 -341 593 -323
rect 559 -391 593 -379
rect 559 -413 593 -391
rect 559 -459 593 -451
rect 559 -485 593 -459
rect -595 -672 -561 -638
<< metal1 >>
rect -599 485 -553 500
rect -599 451 -593 485
rect -559 451 -553 485
rect -599 413 -553 451
rect -599 379 -593 413
rect -559 379 -553 413
rect -599 341 -553 379
rect -599 307 -593 341
rect -559 307 -553 341
rect -599 269 -553 307
rect -599 235 -593 269
rect -559 235 -553 269
rect -599 197 -553 235
rect -599 163 -593 197
rect -559 163 -553 197
rect -599 125 -553 163
rect -599 91 -593 125
rect -559 91 -553 125
rect -599 53 -553 91
rect -599 19 -593 53
rect -559 19 -553 53
rect -599 -19 -553 19
rect -599 -53 -593 -19
rect -559 -53 -553 -19
rect -599 -91 -553 -53
rect -599 -125 -593 -91
rect -559 -125 -553 -91
rect -599 -163 -553 -125
rect -599 -197 -593 -163
rect -559 -197 -553 -163
rect -599 -235 -553 -197
rect -599 -269 -593 -235
rect -559 -269 -553 -235
rect -599 -307 -553 -269
rect -599 -341 -593 -307
rect -559 -341 -553 -307
rect -599 -379 -553 -341
rect -599 -413 -593 -379
rect -559 -413 -553 -379
rect -599 -451 -553 -413
rect -599 -485 -593 -451
rect -559 -485 -553 -451
rect -599 -500 -553 -485
rect -503 485 -457 500
rect -503 451 -497 485
rect -463 451 -457 485
rect -503 413 -457 451
rect -503 379 -497 413
rect -463 379 -457 413
rect -503 341 -457 379
rect -503 307 -497 341
rect -463 307 -457 341
rect -503 269 -457 307
rect -503 235 -497 269
rect -463 235 -457 269
rect -503 197 -457 235
rect -503 163 -497 197
rect -463 163 -457 197
rect -503 125 -457 163
rect -503 91 -497 125
rect -463 91 -457 125
rect -503 53 -457 91
rect -503 19 -497 53
rect -463 19 -457 53
rect -503 -19 -457 19
rect -503 -53 -497 -19
rect -463 -53 -457 -19
rect -503 -91 -457 -53
rect -503 -125 -497 -91
rect -463 -125 -457 -91
rect -503 -163 -457 -125
rect -503 -197 -497 -163
rect -463 -197 -457 -163
rect -503 -235 -457 -197
rect -503 -269 -497 -235
rect -463 -269 -457 -235
rect -503 -307 -457 -269
rect -503 -341 -497 -307
rect -463 -341 -457 -307
rect -503 -379 -457 -341
rect -503 -413 -497 -379
rect -463 -413 -457 -379
rect -503 -451 -457 -413
rect -503 -485 -497 -451
rect -463 -485 -457 -451
rect -503 -500 -457 -485
rect -407 485 -361 500
rect -407 451 -401 485
rect -367 451 -361 485
rect -407 413 -361 451
rect -407 379 -401 413
rect -367 379 -361 413
rect -407 341 -361 379
rect -407 307 -401 341
rect -367 307 -361 341
rect -407 269 -361 307
rect -407 235 -401 269
rect -367 235 -361 269
rect -407 197 -361 235
rect -407 163 -401 197
rect -367 163 -361 197
rect -407 125 -361 163
rect -407 91 -401 125
rect -367 91 -361 125
rect -407 53 -361 91
rect -407 19 -401 53
rect -367 19 -361 53
rect -407 -19 -361 19
rect -407 -53 -401 -19
rect -367 -53 -361 -19
rect -407 -91 -361 -53
rect -407 -125 -401 -91
rect -367 -125 -361 -91
rect -407 -163 -361 -125
rect -407 -197 -401 -163
rect -367 -197 -361 -163
rect -407 -235 -361 -197
rect -407 -269 -401 -235
rect -367 -269 -361 -235
rect -407 -307 -361 -269
rect -407 -341 -401 -307
rect -367 -341 -361 -307
rect -407 -379 -361 -341
rect -407 -413 -401 -379
rect -367 -413 -361 -379
rect -407 -451 -361 -413
rect -407 -485 -401 -451
rect -367 -485 -361 -451
rect -407 -500 -361 -485
rect -311 485 -265 500
rect -311 451 -305 485
rect -271 451 -265 485
rect -311 413 -265 451
rect -311 379 -305 413
rect -271 379 -265 413
rect -311 341 -265 379
rect -311 307 -305 341
rect -271 307 -265 341
rect -311 269 -265 307
rect -311 235 -305 269
rect -271 235 -265 269
rect -311 197 -265 235
rect -311 163 -305 197
rect -271 163 -265 197
rect -311 125 -265 163
rect -311 91 -305 125
rect -271 91 -265 125
rect -311 53 -265 91
rect -311 19 -305 53
rect -271 19 -265 53
rect -311 -19 -265 19
rect -311 -53 -305 -19
rect -271 -53 -265 -19
rect -311 -91 -265 -53
rect -311 -125 -305 -91
rect -271 -125 -265 -91
rect -311 -163 -265 -125
rect -311 -197 -305 -163
rect -271 -197 -265 -163
rect -311 -235 -265 -197
rect -311 -269 -305 -235
rect -271 -269 -265 -235
rect -311 -307 -265 -269
rect -311 -341 -305 -307
rect -271 -341 -265 -307
rect -311 -379 -265 -341
rect -311 -413 -305 -379
rect -271 -413 -265 -379
rect -311 -451 -265 -413
rect -311 -485 -305 -451
rect -271 -485 -265 -451
rect -311 -500 -265 -485
rect -215 485 -169 500
rect -215 451 -209 485
rect -175 451 -169 485
rect -215 413 -169 451
rect -215 379 -209 413
rect -175 379 -169 413
rect -215 341 -169 379
rect -215 307 -209 341
rect -175 307 -169 341
rect -215 269 -169 307
rect -215 235 -209 269
rect -175 235 -169 269
rect -215 197 -169 235
rect -215 163 -209 197
rect -175 163 -169 197
rect -215 125 -169 163
rect -215 91 -209 125
rect -175 91 -169 125
rect -215 53 -169 91
rect -215 19 -209 53
rect -175 19 -169 53
rect -215 -19 -169 19
rect -215 -53 -209 -19
rect -175 -53 -169 -19
rect -215 -91 -169 -53
rect -215 -125 -209 -91
rect -175 -125 -169 -91
rect -215 -163 -169 -125
rect -215 -197 -209 -163
rect -175 -197 -169 -163
rect -215 -235 -169 -197
rect -215 -269 -209 -235
rect -175 -269 -169 -235
rect -215 -307 -169 -269
rect -215 -341 -209 -307
rect -175 -341 -169 -307
rect -215 -379 -169 -341
rect -215 -413 -209 -379
rect -175 -413 -169 -379
rect -215 -451 -169 -413
rect -215 -485 -209 -451
rect -175 -485 -169 -451
rect -215 -500 -169 -485
rect -119 485 -73 500
rect -119 451 -113 485
rect -79 451 -73 485
rect -119 413 -73 451
rect -119 379 -113 413
rect -79 379 -73 413
rect -119 341 -73 379
rect -119 307 -113 341
rect -79 307 -73 341
rect -119 269 -73 307
rect -119 235 -113 269
rect -79 235 -73 269
rect -119 197 -73 235
rect -119 163 -113 197
rect -79 163 -73 197
rect -119 125 -73 163
rect -119 91 -113 125
rect -79 91 -73 125
rect -119 53 -73 91
rect -119 19 -113 53
rect -79 19 -73 53
rect -119 -19 -73 19
rect -119 -53 -113 -19
rect -79 -53 -73 -19
rect -119 -91 -73 -53
rect -119 -125 -113 -91
rect -79 -125 -73 -91
rect -119 -163 -73 -125
rect -119 -197 -113 -163
rect -79 -197 -73 -163
rect -119 -235 -73 -197
rect -119 -269 -113 -235
rect -79 -269 -73 -235
rect -119 -307 -73 -269
rect -119 -341 -113 -307
rect -79 -341 -73 -307
rect -119 -379 -73 -341
rect -119 -413 -113 -379
rect -79 -413 -73 -379
rect -119 -451 -73 -413
rect -119 -485 -113 -451
rect -79 -485 -73 -451
rect -119 -500 -73 -485
rect -23 485 23 500
rect -23 451 -17 485
rect 17 451 23 485
rect -23 413 23 451
rect -23 379 -17 413
rect 17 379 23 413
rect -23 341 23 379
rect -23 307 -17 341
rect 17 307 23 341
rect -23 269 23 307
rect -23 235 -17 269
rect 17 235 23 269
rect -23 197 23 235
rect -23 163 -17 197
rect 17 163 23 197
rect -23 125 23 163
rect -23 91 -17 125
rect 17 91 23 125
rect -23 53 23 91
rect -23 19 -17 53
rect 17 19 23 53
rect -23 -19 23 19
rect -23 -53 -17 -19
rect 17 -53 23 -19
rect -23 -91 23 -53
rect -23 -125 -17 -91
rect 17 -125 23 -91
rect -23 -163 23 -125
rect -23 -197 -17 -163
rect 17 -197 23 -163
rect -23 -235 23 -197
rect -23 -269 -17 -235
rect 17 -269 23 -235
rect -23 -307 23 -269
rect -23 -341 -17 -307
rect 17 -341 23 -307
rect -23 -379 23 -341
rect -23 -413 -17 -379
rect 17 -413 23 -379
rect -23 -451 23 -413
rect -23 -485 -17 -451
rect 17 -485 23 -451
rect -23 -500 23 -485
rect 73 485 119 500
rect 73 451 79 485
rect 113 451 119 485
rect 73 413 119 451
rect 73 379 79 413
rect 113 379 119 413
rect 73 341 119 379
rect 73 307 79 341
rect 113 307 119 341
rect 73 269 119 307
rect 73 235 79 269
rect 113 235 119 269
rect 73 197 119 235
rect 73 163 79 197
rect 113 163 119 197
rect 73 125 119 163
rect 73 91 79 125
rect 113 91 119 125
rect 73 53 119 91
rect 73 19 79 53
rect 113 19 119 53
rect 73 -19 119 19
rect 73 -53 79 -19
rect 113 -53 119 -19
rect 73 -91 119 -53
rect 73 -125 79 -91
rect 113 -125 119 -91
rect 73 -163 119 -125
rect 73 -197 79 -163
rect 113 -197 119 -163
rect 73 -235 119 -197
rect 73 -269 79 -235
rect 113 -269 119 -235
rect 73 -307 119 -269
rect 73 -341 79 -307
rect 113 -341 119 -307
rect 73 -379 119 -341
rect 73 -413 79 -379
rect 113 -413 119 -379
rect 73 -451 119 -413
rect 73 -485 79 -451
rect 113 -485 119 -451
rect 73 -500 119 -485
rect 169 485 215 500
rect 169 451 175 485
rect 209 451 215 485
rect 169 413 215 451
rect 169 379 175 413
rect 209 379 215 413
rect 169 341 215 379
rect 169 307 175 341
rect 209 307 215 341
rect 169 269 215 307
rect 169 235 175 269
rect 209 235 215 269
rect 169 197 215 235
rect 169 163 175 197
rect 209 163 215 197
rect 169 125 215 163
rect 169 91 175 125
rect 209 91 215 125
rect 169 53 215 91
rect 169 19 175 53
rect 209 19 215 53
rect 169 -19 215 19
rect 169 -53 175 -19
rect 209 -53 215 -19
rect 169 -91 215 -53
rect 169 -125 175 -91
rect 209 -125 215 -91
rect 169 -163 215 -125
rect 169 -197 175 -163
rect 209 -197 215 -163
rect 169 -235 215 -197
rect 169 -269 175 -235
rect 209 -269 215 -235
rect 169 -307 215 -269
rect 169 -341 175 -307
rect 209 -341 215 -307
rect 169 -379 215 -341
rect 169 -413 175 -379
rect 209 -413 215 -379
rect 169 -451 215 -413
rect 169 -485 175 -451
rect 209 -485 215 -451
rect 169 -500 215 -485
rect 265 485 311 500
rect 265 451 271 485
rect 305 451 311 485
rect 265 413 311 451
rect 265 379 271 413
rect 305 379 311 413
rect 265 341 311 379
rect 265 307 271 341
rect 305 307 311 341
rect 265 269 311 307
rect 265 235 271 269
rect 305 235 311 269
rect 265 197 311 235
rect 265 163 271 197
rect 305 163 311 197
rect 265 125 311 163
rect 265 91 271 125
rect 305 91 311 125
rect 265 53 311 91
rect 265 19 271 53
rect 305 19 311 53
rect 265 -19 311 19
rect 265 -53 271 -19
rect 305 -53 311 -19
rect 265 -91 311 -53
rect 265 -125 271 -91
rect 305 -125 311 -91
rect 265 -163 311 -125
rect 265 -197 271 -163
rect 305 -197 311 -163
rect 265 -235 311 -197
rect 265 -269 271 -235
rect 305 -269 311 -235
rect 265 -307 311 -269
rect 265 -341 271 -307
rect 305 -341 311 -307
rect 265 -379 311 -341
rect 265 -413 271 -379
rect 305 -413 311 -379
rect 265 -451 311 -413
rect 265 -485 271 -451
rect 305 -485 311 -451
rect 265 -500 311 -485
rect 361 485 407 500
rect 361 451 367 485
rect 401 451 407 485
rect 361 413 407 451
rect 361 379 367 413
rect 401 379 407 413
rect 361 341 407 379
rect 361 307 367 341
rect 401 307 407 341
rect 361 269 407 307
rect 361 235 367 269
rect 401 235 407 269
rect 361 197 407 235
rect 361 163 367 197
rect 401 163 407 197
rect 361 125 407 163
rect 361 91 367 125
rect 401 91 407 125
rect 361 53 407 91
rect 361 19 367 53
rect 401 19 407 53
rect 361 -19 407 19
rect 361 -53 367 -19
rect 401 -53 407 -19
rect 361 -91 407 -53
rect 361 -125 367 -91
rect 401 -125 407 -91
rect 361 -163 407 -125
rect 361 -197 367 -163
rect 401 -197 407 -163
rect 361 -235 407 -197
rect 361 -269 367 -235
rect 401 -269 407 -235
rect 361 -307 407 -269
rect 361 -341 367 -307
rect 401 -341 407 -307
rect 361 -379 407 -341
rect 361 -413 367 -379
rect 401 -413 407 -379
rect 361 -451 407 -413
rect 361 -485 367 -451
rect 401 -485 407 -451
rect 361 -500 407 -485
rect 457 485 503 500
rect 457 451 463 485
rect 497 451 503 485
rect 457 413 503 451
rect 457 379 463 413
rect 497 379 503 413
rect 457 341 503 379
rect 457 307 463 341
rect 497 307 503 341
rect 457 269 503 307
rect 457 235 463 269
rect 497 235 503 269
rect 457 197 503 235
rect 457 163 463 197
rect 497 163 503 197
rect 457 125 503 163
rect 457 91 463 125
rect 497 91 503 125
rect 457 53 503 91
rect 457 19 463 53
rect 497 19 503 53
rect 457 -19 503 19
rect 457 -53 463 -19
rect 497 -53 503 -19
rect 457 -91 503 -53
rect 457 -125 463 -91
rect 497 -125 503 -91
rect 457 -163 503 -125
rect 457 -197 463 -163
rect 497 -197 503 -163
rect 457 -235 503 -197
rect 457 -269 463 -235
rect 497 -269 503 -235
rect 457 -307 503 -269
rect 457 -341 463 -307
rect 497 -341 503 -307
rect 457 -379 503 -341
rect 457 -413 463 -379
rect 497 -413 503 -379
rect 457 -451 503 -413
rect 457 -485 463 -451
rect 497 -485 503 -451
rect 457 -500 503 -485
rect 553 485 599 500
rect 553 451 559 485
rect 593 451 599 485
rect 553 413 599 451
rect 553 379 559 413
rect 593 379 599 413
rect 553 341 599 379
rect 553 307 559 341
rect 593 307 599 341
rect 553 269 599 307
rect 553 235 559 269
rect 593 235 599 269
rect 553 197 599 235
rect 553 163 559 197
rect 593 163 599 197
rect 553 125 599 163
rect 553 91 559 125
rect 593 91 599 125
rect 553 53 599 91
rect 553 19 559 53
rect 593 19 599 53
rect 553 -19 599 19
rect 553 -53 559 -19
rect 593 -53 599 -19
rect 553 -91 599 -53
rect 553 -125 559 -91
rect 593 -125 599 -91
rect 553 -163 599 -125
rect 553 -197 559 -163
rect 593 -197 599 -163
rect 553 -235 599 -197
rect 553 -269 559 -235
rect 593 -269 599 -235
rect 553 -307 599 -269
rect 553 -341 559 -307
rect 593 -341 599 -307
rect 553 -379 599 -341
rect 553 -413 559 -379
rect 593 -413 599 -379
rect 553 -451 599 -413
rect 553 -485 559 -451
rect 593 -485 599 -451
rect 553 -500 599 -485
rect -607 -638 -549 -632
rect -607 -672 -595 -638
rect -561 -672 -549 -638
rect -607 -678 -549 -672
<< end >>
