magic
tech sky130A
magscale 1 2
timestamp 1634821592
<< error_s >>
rect -1176 5049 -1118 5055
rect -1176 5015 -1164 5049
rect 1264 5045 1322 5051
rect -1176 5009 -1118 5015
rect 1264 5011 1276 5045
rect 1264 5005 1322 5011
rect 308 2019 366 2025
rect 308 1985 320 2019
rect 308 1979 366 1985
rect 114 1244 172 1250
rect 114 1210 126 1244
rect 114 1204 172 1210
rect -1308 -1628 -1250 -1622
rect -1308 -1662 -1296 -1628
rect -1308 -1668 -1250 -1662
<< nwell >>
rect -1390 4966 1646 5200
rect -1390 3674 1642 4966
rect -1396 3424 1642 3674
rect -1396 1886 1636 3424
<< locali >>
rect -688 4908 -654 5100
rect 988 4910 1022 4996
rect -572 3648 -538 3792
rect 892 3652 926 3790
rect 128 3236 162 3332
rect 224 1996 258 2128
rect 222 1110 256 1202
rect 126 -62 160 22
rect -718 -446 -684 -334
rect 948 -424 982 -340
rect -622 -1638 -588 -1544
rect 1042 -1612 1076 -1542
<< viali >>
rect -688 5100 -654 5134
rect 988 4996 1022 5030
rect -572 3614 -538 3648
rect 892 3618 926 3652
rect 128 3332 162 3366
rect 224 1962 258 1996
rect 222 1202 256 1236
rect 126 -96 160 -62
rect -718 -334 -684 -300
rect 948 -340 982 -306
rect -622 -1672 -588 -1638
rect 1042 -1646 1076 -1612
<< metal1 >>
rect -700 5134 1036 5148
rect -700 5100 -688 5134
rect -654 5100 1036 5134
rect -700 5090 1036 5100
rect 976 5030 1036 5090
rect 976 4996 988 5030
rect 1022 4996 1036 5030
rect 976 4986 1036 4996
rect -584 3648 -528 3660
rect -584 3614 -572 3648
rect -538 3614 -528 3648
rect -584 3506 -528 3614
rect 876 3652 942 3672
rect 876 3618 892 3652
rect 926 3618 942 3652
rect 876 3506 942 3618
rect -584 3450 942 3506
rect -584 3448 -528 3450
rect 118 3366 172 3450
rect 118 3332 128 3366
rect 162 3332 172 3366
rect 118 3316 172 3332
rect 114 1972 172 2030
rect 210 1996 272 2012
rect 210 1962 224 1996
rect 258 1962 272 1996
rect 210 1236 272 1962
rect 210 1202 222 1236
rect 256 1202 272 1236
rect 210 1190 272 1202
rect 114 -62 172 -50
rect 114 -96 126 -62
rect 160 -96 172 -62
rect 114 -156 172 -96
rect -730 -204 998 -156
rect -730 -300 -672 -204
rect -730 -334 -718 -300
rect -684 -334 -672 -300
rect -730 -346 -672 -334
rect 938 -306 996 -204
rect 938 -340 948 -306
rect 982 -340 996 -306
rect 938 -352 996 -340
rect 1030 -1612 1088 -1598
rect -634 -1638 -576 -1628
rect -634 -1672 -622 -1638
rect -588 -1672 -576 -1638
rect -634 -1718 -576 -1672
rect 1030 -1646 1042 -1612
rect 1076 -1646 1088 -1612
rect 1030 -1718 1088 -1646
rect 1322 -1674 1382 -1618
rect -634 -1778 1092 -1718
use sky130_fd_pr__nfet_01v8_LB5HPE  sky130_fd_pr__nfet_01v8_LB5HPE_0
timestamp 1634821592
transform 1 0 239 0 1 572
box -247 -584 247 688
use sky130_fd_pr__nfet_01v8_Z96LW5  sky130_fd_pr__nfet_01v8_Z96LW5_0
timestamp 1634821592
transform 1 0 1019 0 1 -990
box -583 -688 583 600
use sky130_fd_pr__nfet_01v8_JV9MWK  sky130_fd_pr__nfet_01v8_JV9MWK_0
timestamp 1634821592
transform 1 0 -701 0 1 -990
box -631 -688 631 578
use sky130_fd_pr__pfet_01v8_AWEQDE  sky130_fd_pr__pfet_01v8_AWEQDE_0
timestamp 1634821592
transform 1 0 241 0 1 2686
box -365 -718 257 818
use sky130_fd_pr__pfet_01v8_AWWSCB  sky130_fd_pr__pfet_01v8_AWWSCB_0
timestamp 1634821592
transform 1 0 909 0 1 4344
box -579 -720 449 814
use sky130_fd_pr__pfet_01v8_K2D88D  sky130_fd_pr__pfet_01v8_K2D88D_0
timestamp 1634821592
transform 1 0 -665 0 1 4348
box -803 -742 643 804
<< end >>
