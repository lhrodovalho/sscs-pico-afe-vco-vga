magic
tech sky130A
timestamp 1634782756
<< nwell >>
rect 860 2640 920 2660
rect 860 2610 940 2640
rect 860 -120 920 2610
rect 6580 2600 6630 2650
rect 7430 2640 7480 2650
rect 7500 2640 7560 2660
rect 7430 2610 7560 2640
rect 7430 2600 7480 2610
rect 940 -120 990 -110
rect 860 -160 990 -120
rect 7430 -120 7480 -110
rect 7500 -120 7560 2610
rect 7430 -150 7560 -120
rect 7430 -160 7480 -150
rect 860 -170 940 -160
rect 7500 -170 7560 -150
rect 860 -1340 920 -1320
rect 940 -1340 990 -1330
rect 7430 -1340 7480 -1330
rect 7500 -1340 7560 -1320
rect 860 -1370 7560 -1340
rect 860 -4100 920 -1370
rect 940 -1380 990 -1370
rect 7430 -1380 7480 -1370
rect 940 -4100 990 -4090
rect 1790 -4100 1840 -4090
rect 6580 -4100 6630 -4090
rect 7430 -4100 7480 -4090
rect 7500 -4100 7560 -1370
rect 860 -4130 7560 -4100
rect 860 -4150 920 -4130
rect 940 -4140 990 -4130
rect 1790 -4140 1840 -4130
rect 6580 -4140 6630 -4130
rect 7430 -4140 7480 -4130
rect 7500 -4150 7560 -4130
<< pwell >>
rect 920 2710 7500 2730
rect 2730 2670 2780 2710
rect 2730 -4210 2780 -4160
<< psubdiff >>
rect 810 2680 920 2710
rect 2730 2680 2780 2710
rect 7500 2680 7610 2710
rect 810 -220 7610 -190
rect 810 -1300 860 -1270
rect 7560 -1300 7610 -1270
rect 810 -4200 920 -4170
rect 2730 -4200 2780 -4170
rect 7500 -4200 7610 -4170
<< nsubdiff >>
rect 880 2610 940 2640
rect 6580 2610 6630 2640
rect 7430 2610 7540 2640
rect 880 -150 990 -120
rect 7430 -150 7540 -120
rect 880 -1370 7540 -1340
rect 880 -4130 7540 -4100
<< psubdiffcont >>
rect 810 -190 840 2680
rect 7580 -190 7610 2680
rect 860 -1300 7560 -1270
rect 810 -4170 840 -1300
rect 7580 -4170 7610 -1300
<< nsubdiffcont >>
rect 880 -120 910 2610
rect 7510 -120 7540 2610
rect 880 -4100 910 -1370
rect 7510 -4100 7540 -1370
<< locali >>
rect -1340 -240 -1240 3670
rect -1350 -250 -1240 -240
rect -1350 -280 -1340 -250
rect -1310 -280 -1240 -250
rect -1210 -280 -1040 3670
rect -1010 -280 -840 3670
rect -810 -280 -640 3670
rect -610 -280 -440 3670
rect -410 -280 -240 3670
rect 2730 2710 2780 2720
rect 810 2680 920 2710
rect 2730 2680 2740 2710
rect 2770 2680 2780 2710
rect 2730 2670 2780 2680
rect 5640 2710 5690 2720
rect 5640 2680 5650 2710
rect 5680 2680 5690 2710
rect 7500 2680 7610 2710
rect 5640 2670 5690 2680
rect 940 2640 990 2650
rect 880 2610 950 2640
rect 980 2610 990 2640
rect 940 2600 990 2610
rect 6580 2640 6630 2650
rect 6580 2610 6590 2640
rect 6620 2610 6630 2640
rect 6580 2600 6630 2610
rect 7430 2640 7480 2650
rect 7430 2610 7440 2640
rect 7470 2610 7540 2640
rect 7430 2600 7480 2610
rect 940 -120 990 -110
rect 880 -150 950 -120
rect 980 -150 990 -120
rect 940 -160 990 -150
rect 7430 -120 7480 -110
rect 7430 -150 7440 -120
rect 7470 -150 7540 -120
rect 7430 -160 7480 -150
rect 810 -220 7610 -190
rect -1350 -290 7500 -280
rect -1340 -360 7500 -290
rect -1350 -370 7500 -360
rect -1350 -400 -1340 -370
rect -1310 -400 -1240 -370
rect -1210 -400 -1040 -370
rect -1010 -400 -840 -370
rect -810 -400 -640 -370
rect -610 -400 -440 -370
rect -410 -400 -240 -370
rect -1350 -410 7500 -400
rect -1340 -480 7500 -410
rect -1350 -490 7500 -480
rect -1350 -520 -1340 -490
rect -1310 -520 -1240 -490
rect -1210 -520 -1040 -490
rect -1010 -520 -840 -490
rect -810 -520 -640 -490
rect -610 -520 -440 -490
rect -410 -520 -240 -490
rect -1350 -530 7500 -520
rect -1340 -600 7500 -530
rect -1350 -610 7500 -600
rect -1350 -640 -1340 -610
rect -1310 -640 -1240 -610
rect -1210 -640 -1040 -610
rect -1010 -640 -840 -610
rect -810 -640 -640 -610
rect -610 -640 -440 -610
rect -410 -640 -240 -610
rect -1350 -650 7500 -640
rect -1340 -720 7500 -650
rect -1350 -730 7500 -720
rect -1350 -760 -1340 -730
rect -1310 -760 -1240 -730
rect -1210 -760 -1040 -730
rect -1010 -760 -840 -730
rect -810 -760 -640 -730
rect -610 -760 -440 -730
rect -410 -760 -240 -730
rect -1350 -770 7500 -760
rect -1340 -840 7500 -770
rect -1350 -850 7500 -840
rect -1350 -880 -1340 -850
rect -1310 -880 -1240 -850
rect -1210 -880 -1040 -850
rect -1010 -880 -840 -850
rect -810 -880 -640 -850
rect -610 -880 -440 -850
rect -410 -880 -240 -850
rect -1350 -890 7500 -880
rect -1340 -960 7500 -890
rect -1350 -970 7500 -960
rect -1350 -1000 -1340 -970
rect -1310 -1000 -1240 -970
rect -1210 -1000 -1040 -970
rect -1010 -1000 -840 -970
rect -810 -1000 -640 -970
rect -610 -1000 -440 -970
rect -410 -1000 -240 -970
rect -1350 -1010 7500 -1000
rect -1340 -1080 7500 -1010
rect -1350 -1090 7500 -1080
rect -1350 -1120 -1340 -1090
rect -1310 -1120 -1240 -1090
rect -1210 -1120 -1040 -1090
rect -1010 -1120 -840 -1090
rect -810 -1120 -640 -1090
rect -610 -1120 -440 -1090
rect -410 -1120 -240 -1090
rect -1350 -1130 7500 -1120
rect -1340 -1200 7500 -1130
rect -1350 -1210 7500 -1200
rect -1350 -1240 -1340 -1210
rect -1310 -1240 -1240 -1210
rect -1350 -1250 -1240 -1240
rect -1340 -5160 -1240 -1250
rect -1210 -5160 -1040 -1210
rect -1010 -5160 -840 -1210
rect -810 -5160 -640 -1210
rect -610 -5160 -440 -1210
rect -410 -5160 -240 -1210
rect 810 -1300 860 -1270
rect 7560 -1300 7610 -1270
rect 940 -1340 990 -1330
rect 7430 -1340 7480 -1330
rect 880 -1370 950 -1340
rect 980 -1370 7440 -1340
rect 7470 -1370 7540 -1340
rect 940 -1380 990 -1370
rect 7430 -1380 7480 -1370
rect 940 -4100 990 -4090
rect 1790 -4100 1840 -4090
rect 6580 -4100 6630 -4090
rect 7430 -4100 7480 -4090
rect 880 -4130 950 -4100
rect 980 -4130 1800 -4100
rect 1830 -4130 6590 -4100
rect 6620 -4130 7440 -4100
rect 7470 -4130 7540 -4100
rect 940 -4140 990 -4130
rect 1790 -4140 1840 -4130
rect 6580 -4140 6630 -4130
rect 7430 -4140 7480 -4130
rect 2730 -4170 2780 -4160
rect 810 -4200 920 -4170
rect 2730 -4200 2740 -4170
rect 2770 -4200 2780 -4170
rect 2730 -4210 2780 -4200
rect 5640 -4170 5690 -4160
rect 5640 -4200 5650 -4170
rect 5680 -4200 5690 -4170
rect 7500 -4200 7610 -4170
rect 5640 -4210 5690 -4200
<< viali >>
rect -1340 -280 -1310 -250
rect 2740 2680 2770 2710
rect 5650 2680 5680 2710
rect 950 2610 980 2640
rect 6590 2610 6620 2640
rect 7440 2610 7470 2640
rect 950 -150 980 -120
rect 7440 -150 7470 -120
rect -1340 -400 -1310 -370
rect -1340 -520 -1310 -490
rect -1340 -640 -1310 -610
rect -1340 -760 -1310 -730
rect -1340 -880 -1310 -850
rect -1340 -1000 -1310 -970
rect -1340 -1120 -1310 -1090
rect -1340 -1240 -1310 -1210
rect 950 -1370 980 -1340
rect 7440 -1370 7470 -1340
rect 950 -4130 980 -4100
rect 1800 -4130 1830 -4100
rect 6590 -4130 6620 -4100
rect 7440 -4130 7470 -4100
rect 2740 -4200 2770 -4170
rect 5650 -4200 5680 -4170
<< metal1 >>
rect -1350 -250 -1300 -240
rect -1350 -280 -1340 -250
rect -1310 -280 -1300 -250
rect -1350 -290 -1300 -280
rect -1350 -370 -1300 -360
rect -1350 -400 -1340 -370
rect -1310 -400 -1300 -370
rect -1350 -410 -1300 -400
rect -1350 -490 -1300 -480
rect -1350 -520 -1340 -490
rect -1310 -520 -1300 -490
rect -1350 -530 -1300 -520
rect -1350 -610 -1300 -600
rect -1350 -640 -1340 -610
rect -1310 -640 -1300 -610
rect -1350 -650 -1300 -640
rect -1350 -730 -1300 -720
rect -1350 -760 -1340 -730
rect -1310 -760 -1300 -730
rect -1350 -770 -1300 -760
rect -1350 -850 -1300 -840
rect -1350 -880 -1340 -850
rect -1310 -880 -1300 -850
rect -1350 -890 -1300 -880
rect -1350 -970 -1300 -960
rect -1350 -1000 -1340 -970
rect -1310 -1000 -1300 -970
rect -1350 -1010 -1300 -1000
rect -1350 -1090 -1300 -1080
rect -1350 -1120 -1340 -1090
rect -1310 -1120 -1300 -1090
rect -1350 -1130 -1300 -1120
rect -1350 -1210 -1300 -1200
rect -1350 -1240 -1340 -1210
rect -1310 -1240 -1300 -1210
rect -1350 -1250 -1300 -1240
rect -1240 -5160 -1210 3670
rect -1040 -5160 -1010 3670
rect -840 -5160 -810 3670
rect -640 -5160 -610 3670
rect -440 -5160 -410 3670
rect -240 -5160 -210 3670
rect 950 3660 980 3670
rect 950 2650 980 3520
rect 1800 3660 1830 3670
rect 1800 2730 1830 3520
rect 3680 3660 3710 3670
rect 2740 3020 2770 3030
rect 2740 2730 2770 2880
rect 3680 2730 3710 3520
rect 4620 3660 4650 3670
rect 4620 2730 4650 3520
rect 4710 3660 4740 3670
rect 4710 2730 4740 3520
rect 6590 3660 6620 3670
rect 5650 3020 5680 3030
rect 5650 2730 5680 2880
rect 6590 2730 6620 3520
rect 7440 3660 7470 3670
rect 2730 2710 2780 2720
rect 2730 2680 2740 2710
rect 2770 2680 2780 2710
rect 2730 2670 2780 2680
rect 5640 2710 5690 2720
rect 5640 2680 5650 2710
rect 5680 2680 5690 2710
rect 5640 2670 5690 2680
rect 7440 2650 7470 3520
rect 940 2640 990 2650
rect 940 2610 950 2640
rect 980 2610 990 2640
rect 940 2600 990 2610
rect 6580 2640 6630 2650
rect 6580 2610 6590 2640
rect 6620 2610 6630 2640
rect 6580 2600 6630 2610
rect 7430 2640 7480 2650
rect 7430 2610 7440 2640
rect 7470 2610 7480 2640
rect 7430 2600 7480 2610
rect 950 -110 980 2600
rect 7440 2580 7470 2600
rect 940 -120 990 -110
rect 940 -150 950 -120
rect 980 -150 990 -120
rect 940 -160 990 -150
rect 7430 -120 7480 -110
rect 7430 -150 7440 -120
rect 7470 -150 7480 -120
rect 7430 -160 7480 -150
rect 950 -240 980 -160
rect 1070 -310 1100 -240
rect 1070 -350 1100 -340
rect 1890 -550 1920 -240
rect 1890 -590 1920 -580
rect 1950 -250 1980 -240
rect 1950 -370 1980 -280
rect 1950 -490 1980 -400
rect 2010 -430 2040 -240
rect 2950 -310 2980 -240
rect 2950 -350 2980 -340
rect 2010 -470 2040 -460
rect 1950 -610 1980 -520
rect 3680 -550 3710 -240
rect 3770 -310 3800 -240
rect 3770 -350 3800 -340
rect 3890 -310 3920 -240
rect 3890 -350 3920 -340
rect 3680 -590 3710 -580
rect 1950 -730 1980 -640
rect 1890 -790 1920 -780
rect 1070 -1150 1100 -1140
rect 1070 -1250 1100 -1180
rect 1890 -1250 1920 -820
rect 1950 -850 1980 -760
rect 1950 -970 1980 -880
rect 1950 -1090 1980 -1000
rect 1950 -1210 1980 -1120
rect 1950 -1250 1980 -1240
rect 2010 -670 2040 -660
rect 2010 -1250 2040 -700
rect 3680 -790 3710 -780
rect 2950 -1150 2980 -1140
rect 2950 -1250 2980 -1180
rect 3680 -1250 3710 -820
rect 4710 -790 4740 -240
rect 5440 -310 5470 -240
rect 5440 -350 5470 -340
rect 6380 -670 6410 -240
rect 6380 -710 6410 -700
rect 6440 -250 6470 -240
rect 6440 -370 6470 -280
rect 6440 -490 6470 -400
rect 6440 -610 6470 -520
rect 6440 -730 6470 -640
rect 6440 -770 6470 -760
rect 4710 -830 4740 -820
rect 6500 -790 6530 -240
rect 7320 -310 7350 -240
rect 7320 -350 7350 -340
rect 6500 -830 6530 -820
rect 4710 -910 4740 -900
rect 4500 -1150 4530 -1140
rect 4500 -1250 4530 -1180
rect 4620 -1150 4650 -1140
rect 4620 -1250 4650 -1180
rect 4710 -1250 4740 -940
rect 6500 -910 6530 -900
rect 6440 -970 6470 -960
rect 6380 -1030 6410 -1020
rect 5440 -1150 5470 -1140
rect 5440 -1250 5470 -1180
rect 6380 -1250 6410 -1060
rect 6440 -1090 6470 -1000
rect 6440 -1210 6470 -1120
rect 6440 -1250 6470 -1240
rect 6500 -1250 6530 -940
rect 7320 -1150 7350 -1140
rect 7320 -1250 7350 -1180
rect 940 -1340 990 -1330
rect 940 -1370 950 -1340
rect 980 -1370 990 -1340
rect 940 -1380 990 -1370
rect 7430 -1340 7480 -1330
rect 7430 -1370 7440 -1340
rect 7470 -1370 7480 -1340
rect 7430 -1380 7480 -1370
rect 950 -4090 980 -4070
rect 7440 -4090 7470 -4070
rect 940 -4100 990 -4090
rect 940 -4130 950 -4100
rect 980 -4130 990 -4100
rect 940 -4140 990 -4130
rect 1790 -4100 1840 -4090
rect 1790 -4130 1800 -4100
rect 1830 -4130 1840 -4100
rect 1790 -4140 1840 -4130
rect 6580 -4100 6630 -4090
rect 6580 -4130 6590 -4100
rect 6620 -4130 6630 -4100
rect 6580 -4140 6630 -4130
rect 7430 -4100 7480 -4090
rect 7430 -4130 7440 -4100
rect 7470 -4130 7480 -4100
rect 7430 -4140 7480 -4130
rect 950 -5010 980 -4140
rect 2730 -4170 2780 -4160
rect 2730 -4200 2740 -4170
rect 2770 -4200 2780 -4170
rect 2730 -4210 2780 -4200
rect 5640 -4170 5690 -4160
rect 5640 -4200 5650 -4170
rect 5680 -4200 5690 -4170
rect 5640 -4210 5690 -4200
rect 950 -5160 980 -5150
rect 1800 -5010 1830 -4220
rect 2740 -4370 2770 -4220
rect 2740 -4520 2770 -4510
rect 1800 -5160 1830 -5150
rect 3680 -5010 3710 -4220
rect 3680 -5160 3710 -5150
rect 3770 -5010 3800 -4220
rect 3770 -5160 3800 -5150
rect 4710 -5010 4740 -4220
rect 5650 -4370 5680 -4220
rect 5650 -4520 5680 -4510
rect 4710 -5160 4740 -5150
rect 6590 -5010 6620 -4220
rect 6590 -5160 6620 -5150
rect 7440 -5010 7470 -4140
rect 7440 -5160 7470 -5150
<< via1 >>
rect -1340 -280 -1310 -250
rect -1340 -400 -1310 -370
rect -1340 -520 -1310 -490
rect -1340 -640 -1310 -610
rect -1340 -760 -1310 -730
rect -1340 -880 -1310 -850
rect -1340 -1000 -1310 -970
rect -1340 -1120 -1310 -1090
rect -1340 -1240 -1310 -1210
rect 950 3520 980 3660
rect 1800 3520 1830 3660
rect 3680 3520 3710 3660
rect 2740 2880 2770 3020
rect 4620 3520 4650 3660
rect 4710 3520 4740 3660
rect 6590 3520 6620 3660
rect 5650 2880 5680 3020
rect 7440 3520 7470 3660
rect 1070 -340 1100 -310
rect 1890 -580 1920 -550
rect 1950 -280 1980 -250
rect 1950 -400 1980 -370
rect 2950 -340 2980 -310
rect 2010 -460 2040 -430
rect 1950 -520 1980 -490
rect 3770 -340 3800 -310
rect 3890 -340 3920 -310
rect 3680 -580 3710 -550
rect 1950 -640 1980 -610
rect 1950 -760 1980 -730
rect 1890 -820 1920 -790
rect 1070 -1180 1100 -1150
rect 1950 -880 1980 -850
rect 1950 -1000 1980 -970
rect 1950 -1120 1980 -1090
rect 1950 -1240 1980 -1210
rect 2010 -700 2040 -670
rect 3680 -820 3710 -790
rect 2950 -1180 2980 -1150
rect 5440 -340 5470 -310
rect 6380 -700 6410 -670
rect 6440 -280 6470 -250
rect 6440 -400 6470 -370
rect 6440 -520 6470 -490
rect 6440 -640 6470 -610
rect 6440 -760 6470 -730
rect 4710 -820 4740 -790
rect 7320 -340 7350 -310
rect 6500 -820 6530 -790
rect 4710 -940 4740 -910
rect 4500 -1180 4530 -1150
rect 4620 -1180 4650 -1150
rect 6500 -940 6530 -910
rect 6440 -1000 6470 -970
rect 6380 -1060 6410 -1030
rect 5440 -1180 5470 -1150
rect 6440 -1120 6470 -1090
rect 6440 -1240 6470 -1210
rect 7320 -1180 7350 -1150
rect 950 -5150 980 -5010
rect 2740 -4510 2770 -4370
rect 1800 -5150 1830 -5010
rect 3680 -5150 3710 -5010
rect 3770 -5150 3800 -5010
rect 5650 -4510 5680 -4370
rect 4710 -5150 4740 -5010
rect 6590 -5150 6620 -5010
rect 7440 -5150 7470 -5010
<< metal2 >>
rect -150 3660 8570 3670
rect -150 3520 -140 3660
rect 0 3520 950 3660
rect 980 3520 1800 3660
rect 1830 3520 3680 3660
rect 3710 3520 4620 3660
rect 4650 3520 4710 3660
rect 4740 3520 6590 3660
rect 6620 3520 7440 3660
rect 7470 3520 8420 3660
rect 8560 3520 8570 3660
rect -150 3510 8570 3520
rect 170 3340 8250 3350
rect 170 3200 180 3340
rect 320 3200 8100 3340
rect 8240 3200 8250 3340
rect 170 3190 8250 3200
rect 490 3020 7930 3030
rect 490 2880 500 3020
rect 640 2880 2740 3020
rect 2770 2880 5650 3020
rect 5680 2880 7780 3020
rect 7920 2880 7930 3020
rect 490 2870 7930 2880
rect -1350 -250 -1300 -240
rect -1250 -250 -1200 -240
rect -1050 -250 -1000 -240
rect -850 -250 -800 -240
rect -650 -250 -600 -240
rect -450 -250 -400 -240
rect -250 -250 -200 -240
rect -1350 -280 -1340 -250
rect -1310 -280 -1240 -250
rect -1210 -280 -1040 -250
rect -1010 -280 -840 -250
rect -810 -280 -640 -250
rect -610 -280 -440 -250
rect -410 -280 -240 -250
rect -210 -280 180 -250
rect 320 -280 1950 -250
rect 1980 -280 6440 -250
rect 6470 -280 7500 -250
rect -1350 -290 -1300 -280
rect -1250 -290 -1200 -280
rect -1050 -290 -1000 -280
rect -850 -290 -800 -280
rect -650 -290 -600 -280
rect -450 -290 -400 -280
rect -250 -290 -200 -280
rect -1150 -310 -1100 -300
rect -1340 -340 -1140 -310
rect -1110 -340 1070 -310
rect 1100 -340 2950 -310
rect 2980 -340 3770 -310
rect 3800 -340 3890 -310
rect 3920 -340 5440 -310
rect 5470 -340 7320 -310
rect 7350 -340 7500 -310
rect -1150 -350 -1100 -340
rect -1350 -370 -1300 -360
rect -1250 -370 -1200 -360
rect -1050 -370 -1000 -360
rect -850 -370 -800 -360
rect -650 -370 -600 -360
rect -450 -370 -400 -360
rect -250 -370 -200 -360
rect -1350 -400 -1340 -370
rect -1310 -400 -1240 -370
rect -1210 -400 -1040 -370
rect -1010 -400 -840 -370
rect -810 -400 -640 -370
rect -610 -400 -440 -370
rect -410 -400 -240 -370
rect -210 -400 180 -370
rect 320 -400 1950 -370
rect 1980 -400 6440 -370
rect 6470 -400 7500 -370
rect -1350 -410 -1300 -400
rect -1250 -410 -1200 -400
rect -1050 -410 -1000 -400
rect -850 -410 -800 -400
rect -650 -410 -600 -400
rect -450 -410 -400 -400
rect -250 -410 -200 -400
rect -950 -430 -900 -420
rect -1340 -460 -940 -430
rect -910 -460 2010 -430
rect 2040 -460 7500 -430
rect -950 -470 -900 -460
rect -1350 -490 -1300 -480
rect -1250 -490 -1200 -480
rect -1050 -490 -1000 -480
rect -850 -490 -800 -480
rect -650 -490 -600 -480
rect -450 -490 -400 -480
rect -250 -490 -200 -480
rect -1350 -520 -1340 -490
rect -1310 -520 -1240 -490
rect -1210 -520 -1040 -490
rect -1010 -520 -840 -490
rect -810 -520 -640 -490
rect -610 -520 -440 -490
rect -410 -520 -240 -490
rect -210 -520 180 -490
rect 320 -520 1950 -490
rect 1980 -520 6440 -490
rect 6470 -520 7500 -490
rect -1350 -530 -1300 -520
rect -1250 -530 -1200 -520
rect -1050 -530 -1000 -520
rect -850 -530 -800 -520
rect -650 -530 -600 -520
rect -450 -530 -400 -520
rect -250 -530 -200 -520
rect -750 -550 -700 -540
rect -1340 -580 -740 -550
rect -710 -580 1890 -550
rect 1920 -580 3680 -550
rect 3710 -580 7500 -550
rect -750 -590 -700 -580
rect -1350 -610 -1300 -600
rect -1250 -610 -1200 -600
rect -1050 -610 -1000 -600
rect -850 -610 -800 -600
rect -650 -610 -600 -600
rect -450 -610 -400 -600
rect -250 -610 -200 -600
rect -1350 -640 -1340 -610
rect -1310 -640 -1240 -610
rect -1210 -640 -1040 -610
rect -1010 -640 -840 -610
rect -810 -640 -640 -610
rect -610 -640 -440 -610
rect -410 -640 -240 -610
rect -210 -640 180 -610
rect 320 -640 1950 -610
rect 1980 -640 6440 -610
rect 6470 -640 7500 -610
rect -1350 -650 -1300 -640
rect -1250 -650 -1200 -640
rect -1050 -650 -1000 -640
rect -850 -650 -800 -640
rect -650 -650 -600 -640
rect -450 -650 -400 -640
rect -250 -650 -200 -640
rect -550 -670 -500 -660
rect -1340 -700 -540 -670
rect -510 -700 2010 -670
rect 2040 -700 6380 -670
rect 6410 -700 7500 -670
rect -550 -710 -500 -700
rect -1350 -730 -1300 -720
rect -1250 -730 -1200 -720
rect -1050 -730 -1000 -720
rect -850 -730 -800 -720
rect -650 -730 -600 -720
rect -450 -730 -400 -720
rect -250 -730 -200 -720
rect -1350 -760 -1340 -730
rect -1310 -760 -1240 -730
rect -1210 -760 -1040 -730
rect -1010 -760 -840 -730
rect -810 -760 -640 -730
rect -610 -760 -440 -730
rect -410 -760 -240 -730
rect -210 -760 180 -730
rect 320 -760 1950 -730
rect 1980 -760 6440 -730
rect 6470 -760 7500 -730
rect -1350 -770 -1300 -760
rect -1250 -770 -1200 -760
rect -1050 -770 -1000 -760
rect -850 -770 -800 -760
rect -650 -770 -600 -760
rect -450 -770 -400 -760
rect -250 -770 -200 -760
rect -350 -790 -300 -780
rect -1340 -820 -340 -790
rect -310 -820 1890 -790
rect 1920 -820 3680 -790
rect 3710 -820 4710 -790
rect 4740 -820 6500 -790
rect 6530 -820 7500 -790
rect -350 -830 -300 -820
rect -1350 -850 -1300 -840
rect -1250 -850 -1200 -840
rect -1050 -850 -1000 -840
rect -850 -850 -800 -840
rect -650 -850 -600 -840
rect -450 -850 -400 -840
rect -250 -850 -200 -840
rect -1350 -880 -1340 -850
rect -1310 -880 -1240 -850
rect -1210 -880 -1040 -850
rect -1010 -880 -840 -850
rect -810 -880 -640 -850
rect -610 -880 -440 -850
rect -410 -880 -240 -850
rect -210 -880 180 -850
rect 320 -880 1950 -850
rect 1980 -880 7500 -850
rect -1350 -890 -1300 -880
rect -1250 -890 -1200 -880
rect -1050 -890 -1000 -880
rect -850 -890 -800 -880
rect -650 -890 -600 -880
rect -450 -890 -400 -880
rect -250 -890 -200 -880
rect -750 -910 -700 -900
rect -1340 -940 -740 -910
rect -710 -940 4710 -910
rect 4740 -940 6500 -910
rect 6530 -940 7500 -910
rect -750 -950 -700 -940
rect -1350 -970 -1300 -960
rect -1250 -970 -1200 -960
rect -1050 -970 -1000 -960
rect -850 -970 -800 -960
rect -650 -970 -600 -960
rect -450 -970 -400 -960
rect -250 -970 -200 -960
rect -1350 -1000 -1340 -970
rect -1310 -1000 -1240 -970
rect -1210 -1000 -1040 -970
rect -1010 -1000 -840 -970
rect -810 -1000 -640 -970
rect -610 -1000 -440 -970
rect -410 -1000 -240 -970
rect -210 -1000 180 -970
rect 320 -1000 1950 -970
rect 1980 -1000 6440 -970
rect 6470 -1000 7500 -970
rect -1350 -1010 -1300 -1000
rect -1250 -1010 -1200 -1000
rect -1050 -1010 -1000 -1000
rect -850 -1010 -800 -1000
rect -650 -1010 -600 -1000
rect -450 -1010 -400 -1000
rect -250 -1010 -200 -1000
rect -950 -1030 -900 -1020
rect -1340 -1060 -940 -1030
rect -910 -1060 6380 -1030
rect 6410 -1060 7500 -1030
rect -950 -1070 -900 -1060
rect -1350 -1090 -1300 -1080
rect -1250 -1090 -1200 -1080
rect -1050 -1090 -1000 -1080
rect -850 -1090 -800 -1080
rect -650 -1090 -600 -1080
rect -450 -1090 -400 -1080
rect -250 -1090 -200 -1080
rect -1350 -1120 -1340 -1090
rect -1310 -1120 -1240 -1090
rect -1210 -1120 -1040 -1090
rect -1010 -1120 -840 -1090
rect -810 -1120 -640 -1090
rect -610 -1120 -440 -1090
rect -410 -1120 -240 -1090
rect -210 -1120 180 -1090
rect 320 -1120 1950 -1090
rect 1980 -1120 6440 -1090
rect 6470 -1120 7500 -1090
rect -1350 -1130 -1300 -1120
rect -1250 -1130 -1200 -1120
rect -1050 -1130 -1000 -1120
rect -850 -1130 -800 -1120
rect -650 -1130 -600 -1120
rect -450 -1130 -400 -1120
rect -250 -1130 -200 -1120
rect -1150 -1150 -1100 -1140
rect -1340 -1180 -1140 -1150
rect -1110 -1180 1070 -1150
rect 1100 -1180 2950 -1150
rect 2980 -1180 4500 -1150
rect 4530 -1180 4620 -1150
rect 4650 -1180 5440 -1150
rect 5470 -1180 7320 -1150
rect 7350 -1180 7500 -1150
rect -1150 -1190 -1100 -1180
rect -1350 -1210 -1300 -1200
rect -1250 -1210 -1200 -1200
rect -1050 -1210 -1000 -1200
rect -850 -1210 -800 -1200
rect -650 -1210 -600 -1200
rect -450 -1210 -400 -1200
rect -250 -1210 -200 -1200
rect -1350 -1240 -1340 -1210
rect -1310 -1240 -1240 -1210
rect -1210 -1240 -1040 -1210
rect -1010 -1240 -840 -1210
rect -810 -1240 -640 -1210
rect -610 -1240 -440 -1210
rect -410 -1240 -240 -1210
rect -210 -1240 180 -1210
rect 320 -1240 1950 -1210
rect 1980 -1240 6440 -1210
rect 6470 -1240 7500 -1210
rect -1350 -1250 -1300 -1240
rect -1250 -1250 -1200 -1240
rect -1050 -1250 -1000 -1240
rect -850 -1250 -800 -1240
rect -650 -1250 -600 -1240
rect -450 -1250 -400 -1240
rect -250 -1250 -200 -1240
rect 490 -4370 7930 -4360
rect 490 -4510 500 -4370
rect 640 -4510 2740 -4370
rect 2770 -4510 5650 -4370
rect 5680 -4510 7780 -4370
rect 7920 -4510 7930 -4370
rect 490 -4520 7930 -4510
rect 170 -4690 8250 -4680
rect 170 -4830 180 -4690
rect 320 -4830 8100 -4690
rect 8240 -4830 8250 -4690
rect 170 -4840 8250 -4830
rect -150 -5010 8570 -5000
rect -150 -5150 -140 -5010
rect 0 -5150 950 -5010
rect 980 -5150 1800 -5010
rect 1830 -5150 3680 -5010
rect 3710 -5150 3770 -5010
rect 3800 -5150 4710 -5010
rect 4740 -5150 6590 -5010
rect 6620 -5150 7440 -5010
rect 7470 -5150 8420 -5010
rect 8560 -5150 8570 -5010
rect -150 -5160 8570 -5150
<< via2 >>
rect -140 3520 0 3660
rect 8420 3520 8560 3660
rect 180 3200 320 3340
rect 8100 3200 8240 3340
rect 500 2880 640 3020
rect 7780 2880 7920 3020
rect -1340 -280 -1310 -250
rect -1240 -280 -1210 -250
rect -1040 -280 -1010 -250
rect -840 -280 -810 -250
rect -640 -280 -610 -250
rect -440 -280 -410 -250
rect -240 -280 -210 -250
rect 180 -280 320 -250
rect -1140 -340 -1110 -310
rect -1340 -400 -1310 -370
rect -1240 -400 -1210 -370
rect -1040 -400 -1010 -370
rect -840 -400 -810 -370
rect -640 -400 -610 -370
rect -440 -400 -410 -370
rect -240 -400 -210 -370
rect 180 -400 320 -370
rect -940 -460 -910 -430
rect -1340 -520 -1310 -490
rect -1240 -520 -1210 -490
rect -1040 -520 -1010 -490
rect -840 -520 -810 -490
rect -640 -520 -610 -490
rect -440 -520 -410 -490
rect -240 -520 -210 -490
rect 180 -520 320 -490
rect -740 -580 -710 -550
rect -1340 -640 -1310 -610
rect -1240 -640 -1210 -610
rect -1040 -640 -1010 -610
rect -840 -640 -810 -610
rect -640 -640 -610 -610
rect -440 -640 -410 -610
rect -240 -640 -210 -610
rect 180 -640 320 -610
rect -540 -700 -510 -670
rect -1340 -760 -1310 -730
rect -1240 -760 -1210 -730
rect -1040 -760 -1010 -730
rect -840 -760 -810 -730
rect -640 -760 -610 -730
rect -440 -760 -410 -730
rect -240 -760 -210 -730
rect 180 -760 320 -730
rect -340 -820 -310 -790
rect -1340 -880 -1310 -850
rect -1240 -880 -1210 -850
rect -1040 -880 -1010 -850
rect -840 -880 -810 -850
rect -640 -880 -610 -850
rect -440 -880 -410 -850
rect -240 -880 -210 -850
rect 180 -880 320 -850
rect -740 -940 -710 -910
rect -1340 -1000 -1310 -970
rect -1240 -1000 -1210 -970
rect -1040 -1000 -1010 -970
rect -840 -1000 -810 -970
rect -640 -1000 -610 -970
rect -440 -1000 -410 -970
rect -240 -1000 -210 -970
rect 180 -1000 320 -970
rect -940 -1060 -910 -1030
rect -1340 -1120 -1310 -1090
rect -1240 -1120 -1210 -1090
rect -1040 -1120 -1010 -1090
rect -840 -1120 -810 -1090
rect -640 -1120 -610 -1090
rect -440 -1120 -410 -1090
rect -240 -1120 -210 -1090
rect 180 -1120 320 -1090
rect -1140 -1180 -1110 -1150
rect -1340 -1240 -1310 -1210
rect -1240 -1240 -1210 -1210
rect -1040 -1240 -1010 -1210
rect -840 -1240 -810 -1210
rect -640 -1240 -610 -1210
rect -440 -1240 -410 -1210
rect -240 -1240 -210 -1210
rect 180 -1240 320 -1210
rect 500 -4510 640 -4370
rect 7780 -4510 7920 -4370
rect 180 -4830 320 -4690
rect 8100 -4830 8240 -4690
rect -140 -5150 0 -5010
rect 8420 -5150 8560 -5010
<< metal3 >>
rect -1340 -240 -1310 3670
rect -1240 -240 -1210 3670
rect -1350 -250 -1300 -240
rect -1350 -280 -1340 -250
rect -1310 -280 -1300 -250
rect -1350 -290 -1300 -280
rect -1250 -250 -1200 -240
rect -1250 -280 -1240 -250
rect -1210 -280 -1200 -250
rect -1250 -290 -1200 -280
rect -1340 -360 -1310 -290
rect -1240 -360 -1210 -290
rect -1140 -300 -1110 3700
rect -1040 -240 -1010 3670
rect -1050 -250 -1000 -240
rect -1050 -280 -1040 -250
rect -1010 -280 -1000 -250
rect -1050 -290 -1000 -280
rect -1150 -310 -1100 -300
rect -1150 -340 -1140 -310
rect -1110 -340 -1100 -310
rect -1150 -350 -1100 -340
rect -1350 -370 -1300 -360
rect -1350 -400 -1340 -370
rect -1310 -400 -1300 -370
rect -1350 -410 -1300 -400
rect -1250 -370 -1200 -360
rect -1250 -400 -1240 -370
rect -1210 -400 -1200 -370
rect -1250 -410 -1200 -400
rect -1340 -480 -1310 -410
rect -1240 -480 -1210 -410
rect -1350 -490 -1300 -480
rect -1350 -520 -1340 -490
rect -1310 -520 -1300 -490
rect -1350 -530 -1300 -520
rect -1250 -490 -1200 -480
rect -1250 -520 -1240 -490
rect -1210 -520 -1200 -490
rect -1250 -530 -1200 -520
rect -1340 -600 -1310 -530
rect -1240 -600 -1210 -530
rect -1350 -610 -1300 -600
rect -1350 -640 -1340 -610
rect -1310 -640 -1300 -610
rect -1350 -650 -1300 -640
rect -1250 -610 -1200 -600
rect -1250 -640 -1240 -610
rect -1210 -640 -1200 -610
rect -1250 -650 -1200 -640
rect -1340 -720 -1310 -650
rect -1240 -720 -1210 -650
rect -1350 -730 -1300 -720
rect -1350 -760 -1340 -730
rect -1310 -760 -1300 -730
rect -1350 -770 -1300 -760
rect -1250 -730 -1200 -720
rect -1250 -760 -1240 -730
rect -1210 -760 -1200 -730
rect -1250 -770 -1200 -760
rect -1340 -840 -1310 -770
rect -1240 -840 -1210 -770
rect -1350 -850 -1300 -840
rect -1350 -880 -1340 -850
rect -1310 -880 -1300 -850
rect -1350 -890 -1300 -880
rect -1250 -850 -1200 -840
rect -1250 -880 -1240 -850
rect -1210 -880 -1200 -850
rect -1250 -890 -1200 -880
rect -1340 -960 -1310 -890
rect -1240 -960 -1210 -890
rect -1350 -970 -1300 -960
rect -1350 -1000 -1340 -970
rect -1310 -1000 -1300 -970
rect -1350 -1010 -1300 -1000
rect -1250 -970 -1200 -960
rect -1250 -1000 -1240 -970
rect -1210 -1000 -1200 -970
rect -1250 -1010 -1200 -1000
rect -1340 -1080 -1310 -1010
rect -1240 -1080 -1210 -1010
rect -1350 -1090 -1300 -1080
rect -1350 -1120 -1340 -1090
rect -1310 -1120 -1300 -1090
rect -1350 -1130 -1300 -1120
rect -1250 -1090 -1200 -1080
rect -1250 -1120 -1240 -1090
rect -1210 -1120 -1200 -1090
rect -1250 -1130 -1200 -1120
rect -1340 -1200 -1310 -1130
rect -1240 -1200 -1210 -1130
rect -1140 -1140 -1110 -350
rect -1040 -360 -1010 -290
rect -1050 -370 -1000 -360
rect -1050 -400 -1040 -370
rect -1010 -400 -1000 -370
rect -1050 -410 -1000 -400
rect -1040 -480 -1010 -410
rect -940 -420 -910 3700
rect -840 -240 -810 3670
rect -850 -250 -800 -240
rect -850 -280 -840 -250
rect -810 -280 -800 -250
rect -850 -290 -800 -280
rect -840 -360 -810 -290
rect -850 -370 -800 -360
rect -850 -400 -840 -370
rect -810 -400 -800 -370
rect -850 -410 -800 -400
rect -950 -430 -900 -420
rect -950 -460 -940 -430
rect -910 -460 -900 -430
rect -950 -470 -900 -460
rect -1050 -490 -1000 -480
rect -1050 -520 -1040 -490
rect -1010 -520 -1000 -490
rect -1050 -530 -1000 -520
rect -1040 -600 -1010 -530
rect -1050 -610 -1000 -600
rect -1050 -640 -1040 -610
rect -1010 -640 -1000 -610
rect -1050 -650 -1000 -640
rect -1040 -720 -1010 -650
rect -1050 -730 -1000 -720
rect -1050 -760 -1040 -730
rect -1010 -760 -1000 -730
rect -1050 -770 -1000 -760
rect -1040 -840 -1010 -770
rect -1050 -850 -1000 -840
rect -1050 -880 -1040 -850
rect -1010 -880 -1000 -850
rect -1050 -890 -1000 -880
rect -1040 -960 -1010 -890
rect -1050 -970 -1000 -960
rect -1050 -1000 -1040 -970
rect -1010 -1000 -1000 -970
rect -1050 -1010 -1000 -1000
rect -1040 -1080 -1010 -1010
rect -940 -1020 -910 -470
rect -840 -480 -810 -410
rect -850 -490 -800 -480
rect -850 -520 -840 -490
rect -810 -520 -800 -490
rect -850 -530 -800 -520
rect -840 -600 -810 -530
rect -740 -540 -710 3700
rect -640 -240 -610 3670
rect -650 -250 -600 -240
rect -650 -280 -640 -250
rect -610 -280 -600 -250
rect -650 -290 -600 -280
rect -640 -360 -610 -290
rect -650 -370 -600 -360
rect -650 -400 -640 -370
rect -610 -400 -600 -370
rect -650 -410 -600 -400
rect -640 -480 -610 -410
rect -650 -490 -600 -480
rect -650 -520 -640 -490
rect -610 -520 -600 -490
rect -650 -530 -600 -520
rect -750 -550 -700 -540
rect -750 -580 -740 -550
rect -710 -580 -700 -550
rect -750 -590 -700 -580
rect -850 -610 -800 -600
rect -850 -640 -840 -610
rect -810 -640 -800 -610
rect -850 -650 -800 -640
rect -840 -720 -810 -650
rect -850 -730 -800 -720
rect -850 -760 -840 -730
rect -810 -760 -800 -730
rect -850 -770 -800 -760
rect -840 -840 -810 -770
rect -850 -850 -800 -840
rect -850 -880 -840 -850
rect -810 -880 -800 -850
rect -850 -890 -800 -880
rect -840 -960 -810 -890
rect -740 -900 -710 -590
rect -640 -600 -610 -530
rect -650 -610 -600 -600
rect -650 -640 -640 -610
rect -610 -640 -600 -610
rect -650 -650 -600 -640
rect -640 -720 -610 -650
rect -540 -660 -510 3700
rect -440 -240 -410 3670
rect -450 -250 -400 -240
rect -450 -280 -440 -250
rect -410 -280 -400 -250
rect -450 -290 -400 -280
rect -440 -360 -410 -290
rect -450 -370 -400 -360
rect -450 -400 -440 -370
rect -410 -400 -400 -370
rect -450 -410 -400 -400
rect -440 -480 -410 -410
rect -450 -490 -400 -480
rect -450 -520 -440 -490
rect -410 -520 -400 -490
rect -450 -530 -400 -520
rect -440 -600 -410 -530
rect -450 -610 -400 -600
rect -450 -640 -440 -610
rect -410 -640 -400 -610
rect -450 -650 -400 -640
rect -550 -670 -500 -660
rect -550 -700 -540 -670
rect -510 -700 -500 -670
rect -550 -710 -500 -700
rect -650 -730 -600 -720
rect -650 -760 -640 -730
rect -610 -760 -600 -730
rect -650 -770 -600 -760
rect -640 -840 -610 -770
rect -650 -850 -600 -840
rect -650 -880 -640 -850
rect -610 -880 -600 -850
rect -650 -890 -600 -880
rect -750 -910 -700 -900
rect -750 -940 -740 -910
rect -710 -940 -700 -910
rect -750 -950 -700 -940
rect -850 -970 -800 -960
rect -850 -1000 -840 -970
rect -810 -1000 -800 -970
rect -850 -1010 -800 -1000
rect -950 -1030 -900 -1020
rect -950 -1060 -940 -1030
rect -910 -1060 -900 -1030
rect -950 -1070 -900 -1060
rect -1050 -1090 -1000 -1080
rect -1050 -1120 -1040 -1090
rect -1010 -1120 -1000 -1090
rect -1050 -1130 -1000 -1120
rect -1150 -1150 -1100 -1140
rect -1150 -1180 -1140 -1150
rect -1110 -1180 -1100 -1150
rect -1150 -1190 -1100 -1180
rect -1350 -1210 -1300 -1200
rect -1350 -1240 -1340 -1210
rect -1310 -1240 -1300 -1210
rect -1350 -1250 -1300 -1240
rect -1250 -1210 -1200 -1200
rect -1250 -1240 -1240 -1210
rect -1210 -1240 -1200 -1210
rect -1250 -1250 -1200 -1240
rect -1340 -5160 -1310 -1250
rect -1240 -5160 -1210 -1250
rect -1140 -5160 -1110 -1190
rect -1040 -1200 -1010 -1130
rect -1050 -1210 -1000 -1200
rect -1050 -1240 -1040 -1210
rect -1010 -1240 -1000 -1210
rect -1050 -1250 -1000 -1240
rect -1040 -5160 -1010 -1250
rect -940 -5160 -910 -1070
rect -840 -1080 -810 -1010
rect -850 -1090 -800 -1080
rect -850 -1120 -840 -1090
rect -810 -1120 -800 -1090
rect -850 -1130 -800 -1120
rect -840 -1200 -810 -1130
rect -850 -1210 -800 -1200
rect -850 -1240 -840 -1210
rect -810 -1240 -800 -1210
rect -850 -1250 -800 -1240
rect -840 -5160 -810 -1250
rect -740 -5160 -710 -950
rect -640 -960 -610 -890
rect -650 -970 -600 -960
rect -650 -1000 -640 -970
rect -610 -1000 -600 -970
rect -650 -1010 -600 -1000
rect -640 -1080 -610 -1010
rect -650 -1090 -600 -1080
rect -650 -1120 -640 -1090
rect -610 -1120 -600 -1090
rect -650 -1130 -600 -1120
rect -640 -1200 -610 -1130
rect -650 -1210 -600 -1200
rect -650 -1240 -640 -1210
rect -610 -1240 -600 -1210
rect -650 -1250 -600 -1240
rect -640 -5160 -610 -1250
rect -540 -5160 -510 -710
rect -440 -720 -410 -650
rect -450 -730 -400 -720
rect -450 -760 -440 -730
rect -410 -760 -400 -730
rect -450 -770 -400 -760
rect -440 -840 -410 -770
rect -340 -780 -310 3700
rect -240 -240 -210 3670
rect -150 3660 10 3700
rect -150 3520 -140 3660
rect 0 3520 10 3660
rect -250 -250 -200 -240
rect -250 -280 -240 -250
rect -210 -280 -200 -250
rect -250 -290 -200 -280
rect -240 -360 -210 -290
rect -250 -370 -200 -360
rect -250 -400 -240 -370
rect -210 -400 -200 -370
rect -250 -410 -200 -400
rect -240 -480 -210 -410
rect -250 -490 -200 -480
rect -250 -520 -240 -490
rect -210 -520 -200 -490
rect -250 -530 -200 -520
rect -240 -600 -210 -530
rect -250 -610 -200 -600
rect -250 -640 -240 -610
rect -210 -640 -200 -610
rect -250 -650 -200 -640
rect -240 -720 -210 -650
rect -250 -730 -200 -720
rect -250 -760 -240 -730
rect -210 -760 -200 -730
rect -250 -770 -200 -760
rect -350 -790 -300 -780
rect -350 -820 -340 -790
rect -310 -820 -300 -790
rect -350 -830 -300 -820
rect -450 -850 -400 -840
rect -450 -880 -440 -850
rect -410 -880 -400 -850
rect -450 -890 -400 -880
rect -440 -960 -410 -890
rect -450 -970 -400 -960
rect -450 -1000 -440 -970
rect -410 -1000 -400 -970
rect -450 -1010 -400 -1000
rect -440 -1080 -410 -1010
rect -450 -1090 -400 -1080
rect -450 -1120 -440 -1090
rect -410 -1120 -400 -1090
rect -450 -1130 -400 -1120
rect -440 -1200 -410 -1130
rect -450 -1210 -400 -1200
rect -450 -1240 -440 -1210
rect -410 -1240 -400 -1210
rect -450 -1250 -400 -1240
rect -440 -5160 -410 -1250
rect -340 -5160 -310 -830
rect -240 -840 -210 -770
rect -250 -850 -200 -840
rect -250 -880 -240 -850
rect -210 -880 -200 -850
rect -250 -890 -200 -880
rect -240 -960 -210 -890
rect -250 -970 -200 -960
rect -250 -1000 -240 -970
rect -210 -1000 -200 -970
rect -250 -1010 -200 -1000
rect -240 -1080 -210 -1010
rect -250 -1090 -200 -1080
rect -250 -1120 -240 -1090
rect -210 -1120 -200 -1090
rect -250 -1130 -200 -1120
rect -240 -1200 -210 -1130
rect -250 -1210 -200 -1200
rect -250 -1240 -240 -1210
rect -210 -1240 -200 -1210
rect -250 -1250 -200 -1240
rect -240 -5160 -210 -1250
rect -150 -5010 10 3520
rect -150 -5150 -140 -5010
rect 0 -5150 10 -5010
rect -150 -5160 10 -5150
rect 170 3340 330 3700
rect 170 3200 180 3340
rect 320 3200 330 3340
rect 170 -250 330 3200
rect 170 -280 180 -250
rect 320 -280 330 -250
rect 170 -320 330 -280
rect 170 -450 180 -320
rect 320 -450 330 -320
rect 170 -490 330 -450
rect 170 -520 180 -490
rect 320 -520 330 -490
rect 170 -560 330 -520
rect 170 -690 180 -560
rect 320 -690 330 -560
rect 170 -730 330 -690
rect 170 -760 180 -730
rect 320 -760 330 -730
rect 170 -800 330 -760
rect 170 -930 180 -800
rect 320 -930 330 -800
rect 170 -970 330 -930
rect 170 -1000 180 -970
rect 320 -1000 330 -970
rect 170 -1040 330 -1000
rect 170 -1170 180 -1040
rect 320 -1170 330 -1040
rect 170 -1210 330 -1170
rect 170 -1240 180 -1210
rect 320 -1240 330 -1210
rect 170 -4690 330 -1240
rect 170 -4830 180 -4690
rect 320 -4830 330 -4690
rect 170 -5160 330 -4830
rect 490 3020 650 3700
rect 490 2880 500 3020
rect 640 2880 650 3020
rect 490 -4370 650 2880
rect 490 -4510 500 -4370
rect 640 -4510 650 -4370
rect 490 -5160 650 -4510
rect 7770 3020 7930 3670
rect 7770 2880 7780 3020
rect 7920 2880 7930 3020
rect 7770 -4370 7930 2880
rect 7770 -4510 7780 -4370
rect 7920 -4510 7930 -4370
rect 7770 -5160 7930 -4510
rect 8090 3340 8250 3670
rect 8090 3200 8100 3340
rect 8240 3200 8250 3340
rect 8090 -4690 8250 3200
rect 8090 -4830 8100 -4690
rect 8240 -4830 8250 -4690
rect 8090 -5160 8250 -4830
rect 8410 3660 8570 3670
rect 8410 3520 8420 3660
rect 8560 3520 8570 3660
rect 8410 -5010 8570 3520
rect 8410 -5150 8420 -5010
rect 8560 -5150 8570 -5010
rect 8410 -5160 8570 -5150
<< via3 >>
rect 180 -370 320 -320
rect 180 -400 320 -370
rect 180 -450 320 -400
rect 180 -610 320 -560
rect 180 -640 320 -610
rect 180 -690 320 -640
rect 180 -850 320 -800
rect 180 -880 320 -850
rect 180 -930 320 -880
rect 180 -1090 320 -1040
rect 180 -1120 320 -1090
rect 180 -1170 320 -1120
<< metal4 >>
rect -1340 -320 7500 -310
rect -1340 -450 180 -320
rect 320 -450 7500 -320
rect -1340 -460 7500 -450
rect -1340 -560 7500 -550
rect -1340 -690 180 -560
rect 320 -690 7500 -560
rect -1340 -700 7500 -690
rect -1340 -800 7500 -790
rect -1340 -930 180 -800
rect 320 -930 7500 -800
rect -1340 -940 7500 -930
rect -1340 -1040 7500 -1030
rect -1340 -1170 180 -1040
rect 320 -1170 7500 -1040
rect -1340 -1180 7500 -1170
<< metal5 >>
rect -1340 -5160 -1110 3670
rect -940 -5160 -710 3670
rect -540 -5160 -310 3670
use p8_1  p8_1_6
timestamp 1634440961
transform 1 0 920 0 -1 -1250
box 0 0 940 2970
use p8_1  p8_1_5
timestamp 1634440961
transform 1 0 1860 0 -1 -1250
box 0 0 940 2970
use p1_8  p1_8_2 ota/mag
timestamp 1634440922
transform 1 0 2800 0 -1 -1250
box 0 0 940 2970
use p8_1  p8_1_7
timestamp 1634440961
transform -1 0 4680 0 -1 -1250
box 0 0 940 2970
use p1_8  p1_8_3
timestamp 1634440922
transform -1 0 5620 0 -1 -1250
box 0 0 940 2970
use p8_1  p8_1_8
timestamp 1634440961
transform -1 0 6560 0 -1 -1250
box 0 0 940 2970
use p8_1  p8_1_9
timestamp 1634440961
transform -1 0 7500 0 -1 -1250
box 0 0 940 2970
use p8_1  p8_1_1
timestamp 1634440961
transform 1 0 1860 0 1 -240
box 0 0 940 2970
use p8_1  p8_1_0
timestamp 1634440961
transform 1 0 920 0 1 -240
box 0 0 940 2970
use p1_8  p1_8_0
timestamp 1634440922
transform 1 0 2800 0 1 -240
box 0 0 940 2970
use p8_1  p8_1_2
timestamp 1634440961
transform 1 0 3740 0 1 -240
box 0 0 940 2970
use p1_8  p1_8_1
timestamp 1634440922
transform -1 0 5620 0 1 -240
box 0 0 940 2970
use p8_1  p8_1_3
timestamp 1634440961
transform -1 0 6560 0 1 -240
box 0 0 940 2970
use p8_1  p8_1_4
timestamp 1634440961
transform -1 0 7500 0 1 -240
box 0 0 940 2970
<< labels >>
rlabel metal3 -1140 3670 -1110 3700 1 ib
port 1 n
rlabel metal3 -940 3670 -910 3700 1 xa
port 2 n
rlabel metal3 -740 3670 -710 3700 1 ya
port 3 n
rlabel metal3 -540 3670 -510 3700 1 xb
port 4 n
rlabel metal3 -340 3670 -310 3700 1 yb
port 5 n
rlabel metal3 -150 3670 10 3700 1 vdda
port 6 n
rlabel metal3 170 3670 330 3700 1 gnda
port 7 n
rlabel metal3 490 3670 650 3700 1 vssa
port 8 n
<< end >>
