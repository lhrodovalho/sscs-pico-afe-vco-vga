magic
tech sky130A
magscale 1 2
timestamp 1635533344
<< checkpaint >>
rect 9240 27340 12162 31592
<< pwell >>
rect 13078 29800 13080 30000
rect 7758 27180 7760 27380
rect 13038 25920 13040 26120
rect 7860 25400 11020 25640
rect 7758 24020 7760 24220
rect 7758 21300 7760 21500
rect 13018 19680 13020 19880
rect 7838 17840 7840 18040
<< metal1 >>
rect -2100 17580 -1900 33320
rect 120 21100 320 33360
rect 2280 23780 2480 33360
rect 4500 26920 4700 33360
rect 6740 29880 6940 33360
rect 8880 31246 9080 33360
rect 11140 32760 11340 33360
rect 11140 32560 11960 32760
rect 11760 31600 11960 32560
rect 13340 32080 13540 33360
rect 13340 31960 13380 32080
rect 13500 31960 13540 32080
rect 13340 31920 13540 31960
rect 11760 31480 11800 31600
rect 11920 31480 11960 31600
rect 11760 31420 11960 31480
rect 8880 31240 9620 31246
rect 10260 31240 12720 31246
rect 8880 31200 12720 31240
rect 8880 31080 12580 31200
rect 12700 31080 12720 31200
rect 8880 31060 12720 31080
rect 10788 30530 15316 30532
rect 9040 30346 15316 30530
rect 9040 30344 10810 30346
rect 7520 30300 7720 30340
rect 7520 30160 7560 30300
rect 7680 30160 7720 30300
rect 7520 30140 7720 30160
rect 6740 29680 7740 29880
rect 10598 29766 10810 30344
rect 12880 29960 13080 30000
rect 14406 29972 14610 30346
rect 12880 29820 12920 29960
rect 13040 29820 13080 29960
rect 12880 29800 13080 29820
rect 15120 29698 15312 30346
rect 12580 29480 13100 29540
rect 12700 29360 13100 29480
rect 12580 29340 13100 29360
rect 7800 28580 8060 28620
rect 7800 28420 7840 28580
rect 8020 28420 8060 28580
rect 7800 28380 8060 28420
rect 9046 27572 9386 28826
rect 10598 27572 10818 29182
rect 15110 28484 15298 28576
rect 13120 28220 13380 28260
rect 13120 28060 13160 28220
rect 13340 28060 13380 28220
rect 14400 28184 15298 28484
rect 13120 28020 13380 28060
rect 7560 27340 7760 27380
rect 7560 27200 7600 27340
rect 7720 27200 7760 27340
rect 9046 27296 10818 27572
rect 7560 27180 7760 27200
rect 9090 27154 10818 27296
rect 4500 26720 7780 26920
rect 7860 25600 8120 25640
rect 7860 25440 7900 25600
rect 8080 25440 8120 25600
rect 7860 25400 8120 25440
rect 9108 24396 9452 25838
rect 10598 25776 10818 27154
rect 15110 27080 15298 28184
rect 14290 27078 15298 27080
rect 14286 26860 15298 27078
rect 14286 26198 14558 26860
rect 15110 26262 15298 26860
rect 12840 26080 13040 26120
rect 14354 26100 14558 26198
rect 12840 25940 12880 26080
rect 13000 25940 13040 26080
rect 12840 25920 13040 25940
rect 11760 25620 13060 25660
rect 11760 25500 11780 25620
rect 11900 25500 13060 25620
rect 10606 24396 10798 25480
rect 11760 25460 13060 25500
rect 7560 24180 7760 24220
rect 7560 24040 7600 24180
rect 7720 24040 7760 24180
rect 9108 24056 10798 24396
rect 13100 24360 13360 24400
rect 13100 24200 13140 24360
rect 13320 24200 13360 24360
rect 13100 24160 13360 24200
rect 9190 24052 10798 24056
rect 7560 24020 7760 24040
rect 2280 23560 7860 23780
rect 7960 22440 8220 22480
rect 7960 22280 8000 22440
rect 8180 22280 8220 22440
rect 7960 22240 8220 22280
rect 9194 21680 9460 22698
rect 10606 22636 10798 24052
rect 14356 23516 14616 24596
rect 15106 23516 15306 24082
rect 14356 23438 15306 23516
rect 14356 23296 15310 23438
rect 14358 23294 15310 23296
rect 10620 21680 10784 22490
rect 15102 22400 15310 23294
rect 7560 21460 7900 21520
rect 7560 21320 7600 21460
rect 7720 21320 7900 21460
rect 9194 21438 10784 21680
rect 7560 21300 7900 21320
rect 120 20860 7900 21100
rect 10620 20326 10784 21438
rect 14280 21940 15310 22400
rect 14280 21148 14540 21940
rect 15102 21356 15310 21940
rect 14280 21100 14542 21148
rect 8020 19760 8280 19800
rect 8020 19600 8060 19760
rect 8240 19600 8280 19760
rect 8020 19560 8280 19600
rect 9252 19374 9498 19982
rect 10614 19374 10782 19874
rect 12820 19840 13020 19880
rect 14282 19848 14542 21100
rect 12820 19700 12860 19840
rect 12980 19700 13020 19840
rect 12820 19680 13020 19700
rect 9252 19144 10782 19374
rect 11320 19400 13060 19440
rect 11320 19280 11360 19400
rect 11480 19280 13060 19400
rect 11320 19220 13060 19280
rect 10614 18218 10782 19144
rect 7640 18000 7840 18060
rect 7640 17860 7680 18000
rect 7800 17860 7840 18000
rect 9174 17954 10782 18218
rect 7640 17840 7840 17860
rect -2100 17400 7900 17580
rect 10614 16878 10782 17954
rect 13080 18120 13340 18160
rect 13080 17960 13120 18120
rect 13300 17960 13340 18120
rect 13080 17920 13340 17960
rect 7940 16260 8200 16300
rect 7940 16100 7980 16260
rect 8160 16100 8200 16260
rect 7940 16060 8200 16100
rect 9178 16000 9378 16522
rect 10614 16000 10782 16700
rect 14340 16480 14780 18360
rect 15100 16480 15300 16860
rect 14340 16280 15300 16480
rect -4160 15860 -3140 15900
rect -4160 15740 -3460 15860
rect -3240 15740 -3140 15860
rect -4160 15680 -3140 15740
rect 9178 15840 10782 16000
rect 12500 16060 15300 16280
rect 9178 15720 10780 15840
rect 3880 15400 4080 15440
rect 3880 15260 3920 15400
rect 4040 15260 4080 15400
rect -2220 15080 1220 15120
rect -2220 14920 940 15080
rect 1160 14920 1220 15080
rect -2220 14880 1220 14920
rect -2220 14300 -1900 14880
rect 3880 14300 4080 15260
rect 9180 14300 9440 15720
rect 12500 15100 12700 16060
rect 12500 14920 12520 15100
rect 12660 14920 12700 15100
rect 12500 14860 12700 14920
<< via1 >>
rect 13380 31960 13500 32080
rect 11800 31480 11920 31600
rect 12580 31080 12700 31200
rect 7560 30160 7680 30300
rect 12920 29820 13040 29960
rect 12580 29360 12700 29480
rect 7840 28420 8020 28580
rect 13160 28060 13340 28220
rect 7600 27200 7720 27340
rect 7900 25440 8080 25600
rect 12880 25940 13000 26080
rect 11780 25500 11900 25620
rect 7600 24040 7720 24180
rect 13140 24200 13320 24360
rect 8000 22280 8180 22440
rect 7600 21320 7720 21460
rect 8060 19600 8240 19760
rect 12860 19700 12980 19840
rect 11360 19280 11480 19400
rect 7680 17860 7800 18000
rect 13120 17960 13300 18120
rect 7980 16100 8160 16260
rect -3460 15740 -3240 15860
rect 3920 15260 4040 15400
rect 940 14920 1160 15080
rect 12520 14920 12660 15100
<< metal2 >>
rect 11320 32080 13540 32120
rect 11320 31960 13380 32080
rect 13500 31960 13540 32080
rect 11320 31920 13540 31960
rect 7520 30300 7720 30340
rect 7520 30160 7560 30300
rect 7680 30160 7720 30300
rect 7520 30140 7720 30160
rect 7800 28580 8060 28620
rect 7800 28420 7840 28580
rect 8020 28420 8060 28580
rect 7800 28380 8060 28420
rect 7560 27340 7760 27380
rect 7560 27200 7600 27340
rect 7720 27200 7760 27340
rect 7560 27180 7760 27200
rect 7860 25600 8120 25640
rect 7860 25440 7900 25600
rect 8080 25440 8120 25600
rect 7860 25400 8120 25440
rect 7560 24180 7760 24220
rect 7560 24040 7600 24180
rect 7720 24040 7760 24180
rect 7560 24020 7760 24040
rect 7960 22440 8220 22480
rect 7960 22280 8000 22440
rect 8180 22280 8220 22440
rect 7960 22240 8220 22280
rect 7560 21460 7760 21520
rect 7560 21320 7600 21460
rect 7720 21320 7760 21460
rect 7560 21300 7760 21320
rect 8020 19760 8280 19800
rect 8020 19600 8060 19760
rect 8240 19600 8280 19760
rect 8020 19560 8280 19600
rect 11320 19400 11520 31920
rect 11760 31600 11960 31680
rect 11760 31480 11800 31600
rect 11920 31480 11960 31600
rect 11760 25620 11960 31480
rect 12560 31200 12720 31220
rect 12560 31080 12580 31200
rect 12700 31080 12720 31200
rect 12560 29480 12720 31080
rect 12880 29960 13080 30000
rect 12880 29820 12920 29960
rect 13040 29820 13080 29960
rect 12880 29800 13080 29820
rect 12560 29360 12580 29480
rect 12700 29360 12720 29480
rect 12560 29340 12720 29360
rect 13120 28220 13380 28260
rect 13120 28060 13160 28220
rect 13340 28060 13380 28220
rect 13120 28020 13380 28060
rect 12840 26080 13040 26120
rect 12840 25940 12880 26080
rect 13000 25940 13040 26080
rect 12840 25920 13040 25940
rect 11760 25500 11780 25620
rect 11900 25500 11960 25620
rect 11760 25460 11960 25500
rect 13100 24360 13360 24400
rect 13100 24200 13140 24360
rect 13320 24200 13360 24360
rect 13100 24160 13360 24200
rect 12820 19840 13020 19880
rect 12820 19700 12860 19840
rect 12980 19700 13020 19840
rect 12820 19680 13020 19700
rect 11320 19280 11360 19400
rect 11480 19280 11520 19400
rect 11320 19220 11520 19280
rect 13080 18120 13340 18160
rect 7640 18000 7840 18060
rect 7640 17860 7680 18000
rect 7800 17860 7840 18000
rect 13080 17960 13120 18120
rect 13300 17960 13340 18120
rect 13080 17920 13340 17960
rect 7640 17840 7840 17860
rect 7940 16260 8200 16300
rect 7940 16100 7980 16260
rect 8160 16100 8200 16260
rect 7940 16060 8200 16100
rect -3500 15860 -3180 15900
rect -3500 15740 -3460 15860
rect -3240 15740 -3180 15860
rect -3500 15700 -3180 15740
rect 3880 15400 4080 15440
rect 3880 15260 3920 15400
rect 4040 15260 4080 15400
rect 3880 15220 4080 15260
rect 900 15100 12700 15120
rect 900 15080 12520 15100
rect 900 14920 940 15080
rect 1160 14920 12520 15080
rect 12660 14920 12700 15100
rect 900 14880 12700 14920
<< via2 >>
rect 7560 30160 7680 30300
rect 7840 28420 8020 28580
rect 7600 27200 7720 27340
rect 7900 25440 8080 25600
rect 7600 24040 7720 24180
rect 8000 22280 8180 22440
rect 7600 21320 7720 21460
rect 8060 19600 8240 19760
rect 12920 29820 13040 29960
rect 13160 28060 13340 28220
rect 12880 25940 13000 26080
rect 13140 24200 13320 24360
rect 12860 19700 12980 19840
rect 7680 17860 7800 18000
rect 13120 17960 13300 18120
rect 7980 16100 8160 16260
rect -3460 15740 -3240 15860
rect 3920 15260 4040 15400
<< metal3 >>
rect 7520 30300 13080 30340
rect 7520 30160 7560 30300
rect 7680 30160 13080 30300
rect 7520 30140 13080 30160
rect 7800 28580 8060 28620
rect 7800 28420 7840 28580
rect 8020 28420 8060 28580
rect 7800 28380 8060 28420
rect 11100 27380 11300 30140
rect 12880 29960 13080 30140
rect 12880 29820 12920 29960
rect 13040 29820 13080 29960
rect 12880 29800 13080 29820
rect 13120 28220 13380 28260
rect 13120 28060 13160 28220
rect 13340 28060 13380 28220
rect 13120 28020 13380 28060
rect 7560 27340 11300 27380
rect 7560 27200 7600 27340
rect 7720 27200 11300 27340
rect 7560 27180 11300 27200
rect 11100 26120 11300 27180
rect 11100 26080 13040 26120
rect 11100 25940 12880 26080
rect 13000 25940 13040 26080
rect 7860 25600 8120 25640
rect 7860 25440 7900 25600
rect 8080 25440 8120 25600
rect 7860 25400 8120 25440
rect 11100 24220 11300 25940
rect 12840 25920 13040 25940
rect 7560 24180 11300 24220
rect 7560 24040 7600 24180
rect 7720 24040 11300 24180
rect 13100 24360 13360 24400
rect 13100 24200 13140 24360
rect 13320 24200 13360 24360
rect 13100 24160 13360 24200
rect 7560 24020 11300 24040
rect 7960 22440 8220 22480
rect 7960 22280 8000 22440
rect 8180 22280 8220 22440
rect 7960 22240 8220 22280
rect 11100 21520 11300 24020
rect 7560 21460 11300 21520
rect 7560 21320 7600 21460
rect 7720 21320 11300 21460
rect 7560 21300 11300 21320
rect 11100 19880 11300 21300
rect 11100 19840 13020 19880
rect 8020 19760 8280 19800
rect 8020 19600 8060 19760
rect 8240 19600 8280 19760
rect 8020 19560 8280 19600
rect 11100 19700 12860 19840
rect 12980 19700 13020 19840
rect 11100 18060 11300 19700
rect 12820 19680 13020 19700
rect 7640 18000 11300 18060
rect 7640 17860 7680 18000
rect 7800 17860 11300 18000
rect 13080 18120 13340 18160
rect 13080 17960 13120 18120
rect 13300 17960 13340 18120
rect 13080 17920 13340 17960
rect 7640 17840 11300 17860
rect 7940 16260 8200 16300
rect 7940 16100 7980 16260
rect 8160 16100 8200 16260
rect 7940 16060 8200 16100
rect 11100 15900 11300 17840
rect -3500 15860 11300 15900
rect -3500 15740 -3460 15860
rect -3240 15740 11300 15860
rect -3500 15680 11300 15740
rect 3880 15400 4080 15440
rect 3880 15260 3920 15400
rect 4040 15260 4080 15400
rect 3880 15220 4080 15260
<< via3 >>
rect 7840 28420 8020 28580
rect 13160 28060 13340 28220
rect 7900 25440 8080 25600
rect 13140 24200 13320 24360
rect 8000 22280 8180 22440
rect 8060 19600 8240 19760
rect 13120 17960 13300 18120
rect 7980 16100 8160 16260
rect 3920 15260 4040 15400
<< metal4 >>
rect 7800 28580 8060 28620
rect 7800 28420 7840 28580
rect 8020 28420 11040 28580
rect 7800 28380 11040 28420
rect 10840 28280 11040 28380
rect 10840 28220 13380 28280
rect 10840 28060 13160 28220
rect 13340 28060 13380 28220
rect 10840 28020 13380 28060
rect 10840 25640 11040 28020
rect 7860 25600 11040 25640
rect 7860 25440 7900 25600
rect 8080 25440 11040 25600
rect 7860 25400 11040 25440
rect 10840 24400 11040 25400
rect 10840 24360 13360 24400
rect 10840 24200 13140 24360
rect 13320 24200 13360 24360
rect 10840 24160 13360 24200
rect 10840 22480 11040 24160
rect 7960 22440 11040 22480
rect 7960 22280 8000 22440
rect 8180 22280 11040 22440
rect 7960 22240 11040 22280
rect 10840 19800 11040 22240
rect 8020 19760 11040 19800
rect 8020 19600 8060 19760
rect 8240 19600 11040 19760
rect 8020 19560 11040 19600
rect 10840 18160 11040 19560
rect 10840 18120 13340 18160
rect 10840 17960 13120 18120
rect 13300 17960 13340 18120
rect 10840 17920 13340 17960
rect 10840 16300 11040 17920
rect 3860 16260 11040 16300
rect 3860 16100 7980 16260
rect 8160 16100 11040 16260
rect 3860 16060 11040 16100
rect 3860 15400 4100 16060
rect 3860 15260 3920 15400
rect 4040 15260 4100 15400
rect 3860 15220 4100 15260
use tg  tg_1 ~/sky130_skel/dpga-ieee-sscs-contest-main/magic/digpot/tg/mag
timestamp 1634765323
transform 1 0 7320 0 -1 20198
box 440 -1513 2130 610
use tg  tg_0
timestamp 1634765323
transform 1 0 7248 0 -1 16738
box 440 -1513 2130 610
use sky130_fd_pr__res_high_po_0p35_LN2BL5  XR0
timestamp 1634754066
transform 1 0 10701 0 1 16796
box -201 -696 201 696
use sky130_fd_pr__res_high_po_0p35_QTTEB3  XR1
timestamp 1634590722
transform 1 0 10701 0 1 20105
box -201 -805 201 805
use tg  tg_7
timestamp 1634765323
transform 1 0 12410 0 -1 18572
box 440 -1513 2130 610
use sky130_fd_pr__res_xhigh_po_0p35_QSBVTB  XR7
timestamp 1634590722
transform 1 0 15193 0 1 19096
box -201 -2826 201 2826
use tg  tg_3
timestamp 1634765323
transform 1 0 7160 0 -1 26068
box 440 -1513 2130 610
use tg  tg_2
timestamp 1634765323
transform 1 0 7262 0 -1 22914
box 440 -1513 2130 610
use sky130_fd_pr__res_xhigh_po_0p35_3F46MW  XR3
timestamp 1634590722
transform 1 0 10701 0 1 25626
box -201 -726 201 726
use sky130_fd_pr__res_xhigh_po_0p35_X894K9  XR2
timestamp 1634590722
transform 1 0 10701 0 1 22556
box -201 -656 201 656
use tg  tg_6
timestamp 1634765323
transform 1 0 12424 0 -1 24812
box 440 -1513 2130 610
use sky130_fd_pr__res_xhigh_po_0p35_VTENMF  XR6
timestamp 1634590722
transform 1 0 15201 0 1 25171
box -201 -1671 201 1671
use tg  tg_4
timestamp 1634765323
transform 1 0 7118 0 -1 29032
box 440 -1513 2130 610
use sky130_fd_pr__res_xhigh_po_0p35_378WDC  XR4 VGA/./digpot/mag
timestamp 1635533344
transform 1 0 10701 0 1 29466
box 0 0 1 1
use tg  tg_5
timestamp 1634765323
transform 1 0 12474 0 -1 28694
box 440 -1513 2130 610
use sky130_fd_pr__res_xhigh_po_0p35_XPUJF7  XR5
timestamp 1634590722
transform 1 0 15215 0 1 29144
box -201 -1146 201 1146
<< labels >>
flabel metal1 -2100 33120 -1900 33320 4 FreeSans 3200 0 0 0 c0
port 0 nsew
flabel metal1 120 33160 320 33360 4 FreeSans 3200 0 0 0 c1
port 1 nsew
flabel metal1 2280 33160 2480 33360 4 FreeSans 3200 0 0 0 c2
port 2 nsew
flabel metal1 4500 33160 4700 33360 4 FreeSans 3200 0 0 0 c3
port 3 nsew
flabel metal1 6740 33160 6940 33360 4 FreeSans 3200 0 0 0 c4
port 4 nsew
flabel metal1 8880 33160 9080 33360 4 FreeSans 3200 0 0 0 c5
port 5 nsew
flabel metal1 11140 33160 11340 33360 4 FreeSans 3200 0 0 0 c6
port 6 nsew
flabel metal1 13340 33160 13540 33360 4 FreeSans 3200 0 0 0 c7
port 7 nsew
flabel metal1 -4160 15700 -3960 15900 4 FreeSans 3200 90 0 0 gnd
port 8 nsew
flabel metal1 9200 14312 9400 14512 2 FreeSans 3200 0 0 0 n0
port 10 nsew
flabel metal1 3880 14300 4080 14500 2 FreeSans 3200 0 0 0 vd
port 9 nsew
flabel metal1 -2200 14300 -2000 14500 2 FreeSans 3200 0 0 0 n8
port 11 nsew
<< end >>
