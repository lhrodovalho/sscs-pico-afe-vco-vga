* lna-ota buffer testbench

* Include SkyWater sky130 device models
.lib "/usr/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice" tt
.param mc_mm_switch=0
.include "../mag/lna.spice"


* supply voltages
vdda	vdda 0 1.0
vgnda	gnda 0 0.5
vssa	vssa 0 0.0

* input signals
vin	in gnda dc 0 ac 1 SINE(0 50m 1 0 0 0)
einp	ip gnda in gnda  0.5
einm	im gnda in gnda -0.5

vfsb fsb vssa dc 1.0 pulse(0 1.0 1 10m 1m 10 10)

* DUT
x0 ip im op om fsb ib vdda gnda vssa lna
IB   vdda ib 10n
CLP  op gnda 10p
CLM  om gnda 10p

*.save v(in) v(ip) v(im) v(x0.xp) v(x0.xm) v(op) v(om)
.option gmin=1e-14
*.option NOOPITER
.option NOINIT
.option METHOD=Gear
.control
	op
	print ib i(vdda)
	print ip im x0.xp x0.xm op om
	
	ac dec 10 1m 1Meg
	plot vdb(op,om)

	tran 1m 3 100m uic
	plot ip im x0.xm x0.xp op om
	plot ip-im x0.xm-x0.xp op-om
	wrdata ../data/lna_tb_tran.txt ip im x0.xp x0.xm op om
	
*	noise v(op,om) vin dec 10 1 100
*	print inoise_total onoise_total
*	setplot noise1
*	plot inoise_spectrum loglog
    
.endc

.end
