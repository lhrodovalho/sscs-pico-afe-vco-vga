magic
tech sky130A
timestamp 1638390070
<< locali >>
rect 4240 15710 4440 15720
rect 4240 15690 4250 15710
rect 4270 15690 4330 15710
rect 4350 15690 4410 15710
rect 4430 15690 4440 15710
rect 4240 15680 4440 15690
rect 4480 15710 4680 15720
rect 4480 15690 4490 15710
rect 4510 15690 4570 15710
rect 4590 15690 4650 15710
rect 4670 15690 4680 15710
rect 4480 15680 4680 15690
rect 4720 15710 5720 15720
rect 4720 15690 4730 15710
rect 4750 15690 4810 15710
rect 4830 15690 4890 15710
rect 4910 15690 4970 15710
rect 4990 15690 5050 15710
rect 5070 15690 5130 15710
rect 5150 15690 5210 15710
rect 5230 15690 5290 15710
rect 5310 15690 5370 15710
rect 5390 15690 5450 15710
rect 5470 15690 5530 15710
rect 5550 15690 5610 15710
rect 5630 15690 5690 15710
rect 5710 15690 5720 15710
rect 4720 15680 5720 15690
rect 5760 15710 5960 15720
rect 5760 15690 5770 15710
rect 5790 15690 5850 15710
rect 5870 15690 5930 15710
rect 5950 15690 5960 15710
rect 5760 15680 5960 15690
rect 6000 15710 6200 15720
rect 6000 15690 6010 15710
rect 6030 15690 6090 15710
rect 6110 15690 6170 15710
rect 6190 15690 6200 15710
rect 6000 15680 6200 15690
rect 4240 15630 4440 15640
rect 4240 15610 4250 15630
rect 4270 15610 4330 15630
rect 4350 15610 4410 15630
rect 4430 15610 4440 15630
rect 4240 15600 4440 15610
rect 4480 15630 4680 15640
rect 4480 15610 4490 15630
rect 4510 15610 4570 15630
rect 4590 15610 4650 15630
rect 4670 15610 4680 15630
rect 4480 15600 4680 15610
rect 4720 15630 5720 15640
rect 4720 15610 4730 15630
rect 4750 15610 4810 15630
rect 4830 15610 4890 15630
rect 4910 15610 4970 15630
rect 4990 15610 5050 15630
rect 5070 15610 5130 15630
rect 5150 15610 5210 15630
rect 5230 15610 5290 15630
rect 5310 15610 5370 15630
rect 5390 15610 5450 15630
rect 5470 15610 5530 15630
rect 5550 15610 5610 15630
rect 5630 15610 5690 15630
rect 5710 15610 5720 15630
rect 4720 15600 5720 15610
rect 5760 15630 5960 15640
rect 5760 15610 5770 15630
rect 5790 15610 5850 15630
rect 5870 15610 5930 15630
rect 5950 15610 5960 15630
rect 5760 15600 5960 15610
rect 6000 15630 6200 15640
rect 6000 15610 6010 15630
rect 6030 15610 6090 15630
rect 6110 15610 6170 15630
rect 6190 15610 6200 15630
rect 6000 15600 6200 15610
rect 4240 15550 4440 15560
rect 4240 15530 4250 15550
rect 4270 15530 4330 15550
rect 4350 15530 4410 15550
rect 4430 15530 4440 15550
rect 4240 15520 4440 15530
rect 4480 15550 4680 15560
rect 4480 15530 4490 15550
rect 4510 15530 4570 15550
rect 4590 15530 4650 15550
rect 4670 15530 4680 15550
rect 4480 15520 4680 15530
rect 4720 15550 5720 15560
rect 4720 15530 4730 15550
rect 4750 15530 4810 15550
rect 4830 15530 4890 15550
rect 4910 15530 4970 15550
rect 4990 15530 5050 15550
rect 5070 15530 5130 15550
rect 5150 15530 5210 15550
rect 5230 15530 5290 15550
rect 5310 15530 5370 15550
rect 5390 15530 5450 15550
rect 5470 15530 5530 15550
rect 5550 15530 5610 15550
rect 5630 15530 5690 15550
rect 5710 15530 5720 15550
rect 4720 15520 5720 15530
rect 5760 15550 5960 15560
rect 5760 15530 5770 15550
rect 5790 15530 5850 15550
rect 5870 15530 5930 15550
rect 5950 15530 5960 15550
rect 5760 15520 5960 15530
rect 6000 15550 6200 15560
rect 6000 15530 6010 15550
rect 6030 15530 6090 15550
rect 6110 15530 6170 15550
rect 6190 15530 6200 15550
rect 6000 15520 6200 15530
rect 4240 15470 4440 15480
rect 4240 15450 4250 15470
rect 4270 15450 4330 15470
rect 4350 15450 4410 15470
rect 4430 15450 4440 15470
rect 4240 15440 4440 15450
rect 4480 15470 4680 15480
rect 4480 15450 4490 15470
rect 4510 15450 4570 15470
rect 4590 15450 4650 15470
rect 4670 15450 4680 15470
rect 4480 15440 4680 15450
rect 4720 15470 5720 15480
rect 4720 15450 4730 15470
rect 4750 15450 4810 15470
rect 4830 15450 4890 15470
rect 4910 15450 4970 15470
rect 4990 15450 5050 15470
rect 5070 15450 5130 15470
rect 5150 15450 5210 15470
rect 5230 15450 5290 15470
rect 5310 15450 5370 15470
rect 5390 15450 5450 15470
rect 5470 15450 5530 15470
rect 5550 15450 5610 15470
rect 5630 15450 5690 15470
rect 5710 15450 5720 15470
rect 4720 15440 5720 15450
rect 5760 15470 5960 15480
rect 5760 15450 5770 15470
rect 5790 15450 5850 15470
rect 5870 15450 5930 15470
rect 5950 15450 5960 15470
rect 5760 15440 5960 15450
rect 6000 15470 6200 15480
rect 6000 15450 6010 15470
rect 6030 15450 6090 15470
rect 6110 15450 6170 15470
rect 6190 15450 6200 15470
rect 6000 15440 6200 15450
rect 4240 15390 4440 15400
rect 4240 15370 4250 15390
rect 4270 15370 4330 15390
rect 4350 15370 4410 15390
rect 4430 15370 4440 15390
rect 4240 15360 4440 15370
rect 4480 15390 4680 15400
rect 4480 15370 4490 15390
rect 4510 15370 4570 15390
rect 4590 15370 4650 15390
rect 4670 15370 4680 15390
rect 4480 15360 4680 15370
rect 4720 15390 5720 15400
rect 4720 15370 4730 15390
rect 4750 15370 4810 15390
rect 4830 15370 4890 15390
rect 4910 15370 4970 15390
rect 4990 15370 5050 15390
rect 5070 15370 5130 15390
rect 5150 15370 5210 15390
rect 5230 15370 5290 15390
rect 5310 15370 5370 15390
rect 5390 15370 5450 15390
rect 5470 15370 5530 15390
rect 5550 15370 5610 15390
rect 5630 15370 5690 15390
rect 5710 15370 5720 15390
rect 4720 15360 5720 15370
rect 5760 15390 5960 15400
rect 5760 15370 5770 15390
rect 5790 15370 5850 15390
rect 5870 15370 5930 15390
rect 5950 15370 5960 15390
rect 5760 15360 5960 15370
rect 6000 15390 6200 15400
rect 6000 15370 6010 15390
rect 6030 15370 6090 15390
rect 6110 15370 6170 15390
rect 6190 15370 6200 15390
rect 6000 15360 6200 15370
rect 4240 15310 4440 15320
rect 4240 15290 4250 15310
rect 4270 15290 4330 15310
rect 4350 15290 4410 15310
rect 4430 15290 4440 15310
rect 4240 15280 4440 15290
rect 4480 15310 4680 15320
rect 4480 15290 4490 15310
rect 4510 15290 4570 15310
rect 4590 15290 4650 15310
rect 4670 15290 4680 15310
rect 4480 15280 4680 15290
rect 4720 15310 5720 15320
rect 4720 15290 4730 15310
rect 4750 15290 4810 15310
rect 4830 15290 4890 15310
rect 4910 15290 4970 15310
rect 4990 15290 5050 15310
rect 5070 15290 5130 15310
rect 5150 15290 5210 15310
rect 5230 15290 5290 15310
rect 5310 15290 5370 15310
rect 5390 15290 5450 15310
rect 5470 15290 5530 15310
rect 5550 15290 5610 15310
rect 5630 15290 5690 15310
rect 5710 15290 5720 15310
rect 4720 15280 5720 15290
rect 5760 15310 5960 15320
rect 5760 15290 5770 15310
rect 5790 15290 5850 15310
rect 5870 15290 5930 15310
rect 5950 15290 5960 15310
rect 5760 15280 5960 15290
rect 6000 15310 6200 15320
rect 6000 15290 6010 15310
rect 6030 15290 6090 15310
rect 6110 15290 6170 15310
rect 6190 15290 6200 15310
rect 6000 15280 6200 15290
rect 4240 15230 4440 15240
rect 4240 15210 4250 15230
rect 4270 15210 4330 15230
rect 4350 15210 4410 15230
rect 4430 15210 4440 15230
rect 4240 15200 4440 15210
rect 4480 15230 4680 15240
rect 4480 15210 4490 15230
rect 4510 15210 4570 15230
rect 4590 15210 4650 15230
rect 4670 15210 4680 15230
rect 4480 15200 4680 15210
rect 4720 15230 5720 15240
rect 4720 15210 4730 15230
rect 4750 15210 4810 15230
rect 4830 15210 4890 15230
rect 4910 15210 4970 15230
rect 4990 15210 5050 15230
rect 5070 15210 5130 15230
rect 5150 15210 5210 15230
rect 5230 15210 5290 15230
rect 5310 15210 5370 15230
rect 5390 15210 5450 15230
rect 5470 15210 5530 15230
rect 5550 15210 5610 15230
rect 5630 15210 5690 15230
rect 5710 15210 5720 15230
rect 4720 15200 5720 15210
rect 5760 15230 5960 15240
rect 5760 15210 5770 15230
rect 5790 15210 5850 15230
rect 5870 15210 5930 15230
rect 5950 15210 5960 15230
rect 5760 15200 5960 15210
rect 6000 15230 6200 15240
rect 6000 15210 6010 15230
rect 6030 15210 6090 15230
rect 6110 15210 6170 15230
rect 6190 15210 6200 15230
rect 6000 15200 6200 15210
rect 4240 15150 4440 15160
rect 4240 15130 4250 15150
rect 4270 15130 4330 15150
rect 4350 15130 4410 15150
rect 4430 15130 4440 15150
rect 4240 15120 4440 15130
rect 4480 15150 4680 15160
rect 4480 15130 4490 15150
rect 4510 15130 4570 15150
rect 4590 15130 4650 15150
rect 4670 15130 4680 15150
rect 4480 15120 4680 15130
rect 4720 15150 5720 15160
rect 4720 15130 4730 15150
rect 4750 15130 4810 15150
rect 4830 15130 4890 15150
rect 4910 15130 4970 15150
rect 4990 15130 5050 15150
rect 5070 15130 5130 15150
rect 5150 15130 5210 15150
rect 5230 15130 5290 15150
rect 5310 15130 5370 15150
rect 5390 15130 5450 15150
rect 5470 15130 5530 15150
rect 5550 15130 5610 15150
rect 5630 15130 5690 15150
rect 5710 15130 5720 15150
rect 4720 15120 5720 15130
rect 5760 15150 5960 15160
rect 5760 15130 5770 15150
rect 5790 15130 5850 15150
rect 5870 15130 5930 15150
rect 5950 15130 5960 15150
rect 5760 15120 5960 15130
rect 6000 15150 6200 15160
rect 6000 15130 6010 15150
rect 6030 15130 6090 15150
rect 6110 15130 6170 15150
rect 6190 15130 6200 15150
rect 6000 15120 6200 15130
rect 4240 15070 4440 15080
rect 4240 15050 4250 15070
rect 4270 15050 4330 15070
rect 4350 15050 4410 15070
rect 4430 15050 4440 15070
rect 4240 15040 4440 15050
rect 4480 15070 4680 15080
rect 4480 15050 4490 15070
rect 4510 15050 4570 15070
rect 4590 15050 4650 15070
rect 4670 15050 4680 15070
rect 4480 15040 4680 15050
rect 4720 15070 5720 15080
rect 4720 15050 4730 15070
rect 4750 15050 4810 15070
rect 4830 15050 4890 15070
rect 4910 15050 4970 15070
rect 4990 15050 5050 15070
rect 5070 15050 5130 15070
rect 5150 15050 5210 15070
rect 5230 15050 5290 15070
rect 5310 15050 5370 15070
rect 5390 15050 5450 15070
rect 5470 15050 5530 15070
rect 5550 15050 5610 15070
rect 5630 15050 5690 15070
rect 5710 15050 5720 15070
rect 4720 15040 5720 15050
rect 5760 15070 5960 15080
rect 5760 15050 5770 15070
rect 5790 15050 5850 15070
rect 5870 15050 5930 15070
rect 5950 15050 5960 15070
rect 5760 15040 5960 15050
rect 6000 15070 6200 15080
rect 6000 15050 6010 15070
rect 6030 15050 6090 15070
rect 6110 15050 6170 15070
rect 6190 15050 6200 15070
rect 6000 15040 6200 15050
rect 4240 14990 4440 15000
rect 4240 14970 4250 14990
rect 4270 14970 4330 14990
rect 4350 14970 4410 14990
rect 4430 14970 4440 14990
rect 4240 14960 4440 14970
rect 4480 14990 4680 15000
rect 4480 14970 4490 14990
rect 4510 14970 4570 14990
rect 4590 14970 4650 14990
rect 4670 14970 4680 14990
rect 4480 14960 4680 14970
rect 4720 14990 5720 15000
rect 4720 14970 4730 14990
rect 4750 14970 4810 14990
rect 4830 14970 4890 14990
rect 4910 14970 4970 14990
rect 4990 14970 5050 14990
rect 5070 14970 5130 14990
rect 5150 14970 5210 14990
rect 5230 14970 5290 14990
rect 5310 14970 5370 14990
rect 5390 14970 5450 14990
rect 5470 14970 5530 14990
rect 5550 14970 5610 14990
rect 5630 14970 5690 14990
rect 5710 14970 5720 14990
rect 4720 14960 5720 14970
rect 5760 14990 5960 15000
rect 5760 14970 5770 14990
rect 5790 14970 5850 14990
rect 5870 14970 5930 14990
rect 5950 14970 5960 14990
rect 5760 14960 5960 14970
rect 6000 14990 6200 15000
rect 6000 14970 6010 14990
rect 6030 14970 6090 14990
rect 6110 14970 6170 14990
rect 6190 14970 6200 14990
rect 6000 14960 6200 14970
rect 4240 14910 4440 14920
rect 4240 14890 4250 14910
rect 4270 14890 4330 14910
rect 4350 14890 4410 14910
rect 4430 14890 4440 14910
rect 4240 14880 4440 14890
rect 4480 14910 4680 14920
rect 4480 14890 4490 14910
rect 4510 14890 4570 14910
rect 4590 14890 4650 14910
rect 4670 14890 4680 14910
rect 4480 14880 4680 14890
rect 4720 14910 5720 14920
rect 4720 14890 4730 14910
rect 4750 14890 4810 14910
rect 4830 14890 4890 14910
rect 4910 14890 4970 14910
rect 4990 14890 5050 14910
rect 5070 14890 5130 14910
rect 5150 14890 5210 14910
rect 5230 14890 5290 14910
rect 5310 14890 5370 14910
rect 5390 14890 5450 14910
rect 5470 14890 5530 14910
rect 5550 14890 5610 14910
rect 5630 14890 5690 14910
rect 5710 14890 5720 14910
rect 4720 14880 5720 14890
rect 5760 14910 5960 14920
rect 5760 14890 5770 14910
rect 5790 14890 5850 14910
rect 5870 14890 5930 14910
rect 5950 14890 5960 14910
rect 5760 14880 5960 14890
rect 6000 14910 6200 14920
rect 6000 14890 6010 14910
rect 6030 14890 6090 14910
rect 6110 14890 6170 14910
rect 6190 14890 6200 14910
rect 6000 14880 6200 14890
rect 4240 14830 4440 14840
rect 4240 14810 4250 14830
rect 4270 14810 4330 14830
rect 4350 14810 4410 14830
rect 4430 14810 4440 14830
rect 4240 14800 4440 14810
rect 4480 14830 4680 14840
rect 4480 14810 4490 14830
rect 4510 14810 4570 14830
rect 4590 14810 4650 14830
rect 4670 14810 4680 14830
rect 4480 14800 4680 14810
rect 4720 14830 5720 14840
rect 4720 14810 4730 14830
rect 4750 14810 4810 14830
rect 4830 14810 4890 14830
rect 4910 14810 4970 14830
rect 4990 14810 5050 14830
rect 5070 14810 5130 14830
rect 5150 14810 5210 14830
rect 5230 14810 5290 14830
rect 5310 14810 5370 14830
rect 5390 14810 5450 14830
rect 5470 14810 5530 14830
rect 5550 14810 5610 14830
rect 5630 14810 5690 14830
rect 5710 14810 5720 14830
rect 4720 14800 5720 14810
rect 5760 14830 5960 14840
rect 5760 14810 5770 14830
rect 5790 14810 5850 14830
rect 5870 14810 5930 14830
rect 5950 14810 5960 14830
rect 5760 14800 5960 14810
rect 6000 14830 6200 14840
rect 6000 14810 6010 14830
rect 6030 14810 6090 14830
rect 6110 14810 6170 14830
rect 6190 14810 6200 14830
rect 6000 14800 6200 14810
rect 4240 14750 4440 14760
rect 4240 14730 4250 14750
rect 4270 14730 4330 14750
rect 4350 14730 4410 14750
rect 4430 14730 4440 14750
rect 4240 14720 4440 14730
rect 4480 14750 4680 14760
rect 4480 14730 4490 14750
rect 4510 14730 4570 14750
rect 4590 14730 4650 14750
rect 4670 14730 4680 14750
rect 4480 14720 4680 14730
rect 4720 14750 5720 14760
rect 4720 14730 4730 14750
rect 4750 14730 4810 14750
rect 4830 14730 4890 14750
rect 4910 14730 4970 14750
rect 4990 14730 5050 14750
rect 5070 14730 5130 14750
rect 5150 14730 5210 14750
rect 5230 14730 5290 14750
rect 5310 14730 5370 14750
rect 5390 14730 5450 14750
rect 5470 14730 5530 14750
rect 5550 14730 5610 14750
rect 5630 14730 5690 14750
rect 5710 14730 5720 14750
rect 4720 14720 5720 14730
rect 5760 14750 5960 14760
rect 5760 14730 5770 14750
rect 5790 14730 5850 14750
rect 5870 14730 5930 14750
rect 5950 14730 5960 14750
rect 5760 14720 5960 14730
rect 6000 14750 6200 14760
rect 6000 14730 6010 14750
rect 6030 14730 6090 14750
rect 6110 14730 6170 14750
rect 6190 14730 6200 14750
rect 6000 14720 6200 14730
rect 4240 14670 4440 14680
rect 4240 14650 4250 14670
rect 4270 14650 4330 14670
rect 4350 14650 4410 14670
rect 4430 14650 4440 14670
rect 4240 14640 4440 14650
rect 4480 14670 4680 14680
rect 4480 14650 4490 14670
rect 4510 14650 4570 14670
rect 4590 14650 4650 14670
rect 4670 14650 4680 14670
rect 4480 14640 4680 14650
rect 4720 14670 5720 14680
rect 4720 14650 4730 14670
rect 4750 14650 4810 14670
rect 4830 14650 4890 14670
rect 4910 14650 4970 14670
rect 4990 14650 5050 14670
rect 5070 14650 5130 14670
rect 5150 14650 5210 14670
rect 5230 14650 5290 14670
rect 5310 14650 5370 14670
rect 5390 14650 5450 14670
rect 5470 14650 5530 14670
rect 5550 14650 5610 14670
rect 5630 14650 5690 14670
rect 5710 14650 5720 14670
rect 4720 14640 5720 14650
rect 5760 14670 5960 14680
rect 5760 14650 5770 14670
rect 5790 14650 5850 14670
rect 5870 14650 5930 14670
rect 5950 14650 5960 14670
rect 5760 14640 5960 14650
rect 6000 14670 6200 14680
rect 6000 14650 6010 14670
rect 6030 14650 6090 14670
rect 6110 14650 6170 14670
rect 6190 14650 6200 14670
rect 6000 14640 6200 14650
rect 4240 14590 4440 14600
rect 4240 14570 4250 14590
rect 4270 14570 4330 14590
rect 4350 14570 4410 14590
rect 4430 14570 4440 14590
rect 4240 14560 4440 14570
rect 4480 14590 4680 14600
rect 4480 14570 4490 14590
rect 4510 14570 4570 14590
rect 4590 14570 4650 14590
rect 4670 14570 4680 14590
rect 4480 14560 4680 14570
rect 4720 14590 5720 14600
rect 4720 14570 4730 14590
rect 4750 14570 4810 14590
rect 4830 14570 4890 14590
rect 4910 14570 4970 14590
rect 4990 14570 5050 14590
rect 5070 14570 5130 14590
rect 5150 14570 5210 14590
rect 5230 14570 5290 14590
rect 5310 14570 5370 14590
rect 5390 14570 5450 14590
rect 5470 14570 5530 14590
rect 5550 14570 5610 14590
rect 5630 14570 5690 14590
rect 5710 14570 5720 14590
rect 4720 14560 5720 14570
rect 5760 14590 5960 14600
rect 5760 14570 5770 14590
rect 5790 14570 5850 14590
rect 5870 14570 5930 14590
rect 5950 14570 5960 14590
rect 5760 14560 5960 14570
rect 6000 14590 6200 14600
rect 6000 14570 6010 14590
rect 6030 14570 6090 14590
rect 6110 14570 6170 14590
rect 6190 14570 6200 14590
rect 6000 14560 6200 14570
rect 4240 14510 4440 14520
rect 4240 14490 4250 14510
rect 4270 14490 4330 14510
rect 4350 14490 4410 14510
rect 4430 14490 4440 14510
rect 4240 14480 4440 14490
rect 4480 14510 4680 14520
rect 4480 14490 4490 14510
rect 4510 14490 4570 14510
rect 4590 14490 4650 14510
rect 4670 14490 4680 14510
rect 4480 14480 4680 14490
rect 4720 14510 5720 14520
rect 4720 14490 4730 14510
rect 4750 14490 4810 14510
rect 4830 14490 4890 14510
rect 4910 14490 4970 14510
rect 4990 14490 5050 14510
rect 5070 14490 5130 14510
rect 5150 14490 5210 14510
rect 5230 14490 5290 14510
rect 5310 14490 5370 14510
rect 5390 14490 5450 14510
rect 5470 14490 5530 14510
rect 5550 14490 5610 14510
rect 5630 14490 5690 14510
rect 5710 14490 5720 14510
rect 4720 14480 5720 14490
rect 5760 14510 5960 14520
rect 5760 14490 5770 14510
rect 5790 14490 5850 14510
rect 5870 14490 5930 14510
rect 5950 14490 5960 14510
rect 5760 14480 5960 14490
rect 6000 14510 6200 14520
rect 6000 14490 6010 14510
rect 6030 14490 6090 14510
rect 6110 14490 6170 14510
rect 6190 14490 6200 14510
rect 6000 14480 6200 14490
rect 4240 14430 4440 14440
rect 4240 14410 4250 14430
rect 4270 14410 4330 14430
rect 4350 14410 4410 14430
rect 4430 14410 4440 14430
rect 4240 14400 4440 14410
rect 4480 14430 4680 14440
rect 4480 14410 4490 14430
rect 4510 14410 4570 14430
rect 4590 14410 4650 14430
rect 4670 14410 4680 14430
rect 4480 14400 4680 14410
rect 4720 14430 5720 14440
rect 4720 14410 4730 14430
rect 4750 14410 4810 14430
rect 4830 14410 4890 14430
rect 4910 14410 4970 14430
rect 4990 14410 5050 14430
rect 5070 14410 5130 14430
rect 5150 14410 5210 14430
rect 5230 14410 5290 14430
rect 5310 14410 5370 14430
rect 5390 14410 5450 14430
rect 5470 14410 5530 14430
rect 5550 14410 5610 14430
rect 5630 14410 5690 14430
rect 5710 14410 5720 14430
rect 4720 14400 5720 14410
rect 5760 14430 5960 14440
rect 5760 14410 5770 14430
rect 5790 14410 5850 14430
rect 5870 14410 5930 14430
rect 5950 14410 5960 14430
rect 5760 14400 5960 14410
rect 6000 14430 6200 14440
rect 6000 14410 6010 14430
rect 6030 14410 6090 14430
rect 6110 14410 6170 14430
rect 6190 14410 6200 14430
rect 6000 14400 6200 14410
rect 4240 14350 4440 14360
rect 4240 14330 4250 14350
rect 4270 14330 4330 14350
rect 4350 14330 4410 14350
rect 4430 14330 4440 14350
rect 4240 14320 4440 14330
rect 4480 14350 4680 14360
rect 4480 14330 4490 14350
rect 4510 14330 4570 14350
rect 4590 14330 4650 14350
rect 4670 14330 4680 14350
rect 4480 14320 4680 14330
rect 4720 14350 5720 14360
rect 4720 14330 4730 14350
rect 4750 14330 4810 14350
rect 4830 14330 4890 14350
rect 4910 14330 4970 14350
rect 4990 14330 5050 14350
rect 5070 14330 5130 14350
rect 5150 14330 5210 14350
rect 5230 14330 5290 14350
rect 5310 14330 5370 14350
rect 5390 14330 5450 14350
rect 5470 14330 5530 14350
rect 5550 14330 5610 14350
rect 5630 14330 5690 14350
rect 5710 14330 5720 14350
rect 4720 14320 5720 14330
rect 5760 14350 5960 14360
rect 5760 14330 5770 14350
rect 5790 14330 5850 14350
rect 5870 14330 5930 14350
rect 5950 14330 5960 14350
rect 5760 14320 5960 14330
rect 6000 14350 6200 14360
rect 6000 14330 6010 14350
rect 6030 14330 6090 14350
rect 6110 14330 6170 14350
rect 6190 14330 6200 14350
rect 6000 14320 6200 14330
rect 4240 14270 4440 14280
rect 4240 14250 4250 14270
rect 4270 14250 4330 14270
rect 4350 14250 4410 14270
rect 4430 14250 4440 14270
rect 4240 14240 4440 14250
rect 4480 14270 4680 14280
rect 4480 14250 4490 14270
rect 4510 14250 4570 14270
rect 4590 14250 4650 14270
rect 4670 14250 4680 14270
rect 4480 14240 4680 14250
rect 4720 14270 5720 14280
rect 4720 14250 4730 14270
rect 4750 14250 4810 14270
rect 4830 14250 4890 14270
rect 4910 14250 4970 14270
rect 4990 14250 5050 14270
rect 5070 14250 5130 14270
rect 5150 14250 5210 14270
rect 5230 14250 5290 14270
rect 5310 14250 5370 14270
rect 5390 14250 5450 14270
rect 5470 14250 5530 14270
rect 5550 14250 5610 14270
rect 5630 14250 5690 14270
rect 5710 14250 5720 14270
rect 4720 14240 5720 14250
rect 5760 14270 5960 14280
rect 5760 14250 5770 14270
rect 5790 14250 5850 14270
rect 5870 14250 5930 14270
rect 5950 14250 5960 14270
rect 5760 14240 5960 14250
rect 6000 14270 6200 14280
rect 6000 14250 6010 14270
rect 6030 14250 6090 14270
rect 6110 14250 6170 14270
rect 6190 14250 6200 14270
rect 6000 14240 6200 14250
rect 4240 14190 4440 14200
rect 4240 14170 4250 14190
rect 4270 14170 4330 14190
rect 4350 14170 4410 14190
rect 4430 14170 4440 14190
rect 4240 14160 4440 14170
rect 4480 14190 4680 14200
rect 4480 14170 4490 14190
rect 4510 14170 4570 14190
rect 4590 14170 4650 14190
rect 4670 14170 4680 14190
rect 4480 14160 4680 14170
rect 4720 14190 5720 14200
rect 4720 14170 4730 14190
rect 4750 14170 4810 14190
rect 4830 14170 4890 14190
rect 4910 14170 4970 14190
rect 4990 14170 5050 14190
rect 5070 14170 5130 14190
rect 5150 14170 5210 14190
rect 5230 14170 5290 14190
rect 5310 14170 5370 14190
rect 5390 14170 5450 14190
rect 5470 14170 5530 14190
rect 5550 14170 5610 14190
rect 5630 14170 5690 14190
rect 5710 14170 5720 14190
rect 4720 14160 5720 14170
rect 5760 14190 5960 14200
rect 5760 14170 5770 14190
rect 5790 14170 5850 14190
rect 5870 14170 5930 14190
rect 5950 14170 5960 14190
rect 5760 14160 5960 14170
rect 6000 14190 6200 14200
rect 6000 14170 6010 14190
rect 6030 14170 6090 14190
rect 6110 14170 6170 14190
rect 6190 14170 6200 14190
rect 6000 14160 6200 14170
rect 4240 14110 4440 14120
rect 4240 14090 4250 14110
rect 4270 14090 4330 14110
rect 4350 14090 4410 14110
rect 4430 14090 4440 14110
rect 4240 14080 4440 14090
rect 4480 14110 4680 14120
rect 4480 14090 4490 14110
rect 4510 14090 4570 14110
rect 4590 14090 4650 14110
rect 4670 14090 4680 14110
rect 4480 14080 4680 14090
rect 4720 14110 5720 14120
rect 4720 14090 4730 14110
rect 4750 14090 4810 14110
rect 4830 14090 4890 14110
rect 4910 14090 4970 14110
rect 4990 14090 5050 14110
rect 5070 14090 5130 14110
rect 5150 14090 5210 14110
rect 5230 14090 5290 14110
rect 5310 14090 5370 14110
rect 5390 14090 5450 14110
rect 5470 14090 5530 14110
rect 5550 14090 5610 14110
rect 5630 14090 5690 14110
rect 5710 14090 5720 14110
rect 4720 14080 5720 14090
rect 5760 14110 5960 14120
rect 5760 14090 5770 14110
rect 5790 14090 5850 14110
rect 5870 14090 5930 14110
rect 5950 14090 5960 14110
rect 5760 14080 5960 14090
rect 6000 14110 6200 14120
rect 6000 14090 6010 14110
rect 6030 14090 6090 14110
rect 6110 14090 6170 14110
rect 6190 14090 6200 14110
rect 6000 14080 6200 14090
rect 4240 14030 4440 14040
rect 4240 14010 4250 14030
rect 4270 14010 4330 14030
rect 4350 14010 4410 14030
rect 4430 14010 4440 14030
rect 4240 14000 4440 14010
rect 4480 14030 4680 14040
rect 4480 14010 4490 14030
rect 4510 14010 4570 14030
rect 4590 14010 4650 14030
rect 4670 14010 4680 14030
rect 4480 14000 4680 14010
rect 4720 14030 5720 14040
rect 4720 14010 4730 14030
rect 4750 14010 4810 14030
rect 4830 14010 4890 14030
rect 4910 14010 4970 14030
rect 4990 14010 5050 14030
rect 5070 14010 5130 14030
rect 5150 14010 5210 14030
rect 5230 14010 5290 14030
rect 5310 14010 5370 14030
rect 5390 14010 5450 14030
rect 5470 14010 5530 14030
rect 5550 14010 5610 14030
rect 5630 14010 5690 14030
rect 5710 14010 5720 14030
rect 4720 14000 5720 14010
rect 5760 14030 5960 14040
rect 5760 14010 5770 14030
rect 5790 14010 5850 14030
rect 5870 14010 5930 14030
rect 5950 14010 5960 14030
rect 5760 14000 5960 14010
rect 6000 14030 6200 14040
rect 6000 14010 6010 14030
rect 6030 14010 6090 14030
rect 6110 14010 6170 14030
rect 6190 14010 6200 14030
rect 6000 14000 6200 14010
rect 4240 13950 4440 13960
rect 4240 13930 4250 13950
rect 4270 13930 4330 13950
rect 4350 13930 4410 13950
rect 4430 13930 4440 13950
rect 4240 13920 4440 13930
rect 4480 13950 4680 13960
rect 4480 13930 4490 13950
rect 4510 13930 4570 13950
rect 4590 13930 4650 13950
rect 4670 13930 4680 13950
rect 4480 13920 4680 13930
rect 4720 13950 5720 13960
rect 4720 13930 4730 13950
rect 4750 13930 4810 13950
rect 4830 13930 4890 13950
rect 4910 13930 4970 13950
rect 4990 13930 5050 13950
rect 5070 13930 5130 13950
rect 5150 13930 5210 13950
rect 5230 13930 5290 13950
rect 5310 13930 5370 13950
rect 5390 13930 5450 13950
rect 5470 13930 5530 13950
rect 5550 13930 5610 13950
rect 5630 13930 5690 13950
rect 5710 13930 5720 13950
rect 4720 13920 5720 13930
rect 5760 13950 5960 13960
rect 5760 13930 5770 13950
rect 5790 13930 5850 13950
rect 5870 13930 5930 13950
rect 5950 13930 5960 13950
rect 5760 13920 5960 13930
rect 6000 13950 6200 13960
rect 6000 13930 6010 13950
rect 6030 13930 6090 13950
rect 6110 13930 6170 13950
rect 6190 13930 6200 13950
rect 6000 13920 6200 13930
rect 4240 13870 4440 13880
rect 4240 13850 4250 13870
rect 4270 13850 4330 13870
rect 4350 13850 4410 13870
rect 4430 13850 4440 13870
rect 4240 13840 4440 13850
rect 4480 13870 4680 13880
rect 4480 13850 4490 13870
rect 4510 13850 4570 13870
rect 4590 13850 4650 13870
rect 4670 13850 4680 13870
rect 4480 13840 4680 13850
rect 4720 13870 5720 13880
rect 4720 13850 4730 13870
rect 4750 13850 4810 13870
rect 4830 13850 4890 13870
rect 4910 13850 4970 13870
rect 4990 13850 5050 13870
rect 5070 13850 5130 13870
rect 5150 13850 5210 13870
rect 5230 13850 5290 13870
rect 5310 13850 5370 13870
rect 5390 13850 5450 13870
rect 5470 13850 5530 13870
rect 5550 13850 5610 13870
rect 5630 13850 5690 13870
rect 5710 13850 5720 13870
rect 4720 13840 5720 13850
rect 5760 13870 5960 13880
rect 5760 13850 5770 13870
rect 5790 13850 5850 13870
rect 5870 13850 5930 13870
rect 5950 13850 5960 13870
rect 5760 13840 5960 13850
rect 6000 13870 6200 13880
rect 6000 13850 6010 13870
rect 6030 13850 6090 13870
rect 6110 13850 6170 13870
rect 6190 13850 6200 13870
rect 6000 13840 6200 13850
rect 4240 13790 4440 13800
rect 4240 13770 4250 13790
rect 4270 13770 4330 13790
rect 4350 13770 4410 13790
rect 4430 13770 4440 13790
rect 4240 13760 4440 13770
rect 4480 13790 4680 13800
rect 4480 13770 4490 13790
rect 4510 13770 4570 13790
rect 4590 13770 4650 13790
rect 4670 13770 4680 13790
rect 4480 13760 4680 13770
rect 4720 13790 5720 13800
rect 4720 13770 4730 13790
rect 4750 13770 4810 13790
rect 4830 13770 4890 13790
rect 4910 13770 4970 13790
rect 4990 13770 5050 13790
rect 5070 13770 5130 13790
rect 5150 13770 5210 13790
rect 5230 13770 5290 13790
rect 5310 13770 5370 13790
rect 5390 13770 5450 13790
rect 5470 13770 5530 13790
rect 5550 13770 5610 13790
rect 5630 13770 5690 13790
rect 5710 13770 5720 13790
rect 4720 13760 5720 13770
rect 5760 13790 5960 13800
rect 5760 13770 5770 13790
rect 5790 13770 5850 13790
rect 5870 13770 5930 13790
rect 5950 13770 5960 13790
rect 5760 13760 5960 13770
rect 6000 13790 6200 13800
rect 6000 13770 6010 13790
rect 6030 13770 6090 13790
rect 6110 13770 6170 13790
rect 6190 13770 6200 13790
rect 6000 13760 6200 13770
rect 4240 13710 4440 13720
rect 4240 13690 4250 13710
rect 4270 13690 4330 13710
rect 4350 13690 4410 13710
rect 4430 13690 4440 13710
rect 4240 13680 4440 13690
rect 4480 13710 4680 13720
rect 4480 13690 4490 13710
rect 4510 13690 4570 13710
rect 4590 13690 4650 13710
rect 4670 13690 4680 13710
rect 4480 13680 4680 13690
rect 4720 13710 5720 13720
rect 4720 13690 4730 13710
rect 4750 13690 4810 13710
rect 4830 13690 4890 13710
rect 4910 13690 4970 13710
rect 4990 13690 5050 13710
rect 5070 13690 5130 13710
rect 5150 13690 5210 13710
rect 5230 13690 5290 13710
rect 5310 13690 5370 13710
rect 5390 13690 5450 13710
rect 5470 13690 5530 13710
rect 5550 13690 5610 13710
rect 5630 13690 5690 13710
rect 5710 13690 5720 13710
rect 4720 13680 5720 13690
rect 5760 13710 5960 13720
rect 5760 13690 5770 13710
rect 5790 13690 5850 13710
rect 5870 13690 5930 13710
rect 5950 13690 5960 13710
rect 5760 13680 5960 13690
rect 6000 13710 6200 13720
rect 6000 13690 6010 13710
rect 6030 13690 6090 13710
rect 6110 13690 6170 13710
rect 6190 13690 6200 13710
rect 6000 13680 6200 13690
rect 4240 13630 4440 13640
rect 4240 13610 4250 13630
rect 4270 13610 4330 13630
rect 4350 13610 4410 13630
rect 4430 13610 4440 13630
rect 4240 13600 4440 13610
rect 4480 13630 4680 13640
rect 4480 13610 4490 13630
rect 4510 13610 4570 13630
rect 4590 13610 4650 13630
rect 4670 13610 4680 13630
rect 4480 13600 4680 13610
rect 4720 13630 5720 13640
rect 4720 13610 4730 13630
rect 4750 13610 4810 13630
rect 4830 13610 4890 13630
rect 4910 13610 4970 13630
rect 4990 13610 5050 13630
rect 5070 13610 5130 13630
rect 5150 13610 5210 13630
rect 5230 13610 5290 13630
rect 5310 13610 5370 13630
rect 5390 13610 5450 13630
rect 5470 13610 5530 13630
rect 5550 13610 5610 13630
rect 5630 13610 5690 13630
rect 5710 13610 5720 13630
rect 4720 13600 5720 13610
rect 5760 13630 5960 13640
rect 5760 13610 5770 13630
rect 5790 13610 5850 13630
rect 5870 13610 5930 13630
rect 5950 13610 5960 13630
rect 5760 13600 5960 13610
rect 6000 13630 6200 13640
rect 6000 13610 6010 13630
rect 6030 13610 6090 13630
rect 6110 13610 6170 13630
rect 6190 13610 6200 13630
rect 6000 13600 6200 13610
rect 4240 13550 4440 13560
rect 4240 13530 4250 13550
rect 4270 13530 4330 13550
rect 4350 13530 4410 13550
rect 4430 13530 4440 13550
rect 4240 13520 4440 13530
rect 4480 13550 4680 13560
rect 4480 13530 4490 13550
rect 4510 13530 4570 13550
rect 4590 13530 4650 13550
rect 4670 13530 4680 13550
rect 4480 13520 4680 13530
rect 4720 13550 5720 13560
rect 4720 13530 4730 13550
rect 4750 13530 4810 13550
rect 4830 13530 4890 13550
rect 4910 13530 4970 13550
rect 4990 13530 5050 13550
rect 5070 13530 5130 13550
rect 5150 13530 5210 13550
rect 5230 13530 5290 13550
rect 5310 13530 5370 13550
rect 5390 13530 5450 13550
rect 5470 13530 5530 13550
rect 5550 13530 5610 13550
rect 5630 13530 5690 13550
rect 5710 13530 5720 13550
rect 4720 13520 5720 13530
rect 5760 13550 5960 13560
rect 5760 13530 5770 13550
rect 5790 13530 5850 13550
rect 5870 13530 5930 13550
rect 5950 13530 5960 13550
rect 5760 13520 5960 13530
rect 6000 13550 6200 13560
rect 6000 13530 6010 13550
rect 6030 13530 6090 13550
rect 6110 13530 6170 13550
rect 6190 13530 6200 13550
rect 6000 13520 6200 13530
rect 4240 13470 4440 13480
rect 4240 13450 4250 13470
rect 4270 13450 4330 13470
rect 4350 13450 4410 13470
rect 4430 13450 4440 13470
rect 4240 13440 4440 13450
rect 4480 13470 4680 13480
rect 4480 13450 4490 13470
rect 4510 13450 4570 13470
rect 4590 13450 4650 13470
rect 4670 13450 4680 13470
rect 4480 13440 4680 13450
rect 4720 13470 5720 13480
rect 4720 13450 4730 13470
rect 4750 13450 4810 13470
rect 4830 13450 4890 13470
rect 4910 13450 4970 13470
rect 4990 13450 5050 13470
rect 5070 13450 5130 13470
rect 5150 13450 5210 13470
rect 5230 13450 5290 13470
rect 5310 13450 5370 13470
rect 5390 13450 5450 13470
rect 5470 13450 5530 13470
rect 5550 13450 5610 13470
rect 5630 13450 5690 13470
rect 5710 13450 5720 13470
rect 4720 13440 5720 13450
rect 5760 13470 5960 13480
rect 5760 13450 5770 13470
rect 5790 13450 5850 13470
rect 5870 13450 5930 13470
rect 5950 13450 5960 13470
rect 5760 13440 5960 13450
rect 6000 13470 6200 13480
rect 6000 13450 6010 13470
rect 6030 13450 6090 13470
rect 6110 13450 6170 13470
rect 6190 13450 6200 13470
rect 6000 13440 6200 13450
rect 4240 13390 4440 13400
rect 4240 13370 4250 13390
rect 4270 13370 4330 13390
rect 4350 13370 4410 13390
rect 4430 13370 4440 13390
rect 4240 13360 4440 13370
rect 4480 13390 4680 13400
rect 4480 13370 4490 13390
rect 4510 13370 4570 13390
rect 4590 13370 4650 13390
rect 4670 13370 4680 13390
rect 4480 13360 4680 13370
rect 4720 13390 5720 13400
rect 4720 13370 4730 13390
rect 4750 13370 4810 13390
rect 4830 13370 4890 13390
rect 4910 13370 4970 13390
rect 4990 13370 5050 13390
rect 5070 13370 5130 13390
rect 5150 13370 5210 13390
rect 5230 13370 5290 13390
rect 5310 13370 5370 13390
rect 5390 13370 5450 13390
rect 5470 13370 5530 13390
rect 5550 13370 5610 13390
rect 5630 13370 5690 13390
rect 5710 13370 5720 13390
rect 4720 13360 5720 13370
rect 5760 13390 5960 13400
rect 5760 13370 5770 13390
rect 5790 13370 5850 13390
rect 5870 13370 5930 13390
rect 5950 13370 5960 13390
rect 5760 13360 5960 13370
rect 6000 13390 6200 13400
rect 6000 13370 6010 13390
rect 6030 13370 6090 13390
rect 6110 13370 6170 13390
rect 6190 13370 6200 13390
rect 6000 13360 6200 13370
rect 4240 13310 4440 13320
rect 4240 13290 4250 13310
rect 4270 13290 4330 13310
rect 4350 13290 4410 13310
rect 4430 13290 4440 13310
rect 4240 13280 4440 13290
rect 4480 13310 4680 13320
rect 4480 13290 4490 13310
rect 4510 13290 4570 13310
rect 4590 13290 4650 13310
rect 4670 13290 4680 13310
rect 4480 13280 4680 13290
rect 4720 13310 5720 13320
rect 4720 13290 4730 13310
rect 4750 13290 4810 13310
rect 4830 13290 4890 13310
rect 4910 13290 4970 13310
rect 4990 13290 5050 13310
rect 5070 13290 5130 13310
rect 5150 13290 5210 13310
rect 5230 13290 5290 13310
rect 5310 13290 5370 13310
rect 5390 13290 5450 13310
rect 5470 13290 5530 13310
rect 5550 13290 5610 13310
rect 5630 13290 5690 13310
rect 5710 13290 5720 13310
rect 4720 13280 5720 13290
rect 5760 13310 5960 13320
rect 5760 13290 5770 13310
rect 5790 13290 5850 13310
rect 5870 13290 5930 13310
rect 5950 13290 5960 13310
rect 5760 13280 5960 13290
rect 6000 13310 6200 13320
rect 6000 13290 6010 13310
rect 6030 13290 6090 13310
rect 6110 13290 6170 13310
rect 6190 13290 6200 13310
rect 6000 13280 6200 13290
rect 4240 13230 4440 13240
rect 4240 13210 4250 13230
rect 4270 13210 4330 13230
rect 4350 13210 4410 13230
rect 4430 13210 4440 13230
rect 4240 13200 4440 13210
rect 4480 13230 4680 13240
rect 4480 13210 4490 13230
rect 4510 13210 4570 13230
rect 4590 13210 4650 13230
rect 4670 13210 4680 13230
rect 4480 13200 4680 13210
rect 4720 13230 5720 13240
rect 4720 13210 4730 13230
rect 4750 13210 4810 13230
rect 4830 13210 4890 13230
rect 4910 13210 4970 13230
rect 4990 13210 5050 13230
rect 5070 13210 5130 13230
rect 5150 13210 5210 13230
rect 5230 13210 5290 13230
rect 5310 13210 5370 13230
rect 5390 13210 5450 13230
rect 5470 13210 5530 13230
rect 5550 13210 5610 13230
rect 5630 13210 5690 13230
rect 5710 13210 5720 13230
rect 4720 13200 5720 13210
rect 5760 13230 5960 13240
rect 5760 13210 5770 13230
rect 5790 13210 5850 13230
rect 5870 13210 5930 13230
rect 5950 13210 5960 13230
rect 5760 13200 5960 13210
rect 6000 13230 6200 13240
rect 6000 13210 6010 13230
rect 6030 13210 6090 13230
rect 6110 13210 6170 13230
rect 6190 13210 6200 13230
rect 6000 13200 6200 13210
rect 4240 13150 4440 13160
rect 4240 13130 4250 13150
rect 4270 13130 4330 13150
rect 4350 13130 4410 13150
rect 4430 13130 4440 13150
rect 4240 13120 4440 13130
rect 4480 13150 4680 13160
rect 4480 13130 4490 13150
rect 4510 13130 4570 13150
rect 4590 13130 4650 13150
rect 4670 13130 4680 13150
rect 4480 13120 4680 13130
rect 4720 13150 5720 13160
rect 4720 13130 4730 13150
rect 4750 13130 4810 13150
rect 4830 13130 4890 13150
rect 4910 13130 4970 13150
rect 4990 13130 5050 13150
rect 5070 13130 5130 13150
rect 5150 13130 5210 13150
rect 5230 13130 5290 13150
rect 5310 13130 5370 13150
rect 5390 13130 5450 13150
rect 5470 13130 5530 13150
rect 5550 13130 5610 13150
rect 5630 13130 5690 13150
rect 5710 13130 5720 13150
rect 4720 13120 5720 13130
rect 5760 13150 5960 13160
rect 5760 13130 5770 13150
rect 5790 13130 5850 13150
rect 5870 13130 5930 13150
rect 5950 13130 5960 13150
rect 5760 13120 5960 13130
rect 6000 13150 6200 13160
rect 6000 13130 6010 13150
rect 6030 13130 6090 13150
rect 6110 13130 6170 13150
rect 6190 13130 6200 13150
rect 6000 13120 6200 13130
rect 4240 13070 4440 13080
rect 4240 13050 4250 13070
rect 4270 13050 4330 13070
rect 4350 13050 4410 13070
rect 4430 13050 4440 13070
rect 4240 13040 4440 13050
rect 4480 13070 4680 13080
rect 4480 13050 4490 13070
rect 4510 13050 4570 13070
rect 4590 13050 4650 13070
rect 4670 13050 4680 13070
rect 4480 13040 4680 13050
rect 4720 13070 5720 13080
rect 4720 13050 4730 13070
rect 4750 13050 4810 13070
rect 4830 13050 4890 13070
rect 4910 13050 4970 13070
rect 4990 13050 5050 13070
rect 5070 13050 5130 13070
rect 5150 13050 5210 13070
rect 5230 13050 5290 13070
rect 5310 13050 5370 13070
rect 5390 13050 5450 13070
rect 5470 13050 5530 13070
rect 5550 13050 5610 13070
rect 5630 13050 5690 13070
rect 5710 13050 5720 13070
rect 4720 13040 5720 13050
rect 5760 13070 5960 13080
rect 5760 13050 5770 13070
rect 5790 13050 5850 13070
rect 5870 13050 5930 13070
rect 5950 13050 5960 13070
rect 5760 13040 5960 13050
rect 6000 13070 6200 13080
rect 6000 13050 6010 13070
rect 6030 13050 6090 13070
rect 6110 13050 6170 13070
rect 6190 13050 6200 13070
rect 6000 13040 6200 13050
rect 4240 12990 4440 13000
rect 4240 12970 4250 12990
rect 4270 12970 4330 12990
rect 4350 12970 4410 12990
rect 4430 12970 4440 12990
rect 4240 12960 4440 12970
rect 4480 12990 4680 13000
rect 4480 12970 4490 12990
rect 4510 12970 4570 12990
rect 4590 12970 4650 12990
rect 4670 12970 4680 12990
rect 4480 12960 4680 12970
rect 4720 12990 5720 13000
rect 4720 12970 4730 12990
rect 4750 12970 4810 12990
rect 4830 12970 4890 12990
rect 4910 12970 4970 12990
rect 4990 12970 5050 12990
rect 5070 12970 5130 12990
rect 5150 12970 5210 12990
rect 5230 12970 5290 12990
rect 5310 12970 5370 12990
rect 5390 12970 5450 12990
rect 5470 12970 5530 12990
rect 5550 12970 5610 12990
rect 5630 12970 5690 12990
rect 5710 12970 5720 12990
rect 4720 12960 5720 12970
rect 5760 12990 5960 13000
rect 5760 12970 5770 12990
rect 5790 12970 5850 12990
rect 5870 12970 5930 12990
rect 5950 12970 5960 12990
rect 5760 12960 5960 12970
rect 6000 12990 6200 13000
rect 6000 12970 6010 12990
rect 6030 12970 6090 12990
rect 6110 12970 6170 12990
rect 6190 12970 6200 12990
rect 6000 12960 6200 12970
rect 4240 12910 4440 12920
rect 4240 12890 4250 12910
rect 4270 12890 4330 12910
rect 4350 12890 4410 12910
rect 4430 12890 4440 12910
rect 4240 12880 4440 12890
rect 4480 12910 4680 12920
rect 4480 12890 4490 12910
rect 4510 12890 4570 12910
rect 4590 12890 4650 12910
rect 4670 12890 4680 12910
rect 4480 12880 4680 12890
rect 4720 12910 5720 12920
rect 4720 12890 4730 12910
rect 4750 12890 4810 12910
rect 4830 12890 4890 12910
rect 4910 12890 4970 12910
rect 4990 12890 5050 12910
rect 5070 12890 5130 12910
rect 5150 12890 5210 12910
rect 5230 12890 5290 12910
rect 5310 12890 5370 12910
rect 5390 12890 5450 12910
rect 5470 12890 5530 12910
rect 5550 12890 5610 12910
rect 5630 12890 5690 12910
rect 5710 12890 5720 12910
rect 4720 12880 5720 12890
rect 5760 12910 5960 12920
rect 5760 12890 5770 12910
rect 5790 12890 5850 12910
rect 5870 12890 5930 12910
rect 5950 12890 5960 12910
rect 5760 12880 5960 12890
rect 6000 12910 6200 12920
rect 6000 12890 6010 12910
rect 6030 12890 6090 12910
rect 6110 12890 6170 12910
rect 6190 12890 6200 12910
rect 6000 12880 6200 12890
rect 4240 12830 4440 12840
rect 4240 12810 4250 12830
rect 4270 12810 4330 12830
rect 4350 12810 4410 12830
rect 4430 12810 4440 12830
rect 4240 12800 4440 12810
rect 4480 12830 4680 12840
rect 4480 12810 4490 12830
rect 4510 12810 4570 12830
rect 4590 12810 4650 12830
rect 4670 12810 4680 12830
rect 4480 12800 4680 12810
rect 4720 12830 5720 12840
rect 4720 12810 4730 12830
rect 4750 12810 4810 12830
rect 4830 12810 4890 12830
rect 4910 12810 4970 12830
rect 4990 12810 5050 12830
rect 5070 12810 5130 12830
rect 5150 12810 5210 12830
rect 5230 12810 5290 12830
rect 5310 12810 5370 12830
rect 5390 12810 5450 12830
rect 5470 12810 5530 12830
rect 5550 12810 5610 12830
rect 5630 12810 5690 12830
rect 5710 12810 5720 12830
rect 4720 12800 5720 12810
rect 5760 12830 5960 12840
rect 5760 12810 5770 12830
rect 5790 12810 5850 12830
rect 5870 12810 5930 12830
rect 5950 12810 5960 12830
rect 5760 12800 5960 12810
rect 6000 12830 6200 12840
rect 6000 12810 6010 12830
rect 6030 12810 6090 12830
rect 6110 12810 6170 12830
rect 6190 12810 6200 12830
rect 6000 12800 6200 12810
rect 4240 12750 4440 12760
rect 4240 12730 4250 12750
rect 4270 12730 4330 12750
rect 4350 12730 4410 12750
rect 4430 12730 4440 12750
rect 4240 12720 4440 12730
rect 4480 12750 4680 12760
rect 4480 12730 4490 12750
rect 4510 12730 4570 12750
rect 4590 12730 4650 12750
rect 4670 12730 4680 12750
rect 4480 12720 4680 12730
rect 4720 12750 5720 12760
rect 4720 12730 4730 12750
rect 4750 12730 4810 12750
rect 4830 12730 4890 12750
rect 4910 12730 4970 12750
rect 4990 12730 5050 12750
rect 5070 12730 5130 12750
rect 5150 12730 5210 12750
rect 5230 12730 5290 12750
rect 5310 12730 5370 12750
rect 5390 12730 5450 12750
rect 5470 12730 5530 12750
rect 5550 12730 5610 12750
rect 5630 12730 5690 12750
rect 5710 12730 5720 12750
rect 4720 12720 5720 12730
rect 5760 12750 5960 12760
rect 5760 12730 5770 12750
rect 5790 12730 5850 12750
rect 5870 12730 5930 12750
rect 5950 12730 5960 12750
rect 5760 12720 5960 12730
rect 6000 12750 6200 12760
rect 6000 12730 6010 12750
rect 6030 12730 6090 12750
rect 6110 12730 6170 12750
rect 6190 12730 6200 12750
rect 6000 12720 6200 12730
rect 4240 12670 4440 12680
rect 4240 12650 4250 12670
rect 4270 12650 4330 12670
rect 4350 12650 4410 12670
rect 4430 12650 4440 12670
rect 4240 12640 4440 12650
rect 4480 12670 4680 12680
rect 4480 12650 4490 12670
rect 4510 12650 4570 12670
rect 4590 12650 4650 12670
rect 4670 12650 4680 12670
rect 4480 12640 4680 12650
rect 4720 12670 5720 12680
rect 4720 12650 4730 12670
rect 4750 12650 4810 12670
rect 4830 12650 4890 12670
rect 4910 12650 4970 12670
rect 4990 12650 5050 12670
rect 5070 12650 5130 12670
rect 5150 12650 5210 12670
rect 5230 12650 5290 12670
rect 5310 12650 5370 12670
rect 5390 12650 5450 12670
rect 5470 12650 5530 12670
rect 5550 12650 5610 12670
rect 5630 12650 5690 12670
rect 5710 12650 5720 12670
rect 4720 12640 5720 12650
rect 5760 12670 5960 12680
rect 5760 12650 5770 12670
rect 5790 12650 5850 12670
rect 5870 12650 5930 12670
rect 5950 12650 5960 12670
rect 5760 12640 5960 12650
rect 6000 12670 6200 12680
rect 6000 12650 6010 12670
rect 6030 12650 6090 12670
rect 6110 12650 6170 12670
rect 6190 12650 6200 12670
rect 6000 12640 6200 12650
rect 4240 12590 4440 12600
rect 4240 12570 4250 12590
rect 4270 12570 4330 12590
rect 4350 12570 4410 12590
rect 4430 12570 4440 12590
rect 4240 12560 4440 12570
rect 4480 12590 4680 12600
rect 4480 12570 4490 12590
rect 4510 12570 4570 12590
rect 4590 12570 4650 12590
rect 4670 12570 4680 12590
rect 4480 12560 4680 12570
rect 4720 12590 5720 12600
rect 4720 12570 4730 12590
rect 4750 12570 4810 12590
rect 4830 12570 4890 12590
rect 4910 12570 4970 12590
rect 4990 12570 5050 12590
rect 5070 12570 5130 12590
rect 5150 12570 5210 12590
rect 5230 12570 5290 12590
rect 5310 12570 5370 12590
rect 5390 12570 5450 12590
rect 5470 12570 5530 12590
rect 5550 12570 5610 12590
rect 5630 12570 5690 12590
rect 5710 12570 5720 12590
rect 4720 12560 5720 12570
rect 5760 12590 5960 12600
rect 5760 12570 5770 12590
rect 5790 12570 5850 12590
rect 5870 12570 5930 12590
rect 5950 12570 5960 12590
rect 5760 12560 5960 12570
rect 6000 12590 6200 12600
rect 6000 12570 6010 12590
rect 6030 12570 6090 12590
rect 6110 12570 6170 12590
rect 6190 12570 6200 12590
rect 6000 12560 6200 12570
rect 4240 12510 4440 12520
rect 4240 12490 4250 12510
rect 4270 12490 4330 12510
rect 4350 12490 4410 12510
rect 4430 12490 4440 12510
rect 4240 12480 4440 12490
rect 4480 12510 4680 12520
rect 4480 12490 4490 12510
rect 4510 12490 4570 12510
rect 4590 12490 4650 12510
rect 4670 12490 4680 12510
rect 4480 12480 4680 12490
rect 4720 12510 5720 12520
rect 4720 12490 4730 12510
rect 4750 12490 4810 12510
rect 4830 12490 4890 12510
rect 4910 12490 4970 12510
rect 4990 12490 5050 12510
rect 5070 12490 5130 12510
rect 5150 12490 5210 12510
rect 5230 12490 5290 12510
rect 5310 12490 5370 12510
rect 5390 12490 5450 12510
rect 5470 12490 5530 12510
rect 5550 12490 5610 12510
rect 5630 12490 5690 12510
rect 5710 12490 5720 12510
rect 4720 12480 5720 12490
rect 5760 12510 5960 12520
rect 5760 12490 5770 12510
rect 5790 12490 5850 12510
rect 5870 12490 5930 12510
rect 5950 12490 5960 12510
rect 5760 12480 5960 12490
rect 6000 12510 6200 12520
rect 6000 12490 6010 12510
rect 6030 12490 6090 12510
rect 6110 12490 6170 12510
rect 6190 12490 6200 12510
rect 6000 12480 6200 12490
rect 4240 12430 4440 12440
rect 4240 12410 4250 12430
rect 4270 12410 4330 12430
rect 4350 12410 4410 12430
rect 4430 12410 4440 12430
rect 4240 12400 4440 12410
rect 4480 12430 4680 12440
rect 4480 12410 4490 12430
rect 4510 12410 4570 12430
rect 4590 12410 4650 12430
rect 4670 12410 4680 12430
rect 4480 12400 4680 12410
rect 4720 12430 5720 12440
rect 4720 12410 4730 12430
rect 4750 12410 4810 12430
rect 4830 12410 4890 12430
rect 4910 12410 4970 12430
rect 4990 12410 5050 12430
rect 5070 12410 5130 12430
rect 5150 12410 5210 12430
rect 5230 12410 5290 12430
rect 5310 12410 5370 12430
rect 5390 12410 5450 12430
rect 5470 12410 5530 12430
rect 5550 12410 5610 12430
rect 5630 12410 5690 12430
rect 5710 12410 5720 12430
rect 4720 12400 5720 12410
rect 5760 12430 5960 12440
rect 5760 12410 5770 12430
rect 5790 12410 5850 12430
rect 5870 12410 5930 12430
rect 5950 12410 5960 12430
rect 5760 12400 5960 12410
rect 6000 12430 6200 12440
rect 6000 12410 6010 12430
rect 6030 12410 6090 12430
rect 6110 12410 6170 12430
rect 6190 12410 6200 12430
rect 6000 12400 6200 12410
rect 4240 12350 4440 12360
rect 4240 12330 4250 12350
rect 4270 12330 4330 12350
rect 4350 12330 4410 12350
rect 4430 12330 4440 12350
rect 4240 12320 4440 12330
rect 4480 12350 4680 12360
rect 4480 12330 4490 12350
rect 4510 12330 4570 12350
rect 4590 12330 4650 12350
rect 4670 12330 4680 12350
rect 4480 12320 4680 12330
rect 4720 12350 5720 12360
rect 4720 12330 4730 12350
rect 4750 12330 4810 12350
rect 4830 12330 4890 12350
rect 4910 12330 4970 12350
rect 4990 12330 5050 12350
rect 5070 12330 5130 12350
rect 5150 12330 5210 12350
rect 5230 12330 5290 12350
rect 5310 12330 5370 12350
rect 5390 12330 5450 12350
rect 5470 12330 5530 12350
rect 5550 12330 5610 12350
rect 5630 12330 5690 12350
rect 5710 12330 5720 12350
rect 4720 12320 5720 12330
rect 5760 12350 5960 12360
rect 5760 12330 5770 12350
rect 5790 12330 5850 12350
rect 5870 12330 5930 12350
rect 5950 12330 5960 12350
rect 5760 12320 5960 12330
rect 6000 12350 6200 12360
rect 6000 12330 6010 12350
rect 6030 12330 6090 12350
rect 6110 12330 6170 12350
rect 6190 12330 6200 12350
rect 6000 12320 6200 12330
rect 4240 12270 4440 12280
rect 4240 12250 4250 12270
rect 4270 12250 4330 12270
rect 4350 12250 4410 12270
rect 4430 12250 4440 12270
rect 4240 12240 4440 12250
rect 4480 12270 4680 12280
rect 4480 12250 4490 12270
rect 4510 12250 4570 12270
rect 4590 12250 4650 12270
rect 4670 12250 4680 12270
rect 4480 12240 4680 12250
rect 4720 12270 5720 12280
rect 4720 12250 4730 12270
rect 4750 12250 4810 12270
rect 4830 12250 4890 12270
rect 4910 12250 4970 12270
rect 4990 12250 5050 12270
rect 5070 12250 5130 12270
rect 5150 12250 5210 12270
rect 5230 12250 5290 12270
rect 5310 12250 5370 12270
rect 5390 12250 5450 12270
rect 5470 12250 5530 12270
rect 5550 12250 5610 12270
rect 5630 12250 5690 12270
rect 5710 12250 5720 12270
rect 4720 12240 5720 12250
rect 5760 12270 5960 12280
rect 5760 12250 5770 12270
rect 5790 12250 5850 12270
rect 5870 12250 5930 12270
rect 5950 12250 5960 12270
rect 5760 12240 5960 12250
rect 6000 12270 6200 12280
rect 6000 12250 6010 12270
rect 6030 12250 6090 12270
rect 6110 12250 6170 12270
rect 6190 12250 6200 12270
rect 6000 12240 6200 12250
rect 4240 12190 4440 12200
rect 4240 12170 4250 12190
rect 4270 12170 4330 12190
rect 4350 12170 4410 12190
rect 4430 12170 4440 12190
rect 4240 12160 4440 12170
rect 4480 12190 4680 12200
rect 4480 12170 4490 12190
rect 4510 12170 4570 12190
rect 4590 12170 4650 12190
rect 4670 12170 4680 12190
rect 4480 12160 4680 12170
rect 4720 12190 5720 12200
rect 4720 12170 4730 12190
rect 4750 12170 4810 12190
rect 4830 12170 4890 12190
rect 4910 12170 4970 12190
rect 4990 12170 5050 12190
rect 5070 12170 5130 12190
rect 5150 12170 5210 12190
rect 5230 12170 5290 12190
rect 5310 12170 5370 12190
rect 5390 12170 5450 12190
rect 5470 12170 5530 12190
rect 5550 12170 5610 12190
rect 5630 12170 5690 12190
rect 5710 12170 5720 12190
rect 4720 12160 5720 12170
rect 5760 12190 5960 12200
rect 5760 12170 5770 12190
rect 5790 12170 5850 12190
rect 5870 12170 5930 12190
rect 5950 12170 5960 12190
rect 5760 12160 5960 12170
rect 6000 12190 6200 12200
rect 6000 12170 6010 12190
rect 6030 12170 6090 12190
rect 6110 12170 6170 12190
rect 6190 12170 6200 12190
rect 6000 12160 6200 12170
rect 4240 12110 4440 12120
rect 4240 12090 4250 12110
rect 4270 12090 4330 12110
rect 4350 12090 4410 12110
rect 4430 12090 4440 12110
rect 4240 12080 4440 12090
rect 4480 12110 4680 12120
rect 4480 12090 4490 12110
rect 4510 12090 4570 12110
rect 4590 12090 4650 12110
rect 4670 12090 4680 12110
rect 4480 12080 4680 12090
rect 4720 12110 5720 12120
rect 4720 12090 4730 12110
rect 4750 12090 4810 12110
rect 4830 12090 4890 12110
rect 4910 12090 4970 12110
rect 4990 12090 5050 12110
rect 5070 12090 5130 12110
rect 5150 12090 5210 12110
rect 5230 12090 5290 12110
rect 5310 12090 5370 12110
rect 5390 12090 5450 12110
rect 5470 12090 5530 12110
rect 5550 12090 5610 12110
rect 5630 12090 5690 12110
rect 5710 12090 5720 12110
rect 4720 12080 5720 12090
rect 5760 12110 5960 12120
rect 5760 12090 5770 12110
rect 5790 12090 5850 12110
rect 5870 12090 5930 12110
rect 5950 12090 5960 12110
rect 5760 12080 5960 12090
rect 6000 12110 6200 12120
rect 6000 12090 6010 12110
rect 6030 12090 6090 12110
rect 6110 12090 6170 12110
rect 6190 12090 6200 12110
rect 6000 12080 6200 12090
rect 4240 12030 4440 12040
rect 4240 12010 4250 12030
rect 4270 12010 4330 12030
rect 4350 12010 4410 12030
rect 4430 12010 4440 12030
rect 4240 12000 4440 12010
rect 4480 12030 4680 12040
rect 4480 12010 4490 12030
rect 4510 12010 4570 12030
rect 4590 12010 4650 12030
rect 4670 12010 4680 12030
rect 4480 12000 4680 12010
rect 4720 12030 5720 12040
rect 4720 12010 4730 12030
rect 4750 12010 4810 12030
rect 4830 12010 4890 12030
rect 4910 12010 4970 12030
rect 4990 12010 5050 12030
rect 5070 12010 5130 12030
rect 5150 12010 5210 12030
rect 5230 12010 5290 12030
rect 5310 12010 5370 12030
rect 5390 12010 5450 12030
rect 5470 12010 5530 12030
rect 5550 12010 5610 12030
rect 5630 12010 5690 12030
rect 5710 12010 5720 12030
rect 4720 12000 5720 12010
rect 5760 12030 5960 12040
rect 5760 12010 5770 12030
rect 5790 12010 5850 12030
rect 5870 12010 5930 12030
rect 5950 12010 5960 12030
rect 5760 12000 5960 12010
rect 6000 12030 6200 12040
rect 6000 12010 6010 12030
rect 6030 12010 6090 12030
rect 6110 12010 6170 12030
rect 6190 12010 6200 12030
rect 6000 12000 6200 12010
rect 4240 11950 4440 11960
rect 4240 11930 4250 11950
rect 4270 11930 4330 11950
rect 4350 11930 4410 11950
rect 4430 11930 4440 11950
rect 4240 11920 4440 11930
rect 4480 11950 4680 11960
rect 4480 11930 4490 11950
rect 4510 11930 4570 11950
rect 4590 11930 4650 11950
rect 4670 11930 4680 11950
rect 4480 11920 4680 11930
rect 4720 11950 5720 11960
rect 4720 11930 4730 11950
rect 4750 11930 4810 11950
rect 4830 11930 4890 11950
rect 4910 11930 4970 11950
rect 4990 11930 5050 11950
rect 5070 11930 5130 11950
rect 5150 11930 5210 11950
rect 5230 11930 5290 11950
rect 5310 11930 5370 11950
rect 5390 11930 5450 11950
rect 5470 11930 5530 11950
rect 5550 11930 5610 11950
rect 5630 11930 5690 11950
rect 5710 11930 5720 11950
rect 4720 11920 5720 11930
rect 5760 11950 5960 11960
rect 5760 11930 5770 11950
rect 5790 11930 5850 11950
rect 5870 11930 5930 11950
rect 5950 11930 5960 11950
rect 5760 11920 5960 11930
rect 6000 11950 6200 11960
rect 6000 11930 6010 11950
rect 6030 11930 6090 11950
rect 6110 11930 6170 11950
rect 6190 11930 6200 11950
rect 6000 11920 6200 11930
rect 4240 11870 4440 11880
rect 4240 11850 4250 11870
rect 4270 11850 4330 11870
rect 4350 11850 4410 11870
rect 4430 11850 4440 11870
rect 4240 11840 4440 11850
rect 4480 11870 4680 11880
rect 4480 11850 4490 11870
rect 4510 11850 4570 11870
rect 4590 11850 4650 11870
rect 4670 11850 4680 11870
rect 4480 11840 4680 11850
rect 4720 11870 5720 11880
rect 4720 11850 4730 11870
rect 4750 11850 4810 11870
rect 4830 11850 4890 11870
rect 4910 11850 4970 11870
rect 4990 11850 5050 11870
rect 5070 11850 5130 11870
rect 5150 11850 5210 11870
rect 5230 11850 5290 11870
rect 5310 11850 5370 11870
rect 5390 11850 5450 11870
rect 5470 11850 5530 11870
rect 5550 11850 5610 11870
rect 5630 11850 5690 11870
rect 5710 11850 5720 11870
rect 4720 11840 5720 11850
rect 5760 11870 5960 11880
rect 5760 11850 5770 11870
rect 5790 11850 5850 11870
rect 5870 11850 5930 11870
rect 5950 11850 5960 11870
rect 5760 11840 5960 11850
rect 6000 11870 6200 11880
rect 6000 11850 6010 11870
rect 6030 11850 6090 11870
rect 6110 11850 6170 11870
rect 6190 11850 6200 11870
rect 6000 11840 6200 11850
rect 4240 11790 4440 11800
rect 4240 11770 4250 11790
rect 4270 11770 4330 11790
rect 4350 11770 4410 11790
rect 4430 11770 4440 11790
rect 4240 11760 4440 11770
rect 4480 11790 4680 11800
rect 4480 11770 4490 11790
rect 4510 11770 4570 11790
rect 4590 11770 4650 11790
rect 4670 11770 4680 11790
rect 4480 11760 4680 11770
rect 4720 11790 5720 11800
rect 4720 11770 4730 11790
rect 4750 11770 4810 11790
rect 4830 11770 4890 11790
rect 4910 11770 4970 11790
rect 4990 11770 5050 11790
rect 5070 11770 5130 11790
rect 5150 11770 5210 11790
rect 5230 11770 5290 11790
rect 5310 11770 5370 11790
rect 5390 11770 5450 11790
rect 5470 11770 5530 11790
rect 5550 11770 5610 11790
rect 5630 11770 5690 11790
rect 5710 11770 5720 11790
rect 4720 11760 5720 11770
rect 5760 11790 5960 11800
rect 5760 11770 5770 11790
rect 5790 11770 5850 11790
rect 5870 11770 5930 11790
rect 5950 11770 5960 11790
rect 5760 11760 5960 11770
rect 6000 11790 6200 11800
rect 6000 11770 6010 11790
rect 6030 11770 6090 11790
rect 6110 11770 6170 11790
rect 6190 11770 6200 11790
rect 6000 11760 6200 11770
rect 4240 11710 4440 11720
rect 4240 11690 4250 11710
rect 4270 11690 4330 11710
rect 4350 11690 4410 11710
rect 4430 11690 4440 11710
rect 4240 11680 4440 11690
rect 4480 11710 4680 11720
rect 4480 11690 4490 11710
rect 4510 11690 4570 11710
rect 4590 11690 4650 11710
rect 4670 11690 4680 11710
rect 4480 11680 4680 11690
rect 4720 11710 5720 11720
rect 4720 11690 4730 11710
rect 4750 11690 4810 11710
rect 4830 11690 4890 11710
rect 4910 11690 4970 11710
rect 4990 11690 5050 11710
rect 5070 11690 5130 11710
rect 5150 11690 5210 11710
rect 5230 11690 5290 11710
rect 5310 11690 5370 11710
rect 5390 11690 5450 11710
rect 5470 11690 5530 11710
rect 5550 11690 5610 11710
rect 5630 11690 5690 11710
rect 5710 11690 5720 11710
rect 4720 11680 5720 11690
rect 5760 11710 5960 11720
rect 5760 11690 5770 11710
rect 5790 11690 5850 11710
rect 5870 11690 5930 11710
rect 5950 11690 5960 11710
rect 5760 11680 5960 11690
rect 6000 11710 6200 11720
rect 6000 11690 6010 11710
rect 6030 11690 6090 11710
rect 6110 11690 6170 11710
rect 6190 11690 6200 11710
rect 6000 11680 6200 11690
rect 4240 11630 4440 11640
rect 4240 11610 4250 11630
rect 4270 11610 4330 11630
rect 4350 11610 4410 11630
rect 4430 11610 4440 11630
rect 4240 11600 4440 11610
rect 4480 11630 4680 11640
rect 4480 11610 4490 11630
rect 4510 11610 4570 11630
rect 4590 11610 4650 11630
rect 4670 11610 4680 11630
rect 4480 11600 4680 11610
rect 4720 11630 5720 11640
rect 4720 11610 4730 11630
rect 4750 11610 4810 11630
rect 4830 11610 4890 11630
rect 4910 11610 4970 11630
rect 4990 11610 5050 11630
rect 5070 11610 5130 11630
rect 5150 11610 5210 11630
rect 5230 11610 5290 11630
rect 5310 11610 5370 11630
rect 5390 11610 5450 11630
rect 5470 11610 5530 11630
rect 5550 11610 5610 11630
rect 5630 11610 5690 11630
rect 5710 11610 5720 11630
rect 4720 11600 5720 11610
rect 5760 11630 5960 11640
rect 5760 11610 5770 11630
rect 5790 11610 5850 11630
rect 5870 11610 5930 11630
rect 5950 11610 5960 11630
rect 5760 11600 5960 11610
rect 6000 11630 6200 11640
rect 6000 11610 6010 11630
rect 6030 11610 6090 11630
rect 6110 11610 6170 11630
rect 6190 11610 6200 11630
rect 6000 11600 6200 11610
rect 4240 11550 4440 11560
rect 4240 11530 4250 11550
rect 4270 11530 4330 11550
rect 4350 11530 4410 11550
rect 4430 11530 4440 11550
rect 4240 11520 4440 11530
rect 4480 11550 4680 11560
rect 4480 11530 4490 11550
rect 4510 11530 4570 11550
rect 4590 11530 4650 11550
rect 4670 11530 4680 11550
rect 4480 11520 4680 11530
rect 4720 11550 5720 11560
rect 4720 11530 4730 11550
rect 4750 11530 4810 11550
rect 4830 11530 4890 11550
rect 4910 11530 4970 11550
rect 4990 11530 5050 11550
rect 5070 11530 5130 11550
rect 5150 11530 5210 11550
rect 5230 11530 5290 11550
rect 5310 11530 5370 11550
rect 5390 11530 5450 11550
rect 5470 11530 5530 11550
rect 5550 11530 5610 11550
rect 5630 11530 5690 11550
rect 5710 11530 5720 11550
rect 4720 11520 5720 11530
rect 5760 11550 5960 11560
rect 5760 11530 5770 11550
rect 5790 11530 5850 11550
rect 5870 11530 5930 11550
rect 5950 11530 5960 11550
rect 5760 11520 5960 11530
rect 6000 11550 6200 11560
rect 6000 11530 6010 11550
rect 6030 11530 6090 11550
rect 6110 11530 6170 11550
rect 6190 11530 6200 11550
rect 6000 11520 6200 11530
rect 4240 11470 4440 11480
rect 4240 11450 4250 11470
rect 4270 11450 4330 11470
rect 4350 11450 4410 11470
rect 4430 11450 4440 11470
rect 4240 11440 4440 11450
rect 4480 11470 4680 11480
rect 4480 11450 4490 11470
rect 4510 11450 4570 11470
rect 4590 11450 4650 11470
rect 4670 11450 4680 11470
rect 4480 11440 4680 11450
rect 4720 11470 5720 11480
rect 4720 11450 4730 11470
rect 4750 11450 4810 11470
rect 4830 11450 4890 11470
rect 4910 11450 4970 11470
rect 4990 11450 5050 11470
rect 5070 11450 5130 11470
rect 5150 11450 5210 11470
rect 5230 11450 5290 11470
rect 5310 11450 5370 11470
rect 5390 11450 5450 11470
rect 5470 11450 5530 11470
rect 5550 11450 5610 11470
rect 5630 11450 5690 11470
rect 5710 11450 5720 11470
rect 4720 11440 5720 11450
rect 5760 11470 5960 11480
rect 5760 11450 5770 11470
rect 5790 11450 5850 11470
rect 5870 11450 5930 11470
rect 5950 11450 5960 11470
rect 5760 11440 5960 11450
rect 6000 11470 6200 11480
rect 6000 11450 6010 11470
rect 6030 11450 6090 11470
rect 6110 11450 6170 11470
rect 6190 11450 6200 11470
rect 6000 11440 6200 11450
rect 4240 11390 4440 11400
rect 4240 11370 4250 11390
rect 4270 11370 4330 11390
rect 4350 11370 4410 11390
rect 4430 11370 4440 11390
rect 4240 11360 4440 11370
rect 4480 11390 4680 11400
rect 4480 11370 4490 11390
rect 4510 11370 4570 11390
rect 4590 11370 4650 11390
rect 4670 11370 4680 11390
rect 4480 11360 4680 11370
rect 4720 11390 5720 11400
rect 4720 11370 4730 11390
rect 4750 11370 4810 11390
rect 4830 11370 4890 11390
rect 4910 11370 4970 11390
rect 4990 11370 5050 11390
rect 5070 11370 5130 11390
rect 5150 11370 5210 11390
rect 5230 11370 5290 11390
rect 5310 11370 5370 11390
rect 5390 11370 5450 11390
rect 5470 11370 5530 11390
rect 5550 11370 5610 11390
rect 5630 11370 5690 11390
rect 5710 11370 5720 11390
rect 4720 11360 5720 11370
rect 5760 11390 5960 11400
rect 5760 11370 5770 11390
rect 5790 11370 5850 11390
rect 5870 11370 5930 11390
rect 5950 11370 5960 11390
rect 5760 11360 5960 11370
rect 6000 11390 6200 11400
rect 6000 11370 6010 11390
rect 6030 11370 6090 11390
rect 6110 11370 6170 11390
rect 6190 11370 6200 11390
rect 6000 11360 6200 11370
rect 4240 11310 4440 11320
rect 4240 11290 4250 11310
rect 4270 11290 4330 11310
rect 4350 11290 4410 11310
rect 4430 11290 4440 11310
rect 4240 11280 4440 11290
rect 4480 11310 4680 11320
rect 4480 11290 4490 11310
rect 4510 11290 4570 11310
rect 4590 11290 4650 11310
rect 4670 11290 4680 11310
rect 4480 11280 4680 11290
rect 4720 11310 5720 11320
rect 4720 11290 4730 11310
rect 4750 11290 4810 11310
rect 4830 11290 4890 11310
rect 4910 11290 4970 11310
rect 4990 11290 5050 11310
rect 5070 11290 5130 11310
rect 5150 11290 5210 11310
rect 5230 11290 5290 11310
rect 5310 11290 5370 11310
rect 5390 11290 5450 11310
rect 5470 11290 5530 11310
rect 5550 11290 5610 11310
rect 5630 11290 5690 11310
rect 5710 11290 5720 11310
rect 4720 11280 5720 11290
rect 5760 11310 5960 11320
rect 5760 11290 5770 11310
rect 5790 11290 5850 11310
rect 5870 11290 5930 11310
rect 5950 11290 5960 11310
rect 5760 11280 5960 11290
rect 6000 11310 6200 11320
rect 6000 11290 6010 11310
rect 6030 11290 6090 11310
rect 6110 11290 6170 11310
rect 6190 11290 6200 11310
rect 6000 11280 6200 11290
rect 4240 11230 4440 11240
rect 4240 11210 4250 11230
rect 4270 11210 4330 11230
rect 4350 11210 4410 11230
rect 4430 11210 4440 11230
rect 4240 11200 4440 11210
rect 4480 11230 4680 11240
rect 4480 11210 4490 11230
rect 4510 11210 4570 11230
rect 4590 11210 4650 11230
rect 4670 11210 4680 11230
rect 4480 11200 4680 11210
rect 4720 11230 5720 11240
rect 4720 11210 4730 11230
rect 4750 11210 4810 11230
rect 4830 11210 4890 11230
rect 4910 11210 4970 11230
rect 4990 11210 5050 11230
rect 5070 11210 5130 11230
rect 5150 11210 5210 11230
rect 5230 11210 5290 11230
rect 5310 11210 5370 11230
rect 5390 11210 5450 11230
rect 5470 11210 5530 11230
rect 5550 11210 5610 11230
rect 5630 11210 5690 11230
rect 5710 11210 5720 11230
rect 4720 11200 5720 11210
rect 5760 11230 5960 11240
rect 5760 11210 5770 11230
rect 5790 11210 5850 11230
rect 5870 11210 5930 11230
rect 5950 11210 5960 11230
rect 5760 11200 5960 11210
rect 6000 11230 6200 11240
rect 6000 11210 6010 11230
rect 6030 11210 6090 11230
rect 6110 11210 6170 11230
rect 6190 11210 6200 11230
rect 6000 11200 6200 11210
rect 4240 11150 4440 11160
rect 4240 11130 4250 11150
rect 4270 11130 4330 11150
rect 4350 11130 4410 11150
rect 4430 11130 4440 11150
rect 4240 11120 4440 11130
rect 4480 11150 4680 11160
rect 4480 11130 4490 11150
rect 4510 11130 4570 11150
rect 4590 11130 4650 11150
rect 4670 11130 4680 11150
rect 4480 11120 4680 11130
rect 4720 11150 5720 11160
rect 4720 11130 4730 11150
rect 4750 11130 4810 11150
rect 4830 11130 4890 11150
rect 4910 11130 4970 11150
rect 4990 11130 5050 11150
rect 5070 11130 5130 11150
rect 5150 11130 5210 11150
rect 5230 11130 5290 11150
rect 5310 11130 5370 11150
rect 5390 11130 5450 11150
rect 5470 11130 5530 11150
rect 5550 11130 5610 11150
rect 5630 11130 5690 11150
rect 5710 11130 5720 11150
rect 4720 11120 5720 11130
rect 5760 11150 5960 11160
rect 5760 11130 5770 11150
rect 5790 11130 5850 11150
rect 5870 11130 5930 11150
rect 5950 11130 5960 11150
rect 5760 11120 5960 11130
rect 6000 11150 6200 11160
rect 6000 11130 6010 11150
rect 6030 11130 6090 11150
rect 6110 11130 6170 11150
rect 6190 11130 6200 11150
rect 6000 11120 6200 11130
rect 4240 11070 4440 11080
rect 4240 11050 4250 11070
rect 4270 11050 4330 11070
rect 4350 11050 4410 11070
rect 4430 11050 4440 11070
rect 4240 11040 4440 11050
rect 4480 11070 4680 11080
rect 4480 11050 4490 11070
rect 4510 11050 4570 11070
rect 4590 11050 4650 11070
rect 4670 11050 4680 11070
rect 4480 11040 4680 11050
rect 4720 11070 5720 11080
rect 4720 11050 4730 11070
rect 4750 11050 4810 11070
rect 4830 11050 4890 11070
rect 4910 11050 4970 11070
rect 4990 11050 5050 11070
rect 5070 11050 5130 11070
rect 5150 11050 5210 11070
rect 5230 11050 5290 11070
rect 5310 11050 5370 11070
rect 5390 11050 5450 11070
rect 5470 11050 5530 11070
rect 5550 11050 5610 11070
rect 5630 11050 5690 11070
rect 5710 11050 5720 11070
rect 4720 11040 5720 11050
rect 5760 11070 5960 11080
rect 5760 11050 5770 11070
rect 5790 11050 5850 11070
rect 5870 11050 5930 11070
rect 5950 11050 5960 11070
rect 5760 11040 5960 11050
rect 6000 11070 6200 11080
rect 6000 11050 6010 11070
rect 6030 11050 6090 11070
rect 6110 11050 6170 11070
rect 6190 11050 6200 11070
rect 6000 11040 6200 11050
rect 4240 10990 4440 11000
rect 4240 10970 4250 10990
rect 4270 10970 4330 10990
rect 4350 10970 4410 10990
rect 4430 10970 4440 10990
rect 4240 10960 4440 10970
rect 4480 10990 4680 11000
rect 4480 10970 4490 10990
rect 4510 10970 4570 10990
rect 4590 10970 4650 10990
rect 4670 10970 4680 10990
rect 4480 10960 4680 10970
rect 4720 10990 5720 11000
rect 4720 10970 4730 10990
rect 4750 10970 4810 10990
rect 4830 10970 4890 10990
rect 4910 10970 4970 10990
rect 4990 10970 5050 10990
rect 5070 10970 5130 10990
rect 5150 10970 5210 10990
rect 5230 10970 5290 10990
rect 5310 10970 5370 10990
rect 5390 10970 5450 10990
rect 5470 10970 5530 10990
rect 5550 10970 5610 10990
rect 5630 10970 5690 10990
rect 5710 10970 5720 10990
rect 4720 10960 5720 10970
rect 5760 10990 5960 11000
rect 5760 10970 5770 10990
rect 5790 10970 5850 10990
rect 5870 10970 5930 10990
rect 5950 10970 5960 10990
rect 5760 10960 5960 10970
rect 6000 10990 6200 11000
rect 6000 10970 6010 10990
rect 6030 10970 6090 10990
rect 6110 10970 6170 10990
rect 6190 10970 6200 10990
rect 6000 10960 6200 10970
rect 4240 10910 4440 10920
rect 4240 10890 4250 10910
rect 4270 10890 4330 10910
rect 4350 10890 4410 10910
rect 4430 10890 4440 10910
rect 4240 10880 4440 10890
rect 4480 10910 4680 10920
rect 4480 10890 4490 10910
rect 4510 10890 4570 10910
rect 4590 10890 4650 10910
rect 4670 10890 4680 10910
rect 4480 10880 4680 10890
rect 4720 10910 5720 10920
rect 4720 10890 4730 10910
rect 4750 10890 4810 10910
rect 4830 10890 4890 10910
rect 4910 10890 4970 10910
rect 4990 10890 5050 10910
rect 5070 10890 5130 10910
rect 5150 10890 5210 10910
rect 5230 10890 5290 10910
rect 5310 10890 5370 10910
rect 5390 10890 5450 10910
rect 5470 10890 5530 10910
rect 5550 10890 5610 10910
rect 5630 10890 5690 10910
rect 5710 10890 5720 10910
rect 4720 10880 5720 10890
rect 5760 10910 5960 10920
rect 5760 10890 5770 10910
rect 5790 10890 5850 10910
rect 5870 10890 5930 10910
rect 5950 10890 5960 10910
rect 5760 10880 5960 10890
rect 6000 10910 6200 10920
rect 6000 10890 6010 10910
rect 6030 10890 6090 10910
rect 6110 10890 6170 10910
rect 6190 10890 6200 10910
rect 6000 10880 6200 10890
rect 4240 10830 4440 10840
rect 4240 10810 4250 10830
rect 4270 10810 4330 10830
rect 4350 10810 4410 10830
rect 4430 10810 4440 10830
rect 4240 10800 4440 10810
rect 4480 10830 4680 10840
rect 4480 10810 4490 10830
rect 4510 10810 4570 10830
rect 4590 10810 4650 10830
rect 4670 10810 4680 10830
rect 4480 10800 4680 10810
rect 4720 10830 5720 10840
rect 4720 10810 4730 10830
rect 4750 10810 4810 10830
rect 4830 10810 4890 10830
rect 4910 10810 4970 10830
rect 4990 10810 5050 10830
rect 5070 10810 5130 10830
rect 5150 10810 5210 10830
rect 5230 10810 5290 10830
rect 5310 10810 5370 10830
rect 5390 10810 5450 10830
rect 5470 10810 5530 10830
rect 5550 10810 5610 10830
rect 5630 10810 5690 10830
rect 5710 10810 5720 10830
rect 4720 10800 5720 10810
rect 5760 10830 5960 10840
rect 5760 10810 5770 10830
rect 5790 10810 5850 10830
rect 5870 10810 5930 10830
rect 5950 10810 5960 10830
rect 5760 10800 5960 10810
rect 6000 10830 6200 10840
rect 6000 10810 6010 10830
rect 6030 10810 6090 10830
rect 6110 10810 6170 10830
rect 6190 10810 6200 10830
rect 6000 10800 6200 10810
rect 4240 10750 4440 10760
rect 4240 10730 4250 10750
rect 4270 10730 4330 10750
rect 4350 10730 4410 10750
rect 4430 10730 4440 10750
rect 4240 10720 4440 10730
rect 4480 10750 4680 10760
rect 4480 10730 4490 10750
rect 4510 10730 4570 10750
rect 4590 10730 4650 10750
rect 4670 10730 4680 10750
rect 4480 10720 4680 10730
rect 4720 10750 5720 10760
rect 4720 10730 4730 10750
rect 4750 10730 4810 10750
rect 4830 10730 4890 10750
rect 4910 10730 4970 10750
rect 4990 10730 5050 10750
rect 5070 10730 5130 10750
rect 5150 10730 5210 10750
rect 5230 10730 5290 10750
rect 5310 10730 5370 10750
rect 5390 10730 5450 10750
rect 5470 10730 5530 10750
rect 5550 10730 5610 10750
rect 5630 10730 5690 10750
rect 5710 10730 5720 10750
rect 4720 10720 5720 10730
rect 5760 10750 5960 10760
rect 5760 10730 5770 10750
rect 5790 10730 5850 10750
rect 5870 10730 5930 10750
rect 5950 10730 5960 10750
rect 5760 10720 5960 10730
rect 6000 10750 6200 10760
rect 6000 10730 6010 10750
rect 6030 10730 6090 10750
rect 6110 10730 6170 10750
rect 6190 10730 6200 10750
rect 6000 10720 6200 10730
rect 4240 10670 4440 10680
rect 4240 10650 4250 10670
rect 4270 10650 4330 10670
rect 4350 10650 4410 10670
rect 4430 10650 4440 10670
rect 4240 10640 4440 10650
rect 4480 10670 4680 10680
rect 4480 10650 4490 10670
rect 4510 10650 4570 10670
rect 4590 10650 4650 10670
rect 4670 10650 4680 10670
rect 4480 10640 4680 10650
rect 4720 10670 5720 10680
rect 4720 10650 4730 10670
rect 4750 10650 4810 10670
rect 4830 10650 4890 10670
rect 4910 10650 4970 10670
rect 4990 10650 5050 10670
rect 5070 10650 5130 10670
rect 5150 10650 5210 10670
rect 5230 10650 5290 10670
rect 5310 10650 5370 10670
rect 5390 10650 5450 10670
rect 5470 10650 5530 10670
rect 5550 10650 5610 10670
rect 5630 10650 5690 10670
rect 5710 10650 5720 10670
rect 4720 10640 5720 10650
rect 5760 10670 5960 10680
rect 5760 10650 5770 10670
rect 5790 10650 5850 10670
rect 5870 10650 5930 10670
rect 5950 10650 5960 10670
rect 5760 10640 5960 10650
rect 6000 10670 6200 10680
rect 6000 10650 6010 10670
rect 6030 10650 6090 10670
rect 6110 10650 6170 10670
rect 6190 10650 6200 10670
rect 6000 10640 6200 10650
rect 4240 10590 4440 10600
rect 4240 10570 4250 10590
rect 4270 10570 4330 10590
rect 4350 10570 4410 10590
rect 4430 10570 4440 10590
rect 4240 10560 4440 10570
rect 4480 10590 4680 10600
rect 4480 10570 4490 10590
rect 4510 10570 4570 10590
rect 4590 10570 4650 10590
rect 4670 10570 4680 10590
rect 4480 10560 4680 10570
rect 4720 10590 5720 10600
rect 4720 10570 4730 10590
rect 4750 10570 4810 10590
rect 4830 10570 4890 10590
rect 4910 10570 4970 10590
rect 4990 10570 5050 10590
rect 5070 10570 5130 10590
rect 5150 10570 5210 10590
rect 5230 10570 5290 10590
rect 5310 10570 5370 10590
rect 5390 10570 5450 10590
rect 5470 10570 5530 10590
rect 5550 10570 5610 10590
rect 5630 10570 5690 10590
rect 5710 10570 5720 10590
rect 4720 10560 5720 10570
rect 5760 10590 5960 10600
rect 5760 10570 5770 10590
rect 5790 10570 5850 10590
rect 5870 10570 5930 10590
rect 5950 10570 5960 10590
rect 5760 10560 5960 10570
rect 6000 10590 6200 10600
rect 6000 10570 6010 10590
rect 6030 10570 6090 10590
rect 6110 10570 6170 10590
rect 6190 10570 6200 10590
rect 6000 10560 6200 10570
rect 4240 10510 4440 10520
rect 4240 10490 4250 10510
rect 4270 10490 4330 10510
rect 4350 10490 4410 10510
rect 4430 10490 4440 10510
rect 4240 10480 4440 10490
rect 4480 10510 4680 10520
rect 4480 10490 4490 10510
rect 4510 10490 4570 10510
rect 4590 10490 4650 10510
rect 4670 10490 4680 10510
rect 4480 10480 4680 10490
rect 4720 10510 5720 10520
rect 4720 10490 4730 10510
rect 4750 10490 4810 10510
rect 4830 10490 4890 10510
rect 4910 10490 4970 10510
rect 4990 10490 5050 10510
rect 5070 10490 5130 10510
rect 5150 10490 5210 10510
rect 5230 10490 5290 10510
rect 5310 10490 5370 10510
rect 5390 10490 5450 10510
rect 5470 10490 5530 10510
rect 5550 10490 5610 10510
rect 5630 10490 5690 10510
rect 5710 10490 5720 10510
rect 4720 10480 5720 10490
rect 5760 10510 5960 10520
rect 5760 10490 5770 10510
rect 5790 10490 5850 10510
rect 5870 10490 5930 10510
rect 5950 10490 5960 10510
rect 5760 10480 5960 10490
rect 6000 10510 6200 10520
rect 6000 10490 6010 10510
rect 6030 10490 6090 10510
rect 6110 10490 6170 10510
rect 6190 10490 6200 10510
rect 6000 10480 6200 10490
rect 4240 10430 4440 10440
rect 4240 10410 4250 10430
rect 4270 10410 4330 10430
rect 4350 10410 4410 10430
rect 4430 10410 4440 10430
rect 4240 10400 4440 10410
rect 4480 10430 4680 10440
rect 4480 10410 4490 10430
rect 4510 10410 4570 10430
rect 4590 10410 4650 10430
rect 4670 10410 4680 10430
rect 4480 10400 4680 10410
rect 4720 10430 5720 10440
rect 4720 10410 4730 10430
rect 4750 10410 4810 10430
rect 4830 10410 4890 10430
rect 4910 10410 4970 10430
rect 4990 10410 5050 10430
rect 5070 10410 5130 10430
rect 5150 10410 5210 10430
rect 5230 10410 5290 10430
rect 5310 10410 5370 10430
rect 5390 10410 5450 10430
rect 5470 10410 5530 10430
rect 5550 10410 5610 10430
rect 5630 10410 5690 10430
rect 5710 10410 5720 10430
rect 4720 10400 5720 10410
rect 5760 10430 5960 10440
rect 5760 10410 5770 10430
rect 5790 10410 5850 10430
rect 5870 10410 5930 10430
rect 5950 10410 5960 10430
rect 5760 10400 5960 10410
rect 6000 10430 6200 10440
rect 6000 10410 6010 10430
rect 6030 10410 6090 10430
rect 6110 10410 6170 10430
rect 6190 10410 6200 10430
rect 6000 10400 6200 10410
rect 4240 10350 4440 10360
rect 4240 10330 4250 10350
rect 4270 10330 4330 10350
rect 4350 10330 4410 10350
rect 4430 10330 4440 10350
rect 4240 10320 4440 10330
rect 4480 10350 4680 10360
rect 4480 10330 4490 10350
rect 4510 10330 4570 10350
rect 4590 10330 4650 10350
rect 4670 10330 4680 10350
rect 4480 10320 4680 10330
rect 4720 10350 5720 10360
rect 4720 10330 4730 10350
rect 4750 10330 4810 10350
rect 4830 10330 4890 10350
rect 4910 10330 4970 10350
rect 4990 10330 5050 10350
rect 5070 10330 5130 10350
rect 5150 10330 5210 10350
rect 5230 10330 5290 10350
rect 5310 10330 5370 10350
rect 5390 10330 5450 10350
rect 5470 10330 5530 10350
rect 5550 10330 5610 10350
rect 5630 10330 5690 10350
rect 5710 10330 5720 10350
rect 4720 10320 5720 10330
rect 5760 10350 5960 10360
rect 5760 10330 5770 10350
rect 5790 10330 5850 10350
rect 5870 10330 5930 10350
rect 5950 10330 5960 10350
rect 5760 10320 5960 10330
rect 6000 10350 6200 10360
rect 6000 10330 6010 10350
rect 6030 10330 6090 10350
rect 6110 10330 6170 10350
rect 6190 10330 6200 10350
rect 6000 10320 6200 10330
rect 4240 10270 4440 10280
rect 4240 10250 4250 10270
rect 4270 10250 4330 10270
rect 4350 10250 4410 10270
rect 4430 10250 4440 10270
rect 4240 10240 4440 10250
rect 4480 10270 4680 10280
rect 4480 10250 4490 10270
rect 4510 10250 4570 10270
rect 4590 10250 4650 10270
rect 4670 10250 4680 10270
rect 4480 10240 4680 10250
rect 4720 10270 5720 10280
rect 4720 10250 4730 10270
rect 4750 10250 4810 10270
rect 4830 10250 4890 10270
rect 4910 10250 4970 10270
rect 4990 10250 5050 10270
rect 5070 10250 5130 10270
rect 5150 10250 5210 10270
rect 5230 10250 5290 10270
rect 5310 10250 5370 10270
rect 5390 10250 5450 10270
rect 5470 10250 5530 10270
rect 5550 10250 5610 10270
rect 5630 10250 5690 10270
rect 5710 10250 5720 10270
rect 4720 10240 5720 10250
rect 5760 10270 5960 10280
rect 5760 10250 5770 10270
rect 5790 10250 5850 10270
rect 5870 10250 5930 10270
rect 5950 10250 5960 10270
rect 5760 10240 5960 10250
rect 6000 10270 6200 10280
rect 6000 10250 6010 10270
rect 6030 10250 6090 10270
rect 6110 10250 6170 10270
rect 6190 10250 6200 10270
rect 6000 10240 6200 10250
rect 4240 10190 4440 10200
rect 4240 10170 4250 10190
rect 4270 10170 4330 10190
rect 4350 10170 4410 10190
rect 4430 10170 4440 10190
rect 4240 10160 4440 10170
rect 4480 10190 4680 10200
rect 4480 10170 4490 10190
rect 4510 10170 4570 10190
rect 4590 10170 4650 10190
rect 4670 10170 4680 10190
rect 4480 10160 4680 10170
rect 4720 10190 5720 10200
rect 4720 10170 4730 10190
rect 4750 10170 4810 10190
rect 4830 10170 4890 10190
rect 4910 10170 4970 10190
rect 4990 10170 5050 10190
rect 5070 10170 5130 10190
rect 5150 10170 5210 10190
rect 5230 10170 5290 10190
rect 5310 10170 5370 10190
rect 5390 10170 5450 10190
rect 5470 10170 5530 10190
rect 5550 10170 5610 10190
rect 5630 10170 5690 10190
rect 5710 10170 5720 10190
rect 4720 10160 5720 10170
rect 5760 10190 5960 10200
rect 5760 10170 5770 10190
rect 5790 10170 5850 10190
rect 5870 10170 5930 10190
rect 5950 10170 5960 10190
rect 5760 10160 5960 10170
rect 6000 10190 6200 10200
rect 6000 10170 6010 10190
rect 6030 10170 6090 10190
rect 6110 10170 6170 10190
rect 6190 10170 6200 10190
rect 6000 10160 6200 10170
rect 4240 10110 4440 10120
rect 4240 10090 4250 10110
rect 4270 10090 4330 10110
rect 4350 10090 4410 10110
rect 4430 10090 4440 10110
rect 4240 10080 4440 10090
rect 4480 10110 4680 10120
rect 4480 10090 4490 10110
rect 4510 10090 4570 10110
rect 4590 10090 4650 10110
rect 4670 10090 4680 10110
rect 4480 10080 4680 10090
rect 4720 10110 5720 10120
rect 4720 10090 4730 10110
rect 4750 10090 4810 10110
rect 4830 10090 4890 10110
rect 4910 10090 4970 10110
rect 4990 10090 5050 10110
rect 5070 10090 5130 10110
rect 5150 10090 5210 10110
rect 5230 10090 5290 10110
rect 5310 10090 5370 10110
rect 5390 10090 5450 10110
rect 5470 10090 5530 10110
rect 5550 10090 5610 10110
rect 5630 10090 5690 10110
rect 5710 10090 5720 10110
rect 4720 10080 5720 10090
rect 5760 10110 5960 10120
rect 5760 10090 5770 10110
rect 5790 10090 5850 10110
rect 5870 10090 5930 10110
rect 5950 10090 5960 10110
rect 5760 10080 5960 10090
rect 6000 10110 6200 10120
rect 6000 10090 6010 10110
rect 6030 10090 6090 10110
rect 6110 10090 6170 10110
rect 6190 10090 6200 10110
rect 6000 10080 6200 10090
rect 4240 10030 4440 10040
rect 4240 10010 4250 10030
rect 4270 10010 4330 10030
rect 4350 10010 4410 10030
rect 4430 10010 4440 10030
rect 4240 10000 4440 10010
rect 4480 10030 4680 10040
rect 4480 10010 4490 10030
rect 4510 10010 4570 10030
rect 4590 10010 4650 10030
rect 4670 10010 4680 10030
rect 4480 10000 4680 10010
rect 4720 10030 5720 10040
rect 4720 10010 4730 10030
rect 4750 10010 4810 10030
rect 4830 10010 4890 10030
rect 4910 10010 4970 10030
rect 4990 10010 5050 10030
rect 5070 10010 5130 10030
rect 5150 10010 5210 10030
rect 5230 10010 5290 10030
rect 5310 10010 5370 10030
rect 5390 10010 5450 10030
rect 5470 10010 5530 10030
rect 5550 10010 5610 10030
rect 5630 10010 5690 10030
rect 5710 10010 5720 10030
rect 4720 10000 5720 10010
rect 5760 10030 5960 10040
rect 5760 10010 5770 10030
rect 5790 10010 5850 10030
rect 5870 10010 5930 10030
rect 5950 10010 5960 10030
rect 5760 10000 5960 10010
rect 6000 10030 6200 10040
rect 6000 10010 6010 10030
rect 6030 10010 6090 10030
rect 6110 10010 6170 10030
rect 6190 10010 6200 10030
rect 6000 10000 6200 10010
rect 4240 9950 4440 9960
rect 4240 9930 4250 9950
rect 4270 9930 4330 9950
rect 4350 9930 4410 9950
rect 4430 9930 4440 9950
rect 4240 9920 4440 9930
rect 4480 9950 4680 9960
rect 4480 9930 4490 9950
rect 4510 9930 4570 9950
rect 4590 9930 4650 9950
rect 4670 9930 4680 9950
rect 4480 9920 4680 9930
rect 4720 9950 5720 9960
rect 4720 9930 4730 9950
rect 4750 9930 4810 9950
rect 4830 9930 4890 9950
rect 4910 9930 4970 9950
rect 4990 9930 5050 9950
rect 5070 9930 5130 9950
rect 5150 9930 5210 9950
rect 5230 9930 5290 9950
rect 5310 9930 5370 9950
rect 5390 9930 5450 9950
rect 5470 9930 5530 9950
rect 5550 9930 5610 9950
rect 5630 9930 5690 9950
rect 5710 9930 5720 9950
rect 4720 9920 5720 9930
rect 5760 9950 5960 9960
rect 5760 9930 5770 9950
rect 5790 9930 5850 9950
rect 5870 9930 5930 9950
rect 5950 9930 5960 9950
rect 5760 9920 5960 9930
rect 6000 9950 6200 9960
rect 6000 9930 6010 9950
rect 6030 9930 6090 9950
rect 6110 9930 6170 9950
rect 6190 9930 6200 9950
rect 6000 9920 6200 9930
rect 4240 9870 4440 9880
rect 4240 9850 4250 9870
rect 4270 9850 4330 9870
rect 4350 9850 4410 9870
rect 4430 9850 4440 9870
rect 4240 9840 4440 9850
rect 4480 9870 4680 9880
rect 4480 9850 4490 9870
rect 4510 9850 4570 9870
rect 4590 9850 4650 9870
rect 4670 9850 4680 9870
rect 4480 9840 4680 9850
rect 4720 9870 5720 9880
rect 4720 9850 4730 9870
rect 4750 9850 4810 9870
rect 4830 9850 4890 9870
rect 4910 9850 4970 9870
rect 4990 9850 5050 9870
rect 5070 9850 5130 9870
rect 5150 9850 5210 9870
rect 5230 9850 5290 9870
rect 5310 9850 5370 9870
rect 5390 9850 5450 9870
rect 5470 9850 5530 9870
rect 5550 9850 5610 9870
rect 5630 9850 5690 9870
rect 5710 9850 5720 9870
rect 4720 9840 5720 9850
rect 5760 9870 5960 9880
rect 5760 9850 5770 9870
rect 5790 9850 5850 9870
rect 5870 9850 5930 9870
rect 5950 9850 5960 9870
rect 5760 9840 5960 9850
rect 6000 9870 6200 9880
rect 6000 9850 6010 9870
rect 6030 9850 6090 9870
rect 6110 9850 6170 9870
rect 6190 9850 6200 9870
rect 6000 9840 6200 9850
rect 4240 9790 4440 9800
rect 4240 9770 4250 9790
rect 4270 9770 4330 9790
rect 4350 9770 4410 9790
rect 4430 9770 4440 9790
rect 4240 9760 4440 9770
rect 4480 9790 4680 9800
rect 4480 9770 4490 9790
rect 4510 9770 4570 9790
rect 4590 9770 4650 9790
rect 4670 9770 4680 9790
rect 4480 9760 4680 9770
rect 4720 9790 5720 9800
rect 4720 9770 4730 9790
rect 4750 9770 4810 9790
rect 4830 9770 4890 9790
rect 4910 9770 4970 9790
rect 4990 9770 5050 9790
rect 5070 9770 5130 9790
rect 5150 9770 5210 9790
rect 5230 9770 5290 9790
rect 5310 9770 5370 9790
rect 5390 9770 5450 9790
rect 5470 9770 5530 9790
rect 5550 9770 5610 9790
rect 5630 9770 5690 9790
rect 5710 9770 5720 9790
rect 4720 9760 5720 9770
rect 5760 9790 5960 9800
rect 5760 9770 5770 9790
rect 5790 9770 5850 9790
rect 5870 9770 5930 9790
rect 5950 9770 5960 9790
rect 5760 9760 5960 9770
rect 6000 9790 6200 9800
rect 6000 9770 6010 9790
rect 6030 9770 6090 9790
rect 6110 9770 6170 9790
rect 6190 9770 6200 9790
rect 6000 9760 6200 9770
rect 4240 9710 4440 9720
rect 4240 9690 4250 9710
rect 4270 9690 4330 9710
rect 4350 9690 4410 9710
rect 4430 9690 4440 9710
rect 4240 9680 4440 9690
rect 4480 9710 4680 9720
rect 4480 9690 4490 9710
rect 4510 9690 4570 9710
rect 4590 9690 4650 9710
rect 4670 9690 4680 9710
rect 4480 9680 4680 9690
rect 4720 9710 5720 9720
rect 4720 9690 4730 9710
rect 4750 9690 4810 9710
rect 4830 9690 4890 9710
rect 4910 9690 4970 9710
rect 4990 9690 5050 9710
rect 5070 9690 5130 9710
rect 5150 9690 5210 9710
rect 5230 9690 5290 9710
rect 5310 9690 5370 9710
rect 5390 9690 5450 9710
rect 5470 9690 5530 9710
rect 5550 9690 5610 9710
rect 5630 9690 5690 9710
rect 5710 9690 5720 9710
rect 4720 9680 5720 9690
rect 5760 9710 5960 9720
rect 5760 9690 5770 9710
rect 5790 9690 5850 9710
rect 5870 9690 5930 9710
rect 5950 9690 5960 9710
rect 5760 9680 5960 9690
rect 6000 9710 6200 9720
rect 6000 9690 6010 9710
rect 6030 9690 6090 9710
rect 6110 9690 6170 9710
rect 6190 9690 6200 9710
rect 6000 9680 6200 9690
rect 4240 9630 4440 9640
rect 4240 9610 4250 9630
rect 4270 9610 4330 9630
rect 4350 9610 4410 9630
rect 4430 9610 4440 9630
rect 4240 9600 4440 9610
rect 4480 9630 4680 9640
rect 4480 9610 4490 9630
rect 4510 9610 4570 9630
rect 4590 9610 4650 9630
rect 4670 9610 4680 9630
rect 4480 9600 4680 9610
rect 4720 9630 5720 9640
rect 4720 9610 4730 9630
rect 4750 9610 4810 9630
rect 4830 9610 4890 9630
rect 4910 9610 4970 9630
rect 4990 9610 5050 9630
rect 5070 9610 5130 9630
rect 5150 9610 5210 9630
rect 5230 9610 5290 9630
rect 5310 9610 5370 9630
rect 5390 9610 5450 9630
rect 5470 9610 5530 9630
rect 5550 9610 5610 9630
rect 5630 9610 5690 9630
rect 5710 9610 5720 9630
rect 4720 9600 5720 9610
rect 5760 9630 5960 9640
rect 5760 9610 5770 9630
rect 5790 9610 5850 9630
rect 5870 9610 5930 9630
rect 5950 9610 5960 9630
rect 5760 9600 5960 9610
rect 6000 9630 6200 9640
rect 6000 9610 6010 9630
rect 6030 9610 6090 9630
rect 6110 9610 6170 9630
rect 6190 9610 6200 9630
rect 6000 9600 6200 9610
rect 4240 9550 4440 9560
rect 4240 9530 4250 9550
rect 4270 9530 4330 9550
rect 4350 9530 4410 9550
rect 4430 9530 4440 9550
rect 4240 9520 4440 9530
rect 4480 9550 4680 9560
rect 4480 9530 4490 9550
rect 4510 9530 4570 9550
rect 4590 9530 4650 9550
rect 4670 9530 4680 9550
rect 4480 9520 4680 9530
rect 4720 9550 5720 9560
rect 4720 9530 4730 9550
rect 4750 9530 4810 9550
rect 4830 9530 4890 9550
rect 4910 9530 4970 9550
rect 4990 9530 5050 9550
rect 5070 9530 5130 9550
rect 5150 9530 5210 9550
rect 5230 9530 5290 9550
rect 5310 9530 5370 9550
rect 5390 9530 5450 9550
rect 5470 9530 5530 9550
rect 5550 9530 5610 9550
rect 5630 9530 5690 9550
rect 5710 9530 5720 9550
rect 4720 9520 5720 9530
rect 5760 9550 5960 9560
rect 5760 9530 5770 9550
rect 5790 9530 5850 9550
rect 5870 9530 5930 9550
rect 5950 9530 5960 9550
rect 5760 9520 5960 9530
rect 6000 9550 6200 9560
rect 6000 9530 6010 9550
rect 6030 9530 6090 9550
rect 6110 9530 6170 9550
rect 6190 9530 6200 9550
rect 6000 9520 6200 9530
rect 4240 9470 4440 9480
rect 4240 9450 4250 9470
rect 4270 9450 4330 9470
rect 4350 9450 4410 9470
rect 4430 9450 4440 9470
rect 4240 9440 4440 9450
rect 4480 9470 4680 9480
rect 4480 9450 4490 9470
rect 4510 9450 4570 9470
rect 4590 9450 4650 9470
rect 4670 9450 4680 9470
rect 4480 9440 4680 9450
rect 4720 9470 5720 9480
rect 4720 9450 4730 9470
rect 4750 9450 4810 9470
rect 4830 9450 4890 9470
rect 4910 9450 4970 9470
rect 4990 9450 5050 9470
rect 5070 9450 5130 9470
rect 5150 9450 5210 9470
rect 5230 9450 5290 9470
rect 5310 9450 5370 9470
rect 5390 9450 5450 9470
rect 5470 9450 5530 9470
rect 5550 9450 5610 9470
rect 5630 9450 5690 9470
rect 5710 9450 5720 9470
rect 4720 9440 5720 9450
rect 5760 9470 5960 9480
rect 5760 9450 5770 9470
rect 5790 9450 5850 9470
rect 5870 9450 5930 9470
rect 5950 9450 5960 9470
rect 5760 9440 5960 9450
rect 6000 9470 6200 9480
rect 6000 9450 6010 9470
rect 6030 9450 6090 9470
rect 6110 9450 6170 9470
rect 6190 9450 6200 9470
rect 6000 9440 6200 9450
rect 4240 9390 4440 9400
rect 4240 9370 4250 9390
rect 4270 9370 4330 9390
rect 4350 9370 4410 9390
rect 4430 9370 4440 9390
rect 4240 9360 4440 9370
rect 4480 9390 4680 9400
rect 4480 9370 4490 9390
rect 4510 9370 4570 9390
rect 4590 9370 4650 9390
rect 4670 9370 4680 9390
rect 4480 9360 4680 9370
rect 4720 9390 5720 9400
rect 4720 9370 4730 9390
rect 4750 9370 4810 9390
rect 4830 9370 4890 9390
rect 4910 9370 4970 9390
rect 4990 9370 5050 9390
rect 5070 9370 5130 9390
rect 5150 9370 5210 9390
rect 5230 9370 5290 9390
rect 5310 9370 5370 9390
rect 5390 9370 5450 9390
rect 5470 9370 5530 9390
rect 5550 9370 5610 9390
rect 5630 9370 5690 9390
rect 5710 9370 5720 9390
rect 4720 9360 5720 9370
rect 5760 9390 5960 9400
rect 5760 9370 5770 9390
rect 5790 9370 5850 9390
rect 5870 9370 5930 9390
rect 5950 9370 5960 9390
rect 5760 9360 5960 9370
rect 6000 9390 6200 9400
rect 6000 9370 6010 9390
rect 6030 9370 6090 9390
rect 6110 9370 6170 9390
rect 6190 9370 6200 9390
rect 6000 9360 6200 9370
rect 4240 9310 4440 9320
rect 4240 9290 4250 9310
rect 4270 9290 4330 9310
rect 4350 9290 4410 9310
rect 4430 9290 4440 9310
rect 4240 9280 4440 9290
rect 4480 9310 4680 9320
rect 4480 9290 4490 9310
rect 4510 9290 4570 9310
rect 4590 9290 4650 9310
rect 4670 9290 4680 9310
rect 4480 9280 4680 9290
rect 4720 9310 5720 9320
rect 4720 9290 4730 9310
rect 4750 9290 4810 9310
rect 4830 9290 4890 9310
rect 4910 9290 4970 9310
rect 4990 9290 5050 9310
rect 5070 9290 5130 9310
rect 5150 9290 5210 9310
rect 5230 9290 5290 9310
rect 5310 9290 5370 9310
rect 5390 9290 5450 9310
rect 5470 9290 5530 9310
rect 5550 9290 5610 9310
rect 5630 9290 5690 9310
rect 5710 9290 5720 9310
rect 4720 9280 5720 9290
rect 5760 9310 5960 9320
rect 5760 9290 5770 9310
rect 5790 9290 5850 9310
rect 5870 9290 5930 9310
rect 5950 9290 5960 9310
rect 5760 9280 5960 9290
rect 6000 9310 6200 9320
rect 6000 9290 6010 9310
rect 6030 9290 6090 9310
rect 6110 9290 6170 9310
rect 6190 9290 6200 9310
rect 6000 9280 6200 9290
rect 4240 9230 4440 9240
rect 4240 9210 4250 9230
rect 4270 9210 4330 9230
rect 4350 9210 4410 9230
rect 4430 9210 4440 9230
rect 4240 9200 4440 9210
rect 4480 9230 4680 9240
rect 4480 9210 4490 9230
rect 4510 9210 4570 9230
rect 4590 9210 4650 9230
rect 4670 9210 4680 9230
rect 4480 9200 4680 9210
rect 4720 9230 5720 9240
rect 4720 9210 4730 9230
rect 4750 9210 4810 9230
rect 4830 9210 4890 9230
rect 4910 9210 4970 9230
rect 4990 9210 5050 9230
rect 5070 9210 5130 9230
rect 5150 9210 5210 9230
rect 5230 9210 5290 9230
rect 5310 9210 5370 9230
rect 5390 9210 5450 9230
rect 5470 9210 5530 9230
rect 5550 9210 5610 9230
rect 5630 9210 5690 9230
rect 5710 9210 5720 9230
rect 4720 9200 5720 9210
rect 5760 9230 5960 9240
rect 5760 9210 5770 9230
rect 5790 9210 5850 9230
rect 5870 9210 5930 9230
rect 5950 9210 5960 9230
rect 5760 9200 5960 9210
rect 6000 9230 6200 9240
rect 6000 9210 6010 9230
rect 6030 9210 6090 9230
rect 6110 9210 6170 9230
rect 6190 9210 6200 9230
rect 6000 9200 6200 9210
rect 4240 9150 4440 9160
rect 4240 9130 4250 9150
rect 4270 9130 4330 9150
rect 4350 9130 4410 9150
rect 4430 9130 4440 9150
rect 4240 9120 4440 9130
rect 4480 9150 4680 9160
rect 4480 9130 4490 9150
rect 4510 9130 4570 9150
rect 4590 9130 4650 9150
rect 4670 9130 4680 9150
rect 4480 9120 4680 9130
rect 4720 9150 5720 9160
rect 4720 9130 4730 9150
rect 4750 9130 4810 9150
rect 4830 9130 4890 9150
rect 4910 9130 4970 9150
rect 4990 9130 5050 9150
rect 5070 9130 5130 9150
rect 5150 9130 5210 9150
rect 5230 9130 5290 9150
rect 5310 9130 5370 9150
rect 5390 9130 5450 9150
rect 5470 9130 5530 9150
rect 5550 9130 5610 9150
rect 5630 9130 5690 9150
rect 5710 9130 5720 9150
rect 4720 9120 5720 9130
rect 5760 9150 5960 9160
rect 5760 9130 5770 9150
rect 5790 9130 5850 9150
rect 5870 9130 5930 9150
rect 5950 9130 5960 9150
rect 5760 9120 5960 9130
rect 6000 9150 6200 9160
rect 6000 9130 6010 9150
rect 6030 9130 6090 9150
rect 6110 9130 6170 9150
rect 6190 9130 6200 9150
rect 6000 9120 6200 9130
rect 4240 9070 4440 9080
rect 4240 9050 4250 9070
rect 4270 9050 4330 9070
rect 4350 9050 4410 9070
rect 4430 9050 4440 9070
rect 4240 9040 4440 9050
rect 4480 9070 4680 9080
rect 4480 9050 4490 9070
rect 4510 9050 4570 9070
rect 4590 9050 4650 9070
rect 4670 9050 4680 9070
rect 4480 9040 4680 9050
rect 4720 9070 5720 9080
rect 4720 9050 4730 9070
rect 4750 9050 4810 9070
rect 4830 9050 4890 9070
rect 4910 9050 4970 9070
rect 4990 9050 5050 9070
rect 5070 9050 5130 9070
rect 5150 9050 5210 9070
rect 5230 9050 5290 9070
rect 5310 9050 5370 9070
rect 5390 9050 5450 9070
rect 5470 9050 5530 9070
rect 5550 9050 5610 9070
rect 5630 9050 5690 9070
rect 5710 9050 5720 9070
rect 4720 9040 5720 9050
rect 5760 9070 5960 9080
rect 5760 9050 5770 9070
rect 5790 9050 5850 9070
rect 5870 9050 5930 9070
rect 5950 9050 5960 9070
rect 5760 9040 5960 9050
rect 6000 9070 6200 9080
rect 6000 9050 6010 9070
rect 6030 9050 6090 9070
rect 6110 9050 6170 9070
rect 6190 9050 6200 9070
rect 6000 9040 6200 9050
rect 4240 8990 4440 9000
rect 4240 8970 4250 8990
rect 4270 8970 4330 8990
rect 4350 8970 4410 8990
rect 4430 8970 4440 8990
rect 4240 8960 4440 8970
rect 4480 8990 4680 9000
rect 4480 8970 4490 8990
rect 4510 8970 4570 8990
rect 4590 8970 4650 8990
rect 4670 8970 4680 8990
rect 4480 8960 4680 8970
rect 4720 8990 5720 9000
rect 4720 8970 4730 8990
rect 4750 8970 4810 8990
rect 4830 8970 4890 8990
rect 4910 8970 4970 8990
rect 4990 8970 5050 8990
rect 5070 8970 5130 8990
rect 5150 8970 5210 8990
rect 5230 8970 5290 8990
rect 5310 8970 5370 8990
rect 5390 8970 5450 8990
rect 5470 8970 5530 8990
rect 5550 8970 5610 8990
rect 5630 8970 5690 8990
rect 5710 8970 5720 8990
rect 4720 8960 5720 8970
rect 5760 8990 5960 9000
rect 5760 8970 5770 8990
rect 5790 8970 5850 8990
rect 5870 8970 5930 8990
rect 5950 8970 5960 8990
rect 5760 8960 5960 8970
rect 6000 8990 6200 9000
rect 6000 8970 6010 8990
rect 6030 8970 6090 8990
rect 6110 8970 6170 8990
rect 6190 8970 6200 8990
rect 6000 8960 6200 8970
rect 4240 8910 4440 8920
rect 4240 8890 4250 8910
rect 4270 8890 4330 8910
rect 4350 8890 4410 8910
rect 4430 8890 4440 8910
rect 4240 8880 4440 8890
rect 4480 8910 4680 8920
rect 4480 8890 4490 8910
rect 4510 8890 4570 8910
rect 4590 8890 4650 8910
rect 4670 8890 4680 8910
rect 4480 8880 4680 8890
rect 4720 8910 5720 8920
rect 4720 8890 4730 8910
rect 4750 8890 4810 8910
rect 4830 8890 4890 8910
rect 4910 8890 4970 8910
rect 4990 8890 5050 8910
rect 5070 8890 5130 8910
rect 5150 8890 5210 8910
rect 5230 8890 5290 8910
rect 5310 8890 5370 8910
rect 5390 8890 5450 8910
rect 5470 8890 5530 8910
rect 5550 8890 5610 8910
rect 5630 8890 5690 8910
rect 5710 8890 5720 8910
rect 4720 8880 5720 8890
rect 5760 8910 5960 8920
rect 5760 8890 5770 8910
rect 5790 8890 5850 8910
rect 5870 8890 5930 8910
rect 5950 8890 5960 8910
rect 5760 8880 5960 8890
rect 6000 8910 6200 8920
rect 6000 8890 6010 8910
rect 6030 8890 6090 8910
rect 6110 8890 6170 8910
rect 6190 8890 6200 8910
rect 6000 8880 6200 8890
rect 4240 8830 4440 8840
rect 4240 8810 4250 8830
rect 4270 8810 4330 8830
rect 4350 8810 4410 8830
rect 4430 8810 4440 8830
rect 4240 8800 4440 8810
rect 4480 8830 4680 8840
rect 4480 8810 4490 8830
rect 4510 8810 4570 8830
rect 4590 8810 4650 8830
rect 4670 8810 4680 8830
rect 4480 8800 4680 8810
rect 4720 8830 5720 8840
rect 4720 8810 4730 8830
rect 4750 8810 4810 8830
rect 4830 8810 4890 8830
rect 4910 8810 4970 8830
rect 4990 8810 5050 8830
rect 5070 8810 5130 8830
rect 5150 8810 5210 8830
rect 5230 8810 5290 8830
rect 5310 8810 5370 8830
rect 5390 8810 5450 8830
rect 5470 8810 5530 8830
rect 5550 8810 5610 8830
rect 5630 8810 5690 8830
rect 5710 8810 5720 8830
rect 4720 8800 5720 8810
rect 5760 8830 5960 8840
rect 5760 8810 5770 8830
rect 5790 8810 5850 8830
rect 5870 8810 5930 8830
rect 5950 8810 5960 8830
rect 5760 8800 5960 8810
rect 6000 8830 6200 8840
rect 6000 8810 6010 8830
rect 6030 8810 6090 8830
rect 6110 8810 6170 8830
rect 6190 8810 6200 8830
rect 6000 8800 6200 8810
rect 4240 8750 4440 8760
rect 4240 8730 4250 8750
rect 4270 8730 4330 8750
rect 4350 8730 4410 8750
rect 4430 8730 4440 8750
rect 4240 8720 4440 8730
rect 4480 8750 4680 8760
rect 4480 8730 4490 8750
rect 4510 8730 4570 8750
rect 4590 8730 4650 8750
rect 4670 8730 4680 8750
rect 4480 8720 4680 8730
rect 4720 8750 5720 8760
rect 4720 8730 4730 8750
rect 4750 8730 4810 8750
rect 4830 8730 4890 8750
rect 4910 8730 4970 8750
rect 4990 8730 5050 8750
rect 5070 8730 5130 8750
rect 5150 8730 5210 8750
rect 5230 8730 5290 8750
rect 5310 8730 5370 8750
rect 5390 8730 5450 8750
rect 5470 8730 5530 8750
rect 5550 8730 5610 8750
rect 5630 8730 5690 8750
rect 5710 8730 5720 8750
rect 4720 8720 5720 8730
rect 5760 8750 5960 8760
rect 5760 8730 5770 8750
rect 5790 8730 5850 8750
rect 5870 8730 5930 8750
rect 5950 8730 5960 8750
rect 5760 8720 5960 8730
rect 6000 8750 6200 8760
rect 6000 8730 6010 8750
rect 6030 8730 6090 8750
rect 6110 8730 6170 8750
rect 6190 8730 6200 8750
rect 6000 8720 6200 8730
rect 4240 8670 4440 8680
rect 4240 8650 4250 8670
rect 4270 8650 4330 8670
rect 4350 8650 4410 8670
rect 4430 8650 4440 8670
rect 4240 8640 4440 8650
rect 4480 8670 4680 8680
rect 4480 8650 4490 8670
rect 4510 8650 4570 8670
rect 4590 8650 4650 8670
rect 4670 8650 4680 8670
rect 4480 8640 4680 8650
rect 4720 8670 5720 8680
rect 4720 8650 4730 8670
rect 4750 8650 4810 8670
rect 4830 8650 4890 8670
rect 4910 8650 4970 8670
rect 4990 8650 5050 8670
rect 5070 8650 5130 8670
rect 5150 8650 5210 8670
rect 5230 8650 5290 8670
rect 5310 8650 5370 8670
rect 5390 8650 5450 8670
rect 5470 8650 5530 8670
rect 5550 8650 5610 8670
rect 5630 8650 5690 8670
rect 5710 8650 5720 8670
rect 4720 8640 5720 8650
rect 5760 8670 5960 8680
rect 5760 8650 5770 8670
rect 5790 8650 5850 8670
rect 5870 8650 5930 8670
rect 5950 8650 5960 8670
rect 5760 8640 5960 8650
rect 6000 8670 6200 8680
rect 6000 8650 6010 8670
rect 6030 8650 6090 8670
rect 6110 8650 6170 8670
rect 6190 8650 6200 8670
rect 6000 8640 6200 8650
rect 4240 8590 4440 8600
rect 4240 8570 4250 8590
rect 4270 8570 4330 8590
rect 4350 8570 4410 8590
rect 4430 8570 4440 8590
rect 4240 8560 4440 8570
rect 4480 8590 4680 8600
rect 4480 8570 4490 8590
rect 4510 8570 4570 8590
rect 4590 8570 4650 8590
rect 4670 8570 4680 8590
rect 4480 8560 4680 8570
rect 4720 8590 5720 8600
rect 4720 8570 4730 8590
rect 4750 8570 4810 8590
rect 4830 8570 4890 8590
rect 4910 8570 4970 8590
rect 4990 8570 5050 8590
rect 5070 8570 5130 8590
rect 5150 8570 5210 8590
rect 5230 8570 5290 8590
rect 5310 8570 5370 8590
rect 5390 8570 5450 8590
rect 5470 8570 5530 8590
rect 5550 8570 5610 8590
rect 5630 8570 5690 8590
rect 5710 8570 5720 8590
rect 4720 8560 5720 8570
rect 5760 8590 5960 8600
rect 5760 8570 5770 8590
rect 5790 8570 5850 8590
rect 5870 8570 5930 8590
rect 5950 8570 5960 8590
rect 5760 8560 5960 8570
rect 6000 8590 6200 8600
rect 6000 8570 6010 8590
rect 6030 8570 6090 8590
rect 6110 8570 6170 8590
rect 6190 8570 6200 8590
rect 6000 8560 6200 8570
rect 4240 8510 4440 8520
rect 4240 8490 4250 8510
rect 4270 8490 4330 8510
rect 4350 8490 4410 8510
rect 4430 8490 4440 8510
rect 4240 8480 4440 8490
rect 4480 8510 4680 8520
rect 4480 8490 4490 8510
rect 4510 8490 4570 8510
rect 4590 8490 4650 8510
rect 4670 8490 4680 8510
rect 4480 8480 4680 8490
rect 4720 8510 5720 8520
rect 4720 8490 4730 8510
rect 4750 8490 4810 8510
rect 4830 8490 4890 8510
rect 4910 8490 4970 8510
rect 4990 8490 5050 8510
rect 5070 8490 5130 8510
rect 5150 8490 5210 8510
rect 5230 8490 5290 8510
rect 5310 8490 5370 8510
rect 5390 8490 5450 8510
rect 5470 8490 5530 8510
rect 5550 8490 5610 8510
rect 5630 8490 5690 8510
rect 5710 8490 5720 8510
rect 4720 8480 5720 8490
rect 5760 8510 5960 8520
rect 5760 8490 5770 8510
rect 5790 8490 5850 8510
rect 5870 8490 5930 8510
rect 5950 8490 5960 8510
rect 5760 8480 5960 8490
rect 6000 8510 6200 8520
rect 6000 8490 6010 8510
rect 6030 8490 6090 8510
rect 6110 8490 6170 8510
rect 6190 8490 6200 8510
rect 6000 8480 6200 8490
rect 4240 8430 4440 8440
rect 4240 8410 4250 8430
rect 4270 8410 4330 8430
rect 4350 8410 4410 8430
rect 4430 8410 4440 8430
rect 4240 8400 4440 8410
rect 4480 8430 4680 8440
rect 4480 8410 4490 8430
rect 4510 8410 4570 8430
rect 4590 8410 4650 8430
rect 4670 8410 4680 8430
rect 4480 8400 4680 8410
rect 4720 8430 5720 8440
rect 4720 8410 4730 8430
rect 4750 8410 4810 8430
rect 4830 8410 4890 8430
rect 4910 8410 4970 8430
rect 4990 8410 5050 8430
rect 5070 8410 5130 8430
rect 5150 8410 5210 8430
rect 5230 8410 5290 8430
rect 5310 8410 5370 8430
rect 5390 8410 5450 8430
rect 5470 8410 5530 8430
rect 5550 8410 5610 8430
rect 5630 8410 5690 8430
rect 5710 8410 5720 8430
rect 4720 8400 5720 8410
rect 5760 8430 5960 8440
rect 5760 8410 5770 8430
rect 5790 8410 5850 8430
rect 5870 8410 5930 8430
rect 5950 8410 5960 8430
rect 5760 8400 5960 8410
rect 6000 8430 6200 8440
rect 6000 8410 6010 8430
rect 6030 8410 6090 8430
rect 6110 8410 6170 8430
rect 6190 8410 6200 8430
rect 6000 8400 6200 8410
rect 4240 8350 4440 8360
rect 4240 8330 4250 8350
rect 4270 8330 4330 8350
rect 4350 8330 4410 8350
rect 4430 8330 4440 8350
rect 4240 8320 4440 8330
rect 4480 8350 4680 8360
rect 4480 8330 4490 8350
rect 4510 8330 4570 8350
rect 4590 8330 4650 8350
rect 4670 8330 4680 8350
rect 4480 8320 4680 8330
rect 4720 8350 5720 8360
rect 4720 8330 4730 8350
rect 4750 8330 4810 8350
rect 4830 8330 4890 8350
rect 4910 8330 4970 8350
rect 4990 8330 5050 8350
rect 5070 8330 5130 8350
rect 5150 8330 5210 8350
rect 5230 8330 5290 8350
rect 5310 8330 5370 8350
rect 5390 8330 5450 8350
rect 5470 8330 5530 8350
rect 5550 8330 5610 8350
rect 5630 8330 5690 8350
rect 5710 8330 5720 8350
rect 4720 8320 5720 8330
rect 5760 8350 5960 8360
rect 5760 8330 5770 8350
rect 5790 8330 5850 8350
rect 5870 8330 5930 8350
rect 5950 8330 5960 8350
rect 5760 8320 5960 8330
rect 6000 8350 6200 8360
rect 6000 8330 6010 8350
rect 6030 8330 6090 8350
rect 6110 8330 6170 8350
rect 6190 8330 6200 8350
rect 6000 8320 6200 8330
rect 4240 8270 4440 8280
rect 4240 8250 4250 8270
rect 4270 8250 4330 8270
rect 4350 8250 4410 8270
rect 4430 8250 4440 8270
rect 4240 8240 4440 8250
rect 4480 8270 4680 8280
rect 4480 8250 4490 8270
rect 4510 8250 4570 8270
rect 4590 8250 4650 8270
rect 4670 8250 4680 8270
rect 4480 8240 4680 8250
rect 4720 8270 5720 8280
rect 4720 8250 4730 8270
rect 4750 8250 4810 8270
rect 4830 8250 4890 8270
rect 4910 8250 4970 8270
rect 4990 8250 5050 8270
rect 5070 8250 5130 8270
rect 5150 8250 5210 8270
rect 5230 8250 5290 8270
rect 5310 8250 5370 8270
rect 5390 8250 5450 8270
rect 5470 8250 5530 8270
rect 5550 8250 5610 8270
rect 5630 8250 5690 8270
rect 5710 8250 5720 8270
rect 4720 8240 5720 8250
rect 5760 8270 5960 8280
rect 5760 8250 5770 8270
rect 5790 8250 5850 8270
rect 5870 8250 5930 8270
rect 5950 8250 5960 8270
rect 5760 8240 5960 8250
rect 6000 8270 6200 8280
rect 6000 8250 6010 8270
rect 6030 8250 6090 8270
rect 6110 8250 6170 8270
rect 6190 8250 6200 8270
rect 6000 8240 6200 8250
rect 4240 8190 4440 8200
rect 4240 8170 4250 8190
rect 4270 8170 4330 8190
rect 4350 8170 4410 8190
rect 4430 8170 4440 8190
rect 4240 8160 4440 8170
rect 4480 8190 4680 8200
rect 4480 8170 4490 8190
rect 4510 8170 4570 8190
rect 4590 8170 4650 8190
rect 4670 8170 4680 8190
rect 4480 8160 4680 8170
rect 4720 8190 5720 8200
rect 4720 8170 4730 8190
rect 4750 8170 4810 8190
rect 4830 8170 4890 8190
rect 4910 8170 4970 8190
rect 4990 8170 5050 8190
rect 5070 8170 5130 8190
rect 5150 8170 5210 8190
rect 5230 8170 5290 8190
rect 5310 8170 5370 8190
rect 5390 8170 5450 8190
rect 5470 8170 5530 8190
rect 5550 8170 5610 8190
rect 5630 8170 5690 8190
rect 5710 8170 5720 8190
rect 4720 8160 5720 8170
rect 5760 8190 5960 8200
rect 5760 8170 5770 8190
rect 5790 8170 5850 8190
rect 5870 8170 5930 8190
rect 5950 8170 5960 8190
rect 5760 8160 5960 8170
rect 6000 8190 6200 8200
rect 6000 8170 6010 8190
rect 6030 8170 6090 8190
rect 6110 8170 6170 8190
rect 6190 8170 6200 8190
rect 6000 8160 6200 8170
rect 4240 8110 4440 8120
rect 4240 8090 4250 8110
rect 4270 8090 4330 8110
rect 4350 8090 4410 8110
rect 4430 8090 4440 8110
rect 4240 8080 4440 8090
rect 4480 8110 4680 8120
rect 4480 8090 4490 8110
rect 4510 8090 4570 8110
rect 4590 8090 4650 8110
rect 4670 8090 4680 8110
rect 4480 8080 4680 8090
rect 4720 8110 5720 8120
rect 4720 8090 4730 8110
rect 4750 8090 4810 8110
rect 4830 8090 4890 8110
rect 4910 8090 4970 8110
rect 4990 8090 5050 8110
rect 5070 8090 5130 8110
rect 5150 8090 5210 8110
rect 5230 8090 5290 8110
rect 5310 8090 5370 8110
rect 5390 8090 5450 8110
rect 5470 8090 5530 8110
rect 5550 8090 5610 8110
rect 5630 8090 5690 8110
rect 5710 8090 5720 8110
rect 4720 8080 5720 8090
rect 5760 8110 5960 8120
rect 5760 8090 5770 8110
rect 5790 8090 5850 8110
rect 5870 8090 5930 8110
rect 5950 8090 5960 8110
rect 5760 8080 5960 8090
rect 6000 8110 6200 8120
rect 6000 8090 6010 8110
rect 6030 8090 6090 8110
rect 6110 8090 6170 8110
rect 6190 8090 6200 8110
rect 6000 8080 6200 8090
rect 4240 8030 4440 8040
rect 4240 8010 4250 8030
rect 4270 8010 4330 8030
rect 4350 8010 4410 8030
rect 4430 8010 4440 8030
rect 4240 8000 4440 8010
rect 4480 8030 4680 8040
rect 4480 8010 4490 8030
rect 4510 8010 4570 8030
rect 4590 8010 4650 8030
rect 4670 8010 4680 8030
rect 4480 8000 4680 8010
rect 4720 8030 5720 8040
rect 4720 8010 4730 8030
rect 4750 8010 4810 8030
rect 4830 8010 4890 8030
rect 4910 8010 4970 8030
rect 4990 8010 5050 8030
rect 5070 8010 5130 8030
rect 5150 8010 5210 8030
rect 5230 8010 5290 8030
rect 5310 8010 5370 8030
rect 5390 8010 5450 8030
rect 5470 8010 5530 8030
rect 5550 8010 5610 8030
rect 5630 8010 5690 8030
rect 5710 8010 5720 8030
rect 4720 8000 5720 8010
rect 5760 8030 5960 8040
rect 5760 8010 5770 8030
rect 5790 8010 5850 8030
rect 5870 8010 5930 8030
rect 5950 8010 5960 8030
rect 5760 8000 5960 8010
rect 6000 8030 6200 8040
rect 6000 8010 6010 8030
rect 6030 8010 6090 8030
rect 6110 8010 6170 8030
rect 6190 8010 6200 8030
rect 6000 8000 6200 8010
rect 4240 7950 4440 7960
rect 4240 7930 4250 7950
rect 4270 7930 4330 7950
rect 4350 7930 4410 7950
rect 4430 7930 4440 7950
rect 4240 7920 4440 7930
rect 4480 7950 4680 7960
rect 4480 7930 4490 7950
rect 4510 7930 4570 7950
rect 4590 7930 4650 7950
rect 4670 7930 4680 7950
rect 4480 7920 4680 7930
rect 4720 7950 5720 7960
rect 4720 7930 4730 7950
rect 4750 7930 4810 7950
rect 4830 7930 4890 7950
rect 4910 7930 4970 7950
rect 4990 7930 5050 7950
rect 5070 7930 5130 7950
rect 5150 7930 5210 7950
rect 5230 7930 5290 7950
rect 5310 7930 5370 7950
rect 5390 7930 5450 7950
rect 5470 7930 5530 7950
rect 5550 7930 5610 7950
rect 5630 7930 5690 7950
rect 5710 7930 5720 7950
rect 4720 7920 5720 7930
rect 5760 7950 5960 7960
rect 5760 7930 5770 7950
rect 5790 7930 5850 7950
rect 5870 7930 5930 7950
rect 5950 7930 5960 7950
rect 5760 7920 5960 7930
rect 6000 7950 6200 7960
rect 6000 7930 6010 7950
rect 6030 7930 6090 7950
rect 6110 7930 6170 7950
rect 6190 7930 6200 7950
rect 6000 7920 6200 7930
rect 4240 7870 4440 7880
rect 4240 7850 4250 7870
rect 4270 7850 4330 7870
rect 4350 7850 4410 7870
rect 4430 7850 4440 7870
rect 4240 7840 4440 7850
rect 4480 7870 4680 7880
rect 4480 7850 4490 7870
rect 4510 7850 4570 7870
rect 4590 7850 4650 7870
rect 4670 7850 4680 7870
rect 4480 7840 4680 7850
rect 4720 7870 5720 7880
rect 4720 7850 4730 7870
rect 4750 7850 4810 7870
rect 4830 7850 4890 7870
rect 4910 7850 4970 7870
rect 4990 7850 5050 7870
rect 5070 7850 5130 7870
rect 5150 7850 5210 7870
rect 5230 7850 5290 7870
rect 5310 7850 5370 7870
rect 5390 7850 5450 7870
rect 5470 7850 5530 7870
rect 5550 7850 5610 7870
rect 5630 7850 5690 7870
rect 5710 7850 5720 7870
rect 4720 7840 5720 7850
rect 5760 7870 5960 7880
rect 5760 7850 5770 7870
rect 5790 7850 5850 7870
rect 5870 7850 5930 7870
rect 5950 7850 5960 7870
rect 5760 7840 5960 7850
rect 6000 7870 6200 7880
rect 6000 7850 6010 7870
rect 6030 7850 6090 7870
rect 6110 7850 6170 7870
rect 6190 7850 6200 7870
rect 6000 7840 6200 7850
rect 4240 7790 4440 7800
rect 4240 7770 4250 7790
rect 4270 7770 4330 7790
rect 4350 7770 4410 7790
rect 4430 7770 4440 7790
rect 4240 7760 4440 7770
rect 4480 7790 4680 7800
rect 4480 7770 4490 7790
rect 4510 7770 4570 7790
rect 4590 7770 4650 7790
rect 4670 7770 4680 7790
rect 4480 7760 4680 7770
rect 4720 7790 5720 7800
rect 4720 7770 4730 7790
rect 4750 7770 4810 7790
rect 4830 7770 4890 7790
rect 4910 7770 4970 7790
rect 4990 7770 5050 7790
rect 5070 7770 5130 7790
rect 5150 7770 5210 7790
rect 5230 7770 5290 7790
rect 5310 7770 5370 7790
rect 5390 7770 5450 7790
rect 5470 7770 5530 7790
rect 5550 7770 5610 7790
rect 5630 7770 5690 7790
rect 5710 7770 5720 7790
rect 4720 7760 5720 7770
rect 5760 7790 5960 7800
rect 5760 7770 5770 7790
rect 5790 7770 5850 7790
rect 5870 7770 5930 7790
rect 5950 7770 5960 7790
rect 5760 7760 5960 7770
rect 6000 7790 6200 7800
rect 6000 7770 6010 7790
rect 6030 7770 6090 7790
rect 6110 7770 6170 7790
rect 6190 7770 6200 7790
rect 6000 7760 6200 7770
rect 4240 7710 4440 7720
rect 4240 7690 4250 7710
rect 4270 7690 4330 7710
rect 4350 7690 4410 7710
rect 4430 7690 4440 7710
rect 4240 7680 4440 7690
rect 4480 7710 4680 7720
rect 4480 7690 4490 7710
rect 4510 7690 4570 7710
rect 4590 7690 4650 7710
rect 4670 7690 4680 7710
rect 4480 7680 4680 7690
rect 4720 7710 5720 7720
rect 4720 7690 4730 7710
rect 4750 7690 4810 7710
rect 4830 7690 4890 7710
rect 4910 7690 4970 7710
rect 4990 7690 5050 7710
rect 5070 7690 5130 7710
rect 5150 7690 5210 7710
rect 5230 7690 5290 7710
rect 5310 7690 5370 7710
rect 5390 7690 5450 7710
rect 5470 7690 5530 7710
rect 5550 7690 5610 7710
rect 5630 7690 5690 7710
rect 5710 7690 5720 7710
rect 4720 7680 5720 7690
rect 5760 7710 5960 7720
rect 5760 7690 5770 7710
rect 5790 7690 5850 7710
rect 5870 7690 5930 7710
rect 5950 7690 5960 7710
rect 5760 7680 5960 7690
rect 6000 7710 6200 7720
rect 6000 7690 6010 7710
rect 6030 7690 6090 7710
rect 6110 7690 6170 7710
rect 6190 7690 6200 7710
rect 6000 7680 6200 7690
rect 4240 7630 4440 7640
rect 4240 7610 4250 7630
rect 4270 7610 4330 7630
rect 4350 7610 4410 7630
rect 4430 7610 4440 7630
rect 4240 7600 4440 7610
rect 4480 7630 4680 7640
rect 4480 7610 4490 7630
rect 4510 7610 4570 7630
rect 4590 7610 4650 7630
rect 4670 7610 4680 7630
rect 4480 7600 4680 7610
rect 4720 7630 5720 7640
rect 4720 7610 4730 7630
rect 4750 7610 4810 7630
rect 4830 7610 4890 7630
rect 4910 7610 4970 7630
rect 4990 7610 5050 7630
rect 5070 7610 5130 7630
rect 5150 7610 5210 7630
rect 5230 7610 5290 7630
rect 5310 7610 5370 7630
rect 5390 7610 5450 7630
rect 5470 7610 5530 7630
rect 5550 7610 5610 7630
rect 5630 7610 5690 7630
rect 5710 7610 5720 7630
rect 4720 7600 5720 7610
rect 5760 7630 5960 7640
rect 5760 7610 5770 7630
rect 5790 7610 5850 7630
rect 5870 7610 5930 7630
rect 5950 7610 5960 7630
rect 5760 7600 5960 7610
rect 6000 7630 6200 7640
rect 6000 7610 6010 7630
rect 6030 7610 6090 7630
rect 6110 7610 6170 7630
rect 6190 7610 6200 7630
rect 6000 7600 6200 7610
rect 4240 7550 4440 7560
rect 4240 7530 4250 7550
rect 4270 7530 4330 7550
rect 4350 7530 4410 7550
rect 4430 7530 4440 7550
rect 4240 7520 4440 7530
rect 4480 7550 4680 7560
rect 4480 7530 4490 7550
rect 4510 7530 4570 7550
rect 4590 7530 4650 7550
rect 4670 7530 4680 7550
rect 4480 7520 4680 7530
rect 4720 7550 5720 7560
rect 4720 7530 4730 7550
rect 4750 7530 4810 7550
rect 4830 7530 4890 7550
rect 4910 7530 4970 7550
rect 4990 7530 5050 7550
rect 5070 7530 5130 7550
rect 5150 7530 5210 7550
rect 5230 7530 5290 7550
rect 5310 7530 5370 7550
rect 5390 7530 5450 7550
rect 5470 7530 5530 7550
rect 5550 7530 5610 7550
rect 5630 7530 5690 7550
rect 5710 7530 5720 7550
rect 4720 7520 5720 7530
rect 5760 7550 5960 7560
rect 5760 7530 5770 7550
rect 5790 7530 5850 7550
rect 5870 7530 5930 7550
rect 5950 7530 5960 7550
rect 5760 7520 5960 7530
rect 6000 7550 6200 7560
rect 6000 7530 6010 7550
rect 6030 7530 6090 7550
rect 6110 7530 6170 7550
rect 6190 7530 6200 7550
rect 6000 7520 6200 7530
rect 4240 7470 4440 7480
rect 4240 7450 4250 7470
rect 4270 7450 4330 7470
rect 4350 7450 4410 7470
rect 4430 7450 4440 7470
rect 4240 7440 4440 7450
rect 4480 7470 4680 7480
rect 4480 7450 4490 7470
rect 4510 7450 4570 7470
rect 4590 7450 4650 7470
rect 4670 7450 4680 7470
rect 4480 7440 4680 7450
rect 4720 7470 5720 7480
rect 4720 7450 4730 7470
rect 4750 7450 4810 7470
rect 4830 7450 4890 7470
rect 4910 7450 4970 7470
rect 4990 7450 5050 7470
rect 5070 7450 5130 7470
rect 5150 7450 5210 7470
rect 5230 7450 5290 7470
rect 5310 7450 5370 7470
rect 5390 7450 5450 7470
rect 5470 7450 5530 7470
rect 5550 7450 5610 7470
rect 5630 7450 5690 7470
rect 5710 7450 5720 7470
rect 4720 7440 5720 7450
rect 5760 7470 5960 7480
rect 5760 7450 5770 7470
rect 5790 7450 5850 7470
rect 5870 7450 5930 7470
rect 5950 7450 5960 7470
rect 5760 7440 5960 7450
rect 6000 7470 6200 7480
rect 6000 7450 6010 7470
rect 6030 7450 6090 7470
rect 6110 7450 6170 7470
rect 6190 7450 6200 7470
rect 6000 7440 6200 7450
rect 4240 7390 4440 7400
rect 4240 7370 4250 7390
rect 4270 7370 4330 7390
rect 4350 7370 4410 7390
rect 4430 7370 4440 7390
rect 4240 7360 4440 7370
rect 4480 7390 4680 7400
rect 4480 7370 4490 7390
rect 4510 7370 4570 7390
rect 4590 7370 4650 7390
rect 4670 7370 4680 7390
rect 4480 7360 4680 7370
rect 4720 7390 5720 7400
rect 4720 7370 4730 7390
rect 4750 7370 4810 7390
rect 4830 7370 4890 7390
rect 4910 7370 4970 7390
rect 4990 7370 5050 7390
rect 5070 7370 5130 7390
rect 5150 7370 5210 7390
rect 5230 7370 5290 7390
rect 5310 7370 5370 7390
rect 5390 7370 5450 7390
rect 5470 7370 5530 7390
rect 5550 7370 5610 7390
rect 5630 7370 5690 7390
rect 5710 7370 5720 7390
rect 4720 7360 5720 7370
rect 5760 7390 5960 7400
rect 5760 7370 5770 7390
rect 5790 7370 5850 7390
rect 5870 7370 5930 7390
rect 5950 7370 5960 7390
rect 5760 7360 5960 7370
rect 6000 7390 6200 7400
rect 6000 7370 6010 7390
rect 6030 7370 6090 7390
rect 6110 7370 6170 7390
rect 6190 7370 6200 7390
rect 6000 7360 6200 7370
rect 4240 7310 4440 7320
rect 4240 7290 4250 7310
rect 4270 7290 4330 7310
rect 4350 7290 4410 7310
rect 4430 7290 4440 7310
rect 4240 7280 4440 7290
rect 4480 7310 4680 7320
rect 4480 7290 4490 7310
rect 4510 7290 4570 7310
rect 4590 7290 4650 7310
rect 4670 7290 4680 7310
rect 4480 7280 4680 7290
rect 4720 7310 5720 7320
rect 4720 7290 4730 7310
rect 4750 7290 4810 7310
rect 4830 7290 4890 7310
rect 4910 7290 4970 7310
rect 4990 7290 5050 7310
rect 5070 7290 5130 7310
rect 5150 7290 5210 7310
rect 5230 7290 5290 7310
rect 5310 7290 5370 7310
rect 5390 7290 5450 7310
rect 5470 7290 5530 7310
rect 5550 7290 5610 7310
rect 5630 7290 5690 7310
rect 5710 7290 5720 7310
rect 4720 7280 5720 7290
rect 5760 7310 5960 7320
rect 5760 7290 5770 7310
rect 5790 7290 5850 7310
rect 5870 7290 5930 7310
rect 5950 7290 5960 7310
rect 5760 7280 5960 7290
rect 6000 7310 6200 7320
rect 6000 7290 6010 7310
rect 6030 7290 6090 7310
rect 6110 7290 6170 7310
rect 6190 7290 6200 7310
rect 6000 7280 6200 7290
rect 4240 7230 4440 7240
rect 4240 7210 4250 7230
rect 4270 7210 4330 7230
rect 4350 7210 4410 7230
rect 4430 7210 4440 7230
rect 4240 7200 4440 7210
rect 4480 7230 4680 7240
rect 4480 7210 4490 7230
rect 4510 7210 4570 7230
rect 4590 7210 4650 7230
rect 4670 7210 4680 7230
rect 4480 7200 4680 7210
rect 4720 7230 5720 7240
rect 4720 7210 4730 7230
rect 4750 7210 4810 7230
rect 4830 7210 4890 7230
rect 4910 7210 4970 7230
rect 4990 7210 5050 7230
rect 5070 7210 5130 7230
rect 5150 7210 5210 7230
rect 5230 7210 5290 7230
rect 5310 7210 5370 7230
rect 5390 7210 5450 7230
rect 5470 7210 5530 7230
rect 5550 7210 5610 7230
rect 5630 7210 5690 7230
rect 5710 7210 5720 7230
rect 4720 7200 5720 7210
rect 5760 7230 5960 7240
rect 5760 7210 5770 7230
rect 5790 7210 5850 7230
rect 5870 7210 5930 7230
rect 5950 7210 5960 7230
rect 5760 7200 5960 7210
rect 6000 7230 6200 7240
rect 6000 7210 6010 7230
rect 6030 7210 6090 7230
rect 6110 7210 6170 7230
rect 6190 7210 6200 7230
rect 6000 7200 6200 7210
rect 4240 7150 4440 7160
rect 4240 7130 4250 7150
rect 4270 7130 4330 7150
rect 4350 7130 4410 7150
rect 4430 7130 4440 7150
rect 4240 7120 4440 7130
rect 4480 7150 4680 7160
rect 4480 7130 4490 7150
rect 4510 7130 4570 7150
rect 4590 7130 4650 7150
rect 4670 7130 4680 7150
rect 4480 7120 4680 7130
rect 4720 7150 5720 7160
rect 4720 7130 4730 7150
rect 4750 7130 4810 7150
rect 4830 7130 4890 7150
rect 4910 7130 4970 7150
rect 4990 7130 5050 7150
rect 5070 7130 5130 7150
rect 5150 7130 5210 7150
rect 5230 7130 5290 7150
rect 5310 7130 5370 7150
rect 5390 7130 5450 7150
rect 5470 7130 5530 7150
rect 5550 7130 5610 7150
rect 5630 7130 5690 7150
rect 5710 7130 5720 7150
rect 4720 7120 5720 7130
rect 5760 7150 5960 7160
rect 5760 7130 5770 7150
rect 5790 7130 5850 7150
rect 5870 7130 5930 7150
rect 5950 7130 5960 7150
rect 5760 7120 5960 7130
rect 6000 7150 6200 7160
rect 6000 7130 6010 7150
rect 6030 7130 6090 7150
rect 6110 7130 6170 7150
rect 6190 7130 6200 7150
rect 6000 7120 6200 7130
rect 4240 7070 4440 7080
rect 4240 7050 4250 7070
rect 4270 7050 4330 7070
rect 4350 7050 4410 7070
rect 4430 7050 4440 7070
rect 4240 7040 4440 7050
rect 4480 7070 4680 7080
rect 4480 7050 4490 7070
rect 4510 7050 4570 7070
rect 4590 7050 4650 7070
rect 4670 7050 4680 7070
rect 4480 7040 4680 7050
rect 4720 7070 5720 7080
rect 4720 7050 4730 7070
rect 4750 7050 4810 7070
rect 4830 7050 4890 7070
rect 4910 7050 4970 7070
rect 4990 7050 5050 7070
rect 5070 7050 5130 7070
rect 5150 7050 5210 7070
rect 5230 7050 5290 7070
rect 5310 7050 5370 7070
rect 5390 7050 5450 7070
rect 5470 7050 5530 7070
rect 5550 7050 5610 7070
rect 5630 7050 5690 7070
rect 5710 7050 5720 7070
rect 4720 7040 5720 7050
rect 5760 7070 5960 7080
rect 5760 7050 5770 7070
rect 5790 7050 5850 7070
rect 5870 7050 5930 7070
rect 5950 7050 5960 7070
rect 5760 7040 5960 7050
rect 6000 7070 6200 7080
rect 6000 7050 6010 7070
rect 6030 7050 6090 7070
rect 6110 7050 6170 7070
rect 6190 7050 6200 7070
rect 6000 7040 6200 7050
rect 4240 6990 4440 7000
rect 4240 6970 4250 6990
rect 4270 6970 4330 6990
rect 4350 6970 4410 6990
rect 4430 6970 4440 6990
rect 4240 6960 4440 6970
rect 4480 6990 4680 7000
rect 4480 6970 4490 6990
rect 4510 6970 4570 6990
rect 4590 6970 4650 6990
rect 4670 6970 4680 6990
rect 4480 6960 4680 6970
rect 4720 6990 5720 7000
rect 4720 6970 4730 6990
rect 4750 6970 4810 6990
rect 4830 6970 4890 6990
rect 4910 6970 4970 6990
rect 4990 6970 5050 6990
rect 5070 6970 5130 6990
rect 5150 6970 5210 6990
rect 5230 6970 5290 6990
rect 5310 6970 5370 6990
rect 5390 6970 5450 6990
rect 5470 6970 5530 6990
rect 5550 6970 5610 6990
rect 5630 6970 5690 6990
rect 5710 6970 5720 6990
rect 4720 6960 5720 6970
rect 5760 6990 5960 7000
rect 5760 6970 5770 6990
rect 5790 6970 5850 6990
rect 5870 6970 5930 6990
rect 5950 6970 5960 6990
rect 5760 6960 5960 6970
rect 6000 6990 6200 7000
rect 6000 6970 6010 6990
rect 6030 6970 6090 6990
rect 6110 6970 6170 6990
rect 6190 6970 6200 6990
rect 6000 6960 6200 6970
rect 4240 6910 4440 6920
rect 4240 6890 4250 6910
rect 4270 6890 4330 6910
rect 4350 6890 4410 6910
rect 4430 6890 4440 6910
rect 4240 6880 4440 6890
rect 4480 6910 4680 6920
rect 4480 6890 4490 6910
rect 4510 6890 4570 6910
rect 4590 6890 4650 6910
rect 4670 6890 4680 6910
rect 4480 6880 4680 6890
rect 4720 6910 5720 6920
rect 4720 6890 4730 6910
rect 4750 6890 4810 6910
rect 4830 6890 4890 6910
rect 4910 6890 4970 6910
rect 4990 6890 5050 6910
rect 5070 6890 5130 6910
rect 5150 6890 5210 6910
rect 5230 6890 5290 6910
rect 5310 6890 5370 6910
rect 5390 6890 5450 6910
rect 5470 6890 5530 6910
rect 5550 6890 5610 6910
rect 5630 6890 5690 6910
rect 5710 6890 5720 6910
rect 4720 6880 5720 6890
rect 5760 6910 5960 6920
rect 5760 6890 5770 6910
rect 5790 6890 5850 6910
rect 5870 6890 5930 6910
rect 5950 6890 5960 6910
rect 5760 6880 5960 6890
rect 6000 6910 6200 6920
rect 6000 6890 6010 6910
rect 6030 6890 6090 6910
rect 6110 6890 6170 6910
rect 6190 6890 6200 6910
rect 6000 6880 6200 6890
rect 4240 6830 4440 6840
rect 4240 6810 4250 6830
rect 4270 6810 4330 6830
rect 4350 6810 4410 6830
rect 4430 6810 4440 6830
rect 4240 6800 4440 6810
rect 4480 6830 4680 6840
rect 4480 6810 4490 6830
rect 4510 6810 4570 6830
rect 4590 6810 4650 6830
rect 4670 6810 4680 6830
rect 4480 6800 4680 6810
rect 4720 6830 5720 6840
rect 4720 6810 4730 6830
rect 4750 6810 4810 6830
rect 4830 6810 4890 6830
rect 4910 6810 4970 6830
rect 4990 6810 5050 6830
rect 5070 6810 5130 6830
rect 5150 6810 5210 6830
rect 5230 6810 5290 6830
rect 5310 6810 5370 6830
rect 5390 6810 5450 6830
rect 5470 6810 5530 6830
rect 5550 6810 5610 6830
rect 5630 6810 5690 6830
rect 5710 6810 5720 6830
rect 4720 6800 5720 6810
rect 5760 6830 5960 6840
rect 5760 6810 5770 6830
rect 5790 6810 5850 6830
rect 5870 6810 5930 6830
rect 5950 6810 5960 6830
rect 5760 6800 5960 6810
rect 6000 6830 6200 6840
rect 6000 6810 6010 6830
rect 6030 6810 6090 6830
rect 6110 6810 6170 6830
rect 6190 6810 6200 6830
rect 6000 6800 6200 6810
rect 4240 6750 4440 6760
rect 4240 6730 4250 6750
rect 4270 6730 4330 6750
rect 4350 6730 4410 6750
rect 4430 6730 4440 6750
rect 4240 6720 4440 6730
rect 4480 6750 4680 6760
rect 4480 6730 4490 6750
rect 4510 6730 4570 6750
rect 4590 6730 4650 6750
rect 4670 6730 4680 6750
rect 4480 6720 4680 6730
rect 4720 6750 5720 6760
rect 4720 6730 4730 6750
rect 4750 6730 4810 6750
rect 4830 6730 4890 6750
rect 4910 6730 4970 6750
rect 4990 6730 5050 6750
rect 5070 6730 5130 6750
rect 5150 6730 5210 6750
rect 5230 6730 5290 6750
rect 5310 6730 5370 6750
rect 5390 6730 5450 6750
rect 5470 6730 5530 6750
rect 5550 6730 5610 6750
rect 5630 6730 5690 6750
rect 5710 6730 5720 6750
rect 4720 6720 5720 6730
rect 5760 6750 5960 6760
rect 5760 6730 5770 6750
rect 5790 6730 5850 6750
rect 5870 6730 5930 6750
rect 5950 6730 5960 6750
rect 5760 6720 5960 6730
rect 6000 6750 6200 6760
rect 6000 6730 6010 6750
rect 6030 6730 6090 6750
rect 6110 6730 6170 6750
rect 6190 6730 6200 6750
rect 6000 6720 6200 6730
rect 4240 6670 4440 6680
rect 4240 6650 4250 6670
rect 4270 6650 4330 6670
rect 4350 6650 4410 6670
rect 4430 6650 4440 6670
rect 4240 6640 4440 6650
rect 4480 6670 4680 6680
rect 4480 6650 4490 6670
rect 4510 6650 4570 6670
rect 4590 6650 4650 6670
rect 4670 6650 4680 6670
rect 4480 6640 4680 6650
rect 4720 6670 5720 6680
rect 4720 6650 4730 6670
rect 4750 6650 4810 6670
rect 4830 6650 4890 6670
rect 4910 6650 4970 6670
rect 4990 6650 5050 6670
rect 5070 6650 5130 6670
rect 5150 6650 5210 6670
rect 5230 6650 5290 6670
rect 5310 6650 5370 6670
rect 5390 6650 5450 6670
rect 5470 6650 5530 6670
rect 5550 6650 5610 6670
rect 5630 6650 5690 6670
rect 5710 6650 5720 6670
rect 4720 6640 5720 6650
rect 5760 6670 5960 6680
rect 5760 6650 5770 6670
rect 5790 6650 5850 6670
rect 5870 6650 5930 6670
rect 5950 6650 5960 6670
rect 5760 6640 5960 6650
rect 6000 6670 6200 6680
rect 6000 6650 6010 6670
rect 6030 6650 6090 6670
rect 6110 6650 6170 6670
rect 6190 6650 6200 6670
rect 6000 6640 6200 6650
rect 4240 6590 4440 6600
rect 4240 6570 4250 6590
rect 4270 6570 4330 6590
rect 4350 6570 4410 6590
rect 4430 6570 4440 6590
rect 4240 6560 4440 6570
rect 4480 6590 4680 6600
rect 4480 6570 4490 6590
rect 4510 6570 4570 6590
rect 4590 6570 4650 6590
rect 4670 6570 4680 6590
rect 4480 6560 4680 6570
rect 4720 6590 5720 6600
rect 4720 6570 4730 6590
rect 4750 6570 4810 6590
rect 4830 6570 4890 6590
rect 4910 6570 4970 6590
rect 4990 6570 5050 6590
rect 5070 6570 5130 6590
rect 5150 6570 5210 6590
rect 5230 6570 5290 6590
rect 5310 6570 5370 6590
rect 5390 6570 5450 6590
rect 5470 6570 5530 6590
rect 5550 6570 5610 6590
rect 5630 6570 5690 6590
rect 5710 6570 5720 6590
rect 4720 6560 5720 6570
rect 5760 6590 5960 6600
rect 5760 6570 5770 6590
rect 5790 6570 5850 6590
rect 5870 6570 5930 6590
rect 5950 6570 5960 6590
rect 5760 6560 5960 6570
rect 6000 6590 6200 6600
rect 6000 6570 6010 6590
rect 6030 6570 6090 6590
rect 6110 6570 6170 6590
rect 6190 6570 6200 6590
rect 6000 6560 6200 6570
rect 4240 6510 4440 6520
rect 4240 6490 4250 6510
rect 4270 6490 4330 6510
rect 4350 6490 4410 6510
rect 4430 6490 4440 6510
rect 4240 6480 4440 6490
rect 4480 6510 4680 6520
rect 4480 6490 4490 6510
rect 4510 6490 4570 6510
rect 4590 6490 4650 6510
rect 4670 6490 4680 6510
rect 4480 6480 4680 6490
rect 4720 6510 5720 6520
rect 4720 6490 4730 6510
rect 4750 6490 4810 6510
rect 4830 6490 4890 6510
rect 4910 6490 4970 6510
rect 4990 6490 5050 6510
rect 5070 6490 5130 6510
rect 5150 6490 5210 6510
rect 5230 6490 5290 6510
rect 5310 6490 5370 6510
rect 5390 6490 5450 6510
rect 5470 6490 5530 6510
rect 5550 6490 5610 6510
rect 5630 6490 5690 6510
rect 5710 6490 5720 6510
rect 4720 6480 5720 6490
rect 5760 6510 5960 6520
rect 5760 6490 5770 6510
rect 5790 6490 5850 6510
rect 5870 6490 5930 6510
rect 5950 6490 5960 6510
rect 5760 6480 5960 6490
rect 6000 6510 6200 6520
rect 6000 6490 6010 6510
rect 6030 6490 6090 6510
rect 6110 6490 6170 6510
rect 6190 6490 6200 6510
rect 6000 6480 6200 6490
rect 4240 6430 4440 6440
rect 4240 6410 4250 6430
rect 4270 6410 4330 6430
rect 4350 6410 4410 6430
rect 4430 6410 4440 6430
rect 4240 6400 4440 6410
rect 4480 6430 4680 6440
rect 4480 6410 4490 6430
rect 4510 6410 4570 6430
rect 4590 6410 4650 6430
rect 4670 6410 4680 6430
rect 4480 6400 4680 6410
rect 4720 6430 5720 6440
rect 4720 6410 4730 6430
rect 4750 6410 4810 6430
rect 4830 6410 4890 6430
rect 4910 6410 4970 6430
rect 4990 6410 5050 6430
rect 5070 6410 5130 6430
rect 5150 6410 5210 6430
rect 5230 6410 5290 6430
rect 5310 6410 5370 6430
rect 5390 6410 5450 6430
rect 5470 6410 5530 6430
rect 5550 6410 5610 6430
rect 5630 6410 5690 6430
rect 5710 6410 5720 6430
rect 4720 6400 5720 6410
rect 5760 6430 5960 6440
rect 5760 6410 5770 6430
rect 5790 6410 5850 6430
rect 5870 6410 5930 6430
rect 5950 6410 5960 6430
rect 5760 6400 5960 6410
rect 6000 6430 6200 6440
rect 6000 6410 6010 6430
rect 6030 6410 6090 6430
rect 6110 6410 6170 6430
rect 6190 6410 6200 6430
rect 6000 6400 6200 6410
rect 4240 6350 4440 6360
rect 4240 6330 4250 6350
rect 4270 6330 4330 6350
rect 4350 6330 4410 6350
rect 4430 6330 4440 6350
rect 4240 6320 4440 6330
rect 4480 6350 4680 6360
rect 4480 6330 4490 6350
rect 4510 6330 4570 6350
rect 4590 6330 4650 6350
rect 4670 6330 4680 6350
rect 4480 6320 4680 6330
rect 4720 6350 5720 6360
rect 4720 6330 4730 6350
rect 4750 6330 4810 6350
rect 4830 6330 4890 6350
rect 4910 6330 4970 6350
rect 4990 6330 5050 6350
rect 5070 6330 5130 6350
rect 5150 6330 5210 6350
rect 5230 6330 5290 6350
rect 5310 6330 5370 6350
rect 5390 6330 5450 6350
rect 5470 6330 5530 6350
rect 5550 6330 5610 6350
rect 5630 6330 5690 6350
rect 5710 6330 5720 6350
rect 4720 6320 5720 6330
rect 5760 6350 5960 6360
rect 5760 6330 5770 6350
rect 5790 6330 5850 6350
rect 5870 6330 5930 6350
rect 5950 6330 5960 6350
rect 5760 6320 5960 6330
rect 6000 6350 6200 6360
rect 6000 6330 6010 6350
rect 6030 6330 6090 6350
rect 6110 6330 6170 6350
rect 6190 6330 6200 6350
rect 6000 6320 6200 6330
rect 4240 6270 4440 6280
rect 4240 6250 4250 6270
rect 4270 6250 4330 6270
rect 4350 6250 4410 6270
rect 4430 6250 4440 6270
rect 4240 6240 4440 6250
rect 4480 6270 4680 6280
rect 4480 6250 4490 6270
rect 4510 6250 4570 6270
rect 4590 6250 4650 6270
rect 4670 6250 4680 6270
rect 4480 6240 4680 6250
rect 4720 6270 5720 6280
rect 4720 6250 4730 6270
rect 4750 6250 4810 6270
rect 4830 6250 4890 6270
rect 4910 6250 4970 6270
rect 4990 6250 5050 6270
rect 5070 6250 5130 6270
rect 5150 6250 5210 6270
rect 5230 6250 5290 6270
rect 5310 6250 5370 6270
rect 5390 6250 5450 6270
rect 5470 6250 5530 6270
rect 5550 6250 5610 6270
rect 5630 6250 5690 6270
rect 5710 6250 5720 6270
rect 4720 6240 5720 6250
rect 5760 6270 5960 6280
rect 5760 6250 5770 6270
rect 5790 6250 5850 6270
rect 5870 6250 5930 6270
rect 5950 6250 5960 6270
rect 5760 6240 5960 6250
rect 6000 6270 6200 6280
rect 6000 6250 6010 6270
rect 6030 6250 6090 6270
rect 6110 6250 6170 6270
rect 6190 6250 6200 6270
rect 6000 6240 6200 6250
rect 4240 6190 4440 6200
rect 4240 6170 4250 6190
rect 4270 6170 4330 6190
rect 4350 6170 4410 6190
rect 4430 6170 4440 6190
rect 4240 6160 4440 6170
rect 4480 6190 4680 6200
rect 4480 6170 4490 6190
rect 4510 6170 4570 6190
rect 4590 6170 4650 6190
rect 4670 6170 4680 6190
rect 4480 6160 4680 6170
rect 4720 6190 5720 6200
rect 4720 6170 4730 6190
rect 4750 6170 4810 6190
rect 4830 6170 4890 6190
rect 4910 6170 4970 6190
rect 4990 6170 5050 6190
rect 5070 6170 5130 6190
rect 5150 6170 5210 6190
rect 5230 6170 5290 6190
rect 5310 6170 5370 6190
rect 5390 6170 5450 6190
rect 5470 6170 5530 6190
rect 5550 6170 5610 6190
rect 5630 6170 5690 6190
rect 5710 6170 5720 6190
rect 4720 6160 5720 6170
rect 5760 6190 5960 6200
rect 5760 6170 5770 6190
rect 5790 6170 5850 6190
rect 5870 6170 5930 6190
rect 5950 6170 5960 6190
rect 5760 6160 5960 6170
rect 6000 6190 6200 6200
rect 6000 6170 6010 6190
rect 6030 6170 6090 6190
rect 6110 6170 6170 6190
rect 6190 6170 6200 6190
rect 6000 6160 6200 6170
rect 4240 6110 4440 6120
rect 4240 6090 4250 6110
rect 4270 6090 4330 6110
rect 4350 6090 4410 6110
rect 4430 6090 4440 6110
rect 4240 6080 4440 6090
rect 4480 6110 4680 6120
rect 4480 6090 4490 6110
rect 4510 6090 4570 6110
rect 4590 6090 4650 6110
rect 4670 6090 4680 6110
rect 4480 6080 4680 6090
rect 4720 6110 5720 6120
rect 4720 6090 4730 6110
rect 4750 6090 4810 6110
rect 4830 6090 4890 6110
rect 4910 6090 4970 6110
rect 4990 6090 5050 6110
rect 5070 6090 5130 6110
rect 5150 6090 5210 6110
rect 5230 6090 5290 6110
rect 5310 6090 5370 6110
rect 5390 6090 5450 6110
rect 5470 6090 5530 6110
rect 5550 6090 5610 6110
rect 5630 6090 5690 6110
rect 5710 6090 5720 6110
rect 4720 6080 5720 6090
rect 5760 6110 5960 6120
rect 5760 6090 5770 6110
rect 5790 6090 5850 6110
rect 5870 6090 5930 6110
rect 5950 6090 5960 6110
rect 5760 6080 5960 6090
rect 6000 6110 6200 6120
rect 6000 6090 6010 6110
rect 6030 6090 6090 6110
rect 6110 6090 6170 6110
rect 6190 6090 6200 6110
rect 6000 6080 6200 6090
rect 4240 6030 4440 6040
rect 4240 6010 4250 6030
rect 4270 6010 4330 6030
rect 4350 6010 4410 6030
rect 4430 6010 4440 6030
rect 4240 6000 4440 6010
rect 4480 6030 4680 6040
rect 4480 6010 4490 6030
rect 4510 6010 4570 6030
rect 4590 6010 4650 6030
rect 4670 6010 4680 6030
rect 4480 6000 4680 6010
rect 4720 6030 5720 6040
rect 4720 6010 4730 6030
rect 4750 6010 4810 6030
rect 4830 6010 4890 6030
rect 4910 6010 4970 6030
rect 4990 6010 5050 6030
rect 5070 6010 5130 6030
rect 5150 6010 5210 6030
rect 5230 6010 5290 6030
rect 5310 6010 5370 6030
rect 5390 6010 5450 6030
rect 5470 6010 5530 6030
rect 5550 6010 5610 6030
rect 5630 6010 5690 6030
rect 5710 6010 5720 6030
rect 4720 6000 5720 6010
rect 5760 6030 5960 6040
rect 5760 6010 5770 6030
rect 5790 6010 5850 6030
rect 5870 6010 5930 6030
rect 5950 6010 5960 6030
rect 5760 6000 5960 6010
rect 6000 6030 6200 6040
rect 6000 6010 6010 6030
rect 6030 6010 6090 6030
rect 6110 6010 6170 6030
rect 6190 6010 6200 6030
rect 6000 6000 6200 6010
rect 4240 5950 4440 5960
rect 4240 5930 4250 5950
rect 4270 5930 4330 5950
rect 4350 5930 4410 5950
rect 4430 5930 4440 5950
rect 4240 5920 4440 5930
rect 4480 5950 4680 5960
rect 4480 5930 4490 5950
rect 4510 5930 4570 5950
rect 4590 5930 4650 5950
rect 4670 5930 4680 5950
rect 4480 5920 4680 5930
rect 4720 5950 5720 5960
rect 4720 5930 4730 5950
rect 4750 5930 4810 5950
rect 4830 5930 4890 5950
rect 4910 5930 4970 5950
rect 4990 5930 5050 5950
rect 5070 5930 5130 5950
rect 5150 5930 5210 5950
rect 5230 5930 5290 5950
rect 5310 5930 5370 5950
rect 5390 5930 5450 5950
rect 5470 5930 5530 5950
rect 5550 5930 5610 5950
rect 5630 5930 5690 5950
rect 5710 5930 5720 5950
rect 4720 5920 5720 5930
rect 5760 5950 5960 5960
rect 5760 5930 5770 5950
rect 5790 5930 5850 5950
rect 5870 5930 5930 5950
rect 5950 5930 5960 5950
rect 5760 5920 5960 5930
rect 6000 5950 6200 5960
rect 6000 5930 6010 5950
rect 6030 5930 6090 5950
rect 6110 5930 6170 5950
rect 6190 5930 6200 5950
rect 6000 5920 6200 5930
rect 4240 5870 4440 5880
rect 4240 5850 4250 5870
rect 4270 5850 4330 5870
rect 4350 5850 4410 5870
rect 4430 5850 4440 5870
rect 4240 5840 4440 5850
rect 4480 5870 4680 5880
rect 4480 5850 4490 5870
rect 4510 5850 4570 5870
rect 4590 5850 4650 5870
rect 4670 5850 4680 5870
rect 4480 5840 4680 5850
rect 4720 5870 5720 5880
rect 4720 5850 4730 5870
rect 4750 5850 4810 5870
rect 4830 5850 4890 5870
rect 4910 5850 4970 5870
rect 4990 5850 5050 5870
rect 5070 5850 5130 5870
rect 5150 5850 5210 5870
rect 5230 5850 5290 5870
rect 5310 5850 5370 5870
rect 5390 5850 5450 5870
rect 5470 5850 5530 5870
rect 5550 5850 5610 5870
rect 5630 5850 5690 5870
rect 5710 5850 5720 5870
rect 4720 5840 5720 5850
rect 5760 5870 5960 5880
rect 5760 5850 5770 5870
rect 5790 5850 5850 5870
rect 5870 5850 5930 5870
rect 5950 5850 5960 5870
rect 5760 5840 5960 5850
rect 6000 5870 6200 5880
rect 6000 5850 6010 5870
rect 6030 5850 6090 5870
rect 6110 5850 6170 5870
rect 6190 5850 6200 5870
rect 6000 5840 6200 5850
rect 4240 5790 4440 5800
rect 4240 5770 4250 5790
rect 4270 5770 4330 5790
rect 4350 5770 4410 5790
rect 4430 5770 4440 5790
rect 4240 5760 4440 5770
rect 4480 5790 4680 5800
rect 4480 5770 4490 5790
rect 4510 5770 4570 5790
rect 4590 5770 4650 5790
rect 4670 5770 4680 5790
rect 4480 5760 4680 5770
rect 4720 5790 5720 5800
rect 4720 5770 4730 5790
rect 4750 5770 4810 5790
rect 4830 5770 4890 5790
rect 4910 5770 4970 5790
rect 4990 5770 5050 5790
rect 5070 5770 5130 5790
rect 5150 5770 5210 5790
rect 5230 5770 5290 5790
rect 5310 5770 5370 5790
rect 5390 5770 5450 5790
rect 5470 5770 5530 5790
rect 5550 5770 5610 5790
rect 5630 5770 5690 5790
rect 5710 5770 5720 5790
rect 4720 5760 5720 5770
rect 5760 5790 5960 5800
rect 5760 5770 5770 5790
rect 5790 5770 5850 5790
rect 5870 5770 5930 5790
rect 5950 5770 5960 5790
rect 5760 5760 5960 5770
rect 6000 5790 6200 5800
rect 6000 5770 6010 5790
rect 6030 5770 6090 5790
rect 6110 5770 6170 5790
rect 6190 5770 6200 5790
rect 6000 5760 6200 5770
rect 4240 5710 4440 5720
rect 4240 5690 4250 5710
rect 4270 5690 4330 5710
rect 4350 5690 4410 5710
rect 4430 5690 4440 5710
rect 4240 5680 4440 5690
rect 4480 5710 4680 5720
rect 4480 5690 4490 5710
rect 4510 5690 4570 5710
rect 4590 5690 4650 5710
rect 4670 5690 4680 5710
rect 4480 5680 4680 5690
rect 4720 5710 5720 5720
rect 4720 5690 4730 5710
rect 4750 5690 4810 5710
rect 4830 5690 4890 5710
rect 4910 5690 4970 5710
rect 4990 5690 5050 5710
rect 5070 5690 5130 5710
rect 5150 5690 5210 5710
rect 5230 5690 5290 5710
rect 5310 5690 5370 5710
rect 5390 5690 5450 5710
rect 5470 5690 5530 5710
rect 5550 5690 5610 5710
rect 5630 5690 5690 5710
rect 5710 5690 5720 5710
rect 4720 5680 5720 5690
rect 5760 5710 5960 5720
rect 5760 5690 5770 5710
rect 5790 5690 5850 5710
rect 5870 5690 5930 5710
rect 5950 5690 5960 5710
rect 5760 5680 5960 5690
rect 6000 5710 6200 5720
rect 6000 5690 6010 5710
rect 6030 5690 6090 5710
rect 6110 5690 6170 5710
rect 6190 5690 6200 5710
rect 6000 5680 6200 5690
rect 4240 5630 4440 5640
rect 4240 5610 4250 5630
rect 4270 5610 4330 5630
rect 4350 5610 4410 5630
rect 4430 5610 4440 5630
rect 4240 5600 4440 5610
rect 4480 5630 4680 5640
rect 4480 5610 4490 5630
rect 4510 5610 4570 5630
rect 4590 5610 4650 5630
rect 4670 5610 4680 5630
rect 4480 5600 4680 5610
rect 4720 5630 5720 5640
rect 4720 5610 4730 5630
rect 4750 5610 4810 5630
rect 4830 5610 4890 5630
rect 4910 5610 4970 5630
rect 4990 5610 5050 5630
rect 5070 5610 5130 5630
rect 5150 5610 5210 5630
rect 5230 5610 5290 5630
rect 5310 5610 5370 5630
rect 5390 5610 5450 5630
rect 5470 5610 5530 5630
rect 5550 5610 5610 5630
rect 5630 5610 5690 5630
rect 5710 5610 5720 5630
rect 4720 5600 5720 5610
rect 5760 5630 5960 5640
rect 5760 5610 5770 5630
rect 5790 5610 5850 5630
rect 5870 5610 5930 5630
rect 5950 5610 5960 5630
rect 5760 5600 5960 5610
rect 6000 5630 6200 5640
rect 6000 5610 6010 5630
rect 6030 5610 6090 5630
rect 6110 5610 6170 5630
rect 6190 5610 6200 5630
rect 6000 5600 6200 5610
rect 4240 5550 4440 5560
rect 4240 5530 4250 5550
rect 4270 5530 4330 5550
rect 4350 5530 4410 5550
rect 4430 5530 4440 5550
rect 4240 5520 4440 5530
rect 4480 5550 4680 5560
rect 4480 5530 4490 5550
rect 4510 5530 4570 5550
rect 4590 5530 4650 5550
rect 4670 5530 4680 5550
rect 4480 5520 4680 5530
rect 4720 5550 5720 5560
rect 4720 5530 4730 5550
rect 4750 5530 4810 5550
rect 4830 5530 4890 5550
rect 4910 5530 4970 5550
rect 4990 5530 5050 5550
rect 5070 5530 5130 5550
rect 5150 5530 5210 5550
rect 5230 5530 5290 5550
rect 5310 5530 5370 5550
rect 5390 5530 5450 5550
rect 5470 5530 5530 5550
rect 5550 5530 5610 5550
rect 5630 5530 5690 5550
rect 5710 5530 5720 5550
rect 4720 5520 5720 5530
rect 5760 5550 5960 5560
rect 5760 5530 5770 5550
rect 5790 5530 5850 5550
rect 5870 5530 5930 5550
rect 5950 5530 5960 5550
rect 5760 5520 5960 5530
rect 6000 5550 6200 5560
rect 6000 5530 6010 5550
rect 6030 5530 6090 5550
rect 6110 5530 6170 5550
rect 6190 5530 6200 5550
rect 6000 5520 6200 5530
rect 4240 5470 4440 5480
rect 4240 5450 4250 5470
rect 4270 5450 4330 5470
rect 4350 5450 4410 5470
rect 4430 5450 4440 5470
rect 4240 5440 4440 5450
rect 4480 5470 4680 5480
rect 4480 5450 4490 5470
rect 4510 5450 4570 5470
rect 4590 5450 4650 5470
rect 4670 5450 4680 5470
rect 4480 5440 4680 5450
rect 4720 5470 5720 5480
rect 4720 5450 4730 5470
rect 4750 5450 4810 5470
rect 4830 5450 4890 5470
rect 4910 5450 4970 5470
rect 4990 5450 5050 5470
rect 5070 5450 5130 5470
rect 5150 5450 5210 5470
rect 5230 5450 5290 5470
rect 5310 5450 5370 5470
rect 5390 5450 5450 5470
rect 5470 5450 5530 5470
rect 5550 5450 5610 5470
rect 5630 5450 5690 5470
rect 5710 5450 5720 5470
rect 4720 5440 5720 5450
rect 5760 5470 5960 5480
rect 5760 5450 5770 5470
rect 5790 5450 5850 5470
rect 5870 5450 5930 5470
rect 5950 5450 5960 5470
rect 5760 5440 5960 5450
rect 6000 5470 6200 5480
rect 6000 5450 6010 5470
rect 6030 5450 6090 5470
rect 6110 5450 6170 5470
rect 6190 5450 6200 5470
rect 6000 5440 6200 5450
rect 4240 5390 4440 5400
rect 4240 5370 4250 5390
rect 4270 5370 4330 5390
rect 4350 5370 4410 5390
rect 4430 5370 4440 5390
rect 4240 5360 4440 5370
rect 4480 5390 4680 5400
rect 4480 5370 4490 5390
rect 4510 5370 4570 5390
rect 4590 5370 4650 5390
rect 4670 5370 4680 5390
rect 4480 5360 4680 5370
rect 4720 5390 5720 5400
rect 4720 5370 4730 5390
rect 4750 5370 4810 5390
rect 4830 5370 4890 5390
rect 4910 5370 4970 5390
rect 4990 5370 5050 5390
rect 5070 5370 5130 5390
rect 5150 5370 5210 5390
rect 5230 5370 5290 5390
rect 5310 5370 5370 5390
rect 5390 5370 5450 5390
rect 5470 5370 5530 5390
rect 5550 5370 5610 5390
rect 5630 5370 5690 5390
rect 5710 5370 5720 5390
rect 4720 5360 5720 5370
rect 5760 5390 5960 5400
rect 5760 5370 5770 5390
rect 5790 5370 5850 5390
rect 5870 5370 5930 5390
rect 5950 5370 5960 5390
rect 5760 5360 5960 5370
rect 6000 5390 6200 5400
rect 6000 5370 6010 5390
rect 6030 5370 6090 5390
rect 6110 5370 6170 5390
rect 6190 5370 6200 5390
rect 6000 5360 6200 5370
rect 4240 5310 4440 5320
rect 4240 5290 4250 5310
rect 4270 5290 4330 5310
rect 4350 5290 4410 5310
rect 4430 5290 4440 5310
rect 4240 5280 4440 5290
rect 4480 5310 4680 5320
rect 4480 5290 4490 5310
rect 4510 5290 4570 5310
rect 4590 5290 4650 5310
rect 4670 5290 4680 5310
rect 4480 5280 4680 5290
rect 4720 5310 5720 5320
rect 4720 5290 4730 5310
rect 4750 5290 4810 5310
rect 4830 5290 4890 5310
rect 4910 5290 4970 5310
rect 4990 5290 5050 5310
rect 5070 5290 5130 5310
rect 5150 5290 5210 5310
rect 5230 5290 5290 5310
rect 5310 5290 5370 5310
rect 5390 5290 5450 5310
rect 5470 5290 5530 5310
rect 5550 5290 5610 5310
rect 5630 5290 5690 5310
rect 5710 5290 5720 5310
rect 4720 5280 5720 5290
rect 5760 5310 5960 5320
rect 5760 5290 5770 5310
rect 5790 5290 5850 5310
rect 5870 5290 5930 5310
rect 5950 5290 5960 5310
rect 5760 5280 5960 5290
rect 6000 5310 6200 5320
rect 6000 5290 6010 5310
rect 6030 5290 6090 5310
rect 6110 5290 6170 5310
rect 6190 5290 6200 5310
rect 6000 5280 6200 5290
rect 4240 5230 4440 5240
rect 4240 5210 4250 5230
rect 4270 5210 4330 5230
rect 4350 5210 4410 5230
rect 4430 5210 4440 5230
rect 4240 5200 4440 5210
rect 4480 5230 4680 5240
rect 4480 5210 4490 5230
rect 4510 5210 4570 5230
rect 4590 5210 4650 5230
rect 4670 5210 4680 5230
rect 4480 5200 4680 5210
rect 4720 5230 5720 5240
rect 4720 5210 4730 5230
rect 4750 5210 4810 5230
rect 4830 5210 4890 5230
rect 4910 5210 4970 5230
rect 4990 5210 5050 5230
rect 5070 5210 5130 5230
rect 5150 5210 5210 5230
rect 5230 5210 5290 5230
rect 5310 5210 5370 5230
rect 5390 5210 5450 5230
rect 5470 5210 5530 5230
rect 5550 5210 5610 5230
rect 5630 5210 5690 5230
rect 5710 5210 5720 5230
rect 4720 5200 5720 5210
rect 5760 5230 5960 5240
rect 5760 5210 5770 5230
rect 5790 5210 5850 5230
rect 5870 5210 5930 5230
rect 5950 5210 5960 5230
rect 5760 5200 5960 5210
rect 6000 5230 6200 5240
rect 6000 5210 6010 5230
rect 6030 5210 6090 5230
rect 6110 5210 6170 5230
rect 6190 5210 6200 5230
rect 6000 5200 6200 5210
rect 4240 5150 4440 5160
rect 4240 5130 4250 5150
rect 4270 5130 4330 5150
rect 4350 5130 4410 5150
rect 4430 5130 4440 5150
rect 4240 5120 4440 5130
rect 4480 5150 4680 5160
rect 4480 5130 4490 5150
rect 4510 5130 4570 5150
rect 4590 5130 4650 5150
rect 4670 5130 4680 5150
rect 4480 5120 4680 5130
rect 4720 5150 5720 5160
rect 4720 5130 4730 5150
rect 4750 5130 4810 5150
rect 4830 5130 4890 5150
rect 4910 5130 4970 5150
rect 4990 5130 5050 5150
rect 5070 5130 5130 5150
rect 5150 5130 5210 5150
rect 5230 5130 5290 5150
rect 5310 5130 5370 5150
rect 5390 5130 5450 5150
rect 5470 5130 5530 5150
rect 5550 5130 5610 5150
rect 5630 5130 5690 5150
rect 5710 5130 5720 5150
rect 4720 5120 5720 5130
rect 5760 5150 5960 5160
rect 5760 5130 5770 5150
rect 5790 5130 5850 5150
rect 5870 5130 5930 5150
rect 5950 5130 5960 5150
rect 5760 5120 5960 5130
rect 6000 5150 6200 5160
rect 6000 5130 6010 5150
rect 6030 5130 6090 5150
rect 6110 5130 6170 5150
rect 6190 5130 6200 5150
rect 6000 5120 6200 5130
rect 4240 5070 4440 5080
rect 4240 5050 4250 5070
rect 4270 5050 4330 5070
rect 4350 5050 4410 5070
rect 4430 5050 4440 5070
rect 4240 5040 4440 5050
rect 4480 5070 4680 5080
rect 4480 5050 4490 5070
rect 4510 5050 4570 5070
rect 4590 5050 4650 5070
rect 4670 5050 4680 5070
rect 4480 5040 4680 5050
rect 4720 5070 5720 5080
rect 4720 5050 4730 5070
rect 4750 5050 4810 5070
rect 4830 5050 4890 5070
rect 4910 5050 4970 5070
rect 4990 5050 5050 5070
rect 5070 5050 5130 5070
rect 5150 5050 5210 5070
rect 5230 5050 5290 5070
rect 5310 5050 5370 5070
rect 5390 5050 5450 5070
rect 5470 5050 5530 5070
rect 5550 5050 5610 5070
rect 5630 5050 5690 5070
rect 5710 5050 5720 5070
rect 4720 5040 5720 5050
rect 5760 5070 5960 5080
rect 5760 5050 5770 5070
rect 5790 5050 5850 5070
rect 5870 5050 5930 5070
rect 5950 5050 5960 5070
rect 5760 5040 5960 5050
rect 6000 5070 6200 5080
rect 6000 5050 6010 5070
rect 6030 5050 6090 5070
rect 6110 5050 6170 5070
rect 6190 5050 6200 5070
rect 6000 5040 6200 5050
rect 4240 4990 4440 5000
rect 4240 4970 4250 4990
rect 4270 4970 4330 4990
rect 4350 4970 4410 4990
rect 4430 4970 4440 4990
rect 4240 4960 4440 4970
rect 4480 4990 4680 5000
rect 4480 4970 4490 4990
rect 4510 4970 4570 4990
rect 4590 4970 4650 4990
rect 4670 4970 4680 4990
rect 4480 4960 4680 4970
rect 4720 4990 5720 5000
rect 4720 4970 4730 4990
rect 4750 4970 4810 4990
rect 4830 4970 4890 4990
rect 4910 4970 4970 4990
rect 4990 4970 5050 4990
rect 5070 4970 5130 4990
rect 5150 4970 5210 4990
rect 5230 4970 5290 4990
rect 5310 4970 5370 4990
rect 5390 4970 5450 4990
rect 5470 4970 5530 4990
rect 5550 4970 5610 4990
rect 5630 4970 5690 4990
rect 5710 4970 5720 4990
rect 4720 4960 5720 4970
rect 5760 4990 5960 5000
rect 5760 4970 5770 4990
rect 5790 4970 5850 4990
rect 5870 4970 5930 4990
rect 5950 4970 5960 4990
rect 5760 4960 5960 4970
rect 6000 4990 6200 5000
rect 6000 4970 6010 4990
rect 6030 4970 6090 4990
rect 6110 4970 6170 4990
rect 6190 4970 6200 4990
rect 6000 4960 6200 4970
rect 4240 4910 4440 4920
rect 4240 4890 4250 4910
rect 4270 4890 4330 4910
rect 4350 4890 4410 4910
rect 4430 4890 4440 4910
rect 4240 4880 4440 4890
rect 4480 4910 4680 4920
rect 4480 4890 4490 4910
rect 4510 4890 4570 4910
rect 4590 4890 4650 4910
rect 4670 4890 4680 4910
rect 4480 4880 4680 4890
rect 4720 4910 5720 4920
rect 4720 4890 4730 4910
rect 4750 4890 4810 4910
rect 4830 4890 4890 4910
rect 4910 4890 4970 4910
rect 4990 4890 5050 4910
rect 5070 4890 5130 4910
rect 5150 4890 5210 4910
rect 5230 4890 5290 4910
rect 5310 4890 5370 4910
rect 5390 4890 5450 4910
rect 5470 4890 5530 4910
rect 5550 4890 5610 4910
rect 5630 4890 5690 4910
rect 5710 4890 5720 4910
rect 4720 4880 5720 4890
rect 5760 4910 5960 4920
rect 5760 4890 5770 4910
rect 5790 4890 5850 4910
rect 5870 4890 5930 4910
rect 5950 4890 5960 4910
rect 5760 4880 5960 4890
rect 6000 4910 6200 4920
rect 6000 4890 6010 4910
rect 6030 4890 6090 4910
rect 6110 4890 6170 4910
rect 6190 4890 6200 4910
rect 6000 4880 6200 4890
rect 4240 4830 4440 4840
rect 4240 4810 4250 4830
rect 4270 4810 4330 4830
rect 4350 4810 4410 4830
rect 4430 4810 4440 4830
rect 4240 4800 4440 4810
rect 4480 4830 4680 4840
rect 4480 4810 4490 4830
rect 4510 4810 4570 4830
rect 4590 4810 4650 4830
rect 4670 4810 4680 4830
rect 4480 4800 4680 4810
rect 4720 4830 5720 4840
rect 4720 4810 4730 4830
rect 4750 4810 4810 4830
rect 4830 4810 4890 4830
rect 4910 4810 4970 4830
rect 4990 4810 5050 4830
rect 5070 4810 5130 4830
rect 5150 4810 5210 4830
rect 5230 4810 5290 4830
rect 5310 4810 5370 4830
rect 5390 4810 5450 4830
rect 5470 4810 5530 4830
rect 5550 4810 5610 4830
rect 5630 4810 5690 4830
rect 5710 4810 5720 4830
rect 4720 4800 5720 4810
rect 5760 4830 5960 4840
rect 5760 4810 5770 4830
rect 5790 4810 5850 4830
rect 5870 4810 5930 4830
rect 5950 4810 5960 4830
rect 5760 4800 5960 4810
rect 6000 4830 6200 4840
rect 6000 4810 6010 4830
rect 6030 4810 6090 4830
rect 6110 4810 6170 4830
rect 6190 4810 6200 4830
rect 6000 4800 6200 4810
rect 4240 4750 4440 4760
rect 4240 4730 4250 4750
rect 4270 4730 4330 4750
rect 4350 4730 4410 4750
rect 4430 4730 4440 4750
rect 4240 4720 4440 4730
rect 4480 4750 4680 4760
rect 4480 4730 4490 4750
rect 4510 4730 4570 4750
rect 4590 4730 4650 4750
rect 4670 4730 4680 4750
rect 4480 4720 4680 4730
rect 4720 4750 5720 4760
rect 4720 4730 4730 4750
rect 4750 4730 4810 4750
rect 4830 4730 4890 4750
rect 4910 4730 4970 4750
rect 4990 4730 5050 4750
rect 5070 4730 5130 4750
rect 5150 4730 5210 4750
rect 5230 4730 5290 4750
rect 5310 4730 5370 4750
rect 5390 4730 5450 4750
rect 5470 4730 5530 4750
rect 5550 4730 5610 4750
rect 5630 4730 5690 4750
rect 5710 4730 5720 4750
rect 4720 4720 5720 4730
rect 5760 4750 5960 4760
rect 5760 4730 5770 4750
rect 5790 4730 5850 4750
rect 5870 4730 5930 4750
rect 5950 4730 5960 4750
rect 5760 4720 5960 4730
rect 6000 4750 6200 4760
rect 6000 4730 6010 4750
rect 6030 4730 6090 4750
rect 6110 4730 6170 4750
rect 6190 4730 6200 4750
rect 6000 4720 6200 4730
rect 4240 4670 4440 4680
rect 4240 4650 4250 4670
rect 4270 4650 4330 4670
rect 4350 4650 4410 4670
rect 4430 4650 4440 4670
rect 4240 4640 4440 4650
rect 4480 4670 4680 4680
rect 4480 4650 4490 4670
rect 4510 4650 4570 4670
rect 4590 4650 4650 4670
rect 4670 4650 4680 4670
rect 4480 4640 4680 4650
rect 4720 4670 5720 4680
rect 4720 4650 4730 4670
rect 4750 4650 4810 4670
rect 4830 4650 4890 4670
rect 4910 4650 4970 4670
rect 4990 4650 5050 4670
rect 5070 4650 5130 4670
rect 5150 4650 5210 4670
rect 5230 4650 5290 4670
rect 5310 4650 5370 4670
rect 5390 4650 5450 4670
rect 5470 4650 5530 4670
rect 5550 4650 5610 4670
rect 5630 4650 5690 4670
rect 5710 4650 5720 4670
rect 4720 4640 5720 4650
rect 5760 4670 5960 4680
rect 5760 4650 5770 4670
rect 5790 4650 5850 4670
rect 5870 4650 5930 4670
rect 5950 4650 5960 4670
rect 5760 4640 5960 4650
rect 6000 4670 6200 4680
rect 6000 4650 6010 4670
rect 6030 4650 6090 4670
rect 6110 4650 6170 4670
rect 6190 4650 6200 4670
rect 6000 4640 6200 4650
rect 4240 4590 4440 4600
rect 4240 4570 4250 4590
rect 4270 4570 4330 4590
rect 4350 4570 4410 4590
rect 4430 4570 4440 4590
rect 4240 4560 4440 4570
rect 4480 4590 4680 4600
rect 4480 4570 4490 4590
rect 4510 4570 4570 4590
rect 4590 4570 4650 4590
rect 4670 4570 4680 4590
rect 4480 4560 4680 4570
rect 4720 4590 5720 4600
rect 4720 4570 4730 4590
rect 4750 4570 4810 4590
rect 4830 4570 4890 4590
rect 4910 4570 4970 4590
rect 4990 4570 5050 4590
rect 5070 4570 5130 4590
rect 5150 4570 5210 4590
rect 5230 4570 5290 4590
rect 5310 4570 5370 4590
rect 5390 4570 5450 4590
rect 5470 4570 5530 4590
rect 5550 4570 5610 4590
rect 5630 4570 5690 4590
rect 5710 4570 5720 4590
rect 4720 4560 5720 4570
rect 5760 4590 5960 4600
rect 5760 4570 5770 4590
rect 5790 4570 5850 4590
rect 5870 4570 5930 4590
rect 5950 4570 5960 4590
rect 5760 4560 5960 4570
rect 6000 4590 6200 4600
rect 6000 4570 6010 4590
rect 6030 4570 6090 4590
rect 6110 4570 6170 4590
rect 6190 4570 6200 4590
rect 6000 4560 6200 4570
rect 4240 4510 4440 4520
rect 4240 4490 4250 4510
rect 4270 4490 4330 4510
rect 4350 4490 4410 4510
rect 4430 4490 4440 4510
rect 4240 4480 4440 4490
rect 4480 4510 4680 4520
rect 4480 4490 4490 4510
rect 4510 4490 4570 4510
rect 4590 4490 4650 4510
rect 4670 4490 4680 4510
rect 4480 4480 4680 4490
rect 4720 4510 5720 4520
rect 4720 4490 4730 4510
rect 4750 4490 4810 4510
rect 4830 4490 4890 4510
rect 4910 4490 4970 4510
rect 4990 4490 5050 4510
rect 5070 4490 5130 4510
rect 5150 4490 5210 4510
rect 5230 4490 5290 4510
rect 5310 4490 5370 4510
rect 5390 4490 5450 4510
rect 5470 4490 5530 4510
rect 5550 4490 5610 4510
rect 5630 4490 5690 4510
rect 5710 4490 5720 4510
rect 4720 4480 5720 4490
rect 5760 4510 5960 4520
rect 5760 4490 5770 4510
rect 5790 4490 5850 4510
rect 5870 4490 5930 4510
rect 5950 4490 5960 4510
rect 5760 4480 5960 4490
rect 6000 4510 6200 4520
rect 6000 4490 6010 4510
rect 6030 4490 6090 4510
rect 6110 4490 6170 4510
rect 6190 4490 6200 4510
rect 6000 4480 6200 4490
rect 4240 4430 4440 4440
rect 4240 4410 4250 4430
rect 4270 4410 4330 4430
rect 4350 4410 4410 4430
rect 4430 4410 4440 4430
rect 4240 4400 4440 4410
rect 4480 4430 4680 4440
rect 4480 4410 4490 4430
rect 4510 4410 4570 4430
rect 4590 4410 4650 4430
rect 4670 4410 4680 4430
rect 4480 4400 4680 4410
rect 4720 4430 5720 4440
rect 4720 4410 4730 4430
rect 4750 4410 4810 4430
rect 4830 4410 4890 4430
rect 4910 4410 4970 4430
rect 4990 4410 5050 4430
rect 5070 4410 5130 4430
rect 5150 4410 5210 4430
rect 5230 4410 5290 4430
rect 5310 4410 5370 4430
rect 5390 4410 5450 4430
rect 5470 4410 5530 4430
rect 5550 4410 5610 4430
rect 5630 4410 5690 4430
rect 5710 4410 5720 4430
rect 4720 4400 5720 4410
rect 5760 4430 5960 4440
rect 5760 4410 5770 4430
rect 5790 4410 5850 4430
rect 5870 4410 5930 4430
rect 5950 4410 5960 4430
rect 5760 4400 5960 4410
rect 6000 4430 6200 4440
rect 6000 4410 6010 4430
rect 6030 4410 6090 4430
rect 6110 4410 6170 4430
rect 6190 4410 6200 4430
rect 6000 4400 6200 4410
rect 4240 4350 4440 4360
rect 4240 4330 4250 4350
rect 4270 4330 4330 4350
rect 4350 4330 4410 4350
rect 4430 4330 4440 4350
rect 4240 4320 4440 4330
rect 4480 4350 4680 4360
rect 4480 4330 4490 4350
rect 4510 4330 4570 4350
rect 4590 4330 4650 4350
rect 4670 4330 4680 4350
rect 4480 4320 4680 4330
rect 4720 4350 5720 4360
rect 4720 4330 4730 4350
rect 4750 4330 4810 4350
rect 4830 4330 4890 4350
rect 4910 4330 4970 4350
rect 4990 4330 5050 4350
rect 5070 4330 5130 4350
rect 5150 4330 5210 4350
rect 5230 4330 5290 4350
rect 5310 4330 5370 4350
rect 5390 4330 5450 4350
rect 5470 4330 5530 4350
rect 5550 4330 5610 4350
rect 5630 4330 5690 4350
rect 5710 4330 5720 4350
rect 4720 4320 5720 4330
rect 5760 4350 5960 4360
rect 5760 4330 5770 4350
rect 5790 4330 5850 4350
rect 5870 4330 5930 4350
rect 5950 4330 5960 4350
rect 5760 4320 5960 4330
rect 6000 4350 6200 4360
rect 6000 4330 6010 4350
rect 6030 4330 6090 4350
rect 6110 4330 6170 4350
rect 6190 4330 6200 4350
rect 6000 4320 6200 4330
rect 4240 4270 4440 4280
rect 4240 4250 4250 4270
rect 4270 4250 4330 4270
rect 4350 4250 4410 4270
rect 4430 4250 4440 4270
rect 4240 4240 4440 4250
rect 4480 4270 4680 4280
rect 4480 4250 4490 4270
rect 4510 4250 4570 4270
rect 4590 4250 4650 4270
rect 4670 4250 4680 4270
rect 4480 4240 4680 4250
rect 4720 4270 5720 4280
rect 4720 4250 4730 4270
rect 4750 4250 4810 4270
rect 4830 4250 4890 4270
rect 4910 4250 4970 4270
rect 4990 4250 5050 4270
rect 5070 4250 5130 4270
rect 5150 4250 5210 4270
rect 5230 4250 5290 4270
rect 5310 4250 5370 4270
rect 5390 4250 5450 4270
rect 5470 4250 5530 4270
rect 5550 4250 5610 4270
rect 5630 4250 5690 4270
rect 5710 4250 5720 4270
rect 4720 4240 5720 4250
rect 5760 4270 5960 4280
rect 5760 4250 5770 4270
rect 5790 4250 5850 4270
rect 5870 4250 5930 4270
rect 5950 4250 5960 4270
rect 5760 4240 5960 4250
rect 6000 4270 6200 4280
rect 6000 4250 6010 4270
rect 6030 4250 6090 4270
rect 6110 4250 6170 4270
rect 6190 4250 6200 4270
rect 6000 4240 6200 4250
rect 4240 4190 4440 4200
rect 4240 4170 4250 4190
rect 4270 4170 4330 4190
rect 4350 4170 4410 4190
rect 4430 4170 4440 4190
rect 4240 4160 4440 4170
rect 4480 4190 4680 4200
rect 4480 4170 4490 4190
rect 4510 4170 4570 4190
rect 4590 4170 4650 4190
rect 4670 4170 4680 4190
rect 4480 4160 4680 4170
rect 4720 4190 5720 4200
rect 4720 4170 4730 4190
rect 4750 4170 4810 4190
rect 4830 4170 4890 4190
rect 4910 4170 4970 4190
rect 4990 4170 5050 4190
rect 5070 4170 5130 4190
rect 5150 4170 5210 4190
rect 5230 4170 5290 4190
rect 5310 4170 5370 4190
rect 5390 4170 5450 4190
rect 5470 4170 5530 4190
rect 5550 4170 5610 4190
rect 5630 4170 5690 4190
rect 5710 4170 5720 4190
rect 4720 4160 5720 4170
rect 5760 4190 5960 4200
rect 5760 4170 5770 4190
rect 5790 4170 5850 4190
rect 5870 4170 5930 4190
rect 5950 4170 5960 4190
rect 5760 4160 5960 4170
rect 6000 4190 6200 4200
rect 6000 4170 6010 4190
rect 6030 4170 6090 4190
rect 6110 4170 6170 4190
rect 6190 4170 6200 4190
rect 6000 4160 6200 4170
rect 4240 4110 4440 4120
rect 4240 4090 4250 4110
rect 4270 4090 4330 4110
rect 4350 4090 4410 4110
rect 4430 4090 4440 4110
rect 4240 4080 4440 4090
rect 4480 4110 4680 4120
rect 4480 4090 4490 4110
rect 4510 4090 4570 4110
rect 4590 4090 4650 4110
rect 4670 4090 4680 4110
rect 4480 4080 4680 4090
rect 4720 4110 5720 4120
rect 4720 4090 4730 4110
rect 4750 4090 4810 4110
rect 4830 4090 4890 4110
rect 4910 4090 4970 4110
rect 4990 4090 5050 4110
rect 5070 4090 5130 4110
rect 5150 4090 5210 4110
rect 5230 4090 5290 4110
rect 5310 4090 5370 4110
rect 5390 4090 5450 4110
rect 5470 4090 5530 4110
rect 5550 4090 5610 4110
rect 5630 4090 5690 4110
rect 5710 4090 5720 4110
rect 4720 4080 5720 4090
rect 5760 4110 5960 4120
rect 5760 4090 5770 4110
rect 5790 4090 5850 4110
rect 5870 4090 5930 4110
rect 5950 4090 5960 4110
rect 5760 4080 5960 4090
rect 6000 4110 6200 4120
rect 6000 4090 6010 4110
rect 6030 4090 6090 4110
rect 6110 4090 6170 4110
rect 6190 4090 6200 4110
rect 6000 4080 6200 4090
rect 4240 4030 4440 4040
rect 4240 4010 4250 4030
rect 4270 4010 4330 4030
rect 4350 4010 4410 4030
rect 4430 4010 4440 4030
rect 4240 4000 4440 4010
rect 4480 4030 4680 4040
rect 4480 4010 4490 4030
rect 4510 4010 4570 4030
rect 4590 4010 4650 4030
rect 4670 4010 4680 4030
rect 4480 4000 4680 4010
rect 4720 4030 5720 4040
rect 4720 4010 4730 4030
rect 4750 4010 4810 4030
rect 4830 4010 4890 4030
rect 4910 4010 4970 4030
rect 4990 4010 5050 4030
rect 5070 4010 5130 4030
rect 5150 4010 5210 4030
rect 5230 4010 5290 4030
rect 5310 4010 5370 4030
rect 5390 4010 5450 4030
rect 5470 4010 5530 4030
rect 5550 4010 5610 4030
rect 5630 4010 5690 4030
rect 5710 4010 5720 4030
rect 4720 4000 5720 4010
rect 5760 4030 5960 4040
rect 5760 4010 5770 4030
rect 5790 4010 5850 4030
rect 5870 4010 5930 4030
rect 5950 4010 5960 4030
rect 5760 4000 5960 4010
rect 6000 4030 6200 4040
rect 6000 4010 6010 4030
rect 6030 4010 6090 4030
rect 6110 4010 6170 4030
rect 6190 4010 6200 4030
rect 6000 4000 6200 4010
rect 4240 3950 4440 3960
rect 4240 3930 4250 3950
rect 4270 3930 4330 3950
rect 4350 3930 4410 3950
rect 4430 3930 4440 3950
rect 4240 3920 4440 3930
rect 4480 3950 4680 3960
rect 4480 3930 4490 3950
rect 4510 3930 4570 3950
rect 4590 3930 4650 3950
rect 4670 3930 4680 3950
rect 4480 3920 4680 3930
rect 4720 3950 5720 3960
rect 4720 3930 4730 3950
rect 4750 3930 4810 3950
rect 4830 3930 4890 3950
rect 4910 3930 4970 3950
rect 4990 3930 5050 3950
rect 5070 3930 5130 3950
rect 5150 3930 5210 3950
rect 5230 3930 5290 3950
rect 5310 3930 5370 3950
rect 5390 3930 5450 3950
rect 5470 3930 5530 3950
rect 5550 3930 5610 3950
rect 5630 3930 5690 3950
rect 5710 3930 5720 3950
rect 4720 3920 5720 3930
rect 5760 3950 5960 3960
rect 5760 3930 5770 3950
rect 5790 3930 5850 3950
rect 5870 3930 5930 3950
rect 5950 3930 5960 3950
rect 5760 3920 5960 3930
rect 6000 3950 6200 3960
rect 6000 3930 6010 3950
rect 6030 3930 6090 3950
rect 6110 3930 6170 3950
rect 6190 3930 6200 3950
rect 6000 3920 6200 3930
rect 4240 3870 4440 3880
rect 4240 3850 4250 3870
rect 4270 3850 4330 3870
rect 4350 3850 4410 3870
rect 4430 3850 4440 3870
rect 4240 3840 4440 3850
rect 4480 3870 4680 3880
rect 4480 3850 4490 3870
rect 4510 3850 4570 3870
rect 4590 3850 4650 3870
rect 4670 3850 4680 3870
rect 4480 3840 4680 3850
rect 4720 3870 5720 3880
rect 4720 3850 4730 3870
rect 4750 3850 4810 3870
rect 4830 3850 4890 3870
rect 4910 3850 4970 3870
rect 4990 3850 5050 3870
rect 5070 3850 5130 3870
rect 5150 3850 5210 3870
rect 5230 3850 5290 3870
rect 5310 3850 5370 3870
rect 5390 3850 5450 3870
rect 5470 3850 5530 3870
rect 5550 3850 5610 3870
rect 5630 3850 5690 3870
rect 5710 3850 5720 3870
rect 4720 3840 5720 3850
rect 5760 3870 5960 3880
rect 5760 3850 5770 3870
rect 5790 3850 5850 3870
rect 5870 3850 5930 3870
rect 5950 3850 5960 3870
rect 5760 3840 5960 3850
rect 6000 3870 6200 3880
rect 6000 3850 6010 3870
rect 6030 3850 6090 3870
rect 6110 3850 6170 3870
rect 6190 3850 6200 3870
rect 6000 3840 6200 3850
rect 4240 3790 4440 3800
rect 4240 3770 4250 3790
rect 4270 3770 4330 3790
rect 4350 3770 4410 3790
rect 4430 3770 4440 3790
rect 4240 3760 4440 3770
rect 4480 3790 4680 3800
rect 4480 3770 4490 3790
rect 4510 3770 4570 3790
rect 4590 3770 4650 3790
rect 4670 3770 4680 3790
rect 4480 3760 4680 3770
rect 4720 3790 5720 3800
rect 4720 3770 4730 3790
rect 4750 3770 4810 3790
rect 4830 3770 4890 3790
rect 4910 3770 4970 3790
rect 4990 3770 5050 3790
rect 5070 3770 5130 3790
rect 5150 3770 5210 3790
rect 5230 3770 5290 3790
rect 5310 3770 5370 3790
rect 5390 3770 5450 3790
rect 5470 3770 5530 3790
rect 5550 3770 5610 3790
rect 5630 3770 5690 3790
rect 5710 3770 5720 3790
rect 4720 3760 5720 3770
rect 5760 3790 5960 3800
rect 5760 3770 5770 3790
rect 5790 3770 5850 3790
rect 5870 3770 5930 3790
rect 5950 3770 5960 3790
rect 5760 3760 5960 3770
rect 6000 3790 6200 3800
rect 6000 3770 6010 3790
rect 6030 3770 6090 3790
rect 6110 3770 6170 3790
rect 6190 3770 6200 3790
rect 6000 3760 6200 3770
rect 4240 3710 4440 3720
rect 4240 3690 4250 3710
rect 4270 3690 4330 3710
rect 4350 3690 4410 3710
rect 4430 3690 4440 3710
rect 4240 3680 4440 3690
rect 4480 3710 4680 3720
rect 4480 3690 4490 3710
rect 4510 3690 4570 3710
rect 4590 3690 4650 3710
rect 4670 3690 4680 3710
rect 4480 3680 4680 3690
rect 4720 3710 5720 3720
rect 4720 3690 4730 3710
rect 4750 3690 4810 3710
rect 4830 3690 4890 3710
rect 4910 3690 4970 3710
rect 4990 3690 5050 3710
rect 5070 3690 5130 3710
rect 5150 3690 5210 3710
rect 5230 3690 5290 3710
rect 5310 3690 5370 3710
rect 5390 3690 5450 3710
rect 5470 3690 5530 3710
rect 5550 3690 5610 3710
rect 5630 3690 5690 3710
rect 5710 3690 5720 3710
rect 4720 3680 5720 3690
rect 5760 3710 5960 3720
rect 5760 3690 5770 3710
rect 5790 3690 5850 3710
rect 5870 3690 5930 3710
rect 5950 3690 5960 3710
rect 5760 3680 5960 3690
rect 6000 3710 6200 3720
rect 6000 3690 6010 3710
rect 6030 3690 6090 3710
rect 6110 3690 6170 3710
rect 6190 3690 6200 3710
rect 6000 3680 6200 3690
rect 4240 3630 4440 3640
rect 4240 3610 4250 3630
rect 4270 3610 4330 3630
rect 4350 3610 4410 3630
rect 4430 3610 4440 3630
rect 4240 3600 4440 3610
rect 4480 3630 4680 3640
rect 4480 3610 4490 3630
rect 4510 3610 4570 3630
rect 4590 3610 4650 3630
rect 4670 3610 4680 3630
rect 4480 3600 4680 3610
rect 4720 3630 5720 3640
rect 4720 3610 4730 3630
rect 4750 3610 4810 3630
rect 4830 3610 4890 3630
rect 4910 3610 4970 3630
rect 4990 3610 5050 3630
rect 5070 3610 5130 3630
rect 5150 3610 5210 3630
rect 5230 3610 5290 3630
rect 5310 3610 5370 3630
rect 5390 3610 5450 3630
rect 5470 3610 5530 3630
rect 5550 3610 5610 3630
rect 5630 3610 5690 3630
rect 5710 3610 5720 3630
rect 4720 3600 5720 3610
rect 5760 3630 5960 3640
rect 5760 3610 5770 3630
rect 5790 3610 5850 3630
rect 5870 3610 5930 3630
rect 5950 3610 5960 3630
rect 5760 3600 5960 3610
rect 6000 3630 6200 3640
rect 6000 3610 6010 3630
rect 6030 3610 6090 3630
rect 6110 3610 6170 3630
rect 6190 3610 6200 3630
rect 6000 3600 6200 3610
rect 4240 3550 4440 3560
rect 4240 3530 4250 3550
rect 4270 3530 4330 3550
rect 4350 3530 4410 3550
rect 4430 3530 4440 3550
rect 4240 3520 4440 3530
rect 4480 3550 4680 3560
rect 4480 3530 4490 3550
rect 4510 3530 4570 3550
rect 4590 3530 4650 3550
rect 4670 3530 4680 3550
rect 4480 3520 4680 3530
rect 4720 3550 5720 3560
rect 4720 3530 4730 3550
rect 4750 3530 4810 3550
rect 4830 3530 4890 3550
rect 4910 3530 4970 3550
rect 4990 3530 5050 3550
rect 5070 3530 5130 3550
rect 5150 3530 5210 3550
rect 5230 3530 5290 3550
rect 5310 3530 5370 3550
rect 5390 3530 5450 3550
rect 5470 3530 5530 3550
rect 5550 3530 5610 3550
rect 5630 3530 5690 3550
rect 5710 3530 5720 3550
rect 4720 3520 5720 3530
rect 5760 3550 5960 3560
rect 5760 3530 5770 3550
rect 5790 3530 5850 3550
rect 5870 3530 5930 3550
rect 5950 3530 5960 3550
rect 5760 3520 5960 3530
rect 6000 3550 6200 3560
rect 6000 3530 6010 3550
rect 6030 3530 6090 3550
rect 6110 3530 6170 3550
rect 6190 3530 6200 3550
rect 6000 3520 6200 3530
rect 4240 3470 4440 3480
rect 4240 3450 4250 3470
rect 4270 3450 4330 3470
rect 4350 3450 4410 3470
rect 4430 3450 4440 3470
rect 4240 3440 4440 3450
rect 4480 3470 4680 3480
rect 4480 3450 4490 3470
rect 4510 3450 4570 3470
rect 4590 3450 4650 3470
rect 4670 3450 4680 3470
rect 4480 3440 4680 3450
rect 4720 3470 5720 3480
rect 4720 3450 4730 3470
rect 4750 3450 4810 3470
rect 4830 3450 4890 3470
rect 4910 3450 4970 3470
rect 4990 3450 5050 3470
rect 5070 3450 5130 3470
rect 5150 3450 5210 3470
rect 5230 3450 5290 3470
rect 5310 3450 5370 3470
rect 5390 3450 5450 3470
rect 5470 3450 5530 3470
rect 5550 3450 5610 3470
rect 5630 3450 5690 3470
rect 5710 3450 5720 3470
rect 4720 3440 5720 3450
rect 5760 3470 5960 3480
rect 5760 3450 5770 3470
rect 5790 3450 5850 3470
rect 5870 3450 5930 3470
rect 5950 3450 5960 3470
rect 5760 3440 5960 3450
rect 6000 3470 6200 3480
rect 6000 3450 6010 3470
rect 6030 3450 6090 3470
rect 6110 3450 6170 3470
rect 6190 3450 6200 3470
rect 6000 3440 6200 3450
rect 4240 3390 4440 3400
rect 4240 3370 4250 3390
rect 4270 3370 4330 3390
rect 4350 3370 4410 3390
rect 4430 3370 4440 3390
rect 4240 3360 4440 3370
rect 4480 3390 4680 3400
rect 4480 3370 4490 3390
rect 4510 3370 4570 3390
rect 4590 3370 4650 3390
rect 4670 3370 4680 3390
rect 4480 3360 4680 3370
rect 4720 3390 5720 3400
rect 4720 3370 4730 3390
rect 4750 3370 4810 3390
rect 4830 3370 4890 3390
rect 4910 3370 4970 3390
rect 4990 3370 5050 3390
rect 5070 3370 5130 3390
rect 5150 3370 5210 3390
rect 5230 3370 5290 3390
rect 5310 3370 5370 3390
rect 5390 3370 5450 3390
rect 5470 3370 5530 3390
rect 5550 3370 5610 3390
rect 5630 3370 5690 3390
rect 5710 3370 5720 3390
rect 4720 3360 5720 3370
rect 5760 3390 5960 3400
rect 5760 3370 5770 3390
rect 5790 3370 5850 3390
rect 5870 3370 5930 3390
rect 5950 3370 5960 3390
rect 5760 3360 5960 3370
rect 6000 3390 6200 3400
rect 6000 3370 6010 3390
rect 6030 3370 6090 3390
rect 6110 3370 6170 3390
rect 6190 3370 6200 3390
rect 6000 3360 6200 3370
rect 4240 3310 4440 3320
rect 4240 3290 4250 3310
rect 4270 3290 4330 3310
rect 4350 3290 4410 3310
rect 4430 3290 4440 3310
rect 4240 3280 4440 3290
rect 4480 3310 4680 3320
rect 4480 3290 4490 3310
rect 4510 3290 4570 3310
rect 4590 3290 4650 3310
rect 4670 3290 4680 3310
rect 4480 3280 4680 3290
rect 4720 3310 5720 3320
rect 4720 3290 4730 3310
rect 4750 3290 4810 3310
rect 4830 3290 4890 3310
rect 4910 3290 4970 3310
rect 4990 3290 5050 3310
rect 5070 3290 5130 3310
rect 5150 3290 5210 3310
rect 5230 3290 5290 3310
rect 5310 3290 5370 3310
rect 5390 3290 5450 3310
rect 5470 3290 5530 3310
rect 5550 3290 5610 3310
rect 5630 3290 5690 3310
rect 5710 3290 5720 3310
rect 4720 3280 5720 3290
rect 5760 3310 5960 3320
rect 5760 3290 5770 3310
rect 5790 3290 5850 3310
rect 5870 3290 5930 3310
rect 5950 3290 5960 3310
rect 5760 3280 5960 3290
rect 6000 3310 6200 3320
rect 6000 3290 6010 3310
rect 6030 3290 6090 3310
rect 6110 3290 6170 3310
rect 6190 3290 6200 3310
rect 6000 3280 6200 3290
rect 4240 3230 4440 3240
rect 4240 3210 4250 3230
rect 4270 3210 4330 3230
rect 4350 3210 4410 3230
rect 4430 3210 4440 3230
rect 4240 3200 4440 3210
rect 4480 3230 4680 3240
rect 4480 3210 4490 3230
rect 4510 3210 4570 3230
rect 4590 3210 4650 3230
rect 4670 3210 4680 3230
rect 4480 3200 4680 3210
rect 4720 3230 5720 3240
rect 4720 3210 4730 3230
rect 4750 3210 4810 3230
rect 4830 3210 4890 3230
rect 4910 3210 4970 3230
rect 4990 3210 5050 3230
rect 5070 3210 5130 3230
rect 5150 3210 5210 3230
rect 5230 3210 5290 3230
rect 5310 3210 5370 3230
rect 5390 3210 5450 3230
rect 5470 3210 5530 3230
rect 5550 3210 5610 3230
rect 5630 3210 5690 3230
rect 5710 3210 5720 3230
rect 4720 3200 5720 3210
rect 5760 3230 5960 3240
rect 5760 3210 5770 3230
rect 5790 3210 5850 3230
rect 5870 3210 5930 3230
rect 5950 3210 5960 3230
rect 5760 3200 5960 3210
rect 6000 3230 6200 3240
rect 6000 3210 6010 3230
rect 6030 3210 6090 3230
rect 6110 3210 6170 3230
rect 6190 3210 6200 3230
rect 6000 3200 6200 3210
rect 4240 3150 4440 3160
rect 4240 3130 4250 3150
rect 4270 3130 4330 3150
rect 4350 3130 4410 3150
rect 4430 3130 4440 3150
rect 4240 3120 4440 3130
rect 4480 3150 4680 3160
rect 4480 3130 4490 3150
rect 4510 3130 4570 3150
rect 4590 3130 4650 3150
rect 4670 3130 4680 3150
rect 4480 3120 4680 3130
rect 4720 3150 5720 3160
rect 4720 3130 4730 3150
rect 4750 3130 4810 3150
rect 4830 3130 4890 3150
rect 4910 3130 4970 3150
rect 4990 3130 5050 3150
rect 5070 3130 5130 3150
rect 5150 3130 5210 3150
rect 5230 3130 5290 3150
rect 5310 3130 5370 3150
rect 5390 3130 5450 3150
rect 5470 3130 5530 3150
rect 5550 3130 5610 3150
rect 5630 3130 5690 3150
rect 5710 3130 5720 3150
rect 4720 3120 5720 3130
rect 5760 3150 5960 3160
rect 5760 3130 5770 3150
rect 5790 3130 5850 3150
rect 5870 3130 5930 3150
rect 5950 3130 5960 3150
rect 5760 3120 5960 3130
rect 6000 3150 6200 3160
rect 6000 3130 6010 3150
rect 6030 3130 6090 3150
rect 6110 3130 6170 3150
rect 6190 3130 6200 3150
rect 6000 3120 6200 3130
rect 4240 3070 4440 3080
rect 4240 3050 4250 3070
rect 4270 3050 4330 3070
rect 4350 3050 4410 3070
rect 4430 3050 4440 3070
rect 4240 3040 4440 3050
rect 4480 3070 4680 3080
rect 4480 3050 4490 3070
rect 4510 3050 4570 3070
rect 4590 3050 4650 3070
rect 4670 3050 4680 3070
rect 4480 3040 4680 3050
rect 4720 3070 5720 3080
rect 4720 3050 4730 3070
rect 4750 3050 4810 3070
rect 4830 3050 4890 3070
rect 4910 3050 4970 3070
rect 4990 3050 5050 3070
rect 5070 3050 5130 3070
rect 5150 3050 5210 3070
rect 5230 3050 5290 3070
rect 5310 3050 5370 3070
rect 5390 3050 5450 3070
rect 5470 3050 5530 3070
rect 5550 3050 5610 3070
rect 5630 3050 5690 3070
rect 5710 3050 5720 3070
rect 4720 3040 5720 3050
rect 5760 3070 5960 3080
rect 5760 3050 5770 3070
rect 5790 3050 5850 3070
rect 5870 3050 5930 3070
rect 5950 3050 5960 3070
rect 5760 3040 5960 3050
rect 6000 3070 6200 3080
rect 6000 3050 6010 3070
rect 6030 3050 6090 3070
rect 6110 3050 6170 3070
rect 6190 3050 6200 3070
rect 6000 3040 6200 3050
rect 4240 2990 4440 3000
rect 4240 2970 4250 2990
rect 4270 2970 4330 2990
rect 4350 2970 4410 2990
rect 4430 2970 4440 2990
rect 4240 2960 4440 2970
rect 4480 2990 4680 3000
rect 4480 2970 4490 2990
rect 4510 2970 4570 2990
rect 4590 2970 4650 2990
rect 4670 2970 4680 2990
rect 4480 2960 4680 2970
rect 4720 2990 5720 3000
rect 4720 2970 4730 2990
rect 4750 2970 4810 2990
rect 4830 2970 4890 2990
rect 4910 2970 4970 2990
rect 4990 2970 5050 2990
rect 5070 2970 5130 2990
rect 5150 2970 5210 2990
rect 5230 2970 5290 2990
rect 5310 2970 5370 2990
rect 5390 2970 5450 2990
rect 5470 2970 5530 2990
rect 5550 2970 5610 2990
rect 5630 2970 5690 2990
rect 5710 2970 5720 2990
rect 4720 2960 5720 2970
rect 5760 2990 5960 3000
rect 5760 2970 5770 2990
rect 5790 2970 5850 2990
rect 5870 2970 5930 2990
rect 5950 2970 5960 2990
rect 5760 2960 5960 2970
rect 6000 2990 6200 3000
rect 6000 2970 6010 2990
rect 6030 2970 6090 2990
rect 6110 2970 6170 2990
rect 6190 2970 6200 2990
rect 6000 2960 6200 2970
rect 4240 2910 4440 2920
rect 4240 2890 4250 2910
rect 4270 2890 4330 2910
rect 4350 2890 4410 2910
rect 4430 2890 4440 2910
rect 4240 2880 4440 2890
rect 4480 2910 4680 2920
rect 4480 2890 4490 2910
rect 4510 2890 4570 2910
rect 4590 2890 4650 2910
rect 4670 2890 4680 2910
rect 4480 2880 4680 2890
rect 4720 2910 5720 2920
rect 4720 2890 4730 2910
rect 4750 2890 4810 2910
rect 4830 2890 4890 2910
rect 4910 2890 4970 2910
rect 4990 2890 5050 2910
rect 5070 2890 5130 2910
rect 5150 2890 5210 2910
rect 5230 2890 5290 2910
rect 5310 2890 5370 2910
rect 5390 2890 5450 2910
rect 5470 2890 5530 2910
rect 5550 2890 5610 2910
rect 5630 2890 5690 2910
rect 5710 2890 5720 2910
rect 4720 2880 5720 2890
rect 5760 2910 5960 2920
rect 5760 2890 5770 2910
rect 5790 2890 5850 2910
rect 5870 2890 5930 2910
rect 5950 2890 5960 2910
rect 5760 2880 5960 2890
rect 6000 2910 6200 2920
rect 6000 2890 6010 2910
rect 6030 2890 6090 2910
rect 6110 2890 6170 2910
rect 6190 2890 6200 2910
rect 6000 2880 6200 2890
rect 4240 2830 4440 2840
rect 4240 2810 4250 2830
rect 4270 2810 4330 2830
rect 4350 2810 4410 2830
rect 4430 2810 4440 2830
rect 4240 2800 4440 2810
rect 4480 2830 4680 2840
rect 4480 2810 4490 2830
rect 4510 2810 4570 2830
rect 4590 2810 4650 2830
rect 4670 2810 4680 2830
rect 4480 2800 4680 2810
rect 4720 2830 5720 2840
rect 4720 2810 4730 2830
rect 4750 2810 4810 2830
rect 4830 2810 4890 2830
rect 4910 2810 4970 2830
rect 4990 2810 5050 2830
rect 5070 2810 5130 2830
rect 5150 2810 5210 2830
rect 5230 2810 5290 2830
rect 5310 2810 5370 2830
rect 5390 2810 5450 2830
rect 5470 2810 5530 2830
rect 5550 2810 5610 2830
rect 5630 2810 5690 2830
rect 5710 2810 5720 2830
rect 4720 2800 5720 2810
rect 5760 2830 5960 2840
rect 5760 2810 5770 2830
rect 5790 2810 5850 2830
rect 5870 2810 5930 2830
rect 5950 2810 5960 2830
rect 5760 2800 5960 2810
rect 6000 2830 6200 2840
rect 6000 2810 6010 2830
rect 6030 2810 6090 2830
rect 6110 2810 6170 2830
rect 6190 2810 6200 2830
rect 6000 2800 6200 2810
rect 4240 2750 4440 2760
rect 4240 2730 4250 2750
rect 4270 2730 4330 2750
rect 4350 2730 4410 2750
rect 4430 2730 4440 2750
rect 4240 2720 4440 2730
rect 4480 2750 4680 2760
rect 4480 2730 4490 2750
rect 4510 2730 4570 2750
rect 4590 2730 4650 2750
rect 4670 2730 4680 2750
rect 4480 2720 4680 2730
rect 4720 2750 5720 2760
rect 4720 2730 4730 2750
rect 4750 2730 4810 2750
rect 4830 2730 4890 2750
rect 4910 2730 4970 2750
rect 4990 2730 5050 2750
rect 5070 2730 5130 2750
rect 5150 2730 5210 2750
rect 5230 2730 5290 2750
rect 5310 2730 5370 2750
rect 5390 2730 5450 2750
rect 5470 2730 5530 2750
rect 5550 2730 5610 2750
rect 5630 2730 5690 2750
rect 5710 2730 5720 2750
rect 4720 2720 5720 2730
rect 5760 2750 5960 2760
rect 5760 2730 5770 2750
rect 5790 2730 5850 2750
rect 5870 2730 5930 2750
rect 5950 2730 5960 2750
rect 5760 2720 5960 2730
rect 6000 2750 6200 2760
rect 6000 2730 6010 2750
rect 6030 2730 6090 2750
rect 6110 2730 6170 2750
rect 6190 2730 6200 2750
rect 6000 2720 6200 2730
rect 4240 2670 4440 2680
rect 4240 2650 4250 2670
rect 4270 2650 4330 2670
rect 4350 2650 4410 2670
rect 4430 2650 4440 2670
rect 4240 2640 4440 2650
rect 4480 2670 4680 2680
rect 4480 2650 4490 2670
rect 4510 2650 4570 2670
rect 4590 2650 4650 2670
rect 4670 2650 4680 2670
rect 4480 2640 4680 2650
rect 4720 2670 5720 2680
rect 4720 2650 4730 2670
rect 4750 2650 4810 2670
rect 4830 2650 4890 2670
rect 4910 2650 4970 2670
rect 4990 2650 5050 2670
rect 5070 2650 5130 2670
rect 5150 2650 5210 2670
rect 5230 2650 5290 2670
rect 5310 2650 5370 2670
rect 5390 2650 5450 2670
rect 5470 2650 5530 2670
rect 5550 2650 5610 2670
rect 5630 2650 5690 2670
rect 5710 2650 5720 2670
rect 4720 2640 5720 2650
rect 5760 2670 5960 2680
rect 5760 2650 5770 2670
rect 5790 2650 5850 2670
rect 5870 2650 5930 2670
rect 5950 2650 5960 2670
rect 5760 2640 5960 2650
rect 6000 2670 6200 2680
rect 6000 2650 6010 2670
rect 6030 2650 6090 2670
rect 6110 2650 6170 2670
rect 6190 2650 6200 2670
rect 6000 2640 6200 2650
rect 4240 2590 4440 2600
rect 4240 2570 4250 2590
rect 4270 2570 4330 2590
rect 4350 2570 4410 2590
rect 4430 2570 4440 2590
rect 4240 2560 4440 2570
rect 4480 2590 4680 2600
rect 4480 2570 4490 2590
rect 4510 2570 4570 2590
rect 4590 2570 4650 2590
rect 4670 2570 4680 2590
rect 4480 2560 4680 2570
rect 4720 2590 5720 2600
rect 4720 2570 4730 2590
rect 4750 2570 4810 2590
rect 4830 2570 4890 2590
rect 4910 2570 4970 2590
rect 4990 2570 5050 2590
rect 5070 2570 5130 2590
rect 5150 2570 5210 2590
rect 5230 2570 5290 2590
rect 5310 2570 5370 2590
rect 5390 2570 5450 2590
rect 5470 2570 5530 2590
rect 5550 2570 5610 2590
rect 5630 2570 5690 2590
rect 5710 2570 5720 2590
rect 4720 2560 5720 2570
rect 5760 2590 5960 2600
rect 5760 2570 5770 2590
rect 5790 2570 5850 2590
rect 5870 2570 5930 2590
rect 5950 2570 5960 2590
rect 5760 2560 5960 2570
rect 6000 2590 6200 2600
rect 6000 2570 6010 2590
rect 6030 2570 6090 2590
rect 6110 2570 6170 2590
rect 6190 2570 6200 2590
rect 6000 2560 6200 2570
rect 4240 2510 4440 2520
rect 4240 2490 4250 2510
rect 4270 2490 4330 2510
rect 4350 2490 4410 2510
rect 4430 2490 4440 2510
rect 4240 2480 4440 2490
rect 4480 2510 4680 2520
rect 4480 2490 4490 2510
rect 4510 2490 4570 2510
rect 4590 2490 4650 2510
rect 4670 2490 4680 2510
rect 4480 2480 4680 2490
rect 4720 2510 5720 2520
rect 4720 2490 4730 2510
rect 4750 2490 4810 2510
rect 4830 2490 4890 2510
rect 4910 2490 4970 2510
rect 4990 2490 5050 2510
rect 5070 2490 5130 2510
rect 5150 2490 5210 2510
rect 5230 2490 5290 2510
rect 5310 2490 5370 2510
rect 5390 2490 5450 2510
rect 5470 2490 5530 2510
rect 5550 2490 5610 2510
rect 5630 2490 5690 2510
rect 5710 2490 5720 2510
rect 4720 2480 5720 2490
rect 5760 2510 5960 2520
rect 5760 2490 5770 2510
rect 5790 2490 5850 2510
rect 5870 2490 5930 2510
rect 5950 2490 5960 2510
rect 5760 2480 5960 2490
rect 6000 2510 6200 2520
rect 6000 2490 6010 2510
rect 6030 2490 6090 2510
rect 6110 2490 6170 2510
rect 6190 2490 6200 2510
rect 6000 2480 6200 2490
rect 4240 2430 4440 2440
rect 4240 2410 4250 2430
rect 4270 2410 4330 2430
rect 4350 2410 4410 2430
rect 4430 2410 4440 2430
rect 4240 2400 4440 2410
rect 4480 2430 4680 2440
rect 4480 2410 4490 2430
rect 4510 2410 4570 2430
rect 4590 2410 4650 2430
rect 4670 2410 4680 2430
rect 4480 2400 4680 2410
rect 4720 2430 5720 2440
rect 4720 2410 4730 2430
rect 4750 2410 4810 2430
rect 4830 2410 4890 2430
rect 4910 2410 4970 2430
rect 4990 2410 5050 2430
rect 5070 2410 5130 2430
rect 5150 2410 5210 2430
rect 5230 2410 5290 2430
rect 5310 2410 5370 2430
rect 5390 2410 5450 2430
rect 5470 2410 5530 2430
rect 5550 2410 5610 2430
rect 5630 2410 5690 2430
rect 5710 2410 5720 2430
rect 4720 2400 5720 2410
rect 5760 2430 5960 2440
rect 5760 2410 5770 2430
rect 5790 2410 5850 2430
rect 5870 2410 5930 2430
rect 5950 2410 5960 2430
rect 5760 2400 5960 2410
rect 6000 2430 6200 2440
rect 6000 2410 6010 2430
rect 6030 2410 6090 2430
rect 6110 2410 6170 2430
rect 6190 2410 6200 2430
rect 6000 2400 6200 2410
rect 4240 2350 4440 2360
rect 4240 2330 4250 2350
rect 4270 2330 4330 2350
rect 4350 2330 4410 2350
rect 4430 2330 4440 2350
rect 4240 2320 4440 2330
rect 4480 2350 4680 2360
rect 4480 2330 4490 2350
rect 4510 2330 4570 2350
rect 4590 2330 4650 2350
rect 4670 2330 4680 2350
rect 4480 2320 4680 2330
rect 4720 2350 5720 2360
rect 4720 2330 4730 2350
rect 4750 2330 4810 2350
rect 4830 2330 4890 2350
rect 4910 2330 4970 2350
rect 4990 2330 5050 2350
rect 5070 2330 5130 2350
rect 5150 2330 5210 2350
rect 5230 2330 5290 2350
rect 5310 2330 5370 2350
rect 5390 2330 5450 2350
rect 5470 2330 5530 2350
rect 5550 2330 5610 2350
rect 5630 2330 5690 2350
rect 5710 2330 5720 2350
rect 4720 2320 5720 2330
rect 5760 2350 5960 2360
rect 5760 2330 5770 2350
rect 5790 2330 5850 2350
rect 5870 2330 5930 2350
rect 5950 2330 5960 2350
rect 5760 2320 5960 2330
rect 6000 2350 6200 2360
rect 6000 2330 6010 2350
rect 6030 2330 6090 2350
rect 6110 2330 6170 2350
rect 6190 2330 6200 2350
rect 6000 2320 6200 2330
rect 4240 2270 4440 2280
rect 4240 2250 4250 2270
rect 4270 2250 4330 2270
rect 4350 2250 4410 2270
rect 4430 2250 4440 2270
rect 4240 2240 4440 2250
rect 4480 2270 4680 2280
rect 4480 2250 4490 2270
rect 4510 2250 4570 2270
rect 4590 2250 4650 2270
rect 4670 2250 4680 2270
rect 4480 2240 4680 2250
rect 4720 2270 5720 2280
rect 4720 2250 4730 2270
rect 4750 2250 4810 2270
rect 4830 2250 4890 2270
rect 4910 2250 4970 2270
rect 4990 2250 5050 2270
rect 5070 2250 5130 2270
rect 5150 2250 5210 2270
rect 5230 2250 5290 2270
rect 5310 2250 5370 2270
rect 5390 2250 5450 2270
rect 5470 2250 5530 2270
rect 5550 2250 5610 2270
rect 5630 2250 5690 2270
rect 5710 2250 5720 2270
rect 4720 2240 5720 2250
rect 5760 2270 5960 2280
rect 5760 2250 5770 2270
rect 5790 2250 5850 2270
rect 5870 2250 5930 2270
rect 5950 2250 5960 2270
rect 5760 2240 5960 2250
rect 6000 2270 6200 2280
rect 6000 2250 6010 2270
rect 6030 2250 6090 2270
rect 6110 2250 6170 2270
rect 6190 2250 6200 2270
rect 6000 2240 6200 2250
rect 4240 2190 4440 2200
rect 4240 2170 4250 2190
rect 4270 2170 4330 2190
rect 4350 2170 4410 2190
rect 4430 2170 4440 2190
rect 4240 2160 4440 2170
rect 4480 2190 4680 2200
rect 4480 2170 4490 2190
rect 4510 2170 4570 2190
rect 4590 2170 4650 2190
rect 4670 2170 4680 2190
rect 4480 2160 4680 2170
rect 4720 2190 5720 2200
rect 4720 2170 4730 2190
rect 4750 2170 4810 2190
rect 4830 2170 4890 2190
rect 4910 2170 4970 2190
rect 4990 2170 5050 2190
rect 5070 2170 5130 2190
rect 5150 2170 5210 2190
rect 5230 2170 5290 2190
rect 5310 2170 5370 2190
rect 5390 2170 5450 2190
rect 5470 2170 5530 2190
rect 5550 2170 5610 2190
rect 5630 2170 5690 2190
rect 5710 2170 5720 2190
rect 4720 2160 5720 2170
rect 5760 2190 5960 2200
rect 5760 2170 5770 2190
rect 5790 2170 5850 2190
rect 5870 2170 5930 2190
rect 5950 2170 5960 2190
rect 5760 2160 5960 2170
rect 6000 2190 6200 2200
rect 6000 2170 6010 2190
rect 6030 2170 6090 2190
rect 6110 2170 6170 2190
rect 6190 2170 6200 2190
rect 6000 2160 6200 2170
rect 4240 2110 4440 2120
rect 4240 2090 4250 2110
rect 4270 2090 4330 2110
rect 4350 2090 4410 2110
rect 4430 2090 4440 2110
rect 4240 2080 4440 2090
rect 4480 2110 4680 2120
rect 4480 2090 4490 2110
rect 4510 2090 4570 2110
rect 4590 2090 4650 2110
rect 4670 2090 4680 2110
rect 4480 2080 4680 2090
rect 4720 2110 5720 2120
rect 4720 2090 4730 2110
rect 4750 2090 4810 2110
rect 4830 2090 4890 2110
rect 4910 2090 4970 2110
rect 4990 2090 5050 2110
rect 5070 2090 5130 2110
rect 5150 2090 5210 2110
rect 5230 2090 5290 2110
rect 5310 2090 5370 2110
rect 5390 2090 5450 2110
rect 5470 2090 5530 2110
rect 5550 2090 5610 2110
rect 5630 2090 5690 2110
rect 5710 2090 5720 2110
rect 4720 2080 5720 2090
rect 5760 2110 5960 2120
rect 5760 2090 5770 2110
rect 5790 2090 5850 2110
rect 5870 2090 5930 2110
rect 5950 2090 5960 2110
rect 5760 2080 5960 2090
rect 6000 2110 6200 2120
rect 6000 2090 6010 2110
rect 6030 2090 6090 2110
rect 6110 2090 6170 2110
rect 6190 2090 6200 2110
rect 6000 2080 6200 2090
rect 4240 2030 4440 2040
rect 4240 2010 4250 2030
rect 4270 2010 4330 2030
rect 4350 2010 4410 2030
rect 4430 2010 4440 2030
rect 4240 2000 4440 2010
rect 4480 2030 4680 2040
rect 4480 2010 4490 2030
rect 4510 2010 4570 2030
rect 4590 2010 4650 2030
rect 4670 2010 4680 2030
rect 4480 2000 4680 2010
rect 4720 2030 5720 2040
rect 4720 2010 4730 2030
rect 4750 2010 4810 2030
rect 4830 2010 4890 2030
rect 4910 2010 4970 2030
rect 4990 2010 5050 2030
rect 5070 2010 5130 2030
rect 5150 2010 5210 2030
rect 5230 2010 5290 2030
rect 5310 2010 5370 2030
rect 5390 2010 5450 2030
rect 5470 2010 5530 2030
rect 5550 2010 5610 2030
rect 5630 2010 5690 2030
rect 5710 2010 5720 2030
rect 4720 2000 5720 2010
rect 5760 2030 5960 2040
rect 5760 2010 5770 2030
rect 5790 2010 5850 2030
rect 5870 2010 5930 2030
rect 5950 2010 5960 2030
rect 5760 2000 5960 2010
rect 6000 2030 6200 2040
rect 6000 2010 6010 2030
rect 6030 2010 6090 2030
rect 6110 2010 6170 2030
rect 6190 2010 6200 2030
rect 6000 2000 6200 2010
rect 4240 1950 4440 1960
rect 4240 1930 4250 1950
rect 4270 1930 4330 1950
rect 4350 1930 4410 1950
rect 4430 1930 4440 1950
rect 4240 1920 4440 1930
rect 4480 1950 4680 1960
rect 4480 1930 4490 1950
rect 4510 1930 4570 1950
rect 4590 1930 4650 1950
rect 4670 1930 4680 1950
rect 4480 1920 4680 1930
rect 4720 1950 5720 1960
rect 4720 1930 4730 1950
rect 4750 1930 4810 1950
rect 4830 1930 4890 1950
rect 4910 1930 4970 1950
rect 4990 1930 5050 1950
rect 5070 1930 5130 1950
rect 5150 1930 5210 1950
rect 5230 1930 5290 1950
rect 5310 1930 5370 1950
rect 5390 1930 5450 1950
rect 5470 1930 5530 1950
rect 5550 1930 5610 1950
rect 5630 1930 5690 1950
rect 5710 1930 5720 1950
rect 4720 1920 5720 1930
rect 5760 1950 5960 1960
rect 5760 1930 5770 1950
rect 5790 1930 5850 1950
rect 5870 1930 5930 1950
rect 5950 1930 5960 1950
rect 5760 1920 5960 1930
rect 6000 1950 6200 1960
rect 6000 1930 6010 1950
rect 6030 1930 6090 1950
rect 6110 1930 6170 1950
rect 6190 1930 6200 1950
rect 6000 1920 6200 1930
rect 4240 1870 4440 1880
rect 4240 1850 4250 1870
rect 4270 1850 4330 1870
rect 4350 1850 4410 1870
rect 4430 1850 4440 1870
rect 4240 1840 4440 1850
rect 4480 1870 4680 1880
rect 4480 1850 4490 1870
rect 4510 1850 4570 1870
rect 4590 1850 4650 1870
rect 4670 1850 4680 1870
rect 4480 1840 4680 1850
rect 4720 1870 5720 1880
rect 4720 1850 4730 1870
rect 4750 1850 4810 1870
rect 4830 1850 4890 1870
rect 4910 1850 4970 1870
rect 4990 1850 5050 1870
rect 5070 1850 5130 1870
rect 5150 1850 5210 1870
rect 5230 1850 5290 1870
rect 5310 1850 5370 1870
rect 5390 1850 5450 1870
rect 5470 1850 5530 1870
rect 5550 1850 5610 1870
rect 5630 1850 5690 1870
rect 5710 1850 5720 1870
rect 4720 1840 5720 1850
rect 5760 1870 5960 1880
rect 5760 1850 5770 1870
rect 5790 1850 5850 1870
rect 5870 1850 5930 1870
rect 5950 1850 5960 1870
rect 5760 1840 5960 1850
rect 6000 1870 6200 1880
rect 6000 1850 6010 1870
rect 6030 1850 6090 1870
rect 6110 1850 6170 1870
rect 6190 1850 6200 1870
rect 6000 1840 6200 1850
rect 4240 1790 4440 1800
rect 4240 1770 4250 1790
rect 4270 1770 4330 1790
rect 4350 1770 4410 1790
rect 4430 1770 4440 1790
rect 4240 1760 4440 1770
rect 4480 1790 4680 1800
rect 4480 1770 4490 1790
rect 4510 1770 4570 1790
rect 4590 1770 4650 1790
rect 4670 1770 4680 1790
rect 4480 1760 4680 1770
rect 4720 1790 5720 1800
rect 4720 1770 4730 1790
rect 4750 1770 4810 1790
rect 4830 1770 4890 1790
rect 4910 1770 4970 1790
rect 4990 1770 5050 1790
rect 5070 1770 5130 1790
rect 5150 1770 5210 1790
rect 5230 1770 5290 1790
rect 5310 1770 5370 1790
rect 5390 1770 5450 1790
rect 5470 1770 5530 1790
rect 5550 1770 5610 1790
rect 5630 1770 5690 1790
rect 5710 1770 5720 1790
rect 4720 1760 5720 1770
rect 5760 1790 5960 1800
rect 5760 1770 5770 1790
rect 5790 1770 5850 1790
rect 5870 1770 5930 1790
rect 5950 1770 5960 1790
rect 5760 1760 5960 1770
rect 6000 1790 6200 1800
rect 6000 1770 6010 1790
rect 6030 1770 6090 1790
rect 6110 1770 6170 1790
rect 6190 1770 6200 1790
rect 6000 1760 6200 1770
rect 4240 1710 4440 1720
rect 4240 1690 4250 1710
rect 4270 1690 4330 1710
rect 4350 1690 4410 1710
rect 4430 1690 4440 1710
rect 4240 1680 4440 1690
rect 4480 1710 4680 1720
rect 4480 1690 4490 1710
rect 4510 1690 4570 1710
rect 4590 1690 4650 1710
rect 4670 1690 4680 1710
rect 4480 1680 4680 1690
rect 4720 1710 5720 1720
rect 4720 1690 4730 1710
rect 4750 1690 4810 1710
rect 4830 1690 4890 1710
rect 4910 1690 4970 1710
rect 4990 1690 5050 1710
rect 5070 1690 5130 1710
rect 5150 1690 5210 1710
rect 5230 1690 5290 1710
rect 5310 1690 5370 1710
rect 5390 1690 5450 1710
rect 5470 1690 5530 1710
rect 5550 1690 5610 1710
rect 5630 1690 5690 1710
rect 5710 1690 5720 1710
rect 4720 1680 5720 1690
rect 5760 1710 5960 1720
rect 5760 1690 5770 1710
rect 5790 1690 5850 1710
rect 5870 1690 5930 1710
rect 5950 1690 5960 1710
rect 5760 1680 5960 1690
rect 6000 1710 6200 1720
rect 6000 1690 6010 1710
rect 6030 1690 6090 1710
rect 6110 1690 6170 1710
rect 6190 1690 6200 1710
rect 6000 1680 6200 1690
rect 4240 1630 4440 1640
rect 4240 1610 4250 1630
rect 4270 1610 4330 1630
rect 4350 1610 4410 1630
rect 4430 1610 4440 1630
rect 4240 1600 4440 1610
rect 4480 1630 4680 1640
rect 4480 1610 4490 1630
rect 4510 1610 4570 1630
rect 4590 1610 4650 1630
rect 4670 1610 4680 1630
rect 4480 1600 4680 1610
rect 4720 1630 5720 1640
rect 4720 1610 4730 1630
rect 4750 1610 4810 1630
rect 4830 1610 4890 1630
rect 4910 1610 4970 1630
rect 4990 1610 5050 1630
rect 5070 1610 5130 1630
rect 5150 1610 5210 1630
rect 5230 1610 5290 1630
rect 5310 1610 5370 1630
rect 5390 1610 5450 1630
rect 5470 1610 5530 1630
rect 5550 1610 5610 1630
rect 5630 1610 5690 1630
rect 5710 1610 5720 1630
rect 4720 1600 5720 1610
rect 5760 1630 5960 1640
rect 5760 1610 5770 1630
rect 5790 1610 5850 1630
rect 5870 1610 5930 1630
rect 5950 1610 5960 1630
rect 5760 1600 5960 1610
rect 6000 1630 6200 1640
rect 6000 1610 6010 1630
rect 6030 1610 6090 1630
rect 6110 1610 6170 1630
rect 6190 1610 6200 1630
rect 6000 1600 6200 1610
rect 4240 1550 4440 1560
rect 4240 1530 4250 1550
rect 4270 1530 4330 1550
rect 4350 1530 4410 1550
rect 4430 1530 4440 1550
rect 4240 1520 4440 1530
rect 4480 1550 4680 1560
rect 4480 1530 4490 1550
rect 4510 1530 4570 1550
rect 4590 1530 4650 1550
rect 4670 1530 4680 1550
rect 4480 1520 4680 1530
rect 4720 1550 5720 1560
rect 4720 1530 4730 1550
rect 4750 1530 4810 1550
rect 4830 1530 4890 1550
rect 4910 1530 4970 1550
rect 4990 1530 5050 1550
rect 5070 1530 5130 1550
rect 5150 1530 5210 1550
rect 5230 1530 5290 1550
rect 5310 1530 5370 1550
rect 5390 1530 5450 1550
rect 5470 1530 5530 1550
rect 5550 1530 5610 1550
rect 5630 1530 5690 1550
rect 5710 1530 5720 1550
rect 4720 1520 5720 1530
rect 5760 1550 5960 1560
rect 5760 1530 5770 1550
rect 5790 1530 5850 1550
rect 5870 1530 5930 1550
rect 5950 1530 5960 1550
rect 5760 1520 5960 1530
rect 6000 1550 6200 1560
rect 6000 1530 6010 1550
rect 6030 1530 6090 1550
rect 6110 1530 6170 1550
rect 6190 1530 6200 1550
rect 6000 1520 6200 1530
rect 4240 1470 4440 1480
rect 4240 1450 4250 1470
rect 4270 1450 4330 1470
rect 4350 1450 4410 1470
rect 4430 1450 4440 1470
rect 4240 1440 4440 1450
rect 4480 1470 4680 1480
rect 4480 1450 4490 1470
rect 4510 1450 4570 1470
rect 4590 1450 4650 1470
rect 4670 1450 4680 1470
rect 4480 1440 4680 1450
rect 4720 1470 5720 1480
rect 4720 1450 4730 1470
rect 4750 1450 4810 1470
rect 4830 1450 4890 1470
rect 4910 1450 4970 1470
rect 4990 1450 5050 1470
rect 5070 1450 5130 1470
rect 5150 1450 5210 1470
rect 5230 1450 5290 1470
rect 5310 1450 5370 1470
rect 5390 1450 5450 1470
rect 5470 1450 5530 1470
rect 5550 1450 5610 1470
rect 5630 1450 5690 1470
rect 5710 1450 5720 1470
rect 4720 1440 5720 1450
rect 5760 1470 5960 1480
rect 5760 1450 5770 1470
rect 5790 1450 5850 1470
rect 5870 1450 5930 1470
rect 5950 1450 5960 1470
rect 5760 1440 5960 1450
rect 6000 1470 6200 1480
rect 6000 1450 6010 1470
rect 6030 1450 6090 1470
rect 6110 1450 6170 1470
rect 6190 1450 6200 1470
rect 6000 1440 6200 1450
rect 4240 1390 4440 1400
rect 4240 1370 4250 1390
rect 4270 1370 4330 1390
rect 4350 1370 4410 1390
rect 4430 1370 4440 1390
rect 4240 1360 4440 1370
rect 4480 1390 4680 1400
rect 4480 1370 4490 1390
rect 4510 1370 4570 1390
rect 4590 1370 4650 1390
rect 4670 1370 4680 1390
rect 4480 1360 4680 1370
rect 4720 1390 5720 1400
rect 4720 1370 4730 1390
rect 4750 1370 4810 1390
rect 4830 1370 4890 1390
rect 4910 1370 4970 1390
rect 4990 1370 5050 1390
rect 5070 1370 5130 1390
rect 5150 1370 5210 1390
rect 5230 1370 5290 1390
rect 5310 1370 5370 1390
rect 5390 1370 5450 1390
rect 5470 1370 5530 1390
rect 5550 1370 5610 1390
rect 5630 1370 5690 1390
rect 5710 1370 5720 1390
rect 4720 1360 5720 1370
rect 5760 1390 5960 1400
rect 5760 1370 5770 1390
rect 5790 1370 5850 1390
rect 5870 1370 5930 1390
rect 5950 1370 5960 1390
rect 5760 1360 5960 1370
rect 6000 1390 6200 1400
rect 6000 1370 6010 1390
rect 6030 1370 6090 1390
rect 6110 1370 6170 1390
rect 6190 1370 6200 1390
rect 6000 1360 6200 1370
rect 4240 1310 4440 1320
rect 4240 1290 4250 1310
rect 4270 1290 4330 1310
rect 4350 1290 4410 1310
rect 4430 1290 4440 1310
rect 4240 1280 4440 1290
rect 4480 1310 4680 1320
rect 4480 1290 4490 1310
rect 4510 1290 4570 1310
rect 4590 1290 4650 1310
rect 4670 1290 4680 1310
rect 4480 1280 4680 1290
rect 4720 1310 5720 1320
rect 4720 1290 4730 1310
rect 4750 1290 4810 1310
rect 4830 1290 4890 1310
rect 4910 1290 4970 1310
rect 4990 1290 5050 1310
rect 5070 1290 5130 1310
rect 5150 1290 5210 1310
rect 5230 1290 5290 1310
rect 5310 1290 5370 1310
rect 5390 1290 5450 1310
rect 5470 1290 5530 1310
rect 5550 1290 5610 1310
rect 5630 1290 5690 1310
rect 5710 1290 5720 1310
rect 4720 1280 5720 1290
rect 5760 1310 5960 1320
rect 5760 1290 5770 1310
rect 5790 1290 5850 1310
rect 5870 1290 5930 1310
rect 5950 1290 5960 1310
rect 5760 1280 5960 1290
rect 6000 1310 6200 1320
rect 6000 1290 6010 1310
rect 6030 1290 6090 1310
rect 6110 1290 6170 1310
rect 6190 1290 6200 1310
rect 6000 1280 6200 1290
rect 4240 1230 4440 1240
rect 4240 1210 4250 1230
rect 4270 1210 4330 1230
rect 4350 1210 4410 1230
rect 4430 1210 4440 1230
rect 4240 1200 4440 1210
rect 4480 1230 4680 1240
rect 4480 1210 4490 1230
rect 4510 1210 4570 1230
rect 4590 1210 4650 1230
rect 4670 1210 4680 1230
rect 4480 1200 4680 1210
rect 4720 1230 5720 1240
rect 4720 1210 4730 1230
rect 4750 1210 4810 1230
rect 4830 1210 4890 1230
rect 4910 1210 4970 1230
rect 4990 1210 5050 1230
rect 5070 1210 5130 1230
rect 5150 1210 5210 1230
rect 5230 1210 5290 1230
rect 5310 1210 5370 1230
rect 5390 1210 5450 1230
rect 5470 1210 5530 1230
rect 5550 1210 5610 1230
rect 5630 1210 5690 1230
rect 5710 1210 5720 1230
rect 4720 1200 5720 1210
rect 5760 1230 5960 1240
rect 5760 1210 5770 1230
rect 5790 1210 5850 1230
rect 5870 1210 5930 1230
rect 5950 1210 5960 1230
rect 5760 1200 5960 1210
rect 6000 1230 6200 1240
rect 6000 1210 6010 1230
rect 6030 1210 6090 1230
rect 6110 1210 6170 1230
rect 6190 1210 6200 1230
rect 6000 1200 6200 1210
rect 4240 1150 4440 1160
rect 4240 1130 4250 1150
rect 4270 1130 4330 1150
rect 4350 1130 4410 1150
rect 4430 1130 4440 1150
rect 4240 1120 4440 1130
rect 4480 1150 4680 1160
rect 4480 1130 4490 1150
rect 4510 1130 4570 1150
rect 4590 1130 4650 1150
rect 4670 1130 4680 1150
rect 4480 1120 4680 1130
rect 4720 1150 5720 1160
rect 4720 1130 4730 1150
rect 4750 1130 4810 1150
rect 4830 1130 4890 1150
rect 4910 1130 4970 1150
rect 4990 1130 5050 1150
rect 5070 1130 5130 1150
rect 5150 1130 5210 1150
rect 5230 1130 5290 1150
rect 5310 1130 5370 1150
rect 5390 1130 5450 1150
rect 5470 1130 5530 1150
rect 5550 1130 5610 1150
rect 5630 1130 5690 1150
rect 5710 1130 5720 1150
rect 4720 1120 5720 1130
rect 5760 1150 5960 1160
rect 5760 1130 5770 1150
rect 5790 1130 5850 1150
rect 5870 1130 5930 1150
rect 5950 1130 5960 1150
rect 5760 1120 5960 1130
rect 6000 1150 6200 1160
rect 6000 1130 6010 1150
rect 6030 1130 6090 1150
rect 6110 1130 6170 1150
rect 6190 1130 6200 1150
rect 6000 1120 6200 1130
rect 4240 1070 4440 1080
rect 4240 1050 4250 1070
rect 4270 1050 4330 1070
rect 4350 1050 4410 1070
rect 4430 1050 4440 1070
rect 4240 1040 4440 1050
rect 4480 1070 4680 1080
rect 4480 1050 4490 1070
rect 4510 1050 4570 1070
rect 4590 1050 4650 1070
rect 4670 1050 4680 1070
rect 4480 1040 4680 1050
rect 4720 1070 5720 1080
rect 4720 1050 4730 1070
rect 4750 1050 4810 1070
rect 4830 1050 4890 1070
rect 4910 1050 4970 1070
rect 4990 1050 5050 1070
rect 5070 1050 5130 1070
rect 5150 1050 5210 1070
rect 5230 1050 5290 1070
rect 5310 1050 5370 1070
rect 5390 1050 5450 1070
rect 5470 1050 5530 1070
rect 5550 1050 5610 1070
rect 5630 1050 5690 1070
rect 5710 1050 5720 1070
rect 4720 1040 5720 1050
rect 5760 1070 5960 1080
rect 5760 1050 5770 1070
rect 5790 1050 5850 1070
rect 5870 1050 5930 1070
rect 5950 1050 5960 1070
rect 5760 1040 5960 1050
rect 6000 1070 6200 1080
rect 6000 1050 6010 1070
rect 6030 1050 6090 1070
rect 6110 1050 6170 1070
rect 6190 1050 6200 1070
rect 6000 1040 6200 1050
rect 4240 990 4440 1000
rect 4240 970 4250 990
rect 4270 970 4330 990
rect 4350 970 4410 990
rect 4430 970 4440 990
rect 4240 960 4440 970
rect 4480 990 4680 1000
rect 4480 970 4490 990
rect 4510 970 4570 990
rect 4590 970 4650 990
rect 4670 970 4680 990
rect 4480 960 4680 970
rect 4720 990 5720 1000
rect 4720 970 4730 990
rect 4750 970 4810 990
rect 4830 970 4890 990
rect 4910 970 4970 990
rect 4990 970 5050 990
rect 5070 970 5130 990
rect 5150 970 5210 990
rect 5230 970 5290 990
rect 5310 970 5370 990
rect 5390 970 5450 990
rect 5470 970 5530 990
rect 5550 970 5610 990
rect 5630 970 5690 990
rect 5710 970 5720 990
rect 4720 960 5720 970
rect 5760 990 5960 1000
rect 5760 970 5770 990
rect 5790 970 5850 990
rect 5870 970 5930 990
rect 5950 970 5960 990
rect 5760 960 5960 970
rect 6000 990 6200 1000
rect 6000 970 6010 990
rect 6030 970 6090 990
rect 6110 970 6170 990
rect 6190 970 6200 990
rect 6000 960 6200 970
rect 4240 910 4440 920
rect 4240 890 4250 910
rect 4270 890 4330 910
rect 4350 890 4410 910
rect 4430 890 4440 910
rect 4240 880 4440 890
rect 4480 910 4680 920
rect 4480 890 4490 910
rect 4510 890 4570 910
rect 4590 890 4650 910
rect 4670 890 4680 910
rect 4480 880 4680 890
rect 4720 910 5720 920
rect 4720 890 4730 910
rect 4750 890 4810 910
rect 4830 890 4890 910
rect 4910 890 4970 910
rect 4990 890 5050 910
rect 5070 890 5130 910
rect 5150 890 5210 910
rect 5230 890 5290 910
rect 5310 890 5370 910
rect 5390 890 5450 910
rect 5470 890 5530 910
rect 5550 890 5610 910
rect 5630 890 5690 910
rect 5710 890 5720 910
rect 4720 880 5720 890
rect 5760 910 5960 920
rect 5760 890 5770 910
rect 5790 890 5850 910
rect 5870 890 5930 910
rect 5950 890 5960 910
rect 5760 880 5960 890
rect 6000 910 6200 920
rect 6000 890 6010 910
rect 6030 890 6090 910
rect 6110 890 6170 910
rect 6190 890 6200 910
rect 6000 880 6200 890
rect 4240 830 4440 840
rect 4240 810 4250 830
rect 4270 810 4330 830
rect 4350 810 4410 830
rect 4430 810 4440 830
rect 4240 800 4440 810
rect 4480 830 4680 840
rect 4480 810 4490 830
rect 4510 810 4570 830
rect 4590 810 4650 830
rect 4670 810 4680 830
rect 4480 800 4680 810
rect 4720 830 5720 840
rect 4720 810 4730 830
rect 4750 810 4810 830
rect 4830 810 4890 830
rect 4910 810 4970 830
rect 4990 810 5050 830
rect 5070 810 5130 830
rect 5150 810 5210 830
rect 5230 810 5290 830
rect 5310 810 5370 830
rect 5390 810 5450 830
rect 5470 810 5530 830
rect 5550 810 5610 830
rect 5630 810 5690 830
rect 5710 810 5720 830
rect 4720 800 5720 810
rect 5760 830 5960 840
rect 5760 810 5770 830
rect 5790 810 5850 830
rect 5870 810 5930 830
rect 5950 810 5960 830
rect 5760 800 5960 810
rect 6000 830 6200 840
rect 6000 810 6010 830
rect 6030 810 6090 830
rect 6110 810 6170 830
rect 6190 810 6200 830
rect 6000 800 6200 810
rect 4240 750 4440 760
rect 4240 730 4250 750
rect 4270 730 4330 750
rect 4350 730 4410 750
rect 4430 730 4440 750
rect 4240 720 4440 730
rect 4480 750 4680 760
rect 4480 730 4490 750
rect 4510 730 4570 750
rect 4590 730 4650 750
rect 4670 730 4680 750
rect 4480 720 4680 730
rect 4720 750 5720 760
rect 4720 730 4730 750
rect 4750 730 4810 750
rect 4830 730 4890 750
rect 4910 730 4970 750
rect 4990 730 5050 750
rect 5070 730 5130 750
rect 5150 730 5210 750
rect 5230 730 5290 750
rect 5310 730 5370 750
rect 5390 730 5450 750
rect 5470 730 5530 750
rect 5550 730 5610 750
rect 5630 730 5690 750
rect 5710 730 5720 750
rect 4720 720 5720 730
rect 5760 750 5960 760
rect 5760 730 5770 750
rect 5790 730 5850 750
rect 5870 730 5930 750
rect 5950 730 5960 750
rect 5760 720 5960 730
rect 6000 750 6200 760
rect 6000 730 6010 750
rect 6030 730 6090 750
rect 6110 730 6170 750
rect 6190 730 6200 750
rect 6000 720 6200 730
rect 4240 670 4440 680
rect 4240 650 4250 670
rect 4270 650 4330 670
rect 4350 650 4410 670
rect 4430 650 4440 670
rect 4240 640 4440 650
rect 4480 670 4680 680
rect 4480 650 4490 670
rect 4510 650 4570 670
rect 4590 650 4650 670
rect 4670 650 4680 670
rect 4480 640 4680 650
rect 4720 670 5720 680
rect 4720 650 4730 670
rect 4750 650 4810 670
rect 4830 650 4890 670
rect 4910 650 4970 670
rect 4990 650 5050 670
rect 5070 650 5130 670
rect 5150 650 5210 670
rect 5230 650 5290 670
rect 5310 650 5370 670
rect 5390 650 5450 670
rect 5470 650 5530 670
rect 5550 650 5610 670
rect 5630 650 5690 670
rect 5710 650 5720 670
rect 4720 640 5720 650
rect 5760 670 5960 680
rect 5760 650 5770 670
rect 5790 650 5850 670
rect 5870 650 5930 670
rect 5950 650 5960 670
rect 5760 640 5960 650
rect 6000 670 6200 680
rect 6000 650 6010 670
rect 6030 650 6090 670
rect 6110 650 6170 670
rect 6190 650 6200 670
rect 6000 640 6200 650
rect 4240 590 4440 600
rect 4240 570 4250 590
rect 4270 570 4330 590
rect 4350 570 4410 590
rect 4430 570 4440 590
rect 4240 560 4440 570
rect 4480 590 4680 600
rect 4480 570 4490 590
rect 4510 570 4570 590
rect 4590 570 4650 590
rect 4670 570 4680 590
rect 4480 560 4680 570
rect 4720 590 5720 600
rect 4720 570 4730 590
rect 4750 570 4810 590
rect 4830 570 4890 590
rect 4910 570 4970 590
rect 4990 570 5050 590
rect 5070 570 5130 590
rect 5150 570 5210 590
rect 5230 570 5290 590
rect 5310 570 5370 590
rect 5390 570 5450 590
rect 5470 570 5530 590
rect 5550 570 5610 590
rect 5630 570 5690 590
rect 5710 570 5720 590
rect 4720 560 5720 570
rect 5760 590 5960 600
rect 5760 570 5770 590
rect 5790 570 5850 590
rect 5870 570 5930 590
rect 5950 570 5960 590
rect 5760 560 5960 570
rect 6000 590 6200 600
rect 6000 570 6010 590
rect 6030 570 6090 590
rect 6110 570 6170 590
rect 6190 570 6200 590
rect 6000 560 6200 570
rect 4240 510 4440 520
rect 4240 490 4250 510
rect 4270 490 4330 510
rect 4350 490 4410 510
rect 4430 490 4440 510
rect 4240 480 4440 490
rect 4480 510 4680 520
rect 4480 490 4490 510
rect 4510 490 4570 510
rect 4590 490 4650 510
rect 4670 490 4680 510
rect 4480 480 4680 490
rect 4720 510 5720 520
rect 4720 490 4730 510
rect 4750 490 4810 510
rect 4830 490 4890 510
rect 4910 490 4970 510
rect 4990 490 5050 510
rect 5070 490 5130 510
rect 5150 490 5210 510
rect 5230 490 5290 510
rect 5310 490 5370 510
rect 5390 490 5450 510
rect 5470 490 5530 510
rect 5550 490 5610 510
rect 5630 490 5690 510
rect 5710 490 5720 510
rect 4720 480 5720 490
rect 5760 510 5960 520
rect 5760 490 5770 510
rect 5790 490 5850 510
rect 5870 490 5930 510
rect 5950 490 5960 510
rect 5760 480 5960 490
rect 6000 510 6200 520
rect 6000 490 6010 510
rect 6030 490 6090 510
rect 6110 490 6170 510
rect 6190 490 6200 510
rect 6000 480 6200 490
rect 4240 430 4440 440
rect 4240 410 4250 430
rect 4270 410 4330 430
rect 4350 410 4410 430
rect 4430 410 4440 430
rect 4240 400 4440 410
rect 4480 430 4680 440
rect 4480 410 4490 430
rect 4510 410 4570 430
rect 4590 410 4650 430
rect 4670 410 4680 430
rect 4480 400 4680 410
rect 4720 430 5720 440
rect 4720 410 4730 430
rect 4750 410 4810 430
rect 4830 410 4890 430
rect 4910 410 4970 430
rect 4990 410 5050 430
rect 5070 410 5130 430
rect 5150 410 5210 430
rect 5230 410 5290 430
rect 5310 410 5370 430
rect 5390 410 5450 430
rect 5470 410 5530 430
rect 5550 410 5610 430
rect 5630 410 5690 430
rect 5710 410 5720 430
rect 4720 400 5720 410
rect 5760 430 5960 440
rect 5760 410 5770 430
rect 5790 410 5850 430
rect 5870 410 5930 430
rect 5950 410 5960 430
rect 5760 400 5960 410
rect 6000 430 6200 440
rect 6000 410 6010 430
rect 6030 410 6090 430
rect 6110 410 6170 430
rect 6190 410 6200 430
rect 6000 400 6200 410
rect 4240 350 4440 360
rect 4240 330 4250 350
rect 4270 330 4330 350
rect 4350 330 4410 350
rect 4430 330 4440 350
rect 4240 320 4440 330
rect 4480 350 4680 360
rect 4480 330 4490 350
rect 4510 330 4570 350
rect 4590 330 4650 350
rect 4670 330 4680 350
rect 4480 320 4680 330
rect 4720 350 5720 360
rect 4720 330 4730 350
rect 4750 330 4810 350
rect 4830 330 4890 350
rect 4910 330 4970 350
rect 4990 330 5050 350
rect 5070 330 5130 350
rect 5150 330 5210 350
rect 5230 330 5290 350
rect 5310 330 5370 350
rect 5390 330 5450 350
rect 5470 330 5530 350
rect 5550 330 5610 350
rect 5630 330 5690 350
rect 5710 330 5720 350
rect 4720 320 5720 330
rect 5760 350 5960 360
rect 5760 330 5770 350
rect 5790 330 5850 350
rect 5870 330 5930 350
rect 5950 330 5960 350
rect 5760 320 5960 330
rect 6000 350 6200 360
rect 6000 330 6010 350
rect 6030 330 6090 350
rect 6110 330 6170 350
rect 6190 330 6200 350
rect 6000 320 6200 330
rect 4240 270 4440 280
rect 4240 250 4250 270
rect 4270 250 4330 270
rect 4350 250 4410 270
rect 4430 250 4440 270
rect 4240 240 4440 250
rect 4480 270 4680 280
rect 4480 250 4490 270
rect 4510 250 4570 270
rect 4590 250 4650 270
rect 4670 250 4680 270
rect 4480 240 4680 250
rect 4720 270 5720 280
rect 4720 250 4730 270
rect 4750 250 4810 270
rect 4830 250 4890 270
rect 4910 250 4970 270
rect 4990 250 5050 270
rect 5070 250 5130 270
rect 5150 250 5210 270
rect 5230 250 5290 270
rect 5310 250 5370 270
rect 5390 250 5450 270
rect 5470 250 5530 270
rect 5550 250 5610 270
rect 5630 250 5690 270
rect 5710 250 5720 270
rect 4720 240 5720 250
rect 5760 270 5960 280
rect 5760 250 5770 270
rect 5790 250 5850 270
rect 5870 250 5930 270
rect 5950 250 5960 270
rect 5760 240 5960 250
rect 6000 270 6200 280
rect 6000 250 6010 270
rect 6030 250 6090 270
rect 6110 250 6170 270
rect 6190 250 6200 270
rect 6000 240 6200 250
rect 4240 190 4440 200
rect 4240 170 4250 190
rect 4270 170 4330 190
rect 4350 170 4410 190
rect 4430 170 4440 190
rect 4240 160 4440 170
rect 4480 190 4680 200
rect 4480 170 4490 190
rect 4510 170 4570 190
rect 4590 170 4650 190
rect 4670 170 4680 190
rect 4480 160 4680 170
rect 4720 190 5720 200
rect 4720 170 4730 190
rect 4750 170 4810 190
rect 4830 170 4890 190
rect 4910 170 4970 190
rect 4990 170 5050 190
rect 5070 170 5130 190
rect 5150 170 5210 190
rect 5230 170 5290 190
rect 5310 170 5370 190
rect 5390 170 5450 190
rect 5470 170 5530 190
rect 5550 170 5610 190
rect 5630 170 5690 190
rect 5710 170 5720 190
rect 4720 160 5720 170
rect 5760 190 5960 200
rect 5760 170 5770 190
rect 5790 170 5850 190
rect 5870 170 5930 190
rect 5950 170 5960 190
rect 5760 160 5960 170
rect 6000 190 6200 200
rect 6000 170 6010 190
rect 6030 170 6090 190
rect 6110 170 6170 190
rect 6190 170 6200 190
rect 6000 160 6200 170
rect 4240 110 4440 120
rect 4240 90 4250 110
rect 4270 90 4330 110
rect 4350 90 4410 110
rect 4430 90 4440 110
rect 4240 80 4440 90
rect 4480 110 4680 120
rect 4480 90 4490 110
rect 4510 90 4570 110
rect 4590 90 4650 110
rect 4670 90 4680 110
rect 4480 80 4680 90
rect 4720 110 5720 120
rect 4720 90 4730 110
rect 4750 90 4810 110
rect 4830 90 4890 110
rect 4910 90 4970 110
rect 4990 90 5050 110
rect 5070 90 5130 110
rect 5150 90 5210 110
rect 5230 90 5290 110
rect 5310 90 5370 110
rect 5390 90 5450 110
rect 5470 90 5530 110
rect 5550 90 5610 110
rect 5630 90 5690 110
rect 5710 90 5720 110
rect 4720 80 5720 90
rect 5760 110 5960 120
rect 5760 90 5770 110
rect 5790 90 5850 110
rect 5870 90 5930 110
rect 5950 90 5960 110
rect 5760 80 5960 90
rect 6000 110 6200 120
rect 6000 90 6010 110
rect 6030 90 6090 110
rect 6110 90 6170 110
rect 6190 90 6200 110
rect 6000 80 6200 90
rect 4240 30 4440 40
rect 4240 10 4250 30
rect 4270 10 4330 30
rect 4350 10 4410 30
rect 4430 10 4440 30
rect 4240 0 4440 10
rect 4480 30 4680 40
rect 4480 10 4490 30
rect 4510 10 4570 30
rect 4590 10 4650 30
rect 4670 10 4680 30
rect 4480 0 4680 10
rect 4720 30 5720 40
rect 4720 10 4730 30
rect 4750 10 4810 30
rect 4830 10 4890 30
rect 4910 10 4970 30
rect 4990 10 5050 30
rect 5070 10 5130 30
rect 5150 10 5210 30
rect 5230 10 5290 30
rect 5310 10 5370 30
rect 5390 10 5450 30
rect 5470 10 5530 30
rect 5550 10 5610 30
rect 5630 10 5690 30
rect 5710 10 5720 30
rect 4720 0 5720 10
rect 5760 30 5960 40
rect 5760 10 5770 30
rect 5790 10 5850 30
rect 5870 10 5930 30
rect 5950 10 5960 30
rect 5760 0 5960 10
rect 6000 30 6200 40
rect 6000 10 6010 30
rect 6030 10 6090 30
rect 6110 10 6170 30
rect 6190 10 6200 30
rect 6000 0 6200 10
<< viali >>
rect 4250 15690 4270 15710
rect 4330 15690 4350 15710
rect 4410 15690 4430 15710
rect 4490 15690 4510 15710
rect 4570 15690 4590 15710
rect 4650 15690 4670 15710
rect 4730 15690 4750 15710
rect 4810 15690 4830 15710
rect 4890 15690 4910 15710
rect 4970 15690 4990 15710
rect 5050 15690 5070 15710
rect 5130 15690 5150 15710
rect 5210 15690 5230 15710
rect 5290 15690 5310 15710
rect 5370 15690 5390 15710
rect 5450 15690 5470 15710
rect 5530 15690 5550 15710
rect 5610 15690 5630 15710
rect 5690 15690 5710 15710
rect 5770 15690 5790 15710
rect 5850 15690 5870 15710
rect 5930 15690 5950 15710
rect 6010 15690 6030 15710
rect 6090 15690 6110 15710
rect 6170 15690 6190 15710
rect 4250 15610 4270 15630
rect 4330 15610 4350 15630
rect 4410 15610 4430 15630
rect 4490 15610 4510 15630
rect 4570 15610 4590 15630
rect 4650 15610 4670 15630
rect 4730 15610 4750 15630
rect 4810 15610 4830 15630
rect 4890 15610 4910 15630
rect 4970 15610 4990 15630
rect 5050 15610 5070 15630
rect 5130 15610 5150 15630
rect 5210 15610 5230 15630
rect 5290 15610 5310 15630
rect 5370 15610 5390 15630
rect 5450 15610 5470 15630
rect 5530 15610 5550 15630
rect 5610 15610 5630 15630
rect 5690 15610 5710 15630
rect 5770 15610 5790 15630
rect 5850 15610 5870 15630
rect 5930 15610 5950 15630
rect 6010 15610 6030 15630
rect 6090 15610 6110 15630
rect 6170 15610 6190 15630
rect 4250 15530 4270 15550
rect 4330 15530 4350 15550
rect 4410 15530 4430 15550
rect 4490 15530 4510 15550
rect 4570 15530 4590 15550
rect 4650 15530 4670 15550
rect 4730 15530 4750 15550
rect 4810 15530 4830 15550
rect 4890 15530 4910 15550
rect 4970 15530 4990 15550
rect 5050 15530 5070 15550
rect 5130 15530 5150 15550
rect 5210 15530 5230 15550
rect 5290 15530 5310 15550
rect 5370 15530 5390 15550
rect 5450 15530 5470 15550
rect 5530 15530 5550 15550
rect 5610 15530 5630 15550
rect 5690 15530 5710 15550
rect 5770 15530 5790 15550
rect 5850 15530 5870 15550
rect 5930 15530 5950 15550
rect 6010 15530 6030 15550
rect 6090 15530 6110 15550
rect 6170 15530 6190 15550
rect 4250 15450 4270 15470
rect 4330 15450 4350 15470
rect 4410 15450 4430 15470
rect 4490 15450 4510 15470
rect 4570 15450 4590 15470
rect 4650 15450 4670 15470
rect 4730 15450 4750 15470
rect 4810 15450 4830 15470
rect 4890 15450 4910 15470
rect 4970 15450 4990 15470
rect 5050 15450 5070 15470
rect 5130 15450 5150 15470
rect 5210 15450 5230 15470
rect 5290 15450 5310 15470
rect 5370 15450 5390 15470
rect 5450 15450 5470 15470
rect 5530 15450 5550 15470
rect 5610 15450 5630 15470
rect 5690 15450 5710 15470
rect 5770 15450 5790 15470
rect 5850 15450 5870 15470
rect 5930 15450 5950 15470
rect 6010 15450 6030 15470
rect 6090 15450 6110 15470
rect 6170 15450 6190 15470
rect 4250 15370 4270 15390
rect 4330 15370 4350 15390
rect 4410 15370 4430 15390
rect 4490 15370 4510 15390
rect 4570 15370 4590 15390
rect 4650 15370 4670 15390
rect 4730 15370 4750 15390
rect 4810 15370 4830 15390
rect 4890 15370 4910 15390
rect 4970 15370 4990 15390
rect 5050 15370 5070 15390
rect 5130 15370 5150 15390
rect 5210 15370 5230 15390
rect 5290 15370 5310 15390
rect 5370 15370 5390 15390
rect 5450 15370 5470 15390
rect 5530 15370 5550 15390
rect 5610 15370 5630 15390
rect 5690 15370 5710 15390
rect 5770 15370 5790 15390
rect 5850 15370 5870 15390
rect 5930 15370 5950 15390
rect 6010 15370 6030 15390
rect 6090 15370 6110 15390
rect 6170 15370 6190 15390
rect 4250 15290 4270 15310
rect 4330 15290 4350 15310
rect 4410 15290 4430 15310
rect 4490 15290 4510 15310
rect 4570 15290 4590 15310
rect 4650 15290 4670 15310
rect 4730 15290 4750 15310
rect 4810 15290 4830 15310
rect 4890 15290 4910 15310
rect 4970 15290 4990 15310
rect 5050 15290 5070 15310
rect 5130 15290 5150 15310
rect 5210 15290 5230 15310
rect 5290 15290 5310 15310
rect 5370 15290 5390 15310
rect 5450 15290 5470 15310
rect 5530 15290 5550 15310
rect 5610 15290 5630 15310
rect 5690 15290 5710 15310
rect 5770 15290 5790 15310
rect 5850 15290 5870 15310
rect 5930 15290 5950 15310
rect 6010 15290 6030 15310
rect 6090 15290 6110 15310
rect 6170 15290 6190 15310
rect 4250 15210 4270 15230
rect 4330 15210 4350 15230
rect 4410 15210 4430 15230
rect 4490 15210 4510 15230
rect 4570 15210 4590 15230
rect 4650 15210 4670 15230
rect 4730 15210 4750 15230
rect 4810 15210 4830 15230
rect 4890 15210 4910 15230
rect 4970 15210 4990 15230
rect 5050 15210 5070 15230
rect 5130 15210 5150 15230
rect 5210 15210 5230 15230
rect 5290 15210 5310 15230
rect 5370 15210 5390 15230
rect 5450 15210 5470 15230
rect 5530 15210 5550 15230
rect 5610 15210 5630 15230
rect 5690 15210 5710 15230
rect 5770 15210 5790 15230
rect 5850 15210 5870 15230
rect 5930 15210 5950 15230
rect 6010 15210 6030 15230
rect 6090 15210 6110 15230
rect 6170 15210 6190 15230
rect 4250 15130 4270 15150
rect 4330 15130 4350 15150
rect 4410 15130 4430 15150
rect 4490 15130 4510 15150
rect 4570 15130 4590 15150
rect 4650 15130 4670 15150
rect 4730 15130 4750 15150
rect 4810 15130 4830 15150
rect 4890 15130 4910 15150
rect 4970 15130 4990 15150
rect 5050 15130 5070 15150
rect 5130 15130 5150 15150
rect 5210 15130 5230 15150
rect 5290 15130 5310 15150
rect 5370 15130 5390 15150
rect 5450 15130 5470 15150
rect 5530 15130 5550 15150
rect 5610 15130 5630 15150
rect 5690 15130 5710 15150
rect 5770 15130 5790 15150
rect 5850 15130 5870 15150
rect 5930 15130 5950 15150
rect 6010 15130 6030 15150
rect 6090 15130 6110 15150
rect 6170 15130 6190 15150
rect 4250 15050 4270 15070
rect 4330 15050 4350 15070
rect 4410 15050 4430 15070
rect 4490 15050 4510 15070
rect 4570 15050 4590 15070
rect 4650 15050 4670 15070
rect 4730 15050 4750 15070
rect 4810 15050 4830 15070
rect 4890 15050 4910 15070
rect 4970 15050 4990 15070
rect 5050 15050 5070 15070
rect 5130 15050 5150 15070
rect 5210 15050 5230 15070
rect 5290 15050 5310 15070
rect 5370 15050 5390 15070
rect 5450 15050 5470 15070
rect 5530 15050 5550 15070
rect 5610 15050 5630 15070
rect 5690 15050 5710 15070
rect 5770 15050 5790 15070
rect 5850 15050 5870 15070
rect 5930 15050 5950 15070
rect 6010 15050 6030 15070
rect 6090 15050 6110 15070
rect 6170 15050 6190 15070
rect 4250 14970 4270 14990
rect 4330 14970 4350 14990
rect 4410 14970 4430 14990
rect 4490 14970 4510 14990
rect 4570 14970 4590 14990
rect 4650 14970 4670 14990
rect 4730 14970 4750 14990
rect 4810 14970 4830 14990
rect 4890 14970 4910 14990
rect 4970 14970 4990 14990
rect 5050 14970 5070 14990
rect 5130 14970 5150 14990
rect 5210 14970 5230 14990
rect 5290 14970 5310 14990
rect 5370 14970 5390 14990
rect 5450 14970 5470 14990
rect 5530 14970 5550 14990
rect 5610 14970 5630 14990
rect 5690 14970 5710 14990
rect 5770 14970 5790 14990
rect 5850 14970 5870 14990
rect 5930 14970 5950 14990
rect 6010 14970 6030 14990
rect 6090 14970 6110 14990
rect 6170 14970 6190 14990
rect 4250 14890 4270 14910
rect 4330 14890 4350 14910
rect 4410 14890 4430 14910
rect 4490 14890 4510 14910
rect 4570 14890 4590 14910
rect 4650 14890 4670 14910
rect 4730 14890 4750 14910
rect 4810 14890 4830 14910
rect 4890 14890 4910 14910
rect 4970 14890 4990 14910
rect 5050 14890 5070 14910
rect 5130 14890 5150 14910
rect 5210 14890 5230 14910
rect 5290 14890 5310 14910
rect 5370 14890 5390 14910
rect 5450 14890 5470 14910
rect 5530 14890 5550 14910
rect 5610 14890 5630 14910
rect 5690 14890 5710 14910
rect 5770 14890 5790 14910
rect 5850 14890 5870 14910
rect 5930 14890 5950 14910
rect 6010 14890 6030 14910
rect 6090 14890 6110 14910
rect 6170 14890 6190 14910
rect 4250 14810 4270 14830
rect 4330 14810 4350 14830
rect 4410 14810 4430 14830
rect 4490 14810 4510 14830
rect 4570 14810 4590 14830
rect 4650 14810 4670 14830
rect 4730 14810 4750 14830
rect 4810 14810 4830 14830
rect 4890 14810 4910 14830
rect 4970 14810 4990 14830
rect 5050 14810 5070 14830
rect 5130 14810 5150 14830
rect 5210 14810 5230 14830
rect 5290 14810 5310 14830
rect 5370 14810 5390 14830
rect 5450 14810 5470 14830
rect 5530 14810 5550 14830
rect 5610 14810 5630 14830
rect 5690 14810 5710 14830
rect 5770 14810 5790 14830
rect 5850 14810 5870 14830
rect 5930 14810 5950 14830
rect 6010 14810 6030 14830
rect 6090 14810 6110 14830
rect 6170 14810 6190 14830
rect 4250 14730 4270 14750
rect 4330 14730 4350 14750
rect 4410 14730 4430 14750
rect 4490 14730 4510 14750
rect 4570 14730 4590 14750
rect 4650 14730 4670 14750
rect 4730 14730 4750 14750
rect 4810 14730 4830 14750
rect 4890 14730 4910 14750
rect 4970 14730 4990 14750
rect 5050 14730 5070 14750
rect 5130 14730 5150 14750
rect 5210 14730 5230 14750
rect 5290 14730 5310 14750
rect 5370 14730 5390 14750
rect 5450 14730 5470 14750
rect 5530 14730 5550 14750
rect 5610 14730 5630 14750
rect 5690 14730 5710 14750
rect 5770 14730 5790 14750
rect 5850 14730 5870 14750
rect 5930 14730 5950 14750
rect 6010 14730 6030 14750
rect 6090 14730 6110 14750
rect 6170 14730 6190 14750
rect 4250 14650 4270 14670
rect 4330 14650 4350 14670
rect 4410 14650 4430 14670
rect 4490 14650 4510 14670
rect 4570 14650 4590 14670
rect 4650 14650 4670 14670
rect 4730 14650 4750 14670
rect 4810 14650 4830 14670
rect 4890 14650 4910 14670
rect 4970 14650 4990 14670
rect 5050 14650 5070 14670
rect 5130 14650 5150 14670
rect 5210 14650 5230 14670
rect 5290 14650 5310 14670
rect 5370 14650 5390 14670
rect 5450 14650 5470 14670
rect 5530 14650 5550 14670
rect 5610 14650 5630 14670
rect 5690 14650 5710 14670
rect 5770 14650 5790 14670
rect 5850 14650 5870 14670
rect 5930 14650 5950 14670
rect 6010 14650 6030 14670
rect 6090 14650 6110 14670
rect 6170 14650 6190 14670
rect 4250 14570 4270 14590
rect 4330 14570 4350 14590
rect 4410 14570 4430 14590
rect 4490 14570 4510 14590
rect 4570 14570 4590 14590
rect 4650 14570 4670 14590
rect 4730 14570 4750 14590
rect 4810 14570 4830 14590
rect 4890 14570 4910 14590
rect 4970 14570 4990 14590
rect 5050 14570 5070 14590
rect 5130 14570 5150 14590
rect 5210 14570 5230 14590
rect 5290 14570 5310 14590
rect 5370 14570 5390 14590
rect 5450 14570 5470 14590
rect 5530 14570 5550 14590
rect 5610 14570 5630 14590
rect 5690 14570 5710 14590
rect 5770 14570 5790 14590
rect 5850 14570 5870 14590
rect 5930 14570 5950 14590
rect 6010 14570 6030 14590
rect 6090 14570 6110 14590
rect 6170 14570 6190 14590
rect 4250 14490 4270 14510
rect 4330 14490 4350 14510
rect 4410 14490 4430 14510
rect 4490 14490 4510 14510
rect 4570 14490 4590 14510
rect 4650 14490 4670 14510
rect 4730 14490 4750 14510
rect 4810 14490 4830 14510
rect 4890 14490 4910 14510
rect 4970 14490 4990 14510
rect 5050 14490 5070 14510
rect 5130 14490 5150 14510
rect 5210 14490 5230 14510
rect 5290 14490 5310 14510
rect 5370 14490 5390 14510
rect 5450 14490 5470 14510
rect 5530 14490 5550 14510
rect 5610 14490 5630 14510
rect 5690 14490 5710 14510
rect 5770 14490 5790 14510
rect 5850 14490 5870 14510
rect 5930 14490 5950 14510
rect 6010 14490 6030 14510
rect 6090 14490 6110 14510
rect 6170 14490 6190 14510
rect 4250 14410 4270 14430
rect 4330 14410 4350 14430
rect 4410 14410 4430 14430
rect 4490 14410 4510 14430
rect 4570 14410 4590 14430
rect 4650 14410 4670 14430
rect 4730 14410 4750 14430
rect 4810 14410 4830 14430
rect 4890 14410 4910 14430
rect 4970 14410 4990 14430
rect 5050 14410 5070 14430
rect 5130 14410 5150 14430
rect 5210 14410 5230 14430
rect 5290 14410 5310 14430
rect 5370 14410 5390 14430
rect 5450 14410 5470 14430
rect 5530 14410 5550 14430
rect 5610 14410 5630 14430
rect 5690 14410 5710 14430
rect 5770 14410 5790 14430
rect 5850 14410 5870 14430
rect 5930 14410 5950 14430
rect 6010 14410 6030 14430
rect 6090 14410 6110 14430
rect 6170 14410 6190 14430
rect 4250 14330 4270 14350
rect 4330 14330 4350 14350
rect 4410 14330 4430 14350
rect 4490 14330 4510 14350
rect 4570 14330 4590 14350
rect 4650 14330 4670 14350
rect 4730 14330 4750 14350
rect 4810 14330 4830 14350
rect 4890 14330 4910 14350
rect 4970 14330 4990 14350
rect 5050 14330 5070 14350
rect 5130 14330 5150 14350
rect 5210 14330 5230 14350
rect 5290 14330 5310 14350
rect 5370 14330 5390 14350
rect 5450 14330 5470 14350
rect 5530 14330 5550 14350
rect 5610 14330 5630 14350
rect 5690 14330 5710 14350
rect 5770 14330 5790 14350
rect 5850 14330 5870 14350
rect 5930 14330 5950 14350
rect 6010 14330 6030 14350
rect 6090 14330 6110 14350
rect 6170 14330 6190 14350
rect 4250 14250 4270 14270
rect 4330 14250 4350 14270
rect 4410 14250 4430 14270
rect 4490 14250 4510 14270
rect 4570 14250 4590 14270
rect 4650 14250 4670 14270
rect 4730 14250 4750 14270
rect 4810 14250 4830 14270
rect 4890 14250 4910 14270
rect 4970 14250 4990 14270
rect 5050 14250 5070 14270
rect 5130 14250 5150 14270
rect 5210 14250 5230 14270
rect 5290 14250 5310 14270
rect 5370 14250 5390 14270
rect 5450 14250 5470 14270
rect 5530 14250 5550 14270
rect 5610 14250 5630 14270
rect 5690 14250 5710 14270
rect 5770 14250 5790 14270
rect 5850 14250 5870 14270
rect 5930 14250 5950 14270
rect 6010 14250 6030 14270
rect 6090 14250 6110 14270
rect 6170 14250 6190 14270
rect 4250 14170 4270 14190
rect 4330 14170 4350 14190
rect 4410 14170 4430 14190
rect 4490 14170 4510 14190
rect 4570 14170 4590 14190
rect 4650 14170 4670 14190
rect 4730 14170 4750 14190
rect 4810 14170 4830 14190
rect 4890 14170 4910 14190
rect 4970 14170 4990 14190
rect 5050 14170 5070 14190
rect 5130 14170 5150 14190
rect 5210 14170 5230 14190
rect 5290 14170 5310 14190
rect 5370 14170 5390 14190
rect 5450 14170 5470 14190
rect 5530 14170 5550 14190
rect 5610 14170 5630 14190
rect 5690 14170 5710 14190
rect 5770 14170 5790 14190
rect 5850 14170 5870 14190
rect 5930 14170 5950 14190
rect 6010 14170 6030 14190
rect 6090 14170 6110 14190
rect 6170 14170 6190 14190
rect 4250 14090 4270 14110
rect 4330 14090 4350 14110
rect 4410 14090 4430 14110
rect 4490 14090 4510 14110
rect 4570 14090 4590 14110
rect 4650 14090 4670 14110
rect 4730 14090 4750 14110
rect 4810 14090 4830 14110
rect 4890 14090 4910 14110
rect 4970 14090 4990 14110
rect 5050 14090 5070 14110
rect 5130 14090 5150 14110
rect 5210 14090 5230 14110
rect 5290 14090 5310 14110
rect 5370 14090 5390 14110
rect 5450 14090 5470 14110
rect 5530 14090 5550 14110
rect 5610 14090 5630 14110
rect 5690 14090 5710 14110
rect 5770 14090 5790 14110
rect 5850 14090 5870 14110
rect 5930 14090 5950 14110
rect 6010 14090 6030 14110
rect 6090 14090 6110 14110
rect 6170 14090 6190 14110
rect 4250 14010 4270 14030
rect 4330 14010 4350 14030
rect 4410 14010 4430 14030
rect 4490 14010 4510 14030
rect 4570 14010 4590 14030
rect 4650 14010 4670 14030
rect 4730 14010 4750 14030
rect 4810 14010 4830 14030
rect 4890 14010 4910 14030
rect 4970 14010 4990 14030
rect 5050 14010 5070 14030
rect 5130 14010 5150 14030
rect 5210 14010 5230 14030
rect 5290 14010 5310 14030
rect 5370 14010 5390 14030
rect 5450 14010 5470 14030
rect 5530 14010 5550 14030
rect 5610 14010 5630 14030
rect 5690 14010 5710 14030
rect 5770 14010 5790 14030
rect 5850 14010 5870 14030
rect 5930 14010 5950 14030
rect 6010 14010 6030 14030
rect 6090 14010 6110 14030
rect 6170 14010 6190 14030
rect 4250 13930 4270 13950
rect 4330 13930 4350 13950
rect 4410 13930 4430 13950
rect 4490 13930 4510 13950
rect 4570 13930 4590 13950
rect 4650 13930 4670 13950
rect 4730 13930 4750 13950
rect 4810 13930 4830 13950
rect 4890 13930 4910 13950
rect 4970 13930 4990 13950
rect 5050 13930 5070 13950
rect 5130 13930 5150 13950
rect 5210 13930 5230 13950
rect 5290 13930 5310 13950
rect 5370 13930 5390 13950
rect 5450 13930 5470 13950
rect 5530 13930 5550 13950
rect 5610 13930 5630 13950
rect 5690 13930 5710 13950
rect 5770 13930 5790 13950
rect 5850 13930 5870 13950
rect 5930 13930 5950 13950
rect 6010 13930 6030 13950
rect 6090 13930 6110 13950
rect 6170 13930 6190 13950
rect 4250 13850 4270 13870
rect 4330 13850 4350 13870
rect 4410 13850 4430 13870
rect 4490 13850 4510 13870
rect 4570 13850 4590 13870
rect 4650 13850 4670 13870
rect 4730 13850 4750 13870
rect 4810 13850 4830 13870
rect 4890 13850 4910 13870
rect 4970 13850 4990 13870
rect 5050 13850 5070 13870
rect 5130 13850 5150 13870
rect 5210 13850 5230 13870
rect 5290 13850 5310 13870
rect 5370 13850 5390 13870
rect 5450 13850 5470 13870
rect 5530 13850 5550 13870
rect 5610 13850 5630 13870
rect 5690 13850 5710 13870
rect 5770 13850 5790 13870
rect 5850 13850 5870 13870
rect 5930 13850 5950 13870
rect 6010 13850 6030 13870
rect 6090 13850 6110 13870
rect 6170 13850 6190 13870
rect 4250 13770 4270 13790
rect 4330 13770 4350 13790
rect 4410 13770 4430 13790
rect 4490 13770 4510 13790
rect 4570 13770 4590 13790
rect 4650 13770 4670 13790
rect 4730 13770 4750 13790
rect 4810 13770 4830 13790
rect 4890 13770 4910 13790
rect 4970 13770 4990 13790
rect 5050 13770 5070 13790
rect 5130 13770 5150 13790
rect 5210 13770 5230 13790
rect 5290 13770 5310 13790
rect 5370 13770 5390 13790
rect 5450 13770 5470 13790
rect 5530 13770 5550 13790
rect 5610 13770 5630 13790
rect 5690 13770 5710 13790
rect 5770 13770 5790 13790
rect 5850 13770 5870 13790
rect 5930 13770 5950 13790
rect 6010 13770 6030 13790
rect 6090 13770 6110 13790
rect 6170 13770 6190 13790
rect 4250 13690 4270 13710
rect 4330 13690 4350 13710
rect 4410 13690 4430 13710
rect 4490 13690 4510 13710
rect 4570 13690 4590 13710
rect 4650 13690 4670 13710
rect 4730 13690 4750 13710
rect 4810 13690 4830 13710
rect 4890 13690 4910 13710
rect 4970 13690 4990 13710
rect 5050 13690 5070 13710
rect 5130 13690 5150 13710
rect 5210 13690 5230 13710
rect 5290 13690 5310 13710
rect 5370 13690 5390 13710
rect 5450 13690 5470 13710
rect 5530 13690 5550 13710
rect 5610 13690 5630 13710
rect 5690 13690 5710 13710
rect 5770 13690 5790 13710
rect 5850 13690 5870 13710
rect 5930 13690 5950 13710
rect 6010 13690 6030 13710
rect 6090 13690 6110 13710
rect 6170 13690 6190 13710
rect 4250 13610 4270 13630
rect 4330 13610 4350 13630
rect 4410 13610 4430 13630
rect 4490 13610 4510 13630
rect 4570 13610 4590 13630
rect 4650 13610 4670 13630
rect 4730 13610 4750 13630
rect 4810 13610 4830 13630
rect 4890 13610 4910 13630
rect 4970 13610 4990 13630
rect 5050 13610 5070 13630
rect 5130 13610 5150 13630
rect 5210 13610 5230 13630
rect 5290 13610 5310 13630
rect 5370 13610 5390 13630
rect 5450 13610 5470 13630
rect 5530 13610 5550 13630
rect 5610 13610 5630 13630
rect 5690 13610 5710 13630
rect 5770 13610 5790 13630
rect 5850 13610 5870 13630
rect 5930 13610 5950 13630
rect 6010 13610 6030 13630
rect 6090 13610 6110 13630
rect 6170 13610 6190 13630
rect 4250 13530 4270 13550
rect 4330 13530 4350 13550
rect 4410 13530 4430 13550
rect 4490 13530 4510 13550
rect 4570 13530 4590 13550
rect 4650 13530 4670 13550
rect 4730 13530 4750 13550
rect 4810 13530 4830 13550
rect 4890 13530 4910 13550
rect 4970 13530 4990 13550
rect 5050 13530 5070 13550
rect 5130 13530 5150 13550
rect 5210 13530 5230 13550
rect 5290 13530 5310 13550
rect 5370 13530 5390 13550
rect 5450 13530 5470 13550
rect 5530 13530 5550 13550
rect 5610 13530 5630 13550
rect 5690 13530 5710 13550
rect 5770 13530 5790 13550
rect 5850 13530 5870 13550
rect 5930 13530 5950 13550
rect 6010 13530 6030 13550
rect 6090 13530 6110 13550
rect 6170 13530 6190 13550
rect 4250 13450 4270 13470
rect 4330 13450 4350 13470
rect 4410 13450 4430 13470
rect 4490 13450 4510 13470
rect 4570 13450 4590 13470
rect 4650 13450 4670 13470
rect 4730 13450 4750 13470
rect 4810 13450 4830 13470
rect 4890 13450 4910 13470
rect 4970 13450 4990 13470
rect 5050 13450 5070 13470
rect 5130 13450 5150 13470
rect 5210 13450 5230 13470
rect 5290 13450 5310 13470
rect 5370 13450 5390 13470
rect 5450 13450 5470 13470
rect 5530 13450 5550 13470
rect 5610 13450 5630 13470
rect 5690 13450 5710 13470
rect 5770 13450 5790 13470
rect 5850 13450 5870 13470
rect 5930 13450 5950 13470
rect 6010 13450 6030 13470
rect 6090 13450 6110 13470
rect 6170 13450 6190 13470
rect 4250 13370 4270 13390
rect 4330 13370 4350 13390
rect 4410 13370 4430 13390
rect 4490 13370 4510 13390
rect 4570 13370 4590 13390
rect 4650 13370 4670 13390
rect 4730 13370 4750 13390
rect 4810 13370 4830 13390
rect 4890 13370 4910 13390
rect 4970 13370 4990 13390
rect 5050 13370 5070 13390
rect 5130 13370 5150 13390
rect 5210 13370 5230 13390
rect 5290 13370 5310 13390
rect 5370 13370 5390 13390
rect 5450 13370 5470 13390
rect 5530 13370 5550 13390
rect 5610 13370 5630 13390
rect 5690 13370 5710 13390
rect 5770 13370 5790 13390
rect 5850 13370 5870 13390
rect 5930 13370 5950 13390
rect 6010 13370 6030 13390
rect 6090 13370 6110 13390
rect 6170 13370 6190 13390
rect 4250 13290 4270 13310
rect 4330 13290 4350 13310
rect 4410 13290 4430 13310
rect 4490 13290 4510 13310
rect 4570 13290 4590 13310
rect 4650 13290 4670 13310
rect 4730 13290 4750 13310
rect 4810 13290 4830 13310
rect 4890 13290 4910 13310
rect 4970 13290 4990 13310
rect 5050 13290 5070 13310
rect 5130 13290 5150 13310
rect 5210 13290 5230 13310
rect 5290 13290 5310 13310
rect 5370 13290 5390 13310
rect 5450 13290 5470 13310
rect 5530 13290 5550 13310
rect 5610 13290 5630 13310
rect 5690 13290 5710 13310
rect 5770 13290 5790 13310
rect 5850 13290 5870 13310
rect 5930 13290 5950 13310
rect 6010 13290 6030 13310
rect 6090 13290 6110 13310
rect 6170 13290 6190 13310
rect 4250 13210 4270 13230
rect 4330 13210 4350 13230
rect 4410 13210 4430 13230
rect 4490 13210 4510 13230
rect 4570 13210 4590 13230
rect 4650 13210 4670 13230
rect 4730 13210 4750 13230
rect 4810 13210 4830 13230
rect 4890 13210 4910 13230
rect 4970 13210 4990 13230
rect 5050 13210 5070 13230
rect 5130 13210 5150 13230
rect 5210 13210 5230 13230
rect 5290 13210 5310 13230
rect 5370 13210 5390 13230
rect 5450 13210 5470 13230
rect 5530 13210 5550 13230
rect 5610 13210 5630 13230
rect 5690 13210 5710 13230
rect 5770 13210 5790 13230
rect 5850 13210 5870 13230
rect 5930 13210 5950 13230
rect 6010 13210 6030 13230
rect 6090 13210 6110 13230
rect 6170 13210 6190 13230
rect 4250 13130 4270 13150
rect 4330 13130 4350 13150
rect 4410 13130 4430 13150
rect 4490 13130 4510 13150
rect 4570 13130 4590 13150
rect 4650 13130 4670 13150
rect 4730 13130 4750 13150
rect 4810 13130 4830 13150
rect 4890 13130 4910 13150
rect 4970 13130 4990 13150
rect 5050 13130 5070 13150
rect 5130 13130 5150 13150
rect 5210 13130 5230 13150
rect 5290 13130 5310 13150
rect 5370 13130 5390 13150
rect 5450 13130 5470 13150
rect 5530 13130 5550 13150
rect 5610 13130 5630 13150
rect 5690 13130 5710 13150
rect 5770 13130 5790 13150
rect 5850 13130 5870 13150
rect 5930 13130 5950 13150
rect 6010 13130 6030 13150
rect 6090 13130 6110 13150
rect 6170 13130 6190 13150
rect 4250 13050 4270 13070
rect 4330 13050 4350 13070
rect 4410 13050 4430 13070
rect 4490 13050 4510 13070
rect 4570 13050 4590 13070
rect 4650 13050 4670 13070
rect 4730 13050 4750 13070
rect 4810 13050 4830 13070
rect 4890 13050 4910 13070
rect 4970 13050 4990 13070
rect 5050 13050 5070 13070
rect 5130 13050 5150 13070
rect 5210 13050 5230 13070
rect 5290 13050 5310 13070
rect 5370 13050 5390 13070
rect 5450 13050 5470 13070
rect 5530 13050 5550 13070
rect 5610 13050 5630 13070
rect 5690 13050 5710 13070
rect 5770 13050 5790 13070
rect 5850 13050 5870 13070
rect 5930 13050 5950 13070
rect 6010 13050 6030 13070
rect 6090 13050 6110 13070
rect 6170 13050 6190 13070
rect 4250 12970 4270 12990
rect 4330 12970 4350 12990
rect 4410 12970 4430 12990
rect 4490 12970 4510 12990
rect 4570 12970 4590 12990
rect 4650 12970 4670 12990
rect 4730 12970 4750 12990
rect 4810 12970 4830 12990
rect 4890 12970 4910 12990
rect 4970 12970 4990 12990
rect 5050 12970 5070 12990
rect 5130 12970 5150 12990
rect 5210 12970 5230 12990
rect 5290 12970 5310 12990
rect 5370 12970 5390 12990
rect 5450 12970 5470 12990
rect 5530 12970 5550 12990
rect 5610 12970 5630 12990
rect 5690 12970 5710 12990
rect 5770 12970 5790 12990
rect 5850 12970 5870 12990
rect 5930 12970 5950 12990
rect 6010 12970 6030 12990
rect 6090 12970 6110 12990
rect 6170 12970 6190 12990
rect 4250 12890 4270 12910
rect 4330 12890 4350 12910
rect 4410 12890 4430 12910
rect 4490 12890 4510 12910
rect 4570 12890 4590 12910
rect 4650 12890 4670 12910
rect 4730 12890 4750 12910
rect 4810 12890 4830 12910
rect 4890 12890 4910 12910
rect 4970 12890 4990 12910
rect 5050 12890 5070 12910
rect 5130 12890 5150 12910
rect 5210 12890 5230 12910
rect 5290 12890 5310 12910
rect 5370 12890 5390 12910
rect 5450 12890 5470 12910
rect 5530 12890 5550 12910
rect 5610 12890 5630 12910
rect 5690 12890 5710 12910
rect 5770 12890 5790 12910
rect 5850 12890 5870 12910
rect 5930 12890 5950 12910
rect 6010 12890 6030 12910
rect 6090 12890 6110 12910
rect 6170 12890 6190 12910
rect 4250 12810 4270 12830
rect 4330 12810 4350 12830
rect 4410 12810 4430 12830
rect 4490 12810 4510 12830
rect 4570 12810 4590 12830
rect 4650 12810 4670 12830
rect 4730 12810 4750 12830
rect 4810 12810 4830 12830
rect 4890 12810 4910 12830
rect 4970 12810 4990 12830
rect 5050 12810 5070 12830
rect 5130 12810 5150 12830
rect 5210 12810 5230 12830
rect 5290 12810 5310 12830
rect 5370 12810 5390 12830
rect 5450 12810 5470 12830
rect 5530 12810 5550 12830
rect 5610 12810 5630 12830
rect 5690 12810 5710 12830
rect 5770 12810 5790 12830
rect 5850 12810 5870 12830
rect 5930 12810 5950 12830
rect 6010 12810 6030 12830
rect 6090 12810 6110 12830
rect 6170 12810 6190 12830
rect 4250 12730 4270 12750
rect 4330 12730 4350 12750
rect 4410 12730 4430 12750
rect 4490 12730 4510 12750
rect 4570 12730 4590 12750
rect 4650 12730 4670 12750
rect 4730 12730 4750 12750
rect 4810 12730 4830 12750
rect 4890 12730 4910 12750
rect 4970 12730 4990 12750
rect 5050 12730 5070 12750
rect 5130 12730 5150 12750
rect 5210 12730 5230 12750
rect 5290 12730 5310 12750
rect 5370 12730 5390 12750
rect 5450 12730 5470 12750
rect 5530 12730 5550 12750
rect 5610 12730 5630 12750
rect 5690 12730 5710 12750
rect 5770 12730 5790 12750
rect 5850 12730 5870 12750
rect 5930 12730 5950 12750
rect 6010 12730 6030 12750
rect 6090 12730 6110 12750
rect 6170 12730 6190 12750
rect 4250 12650 4270 12670
rect 4330 12650 4350 12670
rect 4410 12650 4430 12670
rect 4490 12650 4510 12670
rect 4570 12650 4590 12670
rect 4650 12650 4670 12670
rect 4730 12650 4750 12670
rect 4810 12650 4830 12670
rect 4890 12650 4910 12670
rect 4970 12650 4990 12670
rect 5050 12650 5070 12670
rect 5130 12650 5150 12670
rect 5210 12650 5230 12670
rect 5290 12650 5310 12670
rect 5370 12650 5390 12670
rect 5450 12650 5470 12670
rect 5530 12650 5550 12670
rect 5610 12650 5630 12670
rect 5690 12650 5710 12670
rect 5770 12650 5790 12670
rect 5850 12650 5870 12670
rect 5930 12650 5950 12670
rect 6010 12650 6030 12670
rect 6090 12650 6110 12670
rect 6170 12650 6190 12670
rect 4250 12570 4270 12590
rect 4330 12570 4350 12590
rect 4410 12570 4430 12590
rect 4490 12570 4510 12590
rect 4570 12570 4590 12590
rect 4650 12570 4670 12590
rect 4730 12570 4750 12590
rect 4810 12570 4830 12590
rect 4890 12570 4910 12590
rect 4970 12570 4990 12590
rect 5050 12570 5070 12590
rect 5130 12570 5150 12590
rect 5210 12570 5230 12590
rect 5290 12570 5310 12590
rect 5370 12570 5390 12590
rect 5450 12570 5470 12590
rect 5530 12570 5550 12590
rect 5610 12570 5630 12590
rect 5690 12570 5710 12590
rect 5770 12570 5790 12590
rect 5850 12570 5870 12590
rect 5930 12570 5950 12590
rect 6010 12570 6030 12590
rect 6090 12570 6110 12590
rect 6170 12570 6190 12590
rect 4250 12490 4270 12510
rect 4330 12490 4350 12510
rect 4410 12490 4430 12510
rect 4490 12490 4510 12510
rect 4570 12490 4590 12510
rect 4650 12490 4670 12510
rect 4730 12490 4750 12510
rect 4810 12490 4830 12510
rect 4890 12490 4910 12510
rect 4970 12490 4990 12510
rect 5050 12490 5070 12510
rect 5130 12490 5150 12510
rect 5210 12490 5230 12510
rect 5290 12490 5310 12510
rect 5370 12490 5390 12510
rect 5450 12490 5470 12510
rect 5530 12490 5550 12510
rect 5610 12490 5630 12510
rect 5690 12490 5710 12510
rect 5770 12490 5790 12510
rect 5850 12490 5870 12510
rect 5930 12490 5950 12510
rect 6010 12490 6030 12510
rect 6090 12490 6110 12510
rect 6170 12490 6190 12510
rect 4250 12410 4270 12430
rect 4330 12410 4350 12430
rect 4410 12410 4430 12430
rect 4490 12410 4510 12430
rect 4570 12410 4590 12430
rect 4650 12410 4670 12430
rect 4730 12410 4750 12430
rect 4810 12410 4830 12430
rect 4890 12410 4910 12430
rect 4970 12410 4990 12430
rect 5050 12410 5070 12430
rect 5130 12410 5150 12430
rect 5210 12410 5230 12430
rect 5290 12410 5310 12430
rect 5370 12410 5390 12430
rect 5450 12410 5470 12430
rect 5530 12410 5550 12430
rect 5610 12410 5630 12430
rect 5690 12410 5710 12430
rect 5770 12410 5790 12430
rect 5850 12410 5870 12430
rect 5930 12410 5950 12430
rect 6010 12410 6030 12430
rect 6090 12410 6110 12430
rect 6170 12410 6190 12430
rect 4250 12330 4270 12350
rect 4330 12330 4350 12350
rect 4410 12330 4430 12350
rect 4490 12330 4510 12350
rect 4570 12330 4590 12350
rect 4650 12330 4670 12350
rect 4730 12330 4750 12350
rect 4810 12330 4830 12350
rect 4890 12330 4910 12350
rect 4970 12330 4990 12350
rect 5050 12330 5070 12350
rect 5130 12330 5150 12350
rect 5210 12330 5230 12350
rect 5290 12330 5310 12350
rect 5370 12330 5390 12350
rect 5450 12330 5470 12350
rect 5530 12330 5550 12350
rect 5610 12330 5630 12350
rect 5690 12330 5710 12350
rect 5770 12330 5790 12350
rect 5850 12330 5870 12350
rect 5930 12330 5950 12350
rect 6010 12330 6030 12350
rect 6090 12330 6110 12350
rect 6170 12330 6190 12350
rect 4250 12250 4270 12270
rect 4330 12250 4350 12270
rect 4410 12250 4430 12270
rect 4490 12250 4510 12270
rect 4570 12250 4590 12270
rect 4650 12250 4670 12270
rect 4730 12250 4750 12270
rect 4810 12250 4830 12270
rect 4890 12250 4910 12270
rect 4970 12250 4990 12270
rect 5050 12250 5070 12270
rect 5130 12250 5150 12270
rect 5210 12250 5230 12270
rect 5290 12250 5310 12270
rect 5370 12250 5390 12270
rect 5450 12250 5470 12270
rect 5530 12250 5550 12270
rect 5610 12250 5630 12270
rect 5690 12250 5710 12270
rect 5770 12250 5790 12270
rect 5850 12250 5870 12270
rect 5930 12250 5950 12270
rect 6010 12250 6030 12270
rect 6090 12250 6110 12270
rect 6170 12250 6190 12270
rect 4250 12170 4270 12190
rect 4330 12170 4350 12190
rect 4410 12170 4430 12190
rect 4490 12170 4510 12190
rect 4570 12170 4590 12190
rect 4650 12170 4670 12190
rect 4730 12170 4750 12190
rect 4810 12170 4830 12190
rect 4890 12170 4910 12190
rect 4970 12170 4990 12190
rect 5050 12170 5070 12190
rect 5130 12170 5150 12190
rect 5210 12170 5230 12190
rect 5290 12170 5310 12190
rect 5370 12170 5390 12190
rect 5450 12170 5470 12190
rect 5530 12170 5550 12190
rect 5610 12170 5630 12190
rect 5690 12170 5710 12190
rect 5770 12170 5790 12190
rect 5850 12170 5870 12190
rect 5930 12170 5950 12190
rect 6010 12170 6030 12190
rect 6090 12170 6110 12190
rect 6170 12170 6190 12190
rect 4250 12090 4270 12110
rect 4330 12090 4350 12110
rect 4410 12090 4430 12110
rect 4490 12090 4510 12110
rect 4570 12090 4590 12110
rect 4650 12090 4670 12110
rect 4730 12090 4750 12110
rect 4810 12090 4830 12110
rect 4890 12090 4910 12110
rect 4970 12090 4990 12110
rect 5050 12090 5070 12110
rect 5130 12090 5150 12110
rect 5210 12090 5230 12110
rect 5290 12090 5310 12110
rect 5370 12090 5390 12110
rect 5450 12090 5470 12110
rect 5530 12090 5550 12110
rect 5610 12090 5630 12110
rect 5690 12090 5710 12110
rect 5770 12090 5790 12110
rect 5850 12090 5870 12110
rect 5930 12090 5950 12110
rect 6010 12090 6030 12110
rect 6090 12090 6110 12110
rect 6170 12090 6190 12110
rect 4250 12010 4270 12030
rect 4330 12010 4350 12030
rect 4410 12010 4430 12030
rect 4490 12010 4510 12030
rect 4570 12010 4590 12030
rect 4650 12010 4670 12030
rect 4730 12010 4750 12030
rect 4810 12010 4830 12030
rect 4890 12010 4910 12030
rect 4970 12010 4990 12030
rect 5050 12010 5070 12030
rect 5130 12010 5150 12030
rect 5210 12010 5230 12030
rect 5290 12010 5310 12030
rect 5370 12010 5390 12030
rect 5450 12010 5470 12030
rect 5530 12010 5550 12030
rect 5610 12010 5630 12030
rect 5690 12010 5710 12030
rect 5770 12010 5790 12030
rect 5850 12010 5870 12030
rect 5930 12010 5950 12030
rect 6010 12010 6030 12030
rect 6090 12010 6110 12030
rect 6170 12010 6190 12030
rect 4250 11930 4270 11950
rect 4330 11930 4350 11950
rect 4410 11930 4430 11950
rect 4490 11930 4510 11950
rect 4570 11930 4590 11950
rect 4650 11930 4670 11950
rect 4730 11930 4750 11950
rect 4810 11930 4830 11950
rect 4890 11930 4910 11950
rect 4970 11930 4990 11950
rect 5050 11930 5070 11950
rect 5130 11930 5150 11950
rect 5210 11930 5230 11950
rect 5290 11930 5310 11950
rect 5370 11930 5390 11950
rect 5450 11930 5470 11950
rect 5530 11930 5550 11950
rect 5610 11930 5630 11950
rect 5690 11930 5710 11950
rect 5770 11930 5790 11950
rect 5850 11930 5870 11950
rect 5930 11930 5950 11950
rect 6010 11930 6030 11950
rect 6090 11930 6110 11950
rect 6170 11930 6190 11950
rect 4250 11850 4270 11870
rect 4330 11850 4350 11870
rect 4410 11850 4430 11870
rect 4490 11850 4510 11870
rect 4570 11850 4590 11870
rect 4650 11850 4670 11870
rect 4730 11850 4750 11870
rect 4810 11850 4830 11870
rect 4890 11850 4910 11870
rect 4970 11850 4990 11870
rect 5050 11850 5070 11870
rect 5130 11850 5150 11870
rect 5210 11850 5230 11870
rect 5290 11850 5310 11870
rect 5370 11850 5390 11870
rect 5450 11850 5470 11870
rect 5530 11850 5550 11870
rect 5610 11850 5630 11870
rect 5690 11850 5710 11870
rect 5770 11850 5790 11870
rect 5850 11850 5870 11870
rect 5930 11850 5950 11870
rect 6010 11850 6030 11870
rect 6090 11850 6110 11870
rect 6170 11850 6190 11870
rect 4250 11770 4270 11790
rect 4330 11770 4350 11790
rect 4410 11770 4430 11790
rect 4490 11770 4510 11790
rect 4570 11770 4590 11790
rect 4650 11770 4670 11790
rect 4730 11770 4750 11790
rect 4810 11770 4830 11790
rect 4890 11770 4910 11790
rect 4970 11770 4990 11790
rect 5050 11770 5070 11790
rect 5130 11770 5150 11790
rect 5210 11770 5230 11790
rect 5290 11770 5310 11790
rect 5370 11770 5390 11790
rect 5450 11770 5470 11790
rect 5530 11770 5550 11790
rect 5610 11770 5630 11790
rect 5690 11770 5710 11790
rect 5770 11770 5790 11790
rect 5850 11770 5870 11790
rect 5930 11770 5950 11790
rect 6010 11770 6030 11790
rect 6090 11770 6110 11790
rect 6170 11770 6190 11790
rect 4250 11690 4270 11710
rect 4330 11690 4350 11710
rect 4410 11690 4430 11710
rect 4490 11690 4510 11710
rect 4570 11690 4590 11710
rect 4650 11690 4670 11710
rect 4730 11690 4750 11710
rect 4810 11690 4830 11710
rect 4890 11690 4910 11710
rect 4970 11690 4990 11710
rect 5050 11690 5070 11710
rect 5130 11690 5150 11710
rect 5210 11690 5230 11710
rect 5290 11690 5310 11710
rect 5370 11690 5390 11710
rect 5450 11690 5470 11710
rect 5530 11690 5550 11710
rect 5610 11690 5630 11710
rect 5690 11690 5710 11710
rect 5770 11690 5790 11710
rect 5850 11690 5870 11710
rect 5930 11690 5950 11710
rect 6010 11690 6030 11710
rect 6090 11690 6110 11710
rect 6170 11690 6190 11710
rect 4250 11610 4270 11630
rect 4330 11610 4350 11630
rect 4410 11610 4430 11630
rect 4490 11610 4510 11630
rect 4570 11610 4590 11630
rect 4650 11610 4670 11630
rect 4730 11610 4750 11630
rect 4810 11610 4830 11630
rect 4890 11610 4910 11630
rect 4970 11610 4990 11630
rect 5050 11610 5070 11630
rect 5130 11610 5150 11630
rect 5210 11610 5230 11630
rect 5290 11610 5310 11630
rect 5370 11610 5390 11630
rect 5450 11610 5470 11630
rect 5530 11610 5550 11630
rect 5610 11610 5630 11630
rect 5690 11610 5710 11630
rect 5770 11610 5790 11630
rect 5850 11610 5870 11630
rect 5930 11610 5950 11630
rect 6010 11610 6030 11630
rect 6090 11610 6110 11630
rect 6170 11610 6190 11630
rect 4250 11530 4270 11550
rect 4330 11530 4350 11550
rect 4410 11530 4430 11550
rect 4490 11530 4510 11550
rect 4570 11530 4590 11550
rect 4650 11530 4670 11550
rect 4730 11530 4750 11550
rect 4810 11530 4830 11550
rect 4890 11530 4910 11550
rect 4970 11530 4990 11550
rect 5050 11530 5070 11550
rect 5130 11530 5150 11550
rect 5210 11530 5230 11550
rect 5290 11530 5310 11550
rect 5370 11530 5390 11550
rect 5450 11530 5470 11550
rect 5530 11530 5550 11550
rect 5610 11530 5630 11550
rect 5690 11530 5710 11550
rect 5770 11530 5790 11550
rect 5850 11530 5870 11550
rect 5930 11530 5950 11550
rect 6010 11530 6030 11550
rect 6090 11530 6110 11550
rect 6170 11530 6190 11550
rect 4250 11450 4270 11470
rect 4330 11450 4350 11470
rect 4410 11450 4430 11470
rect 4490 11450 4510 11470
rect 4570 11450 4590 11470
rect 4650 11450 4670 11470
rect 4730 11450 4750 11470
rect 4810 11450 4830 11470
rect 4890 11450 4910 11470
rect 4970 11450 4990 11470
rect 5050 11450 5070 11470
rect 5130 11450 5150 11470
rect 5210 11450 5230 11470
rect 5290 11450 5310 11470
rect 5370 11450 5390 11470
rect 5450 11450 5470 11470
rect 5530 11450 5550 11470
rect 5610 11450 5630 11470
rect 5690 11450 5710 11470
rect 5770 11450 5790 11470
rect 5850 11450 5870 11470
rect 5930 11450 5950 11470
rect 6010 11450 6030 11470
rect 6090 11450 6110 11470
rect 6170 11450 6190 11470
rect 4250 11370 4270 11390
rect 4330 11370 4350 11390
rect 4410 11370 4430 11390
rect 4490 11370 4510 11390
rect 4570 11370 4590 11390
rect 4650 11370 4670 11390
rect 4730 11370 4750 11390
rect 4810 11370 4830 11390
rect 4890 11370 4910 11390
rect 4970 11370 4990 11390
rect 5050 11370 5070 11390
rect 5130 11370 5150 11390
rect 5210 11370 5230 11390
rect 5290 11370 5310 11390
rect 5370 11370 5390 11390
rect 5450 11370 5470 11390
rect 5530 11370 5550 11390
rect 5610 11370 5630 11390
rect 5690 11370 5710 11390
rect 5770 11370 5790 11390
rect 5850 11370 5870 11390
rect 5930 11370 5950 11390
rect 6010 11370 6030 11390
rect 6090 11370 6110 11390
rect 6170 11370 6190 11390
rect 4250 11290 4270 11310
rect 4330 11290 4350 11310
rect 4410 11290 4430 11310
rect 4490 11290 4510 11310
rect 4570 11290 4590 11310
rect 4650 11290 4670 11310
rect 4730 11290 4750 11310
rect 4810 11290 4830 11310
rect 4890 11290 4910 11310
rect 4970 11290 4990 11310
rect 5050 11290 5070 11310
rect 5130 11290 5150 11310
rect 5210 11290 5230 11310
rect 5290 11290 5310 11310
rect 5370 11290 5390 11310
rect 5450 11290 5470 11310
rect 5530 11290 5550 11310
rect 5610 11290 5630 11310
rect 5690 11290 5710 11310
rect 5770 11290 5790 11310
rect 5850 11290 5870 11310
rect 5930 11290 5950 11310
rect 6010 11290 6030 11310
rect 6090 11290 6110 11310
rect 6170 11290 6190 11310
rect 4250 11210 4270 11230
rect 4330 11210 4350 11230
rect 4410 11210 4430 11230
rect 4490 11210 4510 11230
rect 4570 11210 4590 11230
rect 4650 11210 4670 11230
rect 4730 11210 4750 11230
rect 4810 11210 4830 11230
rect 4890 11210 4910 11230
rect 4970 11210 4990 11230
rect 5050 11210 5070 11230
rect 5130 11210 5150 11230
rect 5210 11210 5230 11230
rect 5290 11210 5310 11230
rect 5370 11210 5390 11230
rect 5450 11210 5470 11230
rect 5530 11210 5550 11230
rect 5610 11210 5630 11230
rect 5690 11210 5710 11230
rect 5770 11210 5790 11230
rect 5850 11210 5870 11230
rect 5930 11210 5950 11230
rect 6010 11210 6030 11230
rect 6090 11210 6110 11230
rect 6170 11210 6190 11230
rect 4250 11130 4270 11150
rect 4330 11130 4350 11150
rect 4410 11130 4430 11150
rect 4490 11130 4510 11150
rect 4570 11130 4590 11150
rect 4650 11130 4670 11150
rect 4730 11130 4750 11150
rect 4810 11130 4830 11150
rect 4890 11130 4910 11150
rect 4970 11130 4990 11150
rect 5050 11130 5070 11150
rect 5130 11130 5150 11150
rect 5210 11130 5230 11150
rect 5290 11130 5310 11150
rect 5370 11130 5390 11150
rect 5450 11130 5470 11150
rect 5530 11130 5550 11150
rect 5610 11130 5630 11150
rect 5690 11130 5710 11150
rect 5770 11130 5790 11150
rect 5850 11130 5870 11150
rect 5930 11130 5950 11150
rect 6010 11130 6030 11150
rect 6090 11130 6110 11150
rect 6170 11130 6190 11150
rect 4250 11050 4270 11070
rect 4330 11050 4350 11070
rect 4410 11050 4430 11070
rect 4490 11050 4510 11070
rect 4570 11050 4590 11070
rect 4650 11050 4670 11070
rect 4730 11050 4750 11070
rect 4810 11050 4830 11070
rect 4890 11050 4910 11070
rect 4970 11050 4990 11070
rect 5050 11050 5070 11070
rect 5130 11050 5150 11070
rect 5210 11050 5230 11070
rect 5290 11050 5310 11070
rect 5370 11050 5390 11070
rect 5450 11050 5470 11070
rect 5530 11050 5550 11070
rect 5610 11050 5630 11070
rect 5690 11050 5710 11070
rect 5770 11050 5790 11070
rect 5850 11050 5870 11070
rect 5930 11050 5950 11070
rect 6010 11050 6030 11070
rect 6090 11050 6110 11070
rect 6170 11050 6190 11070
rect 4250 10970 4270 10990
rect 4330 10970 4350 10990
rect 4410 10970 4430 10990
rect 4490 10970 4510 10990
rect 4570 10970 4590 10990
rect 4650 10970 4670 10990
rect 4730 10970 4750 10990
rect 4810 10970 4830 10990
rect 4890 10970 4910 10990
rect 4970 10970 4990 10990
rect 5050 10970 5070 10990
rect 5130 10970 5150 10990
rect 5210 10970 5230 10990
rect 5290 10970 5310 10990
rect 5370 10970 5390 10990
rect 5450 10970 5470 10990
rect 5530 10970 5550 10990
rect 5610 10970 5630 10990
rect 5690 10970 5710 10990
rect 5770 10970 5790 10990
rect 5850 10970 5870 10990
rect 5930 10970 5950 10990
rect 6010 10970 6030 10990
rect 6090 10970 6110 10990
rect 6170 10970 6190 10990
rect 4250 10890 4270 10910
rect 4330 10890 4350 10910
rect 4410 10890 4430 10910
rect 4490 10890 4510 10910
rect 4570 10890 4590 10910
rect 4650 10890 4670 10910
rect 4730 10890 4750 10910
rect 4810 10890 4830 10910
rect 4890 10890 4910 10910
rect 4970 10890 4990 10910
rect 5050 10890 5070 10910
rect 5130 10890 5150 10910
rect 5210 10890 5230 10910
rect 5290 10890 5310 10910
rect 5370 10890 5390 10910
rect 5450 10890 5470 10910
rect 5530 10890 5550 10910
rect 5610 10890 5630 10910
rect 5690 10890 5710 10910
rect 5770 10890 5790 10910
rect 5850 10890 5870 10910
rect 5930 10890 5950 10910
rect 6010 10890 6030 10910
rect 6090 10890 6110 10910
rect 6170 10890 6190 10910
rect 4250 10810 4270 10830
rect 4330 10810 4350 10830
rect 4410 10810 4430 10830
rect 4490 10810 4510 10830
rect 4570 10810 4590 10830
rect 4650 10810 4670 10830
rect 4730 10810 4750 10830
rect 4810 10810 4830 10830
rect 4890 10810 4910 10830
rect 4970 10810 4990 10830
rect 5050 10810 5070 10830
rect 5130 10810 5150 10830
rect 5210 10810 5230 10830
rect 5290 10810 5310 10830
rect 5370 10810 5390 10830
rect 5450 10810 5470 10830
rect 5530 10810 5550 10830
rect 5610 10810 5630 10830
rect 5690 10810 5710 10830
rect 5770 10810 5790 10830
rect 5850 10810 5870 10830
rect 5930 10810 5950 10830
rect 6010 10810 6030 10830
rect 6090 10810 6110 10830
rect 6170 10810 6190 10830
rect 4250 10730 4270 10750
rect 4330 10730 4350 10750
rect 4410 10730 4430 10750
rect 4490 10730 4510 10750
rect 4570 10730 4590 10750
rect 4650 10730 4670 10750
rect 4730 10730 4750 10750
rect 4810 10730 4830 10750
rect 4890 10730 4910 10750
rect 4970 10730 4990 10750
rect 5050 10730 5070 10750
rect 5130 10730 5150 10750
rect 5210 10730 5230 10750
rect 5290 10730 5310 10750
rect 5370 10730 5390 10750
rect 5450 10730 5470 10750
rect 5530 10730 5550 10750
rect 5610 10730 5630 10750
rect 5690 10730 5710 10750
rect 5770 10730 5790 10750
rect 5850 10730 5870 10750
rect 5930 10730 5950 10750
rect 6010 10730 6030 10750
rect 6090 10730 6110 10750
rect 6170 10730 6190 10750
rect 4250 10650 4270 10670
rect 4330 10650 4350 10670
rect 4410 10650 4430 10670
rect 4490 10650 4510 10670
rect 4570 10650 4590 10670
rect 4650 10650 4670 10670
rect 4730 10650 4750 10670
rect 4810 10650 4830 10670
rect 4890 10650 4910 10670
rect 4970 10650 4990 10670
rect 5050 10650 5070 10670
rect 5130 10650 5150 10670
rect 5210 10650 5230 10670
rect 5290 10650 5310 10670
rect 5370 10650 5390 10670
rect 5450 10650 5470 10670
rect 5530 10650 5550 10670
rect 5610 10650 5630 10670
rect 5690 10650 5710 10670
rect 5770 10650 5790 10670
rect 5850 10650 5870 10670
rect 5930 10650 5950 10670
rect 6010 10650 6030 10670
rect 6090 10650 6110 10670
rect 6170 10650 6190 10670
rect 4250 10570 4270 10590
rect 4330 10570 4350 10590
rect 4410 10570 4430 10590
rect 4490 10570 4510 10590
rect 4570 10570 4590 10590
rect 4650 10570 4670 10590
rect 4730 10570 4750 10590
rect 4810 10570 4830 10590
rect 4890 10570 4910 10590
rect 4970 10570 4990 10590
rect 5050 10570 5070 10590
rect 5130 10570 5150 10590
rect 5210 10570 5230 10590
rect 5290 10570 5310 10590
rect 5370 10570 5390 10590
rect 5450 10570 5470 10590
rect 5530 10570 5550 10590
rect 5610 10570 5630 10590
rect 5690 10570 5710 10590
rect 5770 10570 5790 10590
rect 5850 10570 5870 10590
rect 5930 10570 5950 10590
rect 6010 10570 6030 10590
rect 6090 10570 6110 10590
rect 6170 10570 6190 10590
rect 4250 10490 4270 10510
rect 4330 10490 4350 10510
rect 4410 10490 4430 10510
rect 4490 10490 4510 10510
rect 4570 10490 4590 10510
rect 4650 10490 4670 10510
rect 4730 10490 4750 10510
rect 4810 10490 4830 10510
rect 4890 10490 4910 10510
rect 4970 10490 4990 10510
rect 5050 10490 5070 10510
rect 5130 10490 5150 10510
rect 5210 10490 5230 10510
rect 5290 10490 5310 10510
rect 5370 10490 5390 10510
rect 5450 10490 5470 10510
rect 5530 10490 5550 10510
rect 5610 10490 5630 10510
rect 5690 10490 5710 10510
rect 5770 10490 5790 10510
rect 5850 10490 5870 10510
rect 5930 10490 5950 10510
rect 6010 10490 6030 10510
rect 6090 10490 6110 10510
rect 6170 10490 6190 10510
rect 4250 10410 4270 10430
rect 4330 10410 4350 10430
rect 4410 10410 4430 10430
rect 4490 10410 4510 10430
rect 4570 10410 4590 10430
rect 4650 10410 4670 10430
rect 4730 10410 4750 10430
rect 4810 10410 4830 10430
rect 4890 10410 4910 10430
rect 4970 10410 4990 10430
rect 5050 10410 5070 10430
rect 5130 10410 5150 10430
rect 5210 10410 5230 10430
rect 5290 10410 5310 10430
rect 5370 10410 5390 10430
rect 5450 10410 5470 10430
rect 5530 10410 5550 10430
rect 5610 10410 5630 10430
rect 5690 10410 5710 10430
rect 5770 10410 5790 10430
rect 5850 10410 5870 10430
rect 5930 10410 5950 10430
rect 6010 10410 6030 10430
rect 6090 10410 6110 10430
rect 6170 10410 6190 10430
rect 4250 10330 4270 10350
rect 4330 10330 4350 10350
rect 4410 10330 4430 10350
rect 4490 10330 4510 10350
rect 4570 10330 4590 10350
rect 4650 10330 4670 10350
rect 4730 10330 4750 10350
rect 4810 10330 4830 10350
rect 4890 10330 4910 10350
rect 4970 10330 4990 10350
rect 5050 10330 5070 10350
rect 5130 10330 5150 10350
rect 5210 10330 5230 10350
rect 5290 10330 5310 10350
rect 5370 10330 5390 10350
rect 5450 10330 5470 10350
rect 5530 10330 5550 10350
rect 5610 10330 5630 10350
rect 5690 10330 5710 10350
rect 5770 10330 5790 10350
rect 5850 10330 5870 10350
rect 5930 10330 5950 10350
rect 6010 10330 6030 10350
rect 6090 10330 6110 10350
rect 6170 10330 6190 10350
rect 4250 10250 4270 10270
rect 4330 10250 4350 10270
rect 4410 10250 4430 10270
rect 4490 10250 4510 10270
rect 4570 10250 4590 10270
rect 4650 10250 4670 10270
rect 4730 10250 4750 10270
rect 4810 10250 4830 10270
rect 4890 10250 4910 10270
rect 4970 10250 4990 10270
rect 5050 10250 5070 10270
rect 5130 10250 5150 10270
rect 5210 10250 5230 10270
rect 5290 10250 5310 10270
rect 5370 10250 5390 10270
rect 5450 10250 5470 10270
rect 5530 10250 5550 10270
rect 5610 10250 5630 10270
rect 5690 10250 5710 10270
rect 5770 10250 5790 10270
rect 5850 10250 5870 10270
rect 5930 10250 5950 10270
rect 6010 10250 6030 10270
rect 6090 10250 6110 10270
rect 6170 10250 6190 10270
rect 4250 10170 4270 10190
rect 4330 10170 4350 10190
rect 4410 10170 4430 10190
rect 4490 10170 4510 10190
rect 4570 10170 4590 10190
rect 4650 10170 4670 10190
rect 4730 10170 4750 10190
rect 4810 10170 4830 10190
rect 4890 10170 4910 10190
rect 4970 10170 4990 10190
rect 5050 10170 5070 10190
rect 5130 10170 5150 10190
rect 5210 10170 5230 10190
rect 5290 10170 5310 10190
rect 5370 10170 5390 10190
rect 5450 10170 5470 10190
rect 5530 10170 5550 10190
rect 5610 10170 5630 10190
rect 5690 10170 5710 10190
rect 5770 10170 5790 10190
rect 5850 10170 5870 10190
rect 5930 10170 5950 10190
rect 6010 10170 6030 10190
rect 6090 10170 6110 10190
rect 6170 10170 6190 10190
rect 4250 10090 4270 10110
rect 4330 10090 4350 10110
rect 4410 10090 4430 10110
rect 4490 10090 4510 10110
rect 4570 10090 4590 10110
rect 4650 10090 4670 10110
rect 4730 10090 4750 10110
rect 4810 10090 4830 10110
rect 4890 10090 4910 10110
rect 4970 10090 4990 10110
rect 5050 10090 5070 10110
rect 5130 10090 5150 10110
rect 5210 10090 5230 10110
rect 5290 10090 5310 10110
rect 5370 10090 5390 10110
rect 5450 10090 5470 10110
rect 5530 10090 5550 10110
rect 5610 10090 5630 10110
rect 5690 10090 5710 10110
rect 5770 10090 5790 10110
rect 5850 10090 5870 10110
rect 5930 10090 5950 10110
rect 6010 10090 6030 10110
rect 6090 10090 6110 10110
rect 6170 10090 6190 10110
rect 4250 10010 4270 10030
rect 4330 10010 4350 10030
rect 4410 10010 4430 10030
rect 4490 10010 4510 10030
rect 4570 10010 4590 10030
rect 4650 10010 4670 10030
rect 4730 10010 4750 10030
rect 4810 10010 4830 10030
rect 4890 10010 4910 10030
rect 4970 10010 4990 10030
rect 5050 10010 5070 10030
rect 5130 10010 5150 10030
rect 5210 10010 5230 10030
rect 5290 10010 5310 10030
rect 5370 10010 5390 10030
rect 5450 10010 5470 10030
rect 5530 10010 5550 10030
rect 5610 10010 5630 10030
rect 5690 10010 5710 10030
rect 5770 10010 5790 10030
rect 5850 10010 5870 10030
rect 5930 10010 5950 10030
rect 6010 10010 6030 10030
rect 6090 10010 6110 10030
rect 6170 10010 6190 10030
rect 4250 9930 4270 9950
rect 4330 9930 4350 9950
rect 4410 9930 4430 9950
rect 4490 9930 4510 9950
rect 4570 9930 4590 9950
rect 4650 9930 4670 9950
rect 4730 9930 4750 9950
rect 4810 9930 4830 9950
rect 4890 9930 4910 9950
rect 4970 9930 4990 9950
rect 5050 9930 5070 9950
rect 5130 9930 5150 9950
rect 5210 9930 5230 9950
rect 5290 9930 5310 9950
rect 5370 9930 5390 9950
rect 5450 9930 5470 9950
rect 5530 9930 5550 9950
rect 5610 9930 5630 9950
rect 5690 9930 5710 9950
rect 5770 9930 5790 9950
rect 5850 9930 5870 9950
rect 5930 9930 5950 9950
rect 6010 9930 6030 9950
rect 6090 9930 6110 9950
rect 6170 9930 6190 9950
rect 4250 9850 4270 9870
rect 4330 9850 4350 9870
rect 4410 9850 4430 9870
rect 4490 9850 4510 9870
rect 4570 9850 4590 9870
rect 4650 9850 4670 9870
rect 4730 9850 4750 9870
rect 4810 9850 4830 9870
rect 4890 9850 4910 9870
rect 4970 9850 4990 9870
rect 5050 9850 5070 9870
rect 5130 9850 5150 9870
rect 5210 9850 5230 9870
rect 5290 9850 5310 9870
rect 5370 9850 5390 9870
rect 5450 9850 5470 9870
rect 5530 9850 5550 9870
rect 5610 9850 5630 9870
rect 5690 9850 5710 9870
rect 5770 9850 5790 9870
rect 5850 9850 5870 9870
rect 5930 9850 5950 9870
rect 6010 9850 6030 9870
rect 6090 9850 6110 9870
rect 6170 9850 6190 9870
rect 4250 9770 4270 9790
rect 4330 9770 4350 9790
rect 4410 9770 4430 9790
rect 4490 9770 4510 9790
rect 4570 9770 4590 9790
rect 4650 9770 4670 9790
rect 4730 9770 4750 9790
rect 4810 9770 4830 9790
rect 4890 9770 4910 9790
rect 4970 9770 4990 9790
rect 5050 9770 5070 9790
rect 5130 9770 5150 9790
rect 5210 9770 5230 9790
rect 5290 9770 5310 9790
rect 5370 9770 5390 9790
rect 5450 9770 5470 9790
rect 5530 9770 5550 9790
rect 5610 9770 5630 9790
rect 5690 9770 5710 9790
rect 5770 9770 5790 9790
rect 5850 9770 5870 9790
rect 5930 9770 5950 9790
rect 6010 9770 6030 9790
rect 6090 9770 6110 9790
rect 6170 9770 6190 9790
rect 4250 9690 4270 9710
rect 4330 9690 4350 9710
rect 4410 9690 4430 9710
rect 4490 9690 4510 9710
rect 4570 9690 4590 9710
rect 4650 9690 4670 9710
rect 4730 9690 4750 9710
rect 4810 9690 4830 9710
rect 4890 9690 4910 9710
rect 4970 9690 4990 9710
rect 5050 9690 5070 9710
rect 5130 9690 5150 9710
rect 5210 9690 5230 9710
rect 5290 9690 5310 9710
rect 5370 9690 5390 9710
rect 5450 9690 5470 9710
rect 5530 9690 5550 9710
rect 5610 9690 5630 9710
rect 5690 9690 5710 9710
rect 5770 9690 5790 9710
rect 5850 9690 5870 9710
rect 5930 9690 5950 9710
rect 6010 9690 6030 9710
rect 6090 9690 6110 9710
rect 6170 9690 6190 9710
rect 4250 9610 4270 9630
rect 4330 9610 4350 9630
rect 4410 9610 4430 9630
rect 4490 9610 4510 9630
rect 4570 9610 4590 9630
rect 4650 9610 4670 9630
rect 4730 9610 4750 9630
rect 4810 9610 4830 9630
rect 4890 9610 4910 9630
rect 4970 9610 4990 9630
rect 5050 9610 5070 9630
rect 5130 9610 5150 9630
rect 5210 9610 5230 9630
rect 5290 9610 5310 9630
rect 5370 9610 5390 9630
rect 5450 9610 5470 9630
rect 5530 9610 5550 9630
rect 5610 9610 5630 9630
rect 5690 9610 5710 9630
rect 5770 9610 5790 9630
rect 5850 9610 5870 9630
rect 5930 9610 5950 9630
rect 6010 9610 6030 9630
rect 6090 9610 6110 9630
rect 6170 9610 6190 9630
rect 4250 9530 4270 9550
rect 4330 9530 4350 9550
rect 4410 9530 4430 9550
rect 4490 9530 4510 9550
rect 4570 9530 4590 9550
rect 4650 9530 4670 9550
rect 4730 9530 4750 9550
rect 4810 9530 4830 9550
rect 4890 9530 4910 9550
rect 4970 9530 4990 9550
rect 5050 9530 5070 9550
rect 5130 9530 5150 9550
rect 5210 9530 5230 9550
rect 5290 9530 5310 9550
rect 5370 9530 5390 9550
rect 5450 9530 5470 9550
rect 5530 9530 5550 9550
rect 5610 9530 5630 9550
rect 5690 9530 5710 9550
rect 5770 9530 5790 9550
rect 5850 9530 5870 9550
rect 5930 9530 5950 9550
rect 6010 9530 6030 9550
rect 6090 9530 6110 9550
rect 6170 9530 6190 9550
rect 4250 9450 4270 9470
rect 4330 9450 4350 9470
rect 4410 9450 4430 9470
rect 4490 9450 4510 9470
rect 4570 9450 4590 9470
rect 4650 9450 4670 9470
rect 4730 9450 4750 9470
rect 4810 9450 4830 9470
rect 4890 9450 4910 9470
rect 4970 9450 4990 9470
rect 5050 9450 5070 9470
rect 5130 9450 5150 9470
rect 5210 9450 5230 9470
rect 5290 9450 5310 9470
rect 5370 9450 5390 9470
rect 5450 9450 5470 9470
rect 5530 9450 5550 9470
rect 5610 9450 5630 9470
rect 5690 9450 5710 9470
rect 5770 9450 5790 9470
rect 5850 9450 5870 9470
rect 5930 9450 5950 9470
rect 6010 9450 6030 9470
rect 6090 9450 6110 9470
rect 6170 9450 6190 9470
rect 4250 9370 4270 9390
rect 4330 9370 4350 9390
rect 4410 9370 4430 9390
rect 4490 9370 4510 9390
rect 4570 9370 4590 9390
rect 4650 9370 4670 9390
rect 4730 9370 4750 9390
rect 4810 9370 4830 9390
rect 4890 9370 4910 9390
rect 4970 9370 4990 9390
rect 5050 9370 5070 9390
rect 5130 9370 5150 9390
rect 5210 9370 5230 9390
rect 5290 9370 5310 9390
rect 5370 9370 5390 9390
rect 5450 9370 5470 9390
rect 5530 9370 5550 9390
rect 5610 9370 5630 9390
rect 5690 9370 5710 9390
rect 5770 9370 5790 9390
rect 5850 9370 5870 9390
rect 5930 9370 5950 9390
rect 6010 9370 6030 9390
rect 6090 9370 6110 9390
rect 6170 9370 6190 9390
rect 4250 9290 4270 9310
rect 4330 9290 4350 9310
rect 4410 9290 4430 9310
rect 4490 9290 4510 9310
rect 4570 9290 4590 9310
rect 4650 9290 4670 9310
rect 4730 9290 4750 9310
rect 4810 9290 4830 9310
rect 4890 9290 4910 9310
rect 4970 9290 4990 9310
rect 5050 9290 5070 9310
rect 5130 9290 5150 9310
rect 5210 9290 5230 9310
rect 5290 9290 5310 9310
rect 5370 9290 5390 9310
rect 5450 9290 5470 9310
rect 5530 9290 5550 9310
rect 5610 9290 5630 9310
rect 5690 9290 5710 9310
rect 5770 9290 5790 9310
rect 5850 9290 5870 9310
rect 5930 9290 5950 9310
rect 6010 9290 6030 9310
rect 6090 9290 6110 9310
rect 6170 9290 6190 9310
rect 4250 9210 4270 9230
rect 4330 9210 4350 9230
rect 4410 9210 4430 9230
rect 4490 9210 4510 9230
rect 4570 9210 4590 9230
rect 4650 9210 4670 9230
rect 4730 9210 4750 9230
rect 4810 9210 4830 9230
rect 4890 9210 4910 9230
rect 4970 9210 4990 9230
rect 5050 9210 5070 9230
rect 5130 9210 5150 9230
rect 5210 9210 5230 9230
rect 5290 9210 5310 9230
rect 5370 9210 5390 9230
rect 5450 9210 5470 9230
rect 5530 9210 5550 9230
rect 5610 9210 5630 9230
rect 5690 9210 5710 9230
rect 5770 9210 5790 9230
rect 5850 9210 5870 9230
rect 5930 9210 5950 9230
rect 6010 9210 6030 9230
rect 6090 9210 6110 9230
rect 6170 9210 6190 9230
rect 4250 9130 4270 9150
rect 4330 9130 4350 9150
rect 4410 9130 4430 9150
rect 4490 9130 4510 9150
rect 4570 9130 4590 9150
rect 4650 9130 4670 9150
rect 4730 9130 4750 9150
rect 4810 9130 4830 9150
rect 4890 9130 4910 9150
rect 4970 9130 4990 9150
rect 5050 9130 5070 9150
rect 5130 9130 5150 9150
rect 5210 9130 5230 9150
rect 5290 9130 5310 9150
rect 5370 9130 5390 9150
rect 5450 9130 5470 9150
rect 5530 9130 5550 9150
rect 5610 9130 5630 9150
rect 5690 9130 5710 9150
rect 5770 9130 5790 9150
rect 5850 9130 5870 9150
rect 5930 9130 5950 9150
rect 6010 9130 6030 9150
rect 6090 9130 6110 9150
rect 6170 9130 6190 9150
rect 4250 9050 4270 9070
rect 4330 9050 4350 9070
rect 4410 9050 4430 9070
rect 4490 9050 4510 9070
rect 4570 9050 4590 9070
rect 4650 9050 4670 9070
rect 4730 9050 4750 9070
rect 4810 9050 4830 9070
rect 4890 9050 4910 9070
rect 4970 9050 4990 9070
rect 5050 9050 5070 9070
rect 5130 9050 5150 9070
rect 5210 9050 5230 9070
rect 5290 9050 5310 9070
rect 5370 9050 5390 9070
rect 5450 9050 5470 9070
rect 5530 9050 5550 9070
rect 5610 9050 5630 9070
rect 5690 9050 5710 9070
rect 5770 9050 5790 9070
rect 5850 9050 5870 9070
rect 5930 9050 5950 9070
rect 6010 9050 6030 9070
rect 6090 9050 6110 9070
rect 6170 9050 6190 9070
rect 4250 8970 4270 8990
rect 4330 8970 4350 8990
rect 4410 8970 4430 8990
rect 4490 8970 4510 8990
rect 4570 8970 4590 8990
rect 4650 8970 4670 8990
rect 4730 8970 4750 8990
rect 4810 8970 4830 8990
rect 4890 8970 4910 8990
rect 4970 8970 4990 8990
rect 5050 8970 5070 8990
rect 5130 8970 5150 8990
rect 5210 8970 5230 8990
rect 5290 8970 5310 8990
rect 5370 8970 5390 8990
rect 5450 8970 5470 8990
rect 5530 8970 5550 8990
rect 5610 8970 5630 8990
rect 5690 8970 5710 8990
rect 5770 8970 5790 8990
rect 5850 8970 5870 8990
rect 5930 8970 5950 8990
rect 6010 8970 6030 8990
rect 6090 8970 6110 8990
rect 6170 8970 6190 8990
rect 4250 8890 4270 8910
rect 4330 8890 4350 8910
rect 4410 8890 4430 8910
rect 4490 8890 4510 8910
rect 4570 8890 4590 8910
rect 4650 8890 4670 8910
rect 4730 8890 4750 8910
rect 4810 8890 4830 8910
rect 4890 8890 4910 8910
rect 4970 8890 4990 8910
rect 5050 8890 5070 8910
rect 5130 8890 5150 8910
rect 5210 8890 5230 8910
rect 5290 8890 5310 8910
rect 5370 8890 5390 8910
rect 5450 8890 5470 8910
rect 5530 8890 5550 8910
rect 5610 8890 5630 8910
rect 5690 8890 5710 8910
rect 5770 8890 5790 8910
rect 5850 8890 5870 8910
rect 5930 8890 5950 8910
rect 6010 8890 6030 8910
rect 6090 8890 6110 8910
rect 6170 8890 6190 8910
rect 4250 8810 4270 8830
rect 4330 8810 4350 8830
rect 4410 8810 4430 8830
rect 4490 8810 4510 8830
rect 4570 8810 4590 8830
rect 4650 8810 4670 8830
rect 4730 8810 4750 8830
rect 4810 8810 4830 8830
rect 4890 8810 4910 8830
rect 4970 8810 4990 8830
rect 5050 8810 5070 8830
rect 5130 8810 5150 8830
rect 5210 8810 5230 8830
rect 5290 8810 5310 8830
rect 5370 8810 5390 8830
rect 5450 8810 5470 8830
rect 5530 8810 5550 8830
rect 5610 8810 5630 8830
rect 5690 8810 5710 8830
rect 5770 8810 5790 8830
rect 5850 8810 5870 8830
rect 5930 8810 5950 8830
rect 6010 8810 6030 8830
rect 6090 8810 6110 8830
rect 6170 8810 6190 8830
rect 4250 8730 4270 8750
rect 4330 8730 4350 8750
rect 4410 8730 4430 8750
rect 4490 8730 4510 8750
rect 4570 8730 4590 8750
rect 4650 8730 4670 8750
rect 4730 8730 4750 8750
rect 4810 8730 4830 8750
rect 4890 8730 4910 8750
rect 4970 8730 4990 8750
rect 5050 8730 5070 8750
rect 5130 8730 5150 8750
rect 5210 8730 5230 8750
rect 5290 8730 5310 8750
rect 5370 8730 5390 8750
rect 5450 8730 5470 8750
rect 5530 8730 5550 8750
rect 5610 8730 5630 8750
rect 5690 8730 5710 8750
rect 5770 8730 5790 8750
rect 5850 8730 5870 8750
rect 5930 8730 5950 8750
rect 6010 8730 6030 8750
rect 6090 8730 6110 8750
rect 6170 8730 6190 8750
rect 4250 8650 4270 8670
rect 4330 8650 4350 8670
rect 4410 8650 4430 8670
rect 4490 8650 4510 8670
rect 4570 8650 4590 8670
rect 4650 8650 4670 8670
rect 4730 8650 4750 8670
rect 4810 8650 4830 8670
rect 4890 8650 4910 8670
rect 4970 8650 4990 8670
rect 5050 8650 5070 8670
rect 5130 8650 5150 8670
rect 5210 8650 5230 8670
rect 5290 8650 5310 8670
rect 5370 8650 5390 8670
rect 5450 8650 5470 8670
rect 5530 8650 5550 8670
rect 5610 8650 5630 8670
rect 5690 8650 5710 8670
rect 5770 8650 5790 8670
rect 5850 8650 5870 8670
rect 5930 8650 5950 8670
rect 6010 8650 6030 8670
rect 6090 8650 6110 8670
rect 6170 8650 6190 8670
rect 4250 8570 4270 8590
rect 4330 8570 4350 8590
rect 4410 8570 4430 8590
rect 4490 8570 4510 8590
rect 4570 8570 4590 8590
rect 4650 8570 4670 8590
rect 4730 8570 4750 8590
rect 4810 8570 4830 8590
rect 4890 8570 4910 8590
rect 4970 8570 4990 8590
rect 5050 8570 5070 8590
rect 5130 8570 5150 8590
rect 5210 8570 5230 8590
rect 5290 8570 5310 8590
rect 5370 8570 5390 8590
rect 5450 8570 5470 8590
rect 5530 8570 5550 8590
rect 5610 8570 5630 8590
rect 5690 8570 5710 8590
rect 5770 8570 5790 8590
rect 5850 8570 5870 8590
rect 5930 8570 5950 8590
rect 6010 8570 6030 8590
rect 6090 8570 6110 8590
rect 6170 8570 6190 8590
rect 4250 8490 4270 8510
rect 4330 8490 4350 8510
rect 4410 8490 4430 8510
rect 4490 8490 4510 8510
rect 4570 8490 4590 8510
rect 4650 8490 4670 8510
rect 4730 8490 4750 8510
rect 4810 8490 4830 8510
rect 4890 8490 4910 8510
rect 4970 8490 4990 8510
rect 5050 8490 5070 8510
rect 5130 8490 5150 8510
rect 5210 8490 5230 8510
rect 5290 8490 5310 8510
rect 5370 8490 5390 8510
rect 5450 8490 5470 8510
rect 5530 8490 5550 8510
rect 5610 8490 5630 8510
rect 5690 8490 5710 8510
rect 5770 8490 5790 8510
rect 5850 8490 5870 8510
rect 5930 8490 5950 8510
rect 6010 8490 6030 8510
rect 6090 8490 6110 8510
rect 6170 8490 6190 8510
rect 4250 8410 4270 8430
rect 4330 8410 4350 8430
rect 4410 8410 4430 8430
rect 4490 8410 4510 8430
rect 4570 8410 4590 8430
rect 4650 8410 4670 8430
rect 4730 8410 4750 8430
rect 4810 8410 4830 8430
rect 4890 8410 4910 8430
rect 4970 8410 4990 8430
rect 5050 8410 5070 8430
rect 5130 8410 5150 8430
rect 5210 8410 5230 8430
rect 5290 8410 5310 8430
rect 5370 8410 5390 8430
rect 5450 8410 5470 8430
rect 5530 8410 5550 8430
rect 5610 8410 5630 8430
rect 5690 8410 5710 8430
rect 5770 8410 5790 8430
rect 5850 8410 5870 8430
rect 5930 8410 5950 8430
rect 6010 8410 6030 8430
rect 6090 8410 6110 8430
rect 6170 8410 6190 8430
rect 4250 8330 4270 8350
rect 4330 8330 4350 8350
rect 4410 8330 4430 8350
rect 4490 8330 4510 8350
rect 4570 8330 4590 8350
rect 4650 8330 4670 8350
rect 4730 8330 4750 8350
rect 4810 8330 4830 8350
rect 4890 8330 4910 8350
rect 4970 8330 4990 8350
rect 5050 8330 5070 8350
rect 5130 8330 5150 8350
rect 5210 8330 5230 8350
rect 5290 8330 5310 8350
rect 5370 8330 5390 8350
rect 5450 8330 5470 8350
rect 5530 8330 5550 8350
rect 5610 8330 5630 8350
rect 5690 8330 5710 8350
rect 5770 8330 5790 8350
rect 5850 8330 5870 8350
rect 5930 8330 5950 8350
rect 6010 8330 6030 8350
rect 6090 8330 6110 8350
rect 6170 8330 6190 8350
rect 4250 8250 4270 8270
rect 4330 8250 4350 8270
rect 4410 8250 4430 8270
rect 4490 8250 4510 8270
rect 4570 8250 4590 8270
rect 4650 8250 4670 8270
rect 4730 8250 4750 8270
rect 4810 8250 4830 8270
rect 4890 8250 4910 8270
rect 4970 8250 4990 8270
rect 5050 8250 5070 8270
rect 5130 8250 5150 8270
rect 5210 8250 5230 8270
rect 5290 8250 5310 8270
rect 5370 8250 5390 8270
rect 5450 8250 5470 8270
rect 5530 8250 5550 8270
rect 5610 8250 5630 8270
rect 5690 8250 5710 8270
rect 5770 8250 5790 8270
rect 5850 8250 5870 8270
rect 5930 8250 5950 8270
rect 6010 8250 6030 8270
rect 6090 8250 6110 8270
rect 6170 8250 6190 8270
rect 4250 8170 4270 8190
rect 4330 8170 4350 8190
rect 4410 8170 4430 8190
rect 4490 8170 4510 8190
rect 4570 8170 4590 8190
rect 4650 8170 4670 8190
rect 4730 8170 4750 8190
rect 4810 8170 4830 8190
rect 4890 8170 4910 8190
rect 4970 8170 4990 8190
rect 5050 8170 5070 8190
rect 5130 8170 5150 8190
rect 5210 8170 5230 8190
rect 5290 8170 5310 8190
rect 5370 8170 5390 8190
rect 5450 8170 5470 8190
rect 5530 8170 5550 8190
rect 5610 8170 5630 8190
rect 5690 8170 5710 8190
rect 5770 8170 5790 8190
rect 5850 8170 5870 8190
rect 5930 8170 5950 8190
rect 6010 8170 6030 8190
rect 6090 8170 6110 8190
rect 6170 8170 6190 8190
rect 4250 8090 4270 8110
rect 4330 8090 4350 8110
rect 4410 8090 4430 8110
rect 4490 8090 4510 8110
rect 4570 8090 4590 8110
rect 4650 8090 4670 8110
rect 4730 8090 4750 8110
rect 4810 8090 4830 8110
rect 4890 8090 4910 8110
rect 4970 8090 4990 8110
rect 5050 8090 5070 8110
rect 5130 8090 5150 8110
rect 5210 8090 5230 8110
rect 5290 8090 5310 8110
rect 5370 8090 5390 8110
rect 5450 8090 5470 8110
rect 5530 8090 5550 8110
rect 5610 8090 5630 8110
rect 5690 8090 5710 8110
rect 5770 8090 5790 8110
rect 5850 8090 5870 8110
rect 5930 8090 5950 8110
rect 6010 8090 6030 8110
rect 6090 8090 6110 8110
rect 6170 8090 6190 8110
rect 4250 8010 4270 8030
rect 4330 8010 4350 8030
rect 4410 8010 4430 8030
rect 4490 8010 4510 8030
rect 4570 8010 4590 8030
rect 4650 8010 4670 8030
rect 4730 8010 4750 8030
rect 4810 8010 4830 8030
rect 4890 8010 4910 8030
rect 4970 8010 4990 8030
rect 5050 8010 5070 8030
rect 5130 8010 5150 8030
rect 5210 8010 5230 8030
rect 5290 8010 5310 8030
rect 5370 8010 5390 8030
rect 5450 8010 5470 8030
rect 5530 8010 5550 8030
rect 5610 8010 5630 8030
rect 5690 8010 5710 8030
rect 5770 8010 5790 8030
rect 5850 8010 5870 8030
rect 5930 8010 5950 8030
rect 6010 8010 6030 8030
rect 6090 8010 6110 8030
rect 6170 8010 6190 8030
rect 4250 7930 4270 7950
rect 4330 7930 4350 7950
rect 4410 7930 4430 7950
rect 4490 7930 4510 7950
rect 4570 7930 4590 7950
rect 4650 7930 4670 7950
rect 4730 7930 4750 7950
rect 4810 7930 4830 7950
rect 4890 7930 4910 7950
rect 4970 7930 4990 7950
rect 5050 7930 5070 7950
rect 5130 7930 5150 7950
rect 5210 7930 5230 7950
rect 5290 7930 5310 7950
rect 5370 7930 5390 7950
rect 5450 7930 5470 7950
rect 5530 7930 5550 7950
rect 5610 7930 5630 7950
rect 5690 7930 5710 7950
rect 5770 7930 5790 7950
rect 5850 7930 5870 7950
rect 5930 7930 5950 7950
rect 6010 7930 6030 7950
rect 6090 7930 6110 7950
rect 6170 7930 6190 7950
rect 4250 7850 4270 7870
rect 4330 7850 4350 7870
rect 4410 7850 4430 7870
rect 4490 7850 4510 7870
rect 4570 7850 4590 7870
rect 4650 7850 4670 7870
rect 4730 7850 4750 7870
rect 4810 7850 4830 7870
rect 4890 7850 4910 7870
rect 4970 7850 4990 7870
rect 5050 7850 5070 7870
rect 5130 7850 5150 7870
rect 5210 7850 5230 7870
rect 5290 7850 5310 7870
rect 5370 7850 5390 7870
rect 5450 7850 5470 7870
rect 5530 7850 5550 7870
rect 5610 7850 5630 7870
rect 5690 7850 5710 7870
rect 5770 7850 5790 7870
rect 5850 7850 5870 7870
rect 5930 7850 5950 7870
rect 6010 7850 6030 7870
rect 6090 7850 6110 7870
rect 6170 7850 6190 7870
rect 4250 7770 4270 7790
rect 4330 7770 4350 7790
rect 4410 7770 4430 7790
rect 4490 7770 4510 7790
rect 4570 7770 4590 7790
rect 4650 7770 4670 7790
rect 4730 7770 4750 7790
rect 4810 7770 4830 7790
rect 4890 7770 4910 7790
rect 4970 7770 4990 7790
rect 5050 7770 5070 7790
rect 5130 7770 5150 7790
rect 5210 7770 5230 7790
rect 5290 7770 5310 7790
rect 5370 7770 5390 7790
rect 5450 7770 5470 7790
rect 5530 7770 5550 7790
rect 5610 7770 5630 7790
rect 5690 7770 5710 7790
rect 5770 7770 5790 7790
rect 5850 7770 5870 7790
rect 5930 7770 5950 7790
rect 6010 7770 6030 7790
rect 6090 7770 6110 7790
rect 6170 7770 6190 7790
rect 4250 7690 4270 7710
rect 4330 7690 4350 7710
rect 4410 7690 4430 7710
rect 4490 7690 4510 7710
rect 4570 7690 4590 7710
rect 4650 7690 4670 7710
rect 4730 7690 4750 7710
rect 4810 7690 4830 7710
rect 4890 7690 4910 7710
rect 4970 7690 4990 7710
rect 5050 7690 5070 7710
rect 5130 7690 5150 7710
rect 5210 7690 5230 7710
rect 5290 7690 5310 7710
rect 5370 7690 5390 7710
rect 5450 7690 5470 7710
rect 5530 7690 5550 7710
rect 5610 7690 5630 7710
rect 5690 7690 5710 7710
rect 5770 7690 5790 7710
rect 5850 7690 5870 7710
rect 5930 7690 5950 7710
rect 6010 7690 6030 7710
rect 6090 7690 6110 7710
rect 6170 7690 6190 7710
rect 4250 7610 4270 7630
rect 4330 7610 4350 7630
rect 4410 7610 4430 7630
rect 4490 7610 4510 7630
rect 4570 7610 4590 7630
rect 4650 7610 4670 7630
rect 4730 7610 4750 7630
rect 4810 7610 4830 7630
rect 4890 7610 4910 7630
rect 4970 7610 4990 7630
rect 5050 7610 5070 7630
rect 5130 7610 5150 7630
rect 5210 7610 5230 7630
rect 5290 7610 5310 7630
rect 5370 7610 5390 7630
rect 5450 7610 5470 7630
rect 5530 7610 5550 7630
rect 5610 7610 5630 7630
rect 5690 7610 5710 7630
rect 5770 7610 5790 7630
rect 5850 7610 5870 7630
rect 5930 7610 5950 7630
rect 6010 7610 6030 7630
rect 6090 7610 6110 7630
rect 6170 7610 6190 7630
rect 4250 7530 4270 7550
rect 4330 7530 4350 7550
rect 4410 7530 4430 7550
rect 4490 7530 4510 7550
rect 4570 7530 4590 7550
rect 4650 7530 4670 7550
rect 4730 7530 4750 7550
rect 4810 7530 4830 7550
rect 4890 7530 4910 7550
rect 4970 7530 4990 7550
rect 5050 7530 5070 7550
rect 5130 7530 5150 7550
rect 5210 7530 5230 7550
rect 5290 7530 5310 7550
rect 5370 7530 5390 7550
rect 5450 7530 5470 7550
rect 5530 7530 5550 7550
rect 5610 7530 5630 7550
rect 5690 7530 5710 7550
rect 5770 7530 5790 7550
rect 5850 7530 5870 7550
rect 5930 7530 5950 7550
rect 6010 7530 6030 7550
rect 6090 7530 6110 7550
rect 6170 7530 6190 7550
rect 4250 7450 4270 7470
rect 4330 7450 4350 7470
rect 4410 7450 4430 7470
rect 4490 7450 4510 7470
rect 4570 7450 4590 7470
rect 4650 7450 4670 7470
rect 4730 7450 4750 7470
rect 4810 7450 4830 7470
rect 4890 7450 4910 7470
rect 4970 7450 4990 7470
rect 5050 7450 5070 7470
rect 5130 7450 5150 7470
rect 5210 7450 5230 7470
rect 5290 7450 5310 7470
rect 5370 7450 5390 7470
rect 5450 7450 5470 7470
rect 5530 7450 5550 7470
rect 5610 7450 5630 7470
rect 5690 7450 5710 7470
rect 5770 7450 5790 7470
rect 5850 7450 5870 7470
rect 5930 7450 5950 7470
rect 6010 7450 6030 7470
rect 6090 7450 6110 7470
rect 6170 7450 6190 7470
rect 4250 7370 4270 7390
rect 4330 7370 4350 7390
rect 4410 7370 4430 7390
rect 4490 7370 4510 7390
rect 4570 7370 4590 7390
rect 4650 7370 4670 7390
rect 4730 7370 4750 7390
rect 4810 7370 4830 7390
rect 4890 7370 4910 7390
rect 4970 7370 4990 7390
rect 5050 7370 5070 7390
rect 5130 7370 5150 7390
rect 5210 7370 5230 7390
rect 5290 7370 5310 7390
rect 5370 7370 5390 7390
rect 5450 7370 5470 7390
rect 5530 7370 5550 7390
rect 5610 7370 5630 7390
rect 5690 7370 5710 7390
rect 5770 7370 5790 7390
rect 5850 7370 5870 7390
rect 5930 7370 5950 7390
rect 6010 7370 6030 7390
rect 6090 7370 6110 7390
rect 6170 7370 6190 7390
rect 4250 7290 4270 7310
rect 4330 7290 4350 7310
rect 4410 7290 4430 7310
rect 4490 7290 4510 7310
rect 4570 7290 4590 7310
rect 4650 7290 4670 7310
rect 4730 7290 4750 7310
rect 4810 7290 4830 7310
rect 4890 7290 4910 7310
rect 4970 7290 4990 7310
rect 5050 7290 5070 7310
rect 5130 7290 5150 7310
rect 5210 7290 5230 7310
rect 5290 7290 5310 7310
rect 5370 7290 5390 7310
rect 5450 7290 5470 7310
rect 5530 7290 5550 7310
rect 5610 7290 5630 7310
rect 5690 7290 5710 7310
rect 5770 7290 5790 7310
rect 5850 7290 5870 7310
rect 5930 7290 5950 7310
rect 6010 7290 6030 7310
rect 6090 7290 6110 7310
rect 6170 7290 6190 7310
rect 4250 7210 4270 7230
rect 4330 7210 4350 7230
rect 4410 7210 4430 7230
rect 4490 7210 4510 7230
rect 4570 7210 4590 7230
rect 4650 7210 4670 7230
rect 4730 7210 4750 7230
rect 4810 7210 4830 7230
rect 4890 7210 4910 7230
rect 4970 7210 4990 7230
rect 5050 7210 5070 7230
rect 5130 7210 5150 7230
rect 5210 7210 5230 7230
rect 5290 7210 5310 7230
rect 5370 7210 5390 7230
rect 5450 7210 5470 7230
rect 5530 7210 5550 7230
rect 5610 7210 5630 7230
rect 5690 7210 5710 7230
rect 5770 7210 5790 7230
rect 5850 7210 5870 7230
rect 5930 7210 5950 7230
rect 6010 7210 6030 7230
rect 6090 7210 6110 7230
rect 6170 7210 6190 7230
rect 4250 7130 4270 7150
rect 4330 7130 4350 7150
rect 4410 7130 4430 7150
rect 4490 7130 4510 7150
rect 4570 7130 4590 7150
rect 4650 7130 4670 7150
rect 4730 7130 4750 7150
rect 4810 7130 4830 7150
rect 4890 7130 4910 7150
rect 4970 7130 4990 7150
rect 5050 7130 5070 7150
rect 5130 7130 5150 7150
rect 5210 7130 5230 7150
rect 5290 7130 5310 7150
rect 5370 7130 5390 7150
rect 5450 7130 5470 7150
rect 5530 7130 5550 7150
rect 5610 7130 5630 7150
rect 5690 7130 5710 7150
rect 5770 7130 5790 7150
rect 5850 7130 5870 7150
rect 5930 7130 5950 7150
rect 6010 7130 6030 7150
rect 6090 7130 6110 7150
rect 6170 7130 6190 7150
rect 4250 7050 4270 7070
rect 4330 7050 4350 7070
rect 4410 7050 4430 7070
rect 4490 7050 4510 7070
rect 4570 7050 4590 7070
rect 4650 7050 4670 7070
rect 4730 7050 4750 7070
rect 4810 7050 4830 7070
rect 4890 7050 4910 7070
rect 4970 7050 4990 7070
rect 5050 7050 5070 7070
rect 5130 7050 5150 7070
rect 5210 7050 5230 7070
rect 5290 7050 5310 7070
rect 5370 7050 5390 7070
rect 5450 7050 5470 7070
rect 5530 7050 5550 7070
rect 5610 7050 5630 7070
rect 5690 7050 5710 7070
rect 5770 7050 5790 7070
rect 5850 7050 5870 7070
rect 5930 7050 5950 7070
rect 6010 7050 6030 7070
rect 6090 7050 6110 7070
rect 6170 7050 6190 7070
rect 4250 6970 4270 6990
rect 4330 6970 4350 6990
rect 4410 6970 4430 6990
rect 4490 6970 4510 6990
rect 4570 6970 4590 6990
rect 4650 6970 4670 6990
rect 4730 6970 4750 6990
rect 4810 6970 4830 6990
rect 4890 6970 4910 6990
rect 4970 6970 4990 6990
rect 5050 6970 5070 6990
rect 5130 6970 5150 6990
rect 5210 6970 5230 6990
rect 5290 6970 5310 6990
rect 5370 6970 5390 6990
rect 5450 6970 5470 6990
rect 5530 6970 5550 6990
rect 5610 6970 5630 6990
rect 5690 6970 5710 6990
rect 5770 6970 5790 6990
rect 5850 6970 5870 6990
rect 5930 6970 5950 6990
rect 6010 6970 6030 6990
rect 6090 6970 6110 6990
rect 6170 6970 6190 6990
rect 4250 6890 4270 6910
rect 4330 6890 4350 6910
rect 4410 6890 4430 6910
rect 4490 6890 4510 6910
rect 4570 6890 4590 6910
rect 4650 6890 4670 6910
rect 4730 6890 4750 6910
rect 4810 6890 4830 6910
rect 4890 6890 4910 6910
rect 4970 6890 4990 6910
rect 5050 6890 5070 6910
rect 5130 6890 5150 6910
rect 5210 6890 5230 6910
rect 5290 6890 5310 6910
rect 5370 6890 5390 6910
rect 5450 6890 5470 6910
rect 5530 6890 5550 6910
rect 5610 6890 5630 6910
rect 5690 6890 5710 6910
rect 5770 6890 5790 6910
rect 5850 6890 5870 6910
rect 5930 6890 5950 6910
rect 6010 6890 6030 6910
rect 6090 6890 6110 6910
rect 6170 6890 6190 6910
rect 4250 6810 4270 6830
rect 4330 6810 4350 6830
rect 4410 6810 4430 6830
rect 4490 6810 4510 6830
rect 4570 6810 4590 6830
rect 4650 6810 4670 6830
rect 4730 6810 4750 6830
rect 4810 6810 4830 6830
rect 4890 6810 4910 6830
rect 4970 6810 4990 6830
rect 5050 6810 5070 6830
rect 5130 6810 5150 6830
rect 5210 6810 5230 6830
rect 5290 6810 5310 6830
rect 5370 6810 5390 6830
rect 5450 6810 5470 6830
rect 5530 6810 5550 6830
rect 5610 6810 5630 6830
rect 5690 6810 5710 6830
rect 5770 6810 5790 6830
rect 5850 6810 5870 6830
rect 5930 6810 5950 6830
rect 6010 6810 6030 6830
rect 6090 6810 6110 6830
rect 6170 6810 6190 6830
rect 4250 6730 4270 6750
rect 4330 6730 4350 6750
rect 4410 6730 4430 6750
rect 4490 6730 4510 6750
rect 4570 6730 4590 6750
rect 4650 6730 4670 6750
rect 4730 6730 4750 6750
rect 4810 6730 4830 6750
rect 4890 6730 4910 6750
rect 4970 6730 4990 6750
rect 5050 6730 5070 6750
rect 5130 6730 5150 6750
rect 5210 6730 5230 6750
rect 5290 6730 5310 6750
rect 5370 6730 5390 6750
rect 5450 6730 5470 6750
rect 5530 6730 5550 6750
rect 5610 6730 5630 6750
rect 5690 6730 5710 6750
rect 5770 6730 5790 6750
rect 5850 6730 5870 6750
rect 5930 6730 5950 6750
rect 6010 6730 6030 6750
rect 6090 6730 6110 6750
rect 6170 6730 6190 6750
rect 4250 6650 4270 6670
rect 4330 6650 4350 6670
rect 4410 6650 4430 6670
rect 4490 6650 4510 6670
rect 4570 6650 4590 6670
rect 4650 6650 4670 6670
rect 4730 6650 4750 6670
rect 4810 6650 4830 6670
rect 4890 6650 4910 6670
rect 4970 6650 4990 6670
rect 5050 6650 5070 6670
rect 5130 6650 5150 6670
rect 5210 6650 5230 6670
rect 5290 6650 5310 6670
rect 5370 6650 5390 6670
rect 5450 6650 5470 6670
rect 5530 6650 5550 6670
rect 5610 6650 5630 6670
rect 5690 6650 5710 6670
rect 5770 6650 5790 6670
rect 5850 6650 5870 6670
rect 5930 6650 5950 6670
rect 6010 6650 6030 6670
rect 6090 6650 6110 6670
rect 6170 6650 6190 6670
rect 4250 6570 4270 6590
rect 4330 6570 4350 6590
rect 4410 6570 4430 6590
rect 4490 6570 4510 6590
rect 4570 6570 4590 6590
rect 4650 6570 4670 6590
rect 4730 6570 4750 6590
rect 4810 6570 4830 6590
rect 4890 6570 4910 6590
rect 4970 6570 4990 6590
rect 5050 6570 5070 6590
rect 5130 6570 5150 6590
rect 5210 6570 5230 6590
rect 5290 6570 5310 6590
rect 5370 6570 5390 6590
rect 5450 6570 5470 6590
rect 5530 6570 5550 6590
rect 5610 6570 5630 6590
rect 5690 6570 5710 6590
rect 5770 6570 5790 6590
rect 5850 6570 5870 6590
rect 5930 6570 5950 6590
rect 6010 6570 6030 6590
rect 6090 6570 6110 6590
rect 6170 6570 6190 6590
rect 4250 6490 4270 6510
rect 4330 6490 4350 6510
rect 4410 6490 4430 6510
rect 4490 6490 4510 6510
rect 4570 6490 4590 6510
rect 4650 6490 4670 6510
rect 4730 6490 4750 6510
rect 4810 6490 4830 6510
rect 4890 6490 4910 6510
rect 4970 6490 4990 6510
rect 5050 6490 5070 6510
rect 5130 6490 5150 6510
rect 5210 6490 5230 6510
rect 5290 6490 5310 6510
rect 5370 6490 5390 6510
rect 5450 6490 5470 6510
rect 5530 6490 5550 6510
rect 5610 6490 5630 6510
rect 5690 6490 5710 6510
rect 5770 6490 5790 6510
rect 5850 6490 5870 6510
rect 5930 6490 5950 6510
rect 6010 6490 6030 6510
rect 6090 6490 6110 6510
rect 6170 6490 6190 6510
rect 4250 6410 4270 6430
rect 4330 6410 4350 6430
rect 4410 6410 4430 6430
rect 4490 6410 4510 6430
rect 4570 6410 4590 6430
rect 4650 6410 4670 6430
rect 4730 6410 4750 6430
rect 4810 6410 4830 6430
rect 4890 6410 4910 6430
rect 4970 6410 4990 6430
rect 5050 6410 5070 6430
rect 5130 6410 5150 6430
rect 5210 6410 5230 6430
rect 5290 6410 5310 6430
rect 5370 6410 5390 6430
rect 5450 6410 5470 6430
rect 5530 6410 5550 6430
rect 5610 6410 5630 6430
rect 5690 6410 5710 6430
rect 5770 6410 5790 6430
rect 5850 6410 5870 6430
rect 5930 6410 5950 6430
rect 6010 6410 6030 6430
rect 6090 6410 6110 6430
rect 6170 6410 6190 6430
rect 4250 6330 4270 6350
rect 4330 6330 4350 6350
rect 4410 6330 4430 6350
rect 4490 6330 4510 6350
rect 4570 6330 4590 6350
rect 4650 6330 4670 6350
rect 4730 6330 4750 6350
rect 4810 6330 4830 6350
rect 4890 6330 4910 6350
rect 4970 6330 4990 6350
rect 5050 6330 5070 6350
rect 5130 6330 5150 6350
rect 5210 6330 5230 6350
rect 5290 6330 5310 6350
rect 5370 6330 5390 6350
rect 5450 6330 5470 6350
rect 5530 6330 5550 6350
rect 5610 6330 5630 6350
rect 5690 6330 5710 6350
rect 5770 6330 5790 6350
rect 5850 6330 5870 6350
rect 5930 6330 5950 6350
rect 6010 6330 6030 6350
rect 6090 6330 6110 6350
rect 6170 6330 6190 6350
rect 4250 6250 4270 6270
rect 4330 6250 4350 6270
rect 4410 6250 4430 6270
rect 4490 6250 4510 6270
rect 4570 6250 4590 6270
rect 4650 6250 4670 6270
rect 4730 6250 4750 6270
rect 4810 6250 4830 6270
rect 4890 6250 4910 6270
rect 4970 6250 4990 6270
rect 5050 6250 5070 6270
rect 5130 6250 5150 6270
rect 5210 6250 5230 6270
rect 5290 6250 5310 6270
rect 5370 6250 5390 6270
rect 5450 6250 5470 6270
rect 5530 6250 5550 6270
rect 5610 6250 5630 6270
rect 5690 6250 5710 6270
rect 5770 6250 5790 6270
rect 5850 6250 5870 6270
rect 5930 6250 5950 6270
rect 6010 6250 6030 6270
rect 6090 6250 6110 6270
rect 6170 6250 6190 6270
rect 4250 6170 4270 6190
rect 4330 6170 4350 6190
rect 4410 6170 4430 6190
rect 4490 6170 4510 6190
rect 4570 6170 4590 6190
rect 4650 6170 4670 6190
rect 4730 6170 4750 6190
rect 4810 6170 4830 6190
rect 4890 6170 4910 6190
rect 4970 6170 4990 6190
rect 5050 6170 5070 6190
rect 5130 6170 5150 6190
rect 5210 6170 5230 6190
rect 5290 6170 5310 6190
rect 5370 6170 5390 6190
rect 5450 6170 5470 6190
rect 5530 6170 5550 6190
rect 5610 6170 5630 6190
rect 5690 6170 5710 6190
rect 5770 6170 5790 6190
rect 5850 6170 5870 6190
rect 5930 6170 5950 6190
rect 6010 6170 6030 6190
rect 6090 6170 6110 6190
rect 6170 6170 6190 6190
rect 4250 6090 4270 6110
rect 4330 6090 4350 6110
rect 4410 6090 4430 6110
rect 4490 6090 4510 6110
rect 4570 6090 4590 6110
rect 4650 6090 4670 6110
rect 4730 6090 4750 6110
rect 4810 6090 4830 6110
rect 4890 6090 4910 6110
rect 4970 6090 4990 6110
rect 5050 6090 5070 6110
rect 5130 6090 5150 6110
rect 5210 6090 5230 6110
rect 5290 6090 5310 6110
rect 5370 6090 5390 6110
rect 5450 6090 5470 6110
rect 5530 6090 5550 6110
rect 5610 6090 5630 6110
rect 5690 6090 5710 6110
rect 5770 6090 5790 6110
rect 5850 6090 5870 6110
rect 5930 6090 5950 6110
rect 6010 6090 6030 6110
rect 6090 6090 6110 6110
rect 6170 6090 6190 6110
rect 4250 6010 4270 6030
rect 4330 6010 4350 6030
rect 4410 6010 4430 6030
rect 4490 6010 4510 6030
rect 4570 6010 4590 6030
rect 4650 6010 4670 6030
rect 4730 6010 4750 6030
rect 4810 6010 4830 6030
rect 4890 6010 4910 6030
rect 4970 6010 4990 6030
rect 5050 6010 5070 6030
rect 5130 6010 5150 6030
rect 5210 6010 5230 6030
rect 5290 6010 5310 6030
rect 5370 6010 5390 6030
rect 5450 6010 5470 6030
rect 5530 6010 5550 6030
rect 5610 6010 5630 6030
rect 5690 6010 5710 6030
rect 5770 6010 5790 6030
rect 5850 6010 5870 6030
rect 5930 6010 5950 6030
rect 6010 6010 6030 6030
rect 6090 6010 6110 6030
rect 6170 6010 6190 6030
rect 4250 5930 4270 5950
rect 4330 5930 4350 5950
rect 4410 5930 4430 5950
rect 4490 5930 4510 5950
rect 4570 5930 4590 5950
rect 4650 5930 4670 5950
rect 4730 5930 4750 5950
rect 4810 5930 4830 5950
rect 4890 5930 4910 5950
rect 4970 5930 4990 5950
rect 5050 5930 5070 5950
rect 5130 5930 5150 5950
rect 5210 5930 5230 5950
rect 5290 5930 5310 5950
rect 5370 5930 5390 5950
rect 5450 5930 5470 5950
rect 5530 5930 5550 5950
rect 5610 5930 5630 5950
rect 5690 5930 5710 5950
rect 5770 5930 5790 5950
rect 5850 5930 5870 5950
rect 5930 5930 5950 5950
rect 6010 5930 6030 5950
rect 6090 5930 6110 5950
rect 6170 5930 6190 5950
rect 4250 5850 4270 5870
rect 4330 5850 4350 5870
rect 4410 5850 4430 5870
rect 4490 5850 4510 5870
rect 4570 5850 4590 5870
rect 4650 5850 4670 5870
rect 4730 5850 4750 5870
rect 4810 5850 4830 5870
rect 4890 5850 4910 5870
rect 4970 5850 4990 5870
rect 5050 5850 5070 5870
rect 5130 5850 5150 5870
rect 5210 5850 5230 5870
rect 5290 5850 5310 5870
rect 5370 5850 5390 5870
rect 5450 5850 5470 5870
rect 5530 5850 5550 5870
rect 5610 5850 5630 5870
rect 5690 5850 5710 5870
rect 5770 5850 5790 5870
rect 5850 5850 5870 5870
rect 5930 5850 5950 5870
rect 6010 5850 6030 5870
rect 6090 5850 6110 5870
rect 6170 5850 6190 5870
rect 4250 5770 4270 5790
rect 4330 5770 4350 5790
rect 4410 5770 4430 5790
rect 4490 5770 4510 5790
rect 4570 5770 4590 5790
rect 4650 5770 4670 5790
rect 4730 5770 4750 5790
rect 4810 5770 4830 5790
rect 4890 5770 4910 5790
rect 4970 5770 4990 5790
rect 5050 5770 5070 5790
rect 5130 5770 5150 5790
rect 5210 5770 5230 5790
rect 5290 5770 5310 5790
rect 5370 5770 5390 5790
rect 5450 5770 5470 5790
rect 5530 5770 5550 5790
rect 5610 5770 5630 5790
rect 5690 5770 5710 5790
rect 5770 5770 5790 5790
rect 5850 5770 5870 5790
rect 5930 5770 5950 5790
rect 6010 5770 6030 5790
rect 6090 5770 6110 5790
rect 6170 5770 6190 5790
rect 4250 5690 4270 5710
rect 4330 5690 4350 5710
rect 4410 5690 4430 5710
rect 4490 5690 4510 5710
rect 4570 5690 4590 5710
rect 4650 5690 4670 5710
rect 4730 5690 4750 5710
rect 4810 5690 4830 5710
rect 4890 5690 4910 5710
rect 4970 5690 4990 5710
rect 5050 5690 5070 5710
rect 5130 5690 5150 5710
rect 5210 5690 5230 5710
rect 5290 5690 5310 5710
rect 5370 5690 5390 5710
rect 5450 5690 5470 5710
rect 5530 5690 5550 5710
rect 5610 5690 5630 5710
rect 5690 5690 5710 5710
rect 5770 5690 5790 5710
rect 5850 5690 5870 5710
rect 5930 5690 5950 5710
rect 6010 5690 6030 5710
rect 6090 5690 6110 5710
rect 6170 5690 6190 5710
rect 4250 5610 4270 5630
rect 4330 5610 4350 5630
rect 4410 5610 4430 5630
rect 4490 5610 4510 5630
rect 4570 5610 4590 5630
rect 4650 5610 4670 5630
rect 4730 5610 4750 5630
rect 4810 5610 4830 5630
rect 4890 5610 4910 5630
rect 4970 5610 4990 5630
rect 5050 5610 5070 5630
rect 5130 5610 5150 5630
rect 5210 5610 5230 5630
rect 5290 5610 5310 5630
rect 5370 5610 5390 5630
rect 5450 5610 5470 5630
rect 5530 5610 5550 5630
rect 5610 5610 5630 5630
rect 5690 5610 5710 5630
rect 5770 5610 5790 5630
rect 5850 5610 5870 5630
rect 5930 5610 5950 5630
rect 6010 5610 6030 5630
rect 6090 5610 6110 5630
rect 6170 5610 6190 5630
rect 4250 5530 4270 5550
rect 4330 5530 4350 5550
rect 4410 5530 4430 5550
rect 4490 5530 4510 5550
rect 4570 5530 4590 5550
rect 4650 5530 4670 5550
rect 4730 5530 4750 5550
rect 4810 5530 4830 5550
rect 4890 5530 4910 5550
rect 4970 5530 4990 5550
rect 5050 5530 5070 5550
rect 5130 5530 5150 5550
rect 5210 5530 5230 5550
rect 5290 5530 5310 5550
rect 5370 5530 5390 5550
rect 5450 5530 5470 5550
rect 5530 5530 5550 5550
rect 5610 5530 5630 5550
rect 5690 5530 5710 5550
rect 5770 5530 5790 5550
rect 5850 5530 5870 5550
rect 5930 5530 5950 5550
rect 6010 5530 6030 5550
rect 6090 5530 6110 5550
rect 6170 5530 6190 5550
rect 4250 5450 4270 5470
rect 4330 5450 4350 5470
rect 4410 5450 4430 5470
rect 4490 5450 4510 5470
rect 4570 5450 4590 5470
rect 4650 5450 4670 5470
rect 4730 5450 4750 5470
rect 4810 5450 4830 5470
rect 4890 5450 4910 5470
rect 4970 5450 4990 5470
rect 5050 5450 5070 5470
rect 5130 5450 5150 5470
rect 5210 5450 5230 5470
rect 5290 5450 5310 5470
rect 5370 5450 5390 5470
rect 5450 5450 5470 5470
rect 5530 5450 5550 5470
rect 5610 5450 5630 5470
rect 5690 5450 5710 5470
rect 5770 5450 5790 5470
rect 5850 5450 5870 5470
rect 5930 5450 5950 5470
rect 6010 5450 6030 5470
rect 6090 5450 6110 5470
rect 6170 5450 6190 5470
rect 4250 5370 4270 5390
rect 4330 5370 4350 5390
rect 4410 5370 4430 5390
rect 4490 5370 4510 5390
rect 4570 5370 4590 5390
rect 4650 5370 4670 5390
rect 4730 5370 4750 5390
rect 4810 5370 4830 5390
rect 4890 5370 4910 5390
rect 4970 5370 4990 5390
rect 5050 5370 5070 5390
rect 5130 5370 5150 5390
rect 5210 5370 5230 5390
rect 5290 5370 5310 5390
rect 5370 5370 5390 5390
rect 5450 5370 5470 5390
rect 5530 5370 5550 5390
rect 5610 5370 5630 5390
rect 5690 5370 5710 5390
rect 5770 5370 5790 5390
rect 5850 5370 5870 5390
rect 5930 5370 5950 5390
rect 6010 5370 6030 5390
rect 6090 5370 6110 5390
rect 6170 5370 6190 5390
rect 4250 5290 4270 5310
rect 4330 5290 4350 5310
rect 4410 5290 4430 5310
rect 4490 5290 4510 5310
rect 4570 5290 4590 5310
rect 4650 5290 4670 5310
rect 4730 5290 4750 5310
rect 4810 5290 4830 5310
rect 4890 5290 4910 5310
rect 4970 5290 4990 5310
rect 5050 5290 5070 5310
rect 5130 5290 5150 5310
rect 5210 5290 5230 5310
rect 5290 5290 5310 5310
rect 5370 5290 5390 5310
rect 5450 5290 5470 5310
rect 5530 5290 5550 5310
rect 5610 5290 5630 5310
rect 5690 5290 5710 5310
rect 5770 5290 5790 5310
rect 5850 5290 5870 5310
rect 5930 5290 5950 5310
rect 6010 5290 6030 5310
rect 6090 5290 6110 5310
rect 6170 5290 6190 5310
rect 4250 5210 4270 5230
rect 4330 5210 4350 5230
rect 4410 5210 4430 5230
rect 4490 5210 4510 5230
rect 4570 5210 4590 5230
rect 4650 5210 4670 5230
rect 4730 5210 4750 5230
rect 4810 5210 4830 5230
rect 4890 5210 4910 5230
rect 4970 5210 4990 5230
rect 5050 5210 5070 5230
rect 5130 5210 5150 5230
rect 5210 5210 5230 5230
rect 5290 5210 5310 5230
rect 5370 5210 5390 5230
rect 5450 5210 5470 5230
rect 5530 5210 5550 5230
rect 5610 5210 5630 5230
rect 5690 5210 5710 5230
rect 5770 5210 5790 5230
rect 5850 5210 5870 5230
rect 5930 5210 5950 5230
rect 6010 5210 6030 5230
rect 6090 5210 6110 5230
rect 6170 5210 6190 5230
rect 4250 5130 4270 5150
rect 4330 5130 4350 5150
rect 4410 5130 4430 5150
rect 4490 5130 4510 5150
rect 4570 5130 4590 5150
rect 4650 5130 4670 5150
rect 4730 5130 4750 5150
rect 4810 5130 4830 5150
rect 4890 5130 4910 5150
rect 4970 5130 4990 5150
rect 5050 5130 5070 5150
rect 5130 5130 5150 5150
rect 5210 5130 5230 5150
rect 5290 5130 5310 5150
rect 5370 5130 5390 5150
rect 5450 5130 5470 5150
rect 5530 5130 5550 5150
rect 5610 5130 5630 5150
rect 5690 5130 5710 5150
rect 5770 5130 5790 5150
rect 5850 5130 5870 5150
rect 5930 5130 5950 5150
rect 6010 5130 6030 5150
rect 6090 5130 6110 5150
rect 6170 5130 6190 5150
rect 4250 5050 4270 5070
rect 4330 5050 4350 5070
rect 4410 5050 4430 5070
rect 4490 5050 4510 5070
rect 4570 5050 4590 5070
rect 4650 5050 4670 5070
rect 4730 5050 4750 5070
rect 4810 5050 4830 5070
rect 4890 5050 4910 5070
rect 4970 5050 4990 5070
rect 5050 5050 5070 5070
rect 5130 5050 5150 5070
rect 5210 5050 5230 5070
rect 5290 5050 5310 5070
rect 5370 5050 5390 5070
rect 5450 5050 5470 5070
rect 5530 5050 5550 5070
rect 5610 5050 5630 5070
rect 5690 5050 5710 5070
rect 5770 5050 5790 5070
rect 5850 5050 5870 5070
rect 5930 5050 5950 5070
rect 6010 5050 6030 5070
rect 6090 5050 6110 5070
rect 6170 5050 6190 5070
rect 4250 4970 4270 4990
rect 4330 4970 4350 4990
rect 4410 4970 4430 4990
rect 4490 4970 4510 4990
rect 4570 4970 4590 4990
rect 4650 4970 4670 4990
rect 4730 4970 4750 4990
rect 4810 4970 4830 4990
rect 4890 4970 4910 4990
rect 4970 4970 4990 4990
rect 5050 4970 5070 4990
rect 5130 4970 5150 4990
rect 5210 4970 5230 4990
rect 5290 4970 5310 4990
rect 5370 4970 5390 4990
rect 5450 4970 5470 4990
rect 5530 4970 5550 4990
rect 5610 4970 5630 4990
rect 5690 4970 5710 4990
rect 5770 4970 5790 4990
rect 5850 4970 5870 4990
rect 5930 4970 5950 4990
rect 6010 4970 6030 4990
rect 6090 4970 6110 4990
rect 6170 4970 6190 4990
rect 4250 4890 4270 4910
rect 4330 4890 4350 4910
rect 4410 4890 4430 4910
rect 4490 4890 4510 4910
rect 4570 4890 4590 4910
rect 4650 4890 4670 4910
rect 4730 4890 4750 4910
rect 4810 4890 4830 4910
rect 4890 4890 4910 4910
rect 4970 4890 4990 4910
rect 5050 4890 5070 4910
rect 5130 4890 5150 4910
rect 5210 4890 5230 4910
rect 5290 4890 5310 4910
rect 5370 4890 5390 4910
rect 5450 4890 5470 4910
rect 5530 4890 5550 4910
rect 5610 4890 5630 4910
rect 5690 4890 5710 4910
rect 5770 4890 5790 4910
rect 5850 4890 5870 4910
rect 5930 4890 5950 4910
rect 6010 4890 6030 4910
rect 6090 4890 6110 4910
rect 6170 4890 6190 4910
rect 4250 4810 4270 4830
rect 4330 4810 4350 4830
rect 4410 4810 4430 4830
rect 4490 4810 4510 4830
rect 4570 4810 4590 4830
rect 4650 4810 4670 4830
rect 4730 4810 4750 4830
rect 4810 4810 4830 4830
rect 4890 4810 4910 4830
rect 4970 4810 4990 4830
rect 5050 4810 5070 4830
rect 5130 4810 5150 4830
rect 5210 4810 5230 4830
rect 5290 4810 5310 4830
rect 5370 4810 5390 4830
rect 5450 4810 5470 4830
rect 5530 4810 5550 4830
rect 5610 4810 5630 4830
rect 5690 4810 5710 4830
rect 5770 4810 5790 4830
rect 5850 4810 5870 4830
rect 5930 4810 5950 4830
rect 6010 4810 6030 4830
rect 6090 4810 6110 4830
rect 6170 4810 6190 4830
rect 4250 4730 4270 4750
rect 4330 4730 4350 4750
rect 4410 4730 4430 4750
rect 4490 4730 4510 4750
rect 4570 4730 4590 4750
rect 4650 4730 4670 4750
rect 4730 4730 4750 4750
rect 4810 4730 4830 4750
rect 4890 4730 4910 4750
rect 4970 4730 4990 4750
rect 5050 4730 5070 4750
rect 5130 4730 5150 4750
rect 5210 4730 5230 4750
rect 5290 4730 5310 4750
rect 5370 4730 5390 4750
rect 5450 4730 5470 4750
rect 5530 4730 5550 4750
rect 5610 4730 5630 4750
rect 5690 4730 5710 4750
rect 5770 4730 5790 4750
rect 5850 4730 5870 4750
rect 5930 4730 5950 4750
rect 6010 4730 6030 4750
rect 6090 4730 6110 4750
rect 6170 4730 6190 4750
rect 4250 4650 4270 4670
rect 4330 4650 4350 4670
rect 4410 4650 4430 4670
rect 4490 4650 4510 4670
rect 4570 4650 4590 4670
rect 4650 4650 4670 4670
rect 4730 4650 4750 4670
rect 4810 4650 4830 4670
rect 4890 4650 4910 4670
rect 4970 4650 4990 4670
rect 5050 4650 5070 4670
rect 5130 4650 5150 4670
rect 5210 4650 5230 4670
rect 5290 4650 5310 4670
rect 5370 4650 5390 4670
rect 5450 4650 5470 4670
rect 5530 4650 5550 4670
rect 5610 4650 5630 4670
rect 5690 4650 5710 4670
rect 5770 4650 5790 4670
rect 5850 4650 5870 4670
rect 5930 4650 5950 4670
rect 6010 4650 6030 4670
rect 6090 4650 6110 4670
rect 6170 4650 6190 4670
rect 4250 4570 4270 4590
rect 4330 4570 4350 4590
rect 4410 4570 4430 4590
rect 4490 4570 4510 4590
rect 4570 4570 4590 4590
rect 4650 4570 4670 4590
rect 4730 4570 4750 4590
rect 4810 4570 4830 4590
rect 4890 4570 4910 4590
rect 4970 4570 4990 4590
rect 5050 4570 5070 4590
rect 5130 4570 5150 4590
rect 5210 4570 5230 4590
rect 5290 4570 5310 4590
rect 5370 4570 5390 4590
rect 5450 4570 5470 4590
rect 5530 4570 5550 4590
rect 5610 4570 5630 4590
rect 5690 4570 5710 4590
rect 5770 4570 5790 4590
rect 5850 4570 5870 4590
rect 5930 4570 5950 4590
rect 6010 4570 6030 4590
rect 6090 4570 6110 4590
rect 6170 4570 6190 4590
rect 4250 4490 4270 4510
rect 4330 4490 4350 4510
rect 4410 4490 4430 4510
rect 4490 4490 4510 4510
rect 4570 4490 4590 4510
rect 4650 4490 4670 4510
rect 4730 4490 4750 4510
rect 4810 4490 4830 4510
rect 4890 4490 4910 4510
rect 4970 4490 4990 4510
rect 5050 4490 5070 4510
rect 5130 4490 5150 4510
rect 5210 4490 5230 4510
rect 5290 4490 5310 4510
rect 5370 4490 5390 4510
rect 5450 4490 5470 4510
rect 5530 4490 5550 4510
rect 5610 4490 5630 4510
rect 5690 4490 5710 4510
rect 5770 4490 5790 4510
rect 5850 4490 5870 4510
rect 5930 4490 5950 4510
rect 6010 4490 6030 4510
rect 6090 4490 6110 4510
rect 6170 4490 6190 4510
rect 4250 4410 4270 4430
rect 4330 4410 4350 4430
rect 4410 4410 4430 4430
rect 4490 4410 4510 4430
rect 4570 4410 4590 4430
rect 4650 4410 4670 4430
rect 4730 4410 4750 4430
rect 4810 4410 4830 4430
rect 4890 4410 4910 4430
rect 4970 4410 4990 4430
rect 5050 4410 5070 4430
rect 5130 4410 5150 4430
rect 5210 4410 5230 4430
rect 5290 4410 5310 4430
rect 5370 4410 5390 4430
rect 5450 4410 5470 4430
rect 5530 4410 5550 4430
rect 5610 4410 5630 4430
rect 5690 4410 5710 4430
rect 5770 4410 5790 4430
rect 5850 4410 5870 4430
rect 5930 4410 5950 4430
rect 6010 4410 6030 4430
rect 6090 4410 6110 4430
rect 6170 4410 6190 4430
rect 4250 4330 4270 4350
rect 4330 4330 4350 4350
rect 4410 4330 4430 4350
rect 4490 4330 4510 4350
rect 4570 4330 4590 4350
rect 4650 4330 4670 4350
rect 4730 4330 4750 4350
rect 4810 4330 4830 4350
rect 4890 4330 4910 4350
rect 4970 4330 4990 4350
rect 5050 4330 5070 4350
rect 5130 4330 5150 4350
rect 5210 4330 5230 4350
rect 5290 4330 5310 4350
rect 5370 4330 5390 4350
rect 5450 4330 5470 4350
rect 5530 4330 5550 4350
rect 5610 4330 5630 4350
rect 5690 4330 5710 4350
rect 5770 4330 5790 4350
rect 5850 4330 5870 4350
rect 5930 4330 5950 4350
rect 6010 4330 6030 4350
rect 6090 4330 6110 4350
rect 6170 4330 6190 4350
rect 4250 4250 4270 4270
rect 4330 4250 4350 4270
rect 4410 4250 4430 4270
rect 4490 4250 4510 4270
rect 4570 4250 4590 4270
rect 4650 4250 4670 4270
rect 4730 4250 4750 4270
rect 4810 4250 4830 4270
rect 4890 4250 4910 4270
rect 4970 4250 4990 4270
rect 5050 4250 5070 4270
rect 5130 4250 5150 4270
rect 5210 4250 5230 4270
rect 5290 4250 5310 4270
rect 5370 4250 5390 4270
rect 5450 4250 5470 4270
rect 5530 4250 5550 4270
rect 5610 4250 5630 4270
rect 5690 4250 5710 4270
rect 5770 4250 5790 4270
rect 5850 4250 5870 4270
rect 5930 4250 5950 4270
rect 6010 4250 6030 4270
rect 6090 4250 6110 4270
rect 6170 4250 6190 4270
rect 4250 4170 4270 4190
rect 4330 4170 4350 4190
rect 4410 4170 4430 4190
rect 4490 4170 4510 4190
rect 4570 4170 4590 4190
rect 4650 4170 4670 4190
rect 4730 4170 4750 4190
rect 4810 4170 4830 4190
rect 4890 4170 4910 4190
rect 4970 4170 4990 4190
rect 5050 4170 5070 4190
rect 5130 4170 5150 4190
rect 5210 4170 5230 4190
rect 5290 4170 5310 4190
rect 5370 4170 5390 4190
rect 5450 4170 5470 4190
rect 5530 4170 5550 4190
rect 5610 4170 5630 4190
rect 5690 4170 5710 4190
rect 5770 4170 5790 4190
rect 5850 4170 5870 4190
rect 5930 4170 5950 4190
rect 6010 4170 6030 4190
rect 6090 4170 6110 4190
rect 6170 4170 6190 4190
rect 4250 4090 4270 4110
rect 4330 4090 4350 4110
rect 4410 4090 4430 4110
rect 4490 4090 4510 4110
rect 4570 4090 4590 4110
rect 4650 4090 4670 4110
rect 4730 4090 4750 4110
rect 4810 4090 4830 4110
rect 4890 4090 4910 4110
rect 4970 4090 4990 4110
rect 5050 4090 5070 4110
rect 5130 4090 5150 4110
rect 5210 4090 5230 4110
rect 5290 4090 5310 4110
rect 5370 4090 5390 4110
rect 5450 4090 5470 4110
rect 5530 4090 5550 4110
rect 5610 4090 5630 4110
rect 5690 4090 5710 4110
rect 5770 4090 5790 4110
rect 5850 4090 5870 4110
rect 5930 4090 5950 4110
rect 6010 4090 6030 4110
rect 6090 4090 6110 4110
rect 6170 4090 6190 4110
rect 4250 4010 4270 4030
rect 4330 4010 4350 4030
rect 4410 4010 4430 4030
rect 4490 4010 4510 4030
rect 4570 4010 4590 4030
rect 4650 4010 4670 4030
rect 4730 4010 4750 4030
rect 4810 4010 4830 4030
rect 4890 4010 4910 4030
rect 4970 4010 4990 4030
rect 5050 4010 5070 4030
rect 5130 4010 5150 4030
rect 5210 4010 5230 4030
rect 5290 4010 5310 4030
rect 5370 4010 5390 4030
rect 5450 4010 5470 4030
rect 5530 4010 5550 4030
rect 5610 4010 5630 4030
rect 5690 4010 5710 4030
rect 5770 4010 5790 4030
rect 5850 4010 5870 4030
rect 5930 4010 5950 4030
rect 6010 4010 6030 4030
rect 6090 4010 6110 4030
rect 6170 4010 6190 4030
rect 4250 3930 4270 3950
rect 4330 3930 4350 3950
rect 4410 3930 4430 3950
rect 4490 3930 4510 3950
rect 4570 3930 4590 3950
rect 4650 3930 4670 3950
rect 4730 3930 4750 3950
rect 4810 3930 4830 3950
rect 4890 3930 4910 3950
rect 4970 3930 4990 3950
rect 5050 3930 5070 3950
rect 5130 3930 5150 3950
rect 5210 3930 5230 3950
rect 5290 3930 5310 3950
rect 5370 3930 5390 3950
rect 5450 3930 5470 3950
rect 5530 3930 5550 3950
rect 5610 3930 5630 3950
rect 5690 3930 5710 3950
rect 5770 3930 5790 3950
rect 5850 3930 5870 3950
rect 5930 3930 5950 3950
rect 6010 3930 6030 3950
rect 6090 3930 6110 3950
rect 6170 3930 6190 3950
rect 4250 3850 4270 3870
rect 4330 3850 4350 3870
rect 4410 3850 4430 3870
rect 4490 3850 4510 3870
rect 4570 3850 4590 3870
rect 4650 3850 4670 3870
rect 4730 3850 4750 3870
rect 4810 3850 4830 3870
rect 4890 3850 4910 3870
rect 4970 3850 4990 3870
rect 5050 3850 5070 3870
rect 5130 3850 5150 3870
rect 5210 3850 5230 3870
rect 5290 3850 5310 3870
rect 5370 3850 5390 3870
rect 5450 3850 5470 3870
rect 5530 3850 5550 3870
rect 5610 3850 5630 3870
rect 5690 3850 5710 3870
rect 5770 3850 5790 3870
rect 5850 3850 5870 3870
rect 5930 3850 5950 3870
rect 6010 3850 6030 3870
rect 6090 3850 6110 3870
rect 6170 3850 6190 3870
rect 4250 3770 4270 3790
rect 4330 3770 4350 3790
rect 4410 3770 4430 3790
rect 4490 3770 4510 3790
rect 4570 3770 4590 3790
rect 4650 3770 4670 3790
rect 4730 3770 4750 3790
rect 4810 3770 4830 3790
rect 4890 3770 4910 3790
rect 4970 3770 4990 3790
rect 5050 3770 5070 3790
rect 5130 3770 5150 3790
rect 5210 3770 5230 3790
rect 5290 3770 5310 3790
rect 5370 3770 5390 3790
rect 5450 3770 5470 3790
rect 5530 3770 5550 3790
rect 5610 3770 5630 3790
rect 5690 3770 5710 3790
rect 5770 3770 5790 3790
rect 5850 3770 5870 3790
rect 5930 3770 5950 3790
rect 6010 3770 6030 3790
rect 6090 3770 6110 3790
rect 6170 3770 6190 3790
rect 4250 3690 4270 3710
rect 4330 3690 4350 3710
rect 4410 3690 4430 3710
rect 4490 3690 4510 3710
rect 4570 3690 4590 3710
rect 4650 3690 4670 3710
rect 4730 3690 4750 3710
rect 4810 3690 4830 3710
rect 4890 3690 4910 3710
rect 4970 3690 4990 3710
rect 5050 3690 5070 3710
rect 5130 3690 5150 3710
rect 5210 3690 5230 3710
rect 5290 3690 5310 3710
rect 5370 3690 5390 3710
rect 5450 3690 5470 3710
rect 5530 3690 5550 3710
rect 5610 3690 5630 3710
rect 5690 3690 5710 3710
rect 5770 3690 5790 3710
rect 5850 3690 5870 3710
rect 5930 3690 5950 3710
rect 6010 3690 6030 3710
rect 6090 3690 6110 3710
rect 6170 3690 6190 3710
rect 4250 3610 4270 3630
rect 4330 3610 4350 3630
rect 4410 3610 4430 3630
rect 4490 3610 4510 3630
rect 4570 3610 4590 3630
rect 4650 3610 4670 3630
rect 4730 3610 4750 3630
rect 4810 3610 4830 3630
rect 4890 3610 4910 3630
rect 4970 3610 4990 3630
rect 5050 3610 5070 3630
rect 5130 3610 5150 3630
rect 5210 3610 5230 3630
rect 5290 3610 5310 3630
rect 5370 3610 5390 3630
rect 5450 3610 5470 3630
rect 5530 3610 5550 3630
rect 5610 3610 5630 3630
rect 5690 3610 5710 3630
rect 5770 3610 5790 3630
rect 5850 3610 5870 3630
rect 5930 3610 5950 3630
rect 6010 3610 6030 3630
rect 6090 3610 6110 3630
rect 6170 3610 6190 3630
rect 4250 3530 4270 3550
rect 4330 3530 4350 3550
rect 4410 3530 4430 3550
rect 4490 3530 4510 3550
rect 4570 3530 4590 3550
rect 4650 3530 4670 3550
rect 4730 3530 4750 3550
rect 4810 3530 4830 3550
rect 4890 3530 4910 3550
rect 4970 3530 4990 3550
rect 5050 3530 5070 3550
rect 5130 3530 5150 3550
rect 5210 3530 5230 3550
rect 5290 3530 5310 3550
rect 5370 3530 5390 3550
rect 5450 3530 5470 3550
rect 5530 3530 5550 3550
rect 5610 3530 5630 3550
rect 5690 3530 5710 3550
rect 5770 3530 5790 3550
rect 5850 3530 5870 3550
rect 5930 3530 5950 3550
rect 6010 3530 6030 3550
rect 6090 3530 6110 3550
rect 6170 3530 6190 3550
rect 4250 3450 4270 3470
rect 4330 3450 4350 3470
rect 4410 3450 4430 3470
rect 4490 3450 4510 3470
rect 4570 3450 4590 3470
rect 4650 3450 4670 3470
rect 4730 3450 4750 3470
rect 4810 3450 4830 3470
rect 4890 3450 4910 3470
rect 4970 3450 4990 3470
rect 5050 3450 5070 3470
rect 5130 3450 5150 3470
rect 5210 3450 5230 3470
rect 5290 3450 5310 3470
rect 5370 3450 5390 3470
rect 5450 3450 5470 3470
rect 5530 3450 5550 3470
rect 5610 3450 5630 3470
rect 5690 3450 5710 3470
rect 5770 3450 5790 3470
rect 5850 3450 5870 3470
rect 5930 3450 5950 3470
rect 6010 3450 6030 3470
rect 6090 3450 6110 3470
rect 6170 3450 6190 3470
rect 4250 3370 4270 3390
rect 4330 3370 4350 3390
rect 4410 3370 4430 3390
rect 4490 3370 4510 3390
rect 4570 3370 4590 3390
rect 4650 3370 4670 3390
rect 4730 3370 4750 3390
rect 4810 3370 4830 3390
rect 4890 3370 4910 3390
rect 4970 3370 4990 3390
rect 5050 3370 5070 3390
rect 5130 3370 5150 3390
rect 5210 3370 5230 3390
rect 5290 3370 5310 3390
rect 5370 3370 5390 3390
rect 5450 3370 5470 3390
rect 5530 3370 5550 3390
rect 5610 3370 5630 3390
rect 5690 3370 5710 3390
rect 5770 3370 5790 3390
rect 5850 3370 5870 3390
rect 5930 3370 5950 3390
rect 6010 3370 6030 3390
rect 6090 3370 6110 3390
rect 6170 3370 6190 3390
rect 4250 3290 4270 3310
rect 4330 3290 4350 3310
rect 4410 3290 4430 3310
rect 4490 3290 4510 3310
rect 4570 3290 4590 3310
rect 4650 3290 4670 3310
rect 4730 3290 4750 3310
rect 4810 3290 4830 3310
rect 4890 3290 4910 3310
rect 4970 3290 4990 3310
rect 5050 3290 5070 3310
rect 5130 3290 5150 3310
rect 5210 3290 5230 3310
rect 5290 3290 5310 3310
rect 5370 3290 5390 3310
rect 5450 3290 5470 3310
rect 5530 3290 5550 3310
rect 5610 3290 5630 3310
rect 5690 3290 5710 3310
rect 5770 3290 5790 3310
rect 5850 3290 5870 3310
rect 5930 3290 5950 3310
rect 6010 3290 6030 3310
rect 6090 3290 6110 3310
rect 6170 3290 6190 3310
rect 4250 3210 4270 3230
rect 4330 3210 4350 3230
rect 4410 3210 4430 3230
rect 4490 3210 4510 3230
rect 4570 3210 4590 3230
rect 4650 3210 4670 3230
rect 4730 3210 4750 3230
rect 4810 3210 4830 3230
rect 4890 3210 4910 3230
rect 4970 3210 4990 3230
rect 5050 3210 5070 3230
rect 5130 3210 5150 3230
rect 5210 3210 5230 3230
rect 5290 3210 5310 3230
rect 5370 3210 5390 3230
rect 5450 3210 5470 3230
rect 5530 3210 5550 3230
rect 5610 3210 5630 3230
rect 5690 3210 5710 3230
rect 5770 3210 5790 3230
rect 5850 3210 5870 3230
rect 5930 3210 5950 3230
rect 6010 3210 6030 3230
rect 6090 3210 6110 3230
rect 6170 3210 6190 3230
rect 4250 3130 4270 3150
rect 4330 3130 4350 3150
rect 4410 3130 4430 3150
rect 4490 3130 4510 3150
rect 4570 3130 4590 3150
rect 4650 3130 4670 3150
rect 4730 3130 4750 3150
rect 4810 3130 4830 3150
rect 4890 3130 4910 3150
rect 4970 3130 4990 3150
rect 5050 3130 5070 3150
rect 5130 3130 5150 3150
rect 5210 3130 5230 3150
rect 5290 3130 5310 3150
rect 5370 3130 5390 3150
rect 5450 3130 5470 3150
rect 5530 3130 5550 3150
rect 5610 3130 5630 3150
rect 5690 3130 5710 3150
rect 5770 3130 5790 3150
rect 5850 3130 5870 3150
rect 5930 3130 5950 3150
rect 6010 3130 6030 3150
rect 6090 3130 6110 3150
rect 6170 3130 6190 3150
rect 4250 3050 4270 3070
rect 4330 3050 4350 3070
rect 4410 3050 4430 3070
rect 4490 3050 4510 3070
rect 4570 3050 4590 3070
rect 4650 3050 4670 3070
rect 4730 3050 4750 3070
rect 4810 3050 4830 3070
rect 4890 3050 4910 3070
rect 4970 3050 4990 3070
rect 5050 3050 5070 3070
rect 5130 3050 5150 3070
rect 5210 3050 5230 3070
rect 5290 3050 5310 3070
rect 5370 3050 5390 3070
rect 5450 3050 5470 3070
rect 5530 3050 5550 3070
rect 5610 3050 5630 3070
rect 5690 3050 5710 3070
rect 5770 3050 5790 3070
rect 5850 3050 5870 3070
rect 5930 3050 5950 3070
rect 6010 3050 6030 3070
rect 6090 3050 6110 3070
rect 6170 3050 6190 3070
rect 4250 2970 4270 2990
rect 4330 2970 4350 2990
rect 4410 2970 4430 2990
rect 4490 2970 4510 2990
rect 4570 2970 4590 2990
rect 4650 2970 4670 2990
rect 4730 2970 4750 2990
rect 4810 2970 4830 2990
rect 4890 2970 4910 2990
rect 4970 2970 4990 2990
rect 5050 2970 5070 2990
rect 5130 2970 5150 2990
rect 5210 2970 5230 2990
rect 5290 2970 5310 2990
rect 5370 2970 5390 2990
rect 5450 2970 5470 2990
rect 5530 2970 5550 2990
rect 5610 2970 5630 2990
rect 5690 2970 5710 2990
rect 5770 2970 5790 2990
rect 5850 2970 5870 2990
rect 5930 2970 5950 2990
rect 6010 2970 6030 2990
rect 6090 2970 6110 2990
rect 6170 2970 6190 2990
rect 4250 2890 4270 2910
rect 4330 2890 4350 2910
rect 4410 2890 4430 2910
rect 4490 2890 4510 2910
rect 4570 2890 4590 2910
rect 4650 2890 4670 2910
rect 4730 2890 4750 2910
rect 4810 2890 4830 2910
rect 4890 2890 4910 2910
rect 4970 2890 4990 2910
rect 5050 2890 5070 2910
rect 5130 2890 5150 2910
rect 5210 2890 5230 2910
rect 5290 2890 5310 2910
rect 5370 2890 5390 2910
rect 5450 2890 5470 2910
rect 5530 2890 5550 2910
rect 5610 2890 5630 2910
rect 5690 2890 5710 2910
rect 5770 2890 5790 2910
rect 5850 2890 5870 2910
rect 5930 2890 5950 2910
rect 6010 2890 6030 2910
rect 6090 2890 6110 2910
rect 6170 2890 6190 2910
rect 4250 2810 4270 2830
rect 4330 2810 4350 2830
rect 4410 2810 4430 2830
rect 4490 2810 4510 2830
rect 4570 2810 4590 2830
rect 4650 2810 4670 2830
rect 4730 2810 4750 2830
rect 4810 2810 4830 2830
rect 4890 2810 4910 2830
rect 4970 2810 4990 2830
rect 5050 2810 5070 2830
rect 5130 2810 5150 2830
rect 5210 2810 5230 2830
rect 5290 2810 5310 2830
rect 5370 2810 5390 2830
rect 5450 2810 5470 2830
rect 5530 2810 5550 2830
rect 5610 2810 5630 2830
rect 5690 2810 5710 2830
rect 5770 2810 5790 2830
rect 5850 2810 5870 2830
rect 5930 2810 5950 2830
rect 6010 2810 6030 2830
rect 6090 2810 6110 2830
rect 6170 2810 6190 2830
rect 4250 2730 4270 2750
rect 4330 2730 4350 2750
rect 4410 2730 4430 2750
rect 4490 2730 4510 2750
rect 4570 2730 4590 2750
rect 4650 2730 4670 2750
rect 4730 2730 4750 2750
rect 4810 2730 4830 2750
rect 4890 2730 4910 2750
rect 4970 2730 4990 2750
rect 5050 2730 5070 2750
rect 5130 2730 5150 2750
rect 5210 2730 5230 2750
rect 5290 2730 5310 2750
rect 5370 2730 5390 2750
rect 5450 2730 5470 2750
rect 5530 2730 5550 2750
rect 5610 2730 5630 2750
rect 5690 2730 5710 2750
rect 5770 2730 5790 2750
rect 5850 2730 5870 2750
rect 5930 2730 5950 2750
rect 6010 2730 6030 2750
rect 6090 2730 6110 2750
rect 6170 2730 6190 2750
rect 4250 2650 4270 2670
rect 4330 2650 4350 2670
rect 4410 2650 4430 2670
rect 4490 2650 4510 2670
rect 4570 2650 4590 2670
rect 4650 2650 4670 2670
rect 4730 2650 4750 2670
rect 4810 2650 4830 2670
rect 4890 2650 4910 2670
rect 4970 2650 4990 2670
rect 5050 2650 5070 2670
rect 5130 2650 5150 2670
rect 5210 2650 5230 2670
rect 5290 2650 5310 2670
rect 5370 2650 5390 2670
rect 5450 2650 5470 2670
rect 5530 2650 5550 2670
rect 5610 2650 5630 2670
rect 5690 2650 5710 2670
rect 5770 2650 5790 2670
rect 5850 2650 5870 2670
rect 5930 2650 5950 2670
rect 6010 2650 6030 2670
rect 6090 2650 6110 2670
rect 6170 2650 6190 2670
rect 4250 2570 4270 2590
rect 4330 2570 4350 2590
rect 4410 2570 4430 2590
rect 4490 2570 4510 2590
rect 4570 2570 4590 2590
rect 4650 2570 4670 2590
rect 4730 2570 4750 2590
rect 4810 2570 4830 2590
rect 4890 2570 4910 2590
rect 4970 2570 4990 2590
rect 5050 2570 5070 2590
rect 5130 2570 5150 2590
rect 5210 2570 5230 2590
rect 5290 2570 5310 2590
rect 5370 2570 5390 2590
rect 5450 2570 5470 2590
rect 5530 2570 5550 2590
rect 5610 2570 5630 2590
rect 5690 2570 5710 2590
rect 5770 2570 5790 2590
rect 5850 2570 5870 2590
rect 5930 2570 5950 2590
rect 6010 2570 6030 2590
rect 6090 2570 6110 2590
rect 6170 2570 6190 2590
rect 4250 2490 4270 2510
rect 4330 2490 4350 2510
rect 4410 2490 4430 2510
rect 4490 2490 4510 2510
rect 4570 2490 4590 2510
rect 4650 2490 4670 2510
rect 4730 2490 4750 2510
rect 4810 2490 4830 2510
rect 4890 2490 4910 2510
rect 4970 2490 4990 2510
rect 5050 2490 5070 2510
rect 5130 2490 5150 2510
rect 5210 2490 5230 2510
rect 5290 2490 5310 2510
rect 5370 2490 5390 2510
rect 5450 2490 5470 2510
rect 5530 2490 5550 2510
rect 5610 2490 5630 2510
rect 5690 2490 5710 2510
rect 5770 2490 5790 2510
rect 5850 2490 5870 2510
rect 5930 2490 5950 2510
rect 6010 2490 6030 2510
rect 6090 2490 6110 2510
rect 6170 2490 6190 2510
rect 4250 2410 4270 2430
rect 4330 2410 4350 2430
rect 4410 2410 4430 2430
rect 4490 2410 4510 2430
rect 4570 2410 4590 2430
rect 4650 2410 4670 2430
rect 4730 2410 4750 2430
rect 4810 2410 4830 2430
rect 4890 2410 4910 2430
rect 4970 2410 4990 2430
rect 5050 2410 5070 2430
rect 5130 2410 5150 2430
rect 5210 2410 5230 2430
rect 5290 2410 5310 2430
rect 5370 2410 5390 2430
rect 5450 2410 5470 2430
rect 5530 2410 5550 2430
rect 5610 2410 5630 2430
rect 5690 2410 5710 2430
rect 5770 2410 5790 2430
rect 5850 2410 5870 2430
rect 5930 2410 5950 2430
rect 6010 2410 6030 2430
rect 6090 2410 6110 2430
rect 6170 2410 6190 2430
rect 4250 2330 4270 2350
rect 4330 2330 4350 2350
rect 4410 2330 4430 2350
rect 4490 2330 4510 2350
rect 4570 2330 4590 2350
rect 4650 2330 4670 2350
rect 4730 2330 4750 2350
rect 4810 2330 4830 2350
rect 4890 2330 4910 2350
rect 4970 2330 4990 2350
rect 5050 2330 5070 2350
rect 5130 2330 5150 2350
rect 5210 2330 5230 2350
rect 5290 2330 5310 2350
rect 5370 2330 5390 2350
rect 5450 2330 5470 2350
rect 5530 2330 5550 2350
rect 5610 2330 5630 2350
rect 5690 2330 5710 2350
rect 5770 2330 5790 2350
rect 5850 2330 5870 2350
rect 5930 2330 5950 2350
rect 6010 2330 6030 2350
rect 6090 2330 6110 2350
rect 6170 2330 6190 2350
rect 4250 2250 4270 2270
rect 4330 2250 4350 2270
rect 4410 2250 4430 2270
rect 4490 2250 4510 2270
rect 4570 2250 4590 2270
rect 4650 2250 4670 2270
rect 4730 2250 4750 2270
rect 4810 2250 4830 2270
rect 4890 2250 4910 2270
rect 4970 2250 4990 2270
rect 5050 2250 5070 2270
rect 5130 2250 5150 2270
rect 5210 2250 5230 2270
rect 5290 2250 5310 2270
rect 5370 2250 5390 2270
rect 5450 2250 5470 2270
rect 5530 2250 5550 2270
rect 5610 2250 5630 2270
rect 5690 2250 5710 2270
rect 5770 2250 5790 2270
rect 5850 2250 5870 2270
rect 5930 2250 5950 2270
rect 6010 2250 6030 2270
rect 6090 2250 6110 2270
rect 6170 2250 6190 2270
rect 4250 2170 4270 2190
rect 4330 2170 4350 2190
rect 4410 2170 4430 2190
rect 4490 2170 4510 2190
rect 4570 2170 4590 2190
rect 4650 2170 4670 2190
rect 4730 2170 4750 2190
rect 4810 2170 4830 2190
rect 4890 2170 4910 2190
rect 4970 2170 4990 2190
rect 5050 2170 5070 2190
rect 5130 2170 5150 2190
rect 5210 2170 5230 2190
rect 5290 2170 5310 2190
rect 5370 2170 5390 2190
rect 5450 2170 5470 2190
rect 5530 2170 5550 2190
rect 5610 2170 5630 2190
rect 5690 2170 5710 2190
rect 5770 2170 5790 2190
rect 5850 2170 5870 2190
rect 5930 2170 5950 2190
rect 6010 2170 6030 2190
rect 6090 2170 6110 2190
rect 6170 2170 6190 2190
rect 4250 2090 4270 2110
rect 4330 2090 4350 2110
rect 4410 2090 4430 2110
rect 4490 2090 4510 2110
rect 4570 2090 4590 2110
rect 4650 2090 4670 2110
rect 4730 2090 4750 2110
rect 4810 2090 4830 2110
rect 4890 2090 4910 2110
rect 4970 2090 4990 2110
rect 5050 2090 5070 2110
rect 5130 2090 5150 2110
rect 5210 2090 5230 2110
rect 5290 2090 5310 2110
rect 5370 2090 5390 2110
rect 5450 2090 5470 2110
rect 5530 2090 5550 2110
rect 5610 2090 5630 2110
rect 5690 2090 5710 2110
rect 5770 2090 5790 2110
rect 5850 2090 5870 2110
rect 5930 2090 5950 2110
rect 6010 2090 6030 2110
rect 6090 2090 6110 2110
rect 6170 2090 6190 2110
rect 4250 2010 4270 2030
rect 4330 2010 4350 2030
rect 4410 2010 4430 2030
rect 4490 2010 4510 2030
rect 4570 2010 4590 2030
rect 4650 2010 4670 2030
rect 4730 2010 4750 2030
rect 4810 2010 4830 2030
rect 4890 2010 4910 2030
rect 4970 2010 4990 2030
rect 5050 2010 5070 2030
rect 5130 2010 5150 2030
rect 5210 2010 5230 2030
rect 5290 2010 5310 2030
rect 5370 2010 5390 2030
rect 5450 2010 5470 2030
rect 5530 2010 5550 2030
rect 5610 2010 5630 2030
rect 5690 2010 5710 2030
rect 5770 2010 5790 2030
rect 5850 2010 5870 2030
rect 5930 2010 5950 2030
rect 6010 2010 6030 2030
rect 6090 2010 6110 2030
rect 6170 2010 6190 2030
rect 4250 1930 4270 1950
rect 4330 1930 4350 1950
rect 4410 1930 4430 1950
rect 4490 1930 4510 1950
rect 4570 1930 4590 1950
rect 4650 1930 4670 1950
rect 4730 1930 4750 1950
rect 4810 1930 4830 1950
rect 4890 1930 4910 1950
rect 4970 1930 4990 1950
rect 5050 1930 5070 1950
rect 5130 1930 5150 1950
rect 5210 1930 5230 1950
rect 5290 1930 5310 1950
rect 5370 1930 5390 1950
rect 5450 1930 5470 1950
rect 5530 1930 5550 1950
rect 5610 1930 5630 1950
rect 5690 1930 5710 1950
rect 5770 1930 5790 1950
rect 5850 1930 5870 1950
rect 5930 1930 5950 1950
rect 6010 1930 6030 1950
rect 6090 1930 6110 1950
rect 6170 1930 6190 1950
rect 4250 1850 4270 1870
rect 4330 1850 4350 1870
rect 4410 1850 4430 1870
rect 4490 1850 4510 1870
rect 4570 1850 4590 1870
rect 4650 1850 4670 1870
rect 4730 1850 4750 1870
rect 4810 1850 4830 1870
rect 4890 1850 4910 1870
rect 4970 1850 4990 1870
rect 5050 1850 5070 1870
rect 5130 1850 5150 1870
rect 5210 1850 5230 1870
rect 5290 1850 5310 1870
rect 5370 1850 5390 1870
rect 5450 1850 5470 1870
rect 5530 1850 5550 1870
rect 5610 1850 5630 1870
rect 5690 1850 5710 1870
rect 5770 1850 5790 1870
rect 5850 1850 5870 1870
rect 5930 1850 5950 1870
rect 6010 1850 6030 1870
rect 6090 1850 6110 1870
rect 6170 1850 6190 1870
rect 4250 1770 4270 1790
rect 4330 1770 4350 1790
rect 4410 1770 4430 1790
rect 4490 1770 4510 1790
rect 4570 1770 4590 1790
rect 4650 1770 4670 1790
rect 4730 1770 4750 1790
rect 4810 1770 4830 1790
rect 4890 1770 4910 1790
rect 4970 1770 4990 1790
rect 5050 1770 5070 1790
rect 5130 1770 5150 1790
rect 5210 1770 5230 1790
rect 5290 1770 5310 1790
rect 5370 1770 5390 1790
rect 5450 1770 5470 1790
rect 5530 1770 5550 1790
rect 5610 1770 5630 1790
rect 5690 1770 5710 1790
rect 5770 1770 5790 1790
rect 5850 1770 5870 1790
rect 5930 1770 5950 1790
rect 6010 1770 6030 1790
rect 6090 1770 6110 1790
rect 6170 1770 6190 1790
rect 4250 1690 4270 1710
rect 4330 1690 4350 1710
rect 4410 1690 4430 1710
rect 4490 1690 4510 1710
rect 4570 1690 4590 1710
rect 4650 1690 4670 1710
rect 4730 1690 4750 1710
rect 4810 1690 4830 1710
rect 4890 1690 4910 1710
rect 4970 1690 4990 1710
rect 5050 1690 5070 1710
rect 5130 1690 5150 1710
rect 5210 1690 5230 1710
rect 5290 1690 5310 1710
rect 5370 1690 5390 1710
rect 5450 1690 5470 1710
rect 5530 1690 5550 1710
rect 5610 1690 5630 1710
rect 5690 1690 5710 1710
rect 5770 1690 5790 1710
rect 5850 1690 5870 1710
rect 5930 1690 5950 1710
rect 6010 1690 6030 1710
rect 6090 1690 6110 1710
rect 6170 1690 6190 1710
rect 4250 1610 4270 1630
rect 4330 1610 4350 1630
rect 4410 1610 4430 1630
rect 4490 1610 4510 1630
rect 4570 1610 4590 1630
rect 4650 1610 4670 1630
rect 4730 1610 4750 1630
rect 4810 1610 4830 1630
rect 4890 1610 4910 1630
rect 4970 1610 4990 1630
rect 5050 1610 5070 1630
rect 5130 1610 5150 1630
rect 5210 1610 5230 1630
rect 5290 1610 5310 1630
rect 5370 1610 5390 1630
rect 5450 1610 5470 1630
rect 5530 1610 5550 1630
rect 5610 1610 5630 1630
rect 5690 1610 5710 1630
rect 5770 1610 5790 1630
rect 5850 1610 5870 1630
rect 5930 1610 5950 1630
rect 6010 1610 6030 1630
rect 6090 1610 6110 1630
rect 6170 1610 6190 1630
rect 4250 1530 4270 1550
rect 4330 1530 4350 1550
rect 4410 1530 4430 1550
rect 4490 1530 4510 1550
rect 4570 1530 4590 1550
rect 4650 1530 4670 1550
rect 4730 1530 4750 1550
rect 4810 1530 4830 1550
rect 4890 1530 4910 1550
rect 4970 1530 4990 1550
rect 5050 1530 5070 1550
rect 5130 1530 5150 1550
rect 5210 1530 5230 1550
rect 5290 1530 5310 1550
rect 5370 1530 5390 1550
rect 5450 1530 5470 1550
rect 5530 1530 5550 1550
rect 5610 1530 5630 1550
rect 5690 1530 5710 1550
rect 5770 1530 5790 1550
rect 5850 1530 5870 1550
rect 5930 1530 5950 1550
rect 6010 1530 6030 1550
rect 6090 1530 6110 1550
rect 6170 1530 6190 1550
rect 4250 1450 4270 1470
rect 4330 1450 4350 1470
rect 4410 1450 4430 1470
rect 4490 1450 4510 1470
rect 4570 1450 4590 1470
rect 4650 1450 4670 1470
rect 4730 1450 4750 1470
rect 4810 1450 4830 1470
rect 4890 1450 4910 1470
rect 4970 1450 4990 1470
rect 5050 1450 5070 1470
rect 5130 1450 5150 1470
rect 5210 1450 5230 1470
rect 5290 1450 5310 1470
rect 5370 1450 5390 1470
rect 5450 1450 5470 1470
rect 5530 1450 5550 1470
rect 5610 1450 5630 1470
rect 5690 1450 5710 1470
rect 5770 1450 5790 1470
rect 5850 1450 5870 1470
rect 5930 1450 5950 1470
rect 6010 1450 6030 1470
rect 6090 1450 6110 1470
rect 6170 1450 6190 1470
rect 4250 1370 4270 1390
rect 4330 1370 4350 1390
rect 4410 1370 4430 1390
rect 4490 1370 4510 1390
rect 4570 1370 4590 1390
rect 4650 1370 4670 1390
rect 4730 1370 4750 1390
rect 4810 1370 4830 1390
rect 4890 1370 4910 1390
rect 4970 1370 4990 1390
rect 5050 1370 5070 1390
rect 5130 1370 5150 1390
rect 5210 1370 5230 1390
rect 5290 1370 5310 1390
rect 5370 1370 5390 1390
rect 5450 1370 5470 1390
rect 5530 1370 5550 1390
rect 5610 1370 5630 1390
rect 5690 1370 5710 1390
rect 5770 1370 5790 1390
rect 5850 1370 5870 1390
rect 5930 1370 5950 1390
rect 6010 1370 6030 1390
rect 6090 1370 6110 1390
rect 6170 1370 6190 1390
rect 4250 1290 4270 1310
rect 4330 1290 4350 1310
rect 4410 1290 4430 1310
rect 4490 1290 4510 1310
rect 4570 1290 4590 1310
rect 4650 1290 4670 1310
rect 4730 1290 4750 1310
rect 4810 1290 4830 1310
rect 4890 1290 4910 1310
rect 4970 1290 4990 1310
rect 5050 1290 5070 1310
rect 5130 1290 5150 1310
rect 5210 1290 5230 1310
rect 5290 1290 5310 1310
rect 5370 1290 5390 1310
rect 5450 1290 5470 1310
rect 5530 1290 5550 1310
rect 5610 1290 5630 1310
rect 5690 1290 5710 1310
rect 5770 1290 5790 1310
rect 5850 1290 5870 1310
rect 5930 1290 5950 1310
rect 6010 1290 6030 1310
rect 6090 1290 6110 1310
rect 6170 1290 6190 1310
rect 4250 1210 4270 1230
rect 4330 1210 4350 1230
rect 4410 1210 4430 1230
rect 4490 1210 4510 1230
rect 4570 1210 4590 1230
rect 4650 1210 4670 1230
rect 4730 1210 4750 1230
rect 4810 1210 4830 1230
rect 4890 1210 4910 1230
rect 4970 1210 4990 1230
rect 5050 1210 5070 1230
rect 5130 1210 5150 1230
rect 5210 1210 5230 1230
rect 5290 1210 5310 1230
rect 5370 1210 5390 1230
rect 5450 1210 5470 1230
rect 5530 1210 5550 1230
rect 5610 1210 5630 1230
rect 5690 1210 5710 1230
rect 5770 1210 5790 1230
rect 5850 1210 5870 1230
rect 5930 1210 5950 1230
rect 6010 1210 6030 1230
rect 6090 1210 6110 1230
rect 6170 1210 6190 1230
rect 4250 1130 4270 1150
rect 4330 1130 4350 1150
rect 4410 1130 4430 1150
rect 4490 1130 4510 1150
rect 4570 1130 4590 1150
rect 4650 1130 4670 1150
rect 4730 1130 4750 1150
rect 4810 1130 4830 1150
rect 4890 1130 4910 1150
rect 4970 1130 4990 1150
rect 5050 1130 5070 1150
rect 5130 1130 5150 1150
rect 5210 1130 5230 1150
rect 5290 1130 5310 1150
rect 5370 1130 5390 1150
rect 5450 1130 5470 1150
rect 5530 1130 5550 1150
rect 5610 1130 5630 1150
rect 5690 1130 5710 1150
rect 5770 1130 5790 1150
rect 5850 1130 5870 1150
rect 5930 1130 5950 1150
rect 6010 1130 6030 1150
rect 6090 1130 6110 1150
rect 6170 1130 6190 1150
rect 4250 1050 4270 1070
rect 4330 1050 4350 1070
rect 4410 1050 4430 1070
rect 4490 1050 4510 1070
rect 4570 1050 4590 1070
rect 4650 1050 4670 1070
rect 4730 1050 4750 1070
rect 4810 1050 4830 1070
rect 4890 1050 4910 1070
rect 4970 1050 4990 1070
rect 5050 1050 5070 1070
rect 5130 1050 5150 1070
rect 5210 1050 5230 1070
rect 5290 1050 5310 1070
rect 5370 1050 5390 1070
rect 5450 1050 5470 1070
rect 5530 1050 5550 1070
rect 5610 1050 5630 1070
rect 5690 1050 5710 1070
rect 5770 1050 5790 1070
rect 5850 1050 5870 1070
rect 5930 1050 5950 1070
rect 6010 1050 6030 1070
rect 6090 1050 6110 1070
rect 6170 1050 6190 1070
rect 4250 970 4270 990
rect 4330 970 4350 990
rect 4410 970 4430 990
rect 4490 970 4510 990
rect 4570 970 4590 990
rect 4650 970 4670 990
rect 4730 970 4750 990
rect 4810 970 4830 990
rect 4890 970 4910 990
rect 4970 970 4990 990
rect 5050 970 5070 990
rect 5130 970 5150 990
rect 5210 970 5230 990
rect 5290 970 5310 990
rect 5370 970 5390 990
rect 5450 970 5470 990
rect 5530 970 5550 990
rect 5610 970 5630 990
rect 5690 970 5710 990
rect 5770 970 5790 990
rect 5850 970 5870 990
rect 5930 970 5950 990
rect 6010 970 6030 990
rect 6090 970 6110 990
rect 6170 970 6190 990
rect 4250 890 4270 910
rect 4330 890 4350 910
rect 4410 890 4430 910
rect 4490 890 4510 910
rect 4570 890 4590 910
rect 4650 890 4670 910
rect 4730 890 4750 910
rect 4810 890 4830 910
rect 4890 890 4910 910
rect 4970 890 4990 910
rect 5050 890 5070 910
rect 5130 890 5150 910
rect 5210 890 5230 910
rect 5290 890 5310 910
rect 5370 890 5390 910
rect 5450 890 5470 910
rect 5530 890 5550 910
rect 5610 890 5630 910
rect 5690 890 5710 910
rect 5770 890 5790 910
rect 5850 890 5870 910
rect 5930 890 5950 910
rect 6010 890 6030 910
rect 6090 890 6110 910
rect 6170 890 6190 910
rect 4250 810 4270 830
rect 4330 810 4350 830
rect 4410 810 4430 830
rect 4490 810 4510 830
rect 4570 810 4590 830
rect 4650 810 4670 830
rect 4730 810 4750 830
rect 4810 810 4830 830
rect 4890 810 4910 830
rect 4970 810 4990 830
rect 5050 810 5070 830
rect 5130 810 5150 830
rect 5210 810 5230 830
rect 5290 810 5310 830
rect 5370 810 5390 830
rect 5450 810 5470 830
rect 5530 810 5550 830
rect 5610 810 5630 830
rect 5690 810 5710 830
rect 5770 810 5790 830
rect 5850 810 5870 830
rect 5930 810 5950 830
rect 6010 810 6030 830
rect 6090 810 6110 830
rect 6170 810 6190 830
rect 4250 730 4270 750
rect 4330 730 4350 750
rect 4410 730 4430 750
rect 4490 730 4510 750
rect 4570 730 4590 750
rect 4650 730 4670 750
rect 4730 730 4750 750
rect 4810 730 4830 750
rect 4890 730 4910 750
rect 4970 730 4990 750
rect 5050 730 5070 750
rect 5130 730 5150 750
rect 5210 730 5230 750
rect 5290 730 5310 750
rect 5370 730 5390 750
rect 5450 730 5470 750
rect 5530 730 5550 750
rect 5610 730 5630 750
rect 5690 730 5710 750
rect 5770 730 5790 750
rect 5850 730 5870 750
rect 5930 730 5950 750
rect 6010 730 6030 750
rect 6090 730 6110 750
rect 6170 730 6190 750
rect 4250 650 4270 670
rect 4330 650 4350 670
rect 4410 650 4430 670
rect 4490 650 4510 670
rect 4570 650 4590 670
rect 4650 650 4670 670
rect 4730 650 4750 670
rect 4810 650 4830 670
rect 4890 650 4910 670
rect 4970 650 4990 670
rect 5050 650 5070 670
rect 5130 650 5150 670
rect 5210 650 5230 670
rect 5290 650 5310 670
rect 5370 650 5390 670
rect 5450 650 5470 670
rect 5530 650 5550 670
rect 5610 650 5630 670
rect 5690 650 5710 670
rect 5770 650 5790 670
rect 5850 650 5870 670
rect 5930 650 5950 670
rect 6010 650 6030 670
rect 6090 650 6110 670
rect 6170 650 6190 670
rect 4250 570 4270 590
rect 4330 570 4350 590
rect 4410 570 4430 590
rect 4490 570 4510 590
rect 4570 570 4590 590
rect 4650 570 4670 590
rect 4730 570 4750 590
rect 4810 570 4830 590
rect 4890 570 4910 590
rect 4970 570 4990 590
rect 5050 570 5070 590
rect 5130 570 5150 590
rect 5210 570 5230 590
rect 5290 570 5310 590
rect 5370 570 5390 590
rect 5450 570 5470 590
rect 5530 570 5550 590
rect 5610 570 5630 590
rect 5690 570 5710 590
rect 5770 570 5790 590
rect 5850 570 5870 590
rect 5930 570 5950 590
rect 6010 570 6030 590
rect 6090 570 6110 590
rect 6170 570 6190 590
rect 4250 490 4270 510
rect 4330 490 4350 510
rect 4410 490 4430 510
rect 4490 490 4510 510
rect 4570 490 4590 510
rect 4650 490 4670 510
rect 4730 490 4750 510
rect 4810 490 4830 510
rect 4890 490 4910 510
rect 4970 490 4990 510
rect 5050 490 5070 510
rect 5130 490 5150 510
rect 5210 490 5230 510
rect 5290 490 5310 510
rect 5370 490 5390 510
rect 5450 490 5470 510
rect 5530 490 5550 510
rect 5610 490 5630 510
rect 5690 490 5710 510
rect 5770 490 5790 510
rect 5850 490 5870 510
rect 5930 490 5950 510
rect 6010 490 6030 510
rect 6090 490 6110 510
rect 6170 490 6190 510
rect 4250 410 4270 430
rect 4330 410 4350 430
rect 4410 410 4430 430
rect 4490 410 4510 430
rect 4570 410 4590 430
rect 4650 410 4670 430
rect 4730 410 4750 430
rect 4810 410 4830 430
rect 4890 410 4910 430
rect 4970 410 4990 430
rect 5050 410 5070 430
rect 5130 410 5150 430
rect 5210 410 5230 430
rect 5290 410 5310 430
rect 5370 410 5390 430
rect 5450 410 5470 430
rect 5530 410 5550 430
rect 5610 410 5630 430
rect 5690 410 5710 430
rect 5770 410 5790 430
rect 5850 410 5870 430
rect 5930 410 5950 430
rect 6010 410 6030 430
rect 6090 410 6110 430
rect 6170 410 6190 430
rect 4250 330 4270 350
rect 4330 330 4350 350
rect 4410 330 4430 350
rect 4490 330 4510 350
rect 4570 330 4590 350
rect 4650 330 4670 350
rect 4730 330 4750 350
rect 4810 330 4830 350
rect 4890 330 4910 350
rect 4970 330 4990 350
rect 5050 330 5070 350
rect 5130 330 5150 350
rect 5210 330 5230 350
rect 5290 330 5310 350
rect 5370 330 5390 350
rect 5450 330 5470 350
rect 5530 330 5550 350
rect 5610 330 5630 350
rect 5690 330 5710 350
rect 5770 330 5790 350
rect 5850 330 5870 350
rect 5930 330 5950 350
rect 6010 330 6030 350
rect 6090 330 6110 350
rect 6170 330 6190 350
rect 4250 250 4270 270
rect 4330 250 4350 270
rect 4410 250 4430 270
rect 4490 250 4510 270
rect 4570 250 4590 270
rect 4650 250 4670 270
rect 4730 250 4750 270
rect 4810 250 4830 270
rect 4890 250 4910 270
rect 4970 250 4990 270
rect 5050 250 5070 270
rect 5130 250 5150 270
rect 5210 250 5230 270
rect 5290 250 5310 270
rect 5370 250 5390 270
rect 5450 250 5470 270
rect 5530 250 5550 270
rect 5610 250 5630 270
rect 5690 250 5710 270
rect 5770 250 5790 270
rect 5850 250 5870 270
rect 5930 250 5950 270
rect 6010 250 6030 270
rect 6090 250 6110 270
rect 6170 250 6190 270
rect 4250 170 4270 190
rect 4330 170 4350 190
rect 4410 170 4430 190
rect 4490 170 4510 190
rect 4570 170 4590 190
rect 4650 170 4670 190
rect 4730 170 4750 190
rect 4810 170 4830 190
rect 4890 170 4910 190
rect 4970 170 4990 190
rect 5050 170 5070 190
rect 5130 170 5150 190
rect 5210 170 5230 190
rect 5290 170 5310 190
rect 5370 170 5390 190
rect 5450 170 5470 190
rect 5530 170 5550 190
rect 5610 170 5630 190
rect 5690 170 5710 190
rect 5770 170 5790 190
rect 5850 170 5870 190
rect 5930 170 5950 190
rect 6010 170 6030 190
rect 6090 170 6110 190
rect 6170 170 6190 190
rect 4250 90 4270 110
rect 4330 90 4350 110
rect 4410 90 4430 110
rect 4490 90 4510 110
rect 4570 90 4590 110
rect 4650 90 4670 110
rect 4730 90 4750 110
rect 4810 90 4830 110
rect 4890 90 4910 110
rect 4970 90 4990 110
rect 5050 90 5070 110
rect 5130 90 5150 110
rect 5210 90 5230 110
rect 5290 90 5310 110
rect 5370 90 5390 110
rect 5450 90 5470 110
rect 5530 90 5550 110
rect 5610 90 5630 110
rect 5690 90 5710 110
rect 5770 90 5790 110
rect 5850 90 5870 110
rect 5930 90 5950 110
rect 6010 90 6030 110
rect 6090 90 6110 110
rect 6170 90 6190 110
rect 4250 10 4270 30
rect 4330 10 4350 30
rect 4410 10 4430 30
rect 4490 10 4510 30
rect 4570 10 4590 30
rect 4650 10 4670 30
rect 4730 10 4750 30
rect 4810 10 4830 30
rect 4890 10 4910 30
rect 4970 10 4990 30
rect 5050 10 5070 30
rect 5130 10 5150 30
rect 5210 10 5230 30
rect 5290 10 5310 30
rect 5370 10 5390 30
rect 5450 10 5470 30
rect 5530 10 5550 30
rect 5610 10 5630 30
rect 5690 10 5710 30
rect 5770 10 5790 30
rect 5850 10 5870 30
rect 5930 10 5950 30
rect 6010 10 6030 30
rect 6090 10 6110 30
rect 6170 10 6190 30
<< metal1 >>
rect 4240 15715 4280 15720
rect 4240 15685 4245 15715
rect 4275 15685 4280 15715
rect 4240 15635 4280 15685
rect 4240 15605 4245 15635
rect 4275 15605 4280 15635
rect 4240 15555 4280 15605
rect 4240 15525 4245 15555
rect 4275 15525 4280 15555
rect 4240 15475 4280 15525
rect 4240 15445 4245 15475
rect 4275 15445 4280 15475
rect 4240 15395 4280 15445
rect 4240 15365 4245 15395
rect 4275 15365 4280 15395
rect 4240 15315 4280 15365
rect 4240 15285 4245 15315
rect 4275 15285 4280 15315
rect 4240 15235 4280 15285
rect 4240 15205 4245 15235
rect 4275 15205 4280 15235
rect 4240 15155 4280 15205
rect 4240 15125 4245 15155
rect 4275 15125 4280 15155
rect 4240 15070 4280 15125
rect 4240 15050 4250 15070
rect 4270 15050 4280 15070
rect 4240 14995 4280 15050
rect 4240 14965 4245 14995
rect 4275 14965 4280 14995
rect 4240 14915 4280 14965
rect 4240 14885 4245 14915
rect 4275 14885 4280 14915
rect 4240 14835 4280 14885
rect 4240 14805 4245 14835
rect 4275 14805 4280 14835
rect 4240 14755 4280 14805
rect 4240 14725 4245 14755
rect 4275 14725 4280 14755
rect 4240 14675 4280 14725
rect 4240 14645 4245 14675
rect 4275 14645 4280 14675
rect 4240 14595 4280 14645
rect 4240 14565 4245 14595
rect 4275 14565 4280 14595
rect 4240 14515 4280 14565
rect 4240 14485 4245 14515
rect 4275 14485 4280 14515
rect 4240 14435 4280 14485
rect 4240 14405 4245 14435
rect 4275 14405 4280 14435
rect 4240 14350 4280 14405
rect 4240 14330 4250 14350
rect 4270 14330 4280 14350
rect 4240 14270 4280 14330
rect 4240 14250 4250 14270
rect 4270 14250 4280 14270
rect 4240 14190 4280 14250
rect 4240 14170 4250 14190
rect 4270 14170 4280 14190
rect 4240 14110 4280 14170
rect 4240 14090 4250 14110
rect 4270 14090 4280 14110
rect 4240 14035 4280 14090
rect 4240 14005 4245 14035
rect 4275 14005 4280 14035
rect 4240 13955 4280 14005
rect 4240 13925 4245 13955
rect 4275 13925 4280 13955
rect 4240 13875 4280 13925
rect 4240 13845 4245 13875
rect 4275 13845 4280 13875
rect 4240 13795 4280 13845
rect 4240 13765 4245 13795
rect 4275 13765 4280 13795
rect 4240 13715 4280 13765
rect 4240 13685 4245 13715
rect 4275 13685 4280 13715
rect 4240 13635 4280 13685
rect 4240 13605 4245 13635
rect 4275 13605 4280 13635
rect 4240 13555 4280 13605
rect 4240 13525 4245 13555
rect 4275 13525 4280 13555
rect 4240 13475 4280 13525
rect 4240 13445 4245 13475
rect 4275 13445 4280 13475
rect 4240 13390 4280 13445
rect 4240 13370 4250 13390
rect 4270 13370 4280 13390
rect 4240 13310 4280 13370
rect 4240 13290 4250 13310
rect 4270 13290 4280 13310
rect 4240 13230 4280 13290
rect 4240 13210 4250 13230
rect 4270 13210 4280 13230
rect 4240 13150 4280 13210
rect 4240 13130 4250 13150
rect 4270 13130 4280 13150
rect 4240 13075 4280 13130
rect 4240 13045 4245 13075
rect 4275 13045 4280 13075
rect 4240 12995 4280 13045
rect 4240 12965 4245 12995
rect 4275 12965 4280 12995
rect 4240 12915 4280 12965
rect 4240 12885 4245 12915
rect 4275 12885 4280 12915
rect 4240 12835 4280 12885
rect 4240 12805 4245 12835
rect 4275 12805 4280 12835
rect 4240 12755 4280 12805
rect 4240 12725 4245 12755
rect 4275 12725 4280 12755
rect 4240 12675 4280 12725
rect 4240 12645 4245 12675
rect 4275 12645 4280 12675
rect 4240 12595 4280 12645
rect 4240 12565 4245 12595
rect 4275 12565 4280 12595
rect 4240 12515 4280 12565
rect 4240 12485 4245 12515
rect 4275 12485 4280 12515
rect 4240 12430 4280 12485
rect 4240 12410 4250 12430
rect 4270 12410 4280 12430
rect 4240 12355 4280 12410
rect 4240 12325 4245 12355
rect 4275 12325 4280 12355
rect 4240 12275 4280 12325
rect 4240 12245 4245 12275
rect 4275 12245 4280 12275
rect 4240 12195 4280 12245
rect 4240 12165 4245 12195
rect 4275 12165 4280 12195
rect 4240 12115 4280 12165
rect 4240 12085 4245 12115
rect 4275 12085 4280 12115
rect 4240 12035 4280 12085
rect 4240 12005 4245 12035
rect 4275 12005 4280 12035
rect 4240 11955 4280 12005
rect 4240 11925 4245 11955
rect 4275 11925 4280 11955
rect 4240 11875 4280 11925
rect 4240 11845 4245 11875
rect 4275 11845 4280 11875
rect 4240 11795 4280 11845
rect 4240 11765 4245 11795
rect 4275 11765 4280 11795
rect 4240 11715 4280 11765
rect 4240 11685 4245 11715
rect 4275 11685 4280 11715
rect 4240 11635 4280 11685
rect 4240 11605 4245 11635
rect 4275 11605 4280 11635
rect 4240 11555 4280 11605
rect 4240 11525 4245 11555
rect 4275 11525 4280 11555
rect 4240 11475 4280 11525
rect 4240 11445 4245 11475
rect 4275 11445 4280 11475
rect 4240 11395 4280 11445
rect 4240 11365 4245 11395
rect 4275 11365 4280 11395
rect 4240 11315 4280 11365
rect 4240 11285 4245 11315
rect 4275 11285 4280 11315
rect 4240 11235 4280 11285
rect 4240 11205 4245 11235
rect 4275 11205 4280 11235
rect 4240 11155 4280 11205
rect 4240 11125 4245 11155
rect 4275 11125 4280 11155
rect 4240 11075 4280 11125
rect 4240 11045 4245 11075
rect 4275 11045 4280 11075
rect 4240 10990 4280 11045
rect 4240 10970 4250 10990
rect 4270 10970 4280 10990
rect 4240 10915 4280 10970
rect 4240 10885 4245 10915
rect 4275 10885 4280 10915
rect 4240 10835 4280 10885
rect 4240 10805 4245 10835
rect 4275 10805 4280 10835
rect 4240 10755 4280 10805
rect 4240 10725 4245 10755
rect 4275 10725 4280 10755
rect 4240 10675 4280 10725
rect 4240 10645 4245 10675
rect 4275 10645 4280 10675
rect 4240 10595 4280 10645
rect 4240 10565 4245 10595
rect 4275 10565 4280 10595
rect 4240 10515 4280 10565
rect 4240 10485 4245 10515
rect 4275 10485 4280 10515
rect 4240 10435 4280 10485
rect 4240 10405 4245 10435
rect 4275 10405 4280 10435
rect 4240 10355 4280 10405
rect 4240 10325 4245 10355
rect 4275 10325 4280 10355
rect 4240 10270 4280 10325
rect 4240 10250 4250 10270
rect 4270 10250 4280 10270
rect 4240 10190 4280 10250
rect 4240 10170 4250 10190
rect 4270 10170 4280 10190
rect 4240 10110 4280 10170
rect 4240 10090 4250 10110
rect 4270 10090 4280 10110
rect 4240 10030 4280 10090
rect 4240 10010 4250 10030
rect 4270 10010 4280 10030
rect 4240 9955 4280 10010
rect 4240 9925 4245 9955
rect 4275 9925 4280 9955
rect 4240 9875 4280 9925
rect 4240 9845 4245 9875
rect 4275 9845 4280 9875
rect 4240 9795 4280 9845
rect 4240 9765 4245 9795
rect 4275 9765 4280 9795
rect 4240 9715 4280 9765
rect 4240 9685 4245 9715
rect 4275 9685 4280 9715
rect 4240 9635 4280 9685
rect 4240 9605 4245 9635
rect 4275 9605 4280 9635
rect 4240 9555 4280 9605
rect 4240 9525 4245 9555
rect 4275 9525 4280 9555
rect 4240 9475 4280 9525
rect 4240 9445 4245 9475
rect 4275 9445 4280 9475
rect 4240 9395 4280 9445
rect 4240 9365 4245 9395
rect 4275 9365 4280 9395
rect 4240 9310 4280 9365
rect 4240 9290 4250 9310
rect 4270 9290 4280 9310
rect 4240 9230 4280 9290
rect 4240 9210 4250 9230
rect 4270 9210 4280 9230
rect 4240 9150 4280 9210
rect 4240 9130 4250 9150
rect 4270 9130 4280 9150
rect 4240 9070 4280 9130
rect 4240 9050 4250 9070
rect 4270 9050 4280 9070
rect 4240 8995 4280 9050
rect 4240 8965 4245 8995
rect 4275 8965 4280 8995
rect 4240 8915 4280 8965
rect 4240 8885 4245 8915
rect 4275 8885 4280 8915
rect 4240 8835 4280 8885
rect 4240 8805 4245 8835
rect 4275 8805 4280 8835
rect 4240 8755 4280 8805
rect 4240 8725 4245 8755
rect 4275 8725 4280 8755
rect 4240 8675 4280 8725
rect 4240 8645 4245 8675
rect 4275 8645 4280 8675
rect 4240 8595 4280 8645
rect 4240 8565 4245 8595
rect 4275 8565 4280 8595
rect 4240 8515 4280 8565
rect 4240 8485 4245 8515
rect 4275 8485 4280 8515
rect 4240 8435 4280 8485
rect 4240 8405 4245 8435
rect 4275 8405 4280 8435
rect 4240 8350 4280 8405
rect 4240 8330 4250 8350
rect 4270 8330 4280 8350
rect 4240 8275 4280 8330
rect 4240 8245 4245 8275
rect 4275 8245 4280 8275
rect 4240 8195 4280 8245
rect 4240 8165 4245 8195
rect 4275 8165 4280 8195
rect 4240 8115 4280 8165
rect 4240 8085 4245 8115
rect 4275 8085 4280 8115
rect 4240 8035 4280 8085
rect 4240 8005 4245 8035
rect 4275 8005 4280 8035
rect 4240 7955 4280 8005
rect 4240 7925 4245 7955
rect 4275 7925 4280 7955
rect 4240 7875 4280 7925
rect 4240 7845 4245 7875
rect 4275 7845 4280 7875
rect 4240 7795 4280 7845
rect 4240 7765 4245 7795
rect 4275 7765 4280 7795
rect 4240 7715 4280 7765
rect 4240 7685 4245 7715
rect 4275 7685 4280 7715
rect 4240 7635 4280 7685
rect 4240 7605 4245 7635
rect 4275 7605 4280 7635
rect 4240 7555 4280 7605
rect 4240 7525 4245 7555
rect 4275 7525 4280 7555
rect 4240 7475 4280 7525
rect 4240 7445 4245 7475
rect 4275 7445 4280 7475
rect 4240 7395 4280 7445
rect 4240 7365 4245 7395
rect 4275 7365 4280 7395
rect 4240 7315 4280 7365
rect 4240 7285 4245 7315
rect 4275 7285 4280 7315
rect 4240 7235 4280 7285
rect 4240 7205 4245 7235
rect 4275 7205 4280 7235
rect 4240 7155 4280 7205
rect 4240 7125 4245 7155
rect 4275 7125 4280 7155
rect 4240 7075 4280 7125
rect 4240 7045 4245 7075
rect 4275 7045 4280 7075
rect 4240 6995 4280 7045
rect 4240 6965 4245 6995
rect 4275 6965 4280 6995
rect 4240 6910 4280 6965
rect 4240 6890 4250 6910
rect 4270 6890 4280 6910
rect 4240 6835 4280 6890
rect 4240 6805 4245 6835
rect 4275 6805 4280 6835
rect 4240 6755 4280 6805
rect 4240 6725 4245 6755
rect 4275 6725 4280 6755
rect 4240 6675 4280 6725
rect 4240 6645 4245 6675
rect 4275 6645 4280 6675
rect 4240 6595 4280 6645
rect 4240 6565 4245 6595
rect 4275 6565 4280 6595
rect 4240 6515 4280 6565
rect 4240 6485 4245 6515
rect 4275 6485 4280 6515
rect 4240 6435 4280 6485
rect 4240 6405 4245 6435
rect 4275 6405 4280 6435
rect 4240 6355 4280 6405
rect 4240 6325 4245 6355
rect 4275 6325 4280 6355
rect 4240 6275 4280 6325
rect 4240 6245 4245 6275
rect 4275 6245 4280 6275
rect 4240 6190 4280 6245
rect 4240 6170 4250 6190
rect 4270 6170 4280 6190
rect 4240 6110 4280 6170
rect 4240 6090 4250 6110
rect 4270 6090 4280 6110
rect 4240 6030 4280 6090
rect 4240 6010 4250 6030
rect 4270 6010 4280 6030
rect 4240 5950 4280 6010
rect 4240 5930 4250 5950
rect 4270 5930 4280 5950
rect 4240 5875 4280 5930
rect 4240 5845 4245 5875
rect 4275 5845 4280 5875
rect 4240 5795 4280 5845
rect 4240 5765 4245 5795
rect 4275 5765 4280 5795
rect 4240 5715 4280 5765
rect 4240 5685 4245 5715
rect 4275 5685 4280 5715
rect 4240 5635 4280 5685
rect 4240 5605 4245 5635
rect 4275 5605 4280 5635
rect 4240 5555 4280 5605
rect 4240 5525 4245 5555
rect 4275 5525 4280 5555
rect 4240 5475 4280 5525
rect 4240 5445 4245 5475
rect 4275 5445 4280 5475
rect 4240 5395 4280 5445
rect 4240 5365 4245 5395
rect 4275 5365 4280 5395
rect 4240 5315 4280 5365
rect 4240 5285 4245 5315
rect 4275 5285 4280 5315
rect 4240 5235 4280 5285
rect 4240 5205 4245 5235
rect 4275 5205 4280 5235
rect 4240 5155 4280 5205
rect 4240 5125 4245 5155
rect 4275 5125 4280 5155
rect 4240 5075 4280 5125
rect 4240 5045 4245 5075
rect 4275 5045 4280 5075
rect 4240 4995 4280 5045
rect 4240 4965 4245 4995
rect 4275 4965 4280 4995
rect 4240 4915 4280 4965
rect 4240 4885 4245 4915
rect 4275 4885 4280 4915
rect 4240 4830 4280 4885
rect 4240 4810 4250 4830
rect 4270 4810 4280 4830
rect 4240 4755 4280 4810
rect 4240 4725 4245 4755
rect 4275 4725 4280 4755
rect 4240 4675 4280 4725
rect 4240 4645 4245 4675
rect 4275 4645 4280 4675
rect 4240 4590 4280 4645
rect 4240 4570 4250 4590
rect 4270 4570 4280 4590
rect 4240 4515 4280 4570
rect 4240 4485 4245 4515
rect 4275 4485 4280 4515
rect 4240 4435 4280 4485
rect 4240 4405 4245 4435
rect 4275 4405 4280 4435
rect 4240 4355 4280 4405
rect 4240 4325 4245 4355
rect 4275 4325 4280 4355
rect 4240 4275 4280 4325
rect 4240 4245 4245 4275
rect 4275 4245 4280 4275
rect 4240 4195 4280 4245
rect 4240 4165 4245 4195
rect 4275 4165 4280 4195
rect 4240 4115 4280 4165
rect 4240 4085 4245 4115
rect 4275 4085 4280 4115
rect 4240 4035 4280 4085
rect 4240 4005 4245 4035
rect 4275 4005 4280 4035
rect 4240 3955 4280 4005
rect 4240 3925 4245 3955
rect 4275 3925 4280 3955
rect 4240 3875 4280 3925
rect 4240 3845 4245 3875
rect 4275 3845 4280 3875
rect 4240 3790 4280 3845
rect 4240 3770 4250 3790
rect 4270 3770 4280 3790
rect 4240 3715 4280 3770
rect 4240 3685 4245 3715
rect 4275 3685 4280 3715
rect 4240 3635 4280 3685
rect 4240 3605 4245 3635
rect 4275 3605 4280 3635
rect 4240 3550 4280 3605
rect 4240 3530 4250 3550
rect 4270 3530 4280 3550
rect 4240 3475 4280 3530
rect 4240 3445 4245 3475
rect 4275 3445 4280 3475
rect 4240 3395 4280 3445
rect 4240 3365 4245 3395
rect 4275 3365 4280 3395
rect 4240 3310 4280 3365
rect 4240 3290 4250 3310
rect 4270 3290 4280 3310
rect 4240 3235 4280 3290
rect 4240 3205 4245 3235
rect 4275 3205 4280 3235
rect 4240 3155 4280 3205
rect 4240 3125 4245 3155
rect 4275 3125 4280 3155
rect 4240 3075 4280 3125
rect 4240 3045 4245 3075
rect 4275 3045 4280 3075
rect 4240 2995 4280 3045
rect 4240 2965 4245 2995
rect 4275 2965 4280 2995
rect 4240 2915 4280 2965
rect 4240 2885 4245 2915
rect 4275 2885 4280 2915
rect 4240 2835 4280 2885
rect 4240 2805 4245 2835
rect 4275 2805 4280 2835
rect 4240 2755 4280 2805
rect 4240 2725 4245 2755
rect 4275 2725 4280 2755
rect 4240 2675 4280 2725
rect 4240 2645 4245 2675
rect 4275 2645 4280 2675
rect 4240 2595 4280 2645
rect 4240 2565 4245 2595
rect 4275 2565 4280 2595
rect 4240 2515 4280 2565
rect 4240 2485 4245 2515
rect 4275 2485 4280 2515
rect 4240 2435 4280 2485
rect 4240 2405 4245 2435
rect 4275 2405 4280 2435
rect 4240 2355 4280 2405
rect 4240 2325 4245 2355
rect 4275 2325 4280 2355
rect 4240 2275 4280 2325
rect 4240 2245 4245 2275
rect 4275 2245 4280 2275
rect 4240 2195 4280 2245
rect 4240 2165 4245 2195
rect 4275 2165 4280 2195
rect 4240 2115 4280 2165
rect 4240 2085 4245 2115
rect 4275 2085 4280 2115
rect 4240 2035 4280 2085
rect 4240 2005 4245 2035
rect 4275 2005 4280 2035
rect 4240 1955 4280 2005
rect 4240 1925 4245 1955
rect 4275 1925 4280 1955
rect 4240 1870 4280 1925
rect 4240 1850 4250 1870
rect 4270 1850 4280 1870
rect 4240 1790 4280 1850
rect 4240 1770 4250 1790
rect 4270 1770 4280 1790
rect 4240 1715 4280 1770
rect 4240 1685 4245 1715
rect 4275 1685 4280 1715
rect 4240 1635 4280 1685
rect 4240 1605 4245 1635
rect 4275 1605 4280 1635
rect 4240 1555 4280 1605
rect 4240 1525 4245 1555
rect 4275 1525 4280 1555
rect 4240 1475 4280 1525
rect 4240 1445 4245 1475
rect 4275 1445 4280 1475
rect 4240 1395 4280 1445
rect 4240 1365 4245 1395
rect 4275 1365 4280 1395
rect 4240 1315 4280 1365
rect 4240 1285 4245 1315
rect 4275 1285 4280 1315
rect 4240 1235 4280 1285
rect 4240 1205 4245 1235
rect 4275 1205 4280 1235
rect 4240 1155 4280 1205
rect 4240 1125 4245 1155
rect 4275 1125 4280 1155
rect 4240 1075 4280 1125
rect 4240 1045 4245 1075
rect 4275 1045 4280 1075
rect 4240 995 4280 1045
rect 4240 965 4245 995
rect 4275 965 4280 995
rect 4240 910 4280 965
rect 4240 890 4250 910
rect 4270 890 4280 910
rect 4240 835 4280 890
rect 4240 805 4245 835
rect 4275 805 4280 835
rect 4240 755 4280 805
rect 4240 725 4245 755
rect 4275 725 4280 755
rect 4240 675 4280 725
rect 4240 645 4245 675
rect 4275 645 4280 675
rect 4240 595 4280 645
rect 4240 565 4245 595
rect 4275 565 4280 595
rect 4240 515 4280 565
rect 4240 485 4245 515
rect 4275 485 4280 515
rect 4240 430 4280 485
rect 4240 410 4250 430
rect 4270 410 4280 430
rect 4240 350 4280 410
rect 4240 330 4250 350
rect 4270 330 4280 350
rect 4240 275 4280 330
rect 4240 245 4245 275
rect 4275 245 4280 275
rect 4240 195 4280 245
rect 4240 165 4245 195
rect 4275 165 4280 195
rect 4240 115 4280 165
rect 4240 85 4245 115
rect 4275 85 4280 115
rect 4240 35 4280 85
rect 4240 5 4245 35
rect 4275 5 4280 35
rect 4240 0 4280 5
rect 4320 15710 4360 15720
rect 4320 15690 4330 15710
rect 4350 15690 4360 15710
rect 4320 15630 4360 15690
rect 4320 15610 4330 15630
rect 4350 15610 4360 15630
rect 4320 15550 4360 15610
rect 4320 15530 4330 15550
rect 4350 15530 4360 15550
rect 4320 15470 4360 15530
rect 4320 15450 4330 15470
rect 4350 15450 4360 15470
rect 4320 15390 4360 15450
rect 4320 15370 4330 15390
rect 4350 15370 4360 15390
rect 4320 15310 4360 15370
rect 4320 15290 4330 15310
rect 4350 15290 4360 15310
rect 4320 15230 4360 15290
rect 4320 15210 4330 15230
rect 4350 15210 4360 15230
rect 4320 15150 4360 15210
rect 4320 15130 4330 15150
rect 4350 15130 4360 15150
rect 4320 15070 4360 15130
rect 4320 15050 4330 15070
rect 4350 15050 4360 15070
rect 4320 14990 4360 15050
rect 4320 14970 4330 14990
rect 4350 14970 4360 14990
rect 4320 14910 4360 14970
rect 4320 14890 4330 14910
rect 4350 14890 4360 14910
rect 4320 14830 4360 14890
rect 4320 14810 4330 14830
rect 4350 14810 4360 14830
rect 4320 14750 4360 14810
rect 4320 14730 4330 14750
rect 4350 14730 4360 14750
rect 4320 14670 4360 14730
rect 4320 14650 4330 14670
rect 4350 14650 4360 14670
rect 4320 14590 4360 14650
rect 4320 14570 4330 14590
rect 4350 14570 4360 14590
rect 4320 14510 4360 14570
rect 4320 14490 4330 14510
rect 4350 14490 4360 14510
rect 4320 14430 4360 14490
rect 4320 14410 4330 14430
rect 4350 14410 4360 14430
rect 4320 14350 4360 14410
rect 4320 14330 4330 14350
rect 4350 14330 4360 14350
rect 4320 14270 4360 14330
rect 4320 14250 4330 14270
rect 4350 14250 4360 14270
rect 4320 14190 4360 14250
rect 4320 14170 4330 14190
rect 4350 14170 4360 14190
rect 4320 14110 4360 14170
rect 4320 14090 4330 14110
rect 4350 14090 4360 14110
rect 4320 14030 4360 14090
rect 4320 14010 4330 14030
rect 4350 14010 4360 14030
rect 4320 13950 4360 14010
rect 4320 13930 4330 13950
rect 4350 13930 4360 13950
rect 4320 13870 4360 13930
rect 4320 13850 4330 13870
rect 4350 13850 4360 13870
rect 4320 13790 4360 13850
rect 4320 13770 4330 13790
rect 4350 13770 4360 13790
rect 4320 13710 4360 13770
rect 4320 13690 4330 13710
rect 4350 13690 4360 13710
rect 4320 13630 4360 13690
rect 4320 13610 4330 13630
rect 4350 13610 4360 13630
rect 4320 13550 4360 13610
rect 4320 13530 4330 13550
rect 4350 13530 4360 13550
rect 4320 13470 4360 13530
rect 4320 13450 4330 13470
rect 4350 13450 4360 13470
rect 4320 13390 4360 13450
rect 4320 13370 4330 13390
rect 4350 13370 4360 13390
rect 4320 13310 4360 13370
rect 4320 13290 4330 13310
rect 4350 13290 4360 13310
rect 4320 13230 4360 13290
rect 4320 13210 4330 13230
rect 4350 13210 4360 13230
rect 4320 13150 4360 13210
rect 4320 13130 4330 13150
rect 4350 13130 4360 13150
rect 4320 13070 4360 13130
rect 4320 13050 4330 13070
rect 4350 13050 4360 13070
rect 4320 12990 4360 13050
rect 4320 12970 4330 12990
rect 4350 12970 4360 12990
rect 4320 12910 4360 12970
rect 4320 12890 4330 12910
rect 4350 12890 4360 12910
rect 4320 12830 4360 12890
rect 4320 12810 4330 12830
rect 4350 12810 4360 12830
rect 4320 12750 4360 12810
rect 4320 12730 4330 12750
rect 4350 12730 4360 12750
rect 4320 12670 4360 12730
rect 4320 12650 4330 12670
rect 4350 12650 4360 12670
rect 4320 12590 4360 12650
rect 4320 12570 4330 12590
rect 4350 12570 4360 12590
rect 4320 12510 4360 12570
rect 4320 12490 4330 12510
rect 4350 12490 4360 12510
rect 4320 12430 4360 12490
rect 4320 12410 4330 12430
rect 4350 12410 4360 12430
rect 4320 12350 4360 12410
rect 4320 12330 4330 12350
rect 4350 12330 4360 12350
rect 4320 12270 4360 12330
rect 4320 12250 4330 12270
rect 4350 12250 4360 12270
rect 4320 12190 4360 12250
rect 4320 12170 4330 12190
rect 4350 12170 4360 12190
rect 4320 12110 4360 12170
rect 4320 12090 4330 12110
rect 4350 12090 4360 12110
rect 4320 12030 4360 12090
rect 4320 12010 4330 12030
rect 4350 12010 4360 12030
rect 4320 11950 4360 12010
rect 4320 11930 4330 11950
rect 4350 11930 4360 11950
rect 4320 11870 4360 11930
rect 4320 11850 4330 11870
rect 4350 11850 4360 11870
rect 4320 11790 4360 11850
rect 4320 11770 4330 11790
rect 4350 11770 4360 11790
rect 4320 11710 4360 11770
rect 4320 11690 4330 11710
rect 4350 11690 4360 11710
rect 4320 11630 4360 11690
rect 4320 11610 4330 11630
rect 4350 11610 4360 11630
rect 4320 11550 4360 11610
rect 4320 11530 4330 11550
rect 4350 11530 4360 11550
rect 4320 11470 4360 11530
rect 4320 11450 4330 11470
rect 4350 11450 4360 11470
rect 4320 11390 4360 11450
rect 4320 11370 4330 11390
rect 4350 11370 4360 11390
rect 4320 11310 4360 11370
rect 4320 11290 4330 11310
rect 4350 11290 4360 11310
rect 4320 11230 4360 11290
rect 4320 11210 4330 11230
rect 4350 11210 4360 11230
rect 4320 11150 4360 11210
rect 4320 11130 4330 11150
rect 4350 11130 4360 11150
rect 4320 11070 4360 11130
rect 4320 11050 4330 11070
rect 4350 11050 4360 11070
rect 4320 10990 4360 11050
rect 4320 10970 4330 10990
rect 4350 10970 4360 10990
rect 4320 10910 4360 10970
rect 4320 10890 4330 10910
rect 4350 10890 4360 10910
rect 4320 10830 4360 10890
rect 4320 10810 4330 10830
rect 4350 10810 4360 10830
rect 4320 10750 4360 10810
rect 4320 10730 4330 10750
rect 4350 10730 4360 10750
rect 4320 10670 4360 10730
rect 4320 10650 4330 10670
rect 4350 10650 4360 10670
rect 4320 10590 4360 10650
rect 4320 10570 4330 10590
rect 4350 10570 4360 10590
rect 4320 10510 4360 10570
rect 4320 10490 4330 10510
rect 4350 10490 4360 10510
rect 4320 10430 4360 10490
rect 4320 10410 4330 10430
rect 4350 10410 4360 10430
rect 4320 10350 4360 10410
rect 4320 10330 4330 10350
rect 4350 10330 4360 10350
rect 4320 10270 4360 10330
rect 4320 10250 4330 10270
rect 4350 10250 4360 10270
rect 4320 10190 4360 10250
rect 4320 10170 4330 10190
rect 4350 10170 4360 10190
rect 4320 10110 4360 10170
rect 4320 10090 4330 10110
rect 4350 10090 4360 10110
rect 4320 10030 4360 10090
rect 4320 10010 4330 10030
rect 4350 10010 4360 10030
rect 4320 9950 4360 10010
rect 4320 9930 4330 9950
rect 4350 9930 4360 9950
rect 4320 9870 4360 9930
rect 4320 9850 4330 9870
rect 4350 9850 4360 9870
rect 4320 9790 4360 9850
rect 4320 9770 4330 9790
rect 4350 9770 4360 9790
rect 4320 9710 4360 9770
rect 4320 9690 4330 9710
rect 4350 9690 4360 9710
rect 4320 9630 4360 9690
rect 4320 9610 4330 9630
rect 4350 9610 4360 9630
rect 4320 9550 4360 9610
rect 4320 9530 4330 9550
rect 4350 9530 4360 9550
rect 4320 9470 4360 9530
rect 4320 9450 4330 9470
rect 4350 9450 4360 9470
rect 4320 9390 4360 9450
rect 4320 9370 4330 9390
rect 4350 9370 4360 9390
rect 4320 9310 4360 9370
rect 4320 9290 4330 9310
rect 4350 9290 4360 9310
rect 4320 9230 4360 9290
rect 4320 9210 4330 9230
rect 4350 9210 4360 9230
rect 4320 9150 4360 9210
rect 4320 9130 4330 9150
rect 4350 9130 4360 9150
rect 4320 9070 4360 9130
rect 4320 9050 4330 9070
rect 4350 9050 4360 9070
rect 4320 8990 4360 9050
rect 4320 8970 4330 8990
rect 4350 8970 4360 8990
rect 4320 8910 4360 8970
rect 4320 8890 4330 8910
rect 4350 8890 4360 8910
rect 4320 8830 4360 8890
rect 4320 8810 4330 8830
rect 4350 8810 4360 8830
rect 4320 8750 4360 8810
rect 4320 8730 4330 8750
rect 4350 8730 4360 8750
rect 4320 8670 4360 8730
rect 4320 8650 4330 8670
rect 4350 8650 4360 8670
rect 4320 8590 4360 8650
rect 4320 8570 4330 8590
rect 4350 8570 4360 8590
rect 4320 8510 4360 8570
rect 4320 8490 4330 8510
rect 4350 8490 4360 8510
rect 4320 8430 4360 8490
rect 4320 8410 4330 8430
rect 4350 8410 4360 8430
rect 4320 8350 4360 8410
rect 4320 8330 4330 8350
rect 4350 8330 4360 8350
rect 4320 8270 4360 8330
rect 4320 8250 4330 8270
rect 4350 8250 4360 8270
rect 4320 8190 4360 8250
rect 4320 8170 4330 8190
rect 4350 8170 4360 8190
rect 4320 8110 4360 8170
rect 4320 8090 4330 8110
rect 4350 8090 4360 8110
rect 4320 8030 4360 8090
rect 4320 8010 4330 8030
rect 4350 8010 4360 8030
rect 4320 7950 4360 8010
rect 4320 7930 4330 7950
rect 4350 7930 4360 7950
rect 4320 7870 4360 7930
rect 4320 7850 4330 7870
rect 4350 7850 4360 7870
rect 4320 7790 4360 7850
rect 4320 7770 4330 7790
rect 4350 7770 4360 7790
rect 4320 7710 4360 7770
rect 4320 7690 4330 7710
rect 4350 7690 4360 7710
rect 4320 7630 4360 7690
rect 4320 7610 4330 7630
rect 4350 7610 4360 7630
rect 4320 7550 4360 7610
rect 4320 7530 4330 7550
rect 4350 7530 4360 7550
rect 4320 7470 4360 7530
rect 4320 7450 4330 7470
rect 4350 7450 4360 7470
rect 4320 7390 4360 7450
rect 4320 7370 4330 7390
rect 4350 7370 4360 7390
rect 4320 7310 4360 7370
rect 4320 7290 4330 7310
rect 4350 7290 4360 7310
rect 4320 7230 4360 7290
rect 4320 7210 4330 7230
rect 4350 7210 4360 7230
rect 4320 7150 4360 7210
rect 4320 7130 4330 7150
rect 4350 7130 4360 7150
rect 4320 7070 4360 7130
rect 4320 7050 4330 7070
rect 4350 7050 4360 7070
rect 4320 6990 4360 7050
rect 4320 6970 4330 6990
rect 4350 6970 4360 6990
rect 4320 6910 4360 6970
rect 4320 6890 4330 6910
rect 4350 6890 4360 6910
rect 4320 6830 4360 6890
rect 4320 6810 4330 6830
rect 4350 6810 4360 6830
rect 4320 6750 4360 6810
rect 4320 6730 4330 6750
rect 4350 6730 4360 6750
rect 4320 6670 4360 6730
rect 4320 6650 4330 6670
rect 4350 6650 4360 6670
rect 4320 6590 4360 6650
rect 4320 6570 4330 6590
rect 4350 6570 4360 6590
rect 4320 6510 4360 6570
rect 4320 6490 4330 6510
rect 4350 6490 4360 6510
rect 4320 6430 4360 6490
rect 4320 6410 4330 6430
rect 4350 6410 4360 6430
rect 4320 6350 4360 6410
rect 4320 6330 4330 6350
rect 4350 6330 4360 6350
rect 4320 6270 4360 6330
rect 4320 6250 4330 6270
rect 4350 6250 4360 6270
rect 4320 6190 4360 6250
rect 4320 6170 4330 6190
rect 4350 6170 4360 6190
rect 4320 6110 4360 6170
rect 4320 6090 4330 6110
rect 4350 6090 4360 6110
rect 4320 6030 4360 6090
rect 4320 6010 4330 6030
rect 4350 6010 4360 6030
rect 4320 5950 4360 6010
rect 4320 5930 4330 5950
rect 4350 5930 4360 5950
rect 4320 5870 4360 5930
rect 4320 5850 4330 5870
rect 4350 5850 4360 5870
rect 4320 5790 4360 5850
rect 4320 5770 4330 5790
rect 4350 5770 4360 5790
rect 4320 5710 4360 5770
rect 4320 5690 4330 5710
rect 4350 5690 4360 5710
rect 4320 5630 4360 5690
rect 4320 5610 4330 5630
rect 4350 5610 4360 5630
rect 4320 5550 4360 5610
rect 4320 5530 4330 5550
rect 4350 5530 4360 5550
rect 4320 5470 4360 5530
rect 4320 5450 4330 5470
rect 4350 5450 4360 5470
rect 4320 5390 4360 5450
rect 4320 5370 4330 5390
rect 4350 5370 4360 5390
rect 4320 5310 4360 5370
rect 4320 5290 4330 5310
rect 4350 5290 4360 5310
rect 4320 5230 4360 5290
rect 4320 5210 4330 5230
rect 4350 5210 4360 5230
rect 4320 5150 4360 5210
rect 4320 5130 4330 5150
rect 4350 5130 4360 5150
rect 4320 5070 4360 5130
rect 4320 5050 4330 5070
rect 4350 5050 4360 5070
rect 4320 4990 4360 5050
rect 4320 4970 4330 4990
rect 4350 4970 4360 4990
rect 4320 4910 4360 4970
rect 4320 4890 4330 4910
rect 4350 4890 4360 4910
rect 4320 4830 4360 4890
rect 4320 4810 4330 4830
rect 4350 4810 4360 4830
rect 4320 4750 4360 4810
rect 4320 4730 4330 4750
rect 4350 4730 4360 4750
rect 4320 4670 4360 4730
rect 4320 4650 4330 4670
rect 4350 4650 4360 4670
rect 4320 4590 4360 4650
rect 4320 4570 4330 4590
rect 4350 4570 4360 4590
rect 4320 4510 4360 4570
rect 4320 4490 4330 4510
rect 4350 4490 4360 4510
rect 4320 4430 4360 4490
rect 4320 4410 4330 4430
rect 4350 4410 4360 4430
rect 4320 4350 4360 4410
rect 4320 4330 4330 4350
rect 4350 4330 4360 4350
rect 4320 4270 4360 4330
rect 4320 4250 4330 4270
rect 4350 4250 4360 4270
rect 4320 4190 4360 4250
rect 4320 4170 4330 4190
rect 4350 4170 4360 4190
rect 4320 4110 4360 4170
rect 4320 4090 4330 4110
rect 4350 4090 4360 4110
rect 4320 4030 4360 4090
rect 4320 4010 4330 4030
rect 4350 4010 4360 4030
rect 4320 3950 4360 4010
rect 4320 3930 4330 3950
rect 4350 3930 4360 3950
rect 4320 3870 4360 3930
rect 4320 3850 4330 3870
rect 4350 3850 4360 3870
rect 4320 3790 4360 3850
rect 4320 3770 4330 3790
rect 4350 3770 4360 3790
rect 4320 3710 4360 3770
rect 4320 3690 4330 3710
rect 4350 3690 4360 3710
rect 4320 3630 4360 3690
rect 4320 3610 4330 3630
rect 4350 3610 4360 3630
rect 4320 3550 4360 3610
rect 4320 3530 4330 3550
rect 4350 3530 4360 3550
rect 4320 3470 4360 3530
rect 4320 3450 4330 3470
rect 4350 3450 4360 3470
rect 4320 3390 4360 3450
rect 4320 3370 4330 3390
rect 4350 3370 4360 3390
rect 4320 3310 4360 3370
rect 4320 3290 4330 3310
rect 4350 3290 4360 3310
rect 4320 3230 4360 3290
rect 4320 3210 4330 3230
rect 4350 3210 4360 3230
rect 4320 3150 4360 3210
rect 4320 3130 4330 3150
rect 4350 3130 4360 3150
rect 4320 3070 4360 3130
rect 4320 3050 4330 3070
rect 4350 3050 4360 3070
rect 4320 2990 4360 3050
rect 4320 2970 4330 2990
rect 4350 2970 4360 2990
rect 4320 2910 4360 2970
rect 4320 2890 4330 2910
rect 4350 2890 4360 2910
rect 4320 2830 4360 2890
rect 4320 2810 4330 2830
rect 4350 2810 4360 2830
rect 4320 2750 4360 2810
rect 4320 2730 4330 2750
rect 4350 2730 4360 2750
rect 4320 2670 4360 2730
rect 4320 2650 4330 2670
rect 4350 2650 4360 2670
rect 4320 2590 4360 2650
rect 4320 2570 4330 2590
rect 4350 2570 4360 2590
rect 4320 2510 4360 2570
rect 4320 2490 4330 2510
rect 4350 2490 4360 2510
rect 4320 2430 4360 2490
rect 4320 2410 4330 2430
rect 4350 2410 4360 2430
rect 4320 2350 4360 2410
rect 4320 2330 4330 2350
rect 4350 2330 4360 2350
rect 4320 2270 4360 2330
rect 4320 2250 4330 2270
rect 4350 2250 4360 2270
rect 4320 2190 4360 2250
rect 4320 2170 4330 2190
rect 4350 2170 4360 2190
rect 4320 2110 4360 2170
rect 4320 2090 4330 2110
rect 4350 2090 4360 2110
rect 4320 2030 4360 2090
rect 4320 2010 4330 2030
rect 4350 2010 4360 2030
rect 4320 1950 4360 2010
rect 4320 1930 4330 1950
rect 4350 1930 4360 1950
rect 4320 1870 4360 1930
rect 4320 1850 4330 1870
rect 4350 1850 4360 1870
rect 4320 1790 4360 1850
rect 4320 1770 4330 1790
rect 4350 1770 4360 1790
rect 4320 1710 4360 1770
rect 4320 1690 4330 1710
rect 4350 1690 4360 1710
rect 4320 1630 4360 1690
rect 4320 1610 4330 1630
rect 4350 1610 4360 1630
rect 4320 1550 4360 1610
rect 4320 1530 4330 1550
rect 4350 1530 4360 1550
rect 4320 1470 4360 1530
rect 4320 1450 4330 1470
rect 4350 1450 4360 1470
rect 4320 1390 4360 1450
rect 4320 1370 4330 1390
rect 4350 1370 4360 1390
rect 4320 1310 4360 1370
rect 4320 1290 4330 1310
rect 4350 1290 4360 1310
rect 4320 1230 4360 1290
rect 4320 1210 4330 1230
rect 4350 1210 4360 1230
rect 4320 1150 4360 1210
rect 4320 1130 4330 1150
rect 4350 1130 4360 1150
rect 4320 1070 4360 1130
rect 4320 1050 4330 1070
rect 4350 1050 4360 1070
rect 4320 990 4360 1050
rect 4320 970 4330 990
rect 4350 970 4360 990
rect 4320 910 4360 970
rect 4320 890 4330 910
rect 4350 890 4360 910
rect 4320 830 4360 890
rect 4320 810 4330 830
rect 4350 810 4360 830
rect 4320 750 4360 810
rect 4320 730 4330 750
rect 4350 730 4360 750
rect 4320 670 4360 730
rect 4320 650 4330 670
rect 4350 650 4360 670
rect 4320 590 4360 650
rect 4320 570 4330 590
rect 4350 570 4360 590
rect 4320 510 4360 570
rect 4320 490 4330 510
rect 4350 490 4360 510
rect 4320 430 4360 490
rect 4320 410 4330 430
rect 4350 410 4360 430
rect 4320 350 4360 410
rect 4320 330 4330 350
rect 4350 330 4360 350
rect 4320 270 4360 330
rect 4320 250 4330 270
rect 4350 250 4360 270
rect 4320 190 4360 250
rect 4320 170 4330 190
rect 4350 170 4360 190
rect 4320 110 4360 170
rect 4320 90 4330 110
rect 4350 90 4360 110
rect 4320 30 4360 90
rect 4320 10 4330 30
rect 4350 10 4360 30
rect 4320 0 4360 10
rect 4400 15715 4440 15720
rect 4400 15685 4405 15715
rect 4435 15685 4440 15715
rect 4400 15635 4440 15685
rect 4400 15605 4405 15635
rect 4435 15605 4440 15635
rect 4400 15555 4440 15605
rect 4400 15525 4405 15555
rect 4435 15525 4440 15555
rect 4400 15475 4440 15525
rect 4400 15445 4405 15475
rect 4435 15445 4440 15475
rect 4400 15395 4440 15445
rect 4400 15365 4405 15395
rect 4435 15365 4440 15395
rect 4400 15315 4440 15365
rect 4400 15285 4405 15315
rect 4435 15285 4440 15315
rect 4400 15235 4440 15285
rect 4400 15205 4405 15235
rect 4435 15205 4440 15235
rect 4400 15155 4440 15205
rect 4400 15125 4405 15155
rect 4435 15125 4440 15155
rect 4400 15070 4440 15125
rect 4400 15050 4410 15070
rect 4430 15050 4440 15070
rect 4400 14995 4440 15050
rect 4400 14965 4405 14995
rect 4435 14965 4440 14995
rect 4400 14915 4440 14965
rect 4400 14885 4405 14915
rect 4435 14885 4440 14915
rect 4400 14835 4440 14885
rect 4400 14805 4405 14835
rect 4435 14805 4440 14835
rect 4400 14755 4440 14805
rect 4400 14725 4405 14755
rect 4435 14725 4440 14755
rect 4400 14675 4440 14725
rect 4400 14645 4405 14675
rect 4435 14645 4440 14675
rect 4400 14595 4440 14645
rect 4400 14565 4405 14595
rect 4435 14565 4440 14595
rect 4400 14515 4440 14565
rect 4400 14485 4405 14515
rect 4435 14485 4440 14515
rect 4400 14435 4440 14485
rect 4400 14405 4405 14435
rect 4435 14405 4440 14435
rect 4400 14350 4440 14405
rect 4400 14330 4410 14350
rect 4430 14330 4440 14350
rect 4400 14270 4440 14330
rect 4400 14250 4410 14270
rect 4430 14250 4440 14270
rect 4400 14190 4440 14250
rect 4400 14170 4410 14190
rect 4430 14170 4440 14190
rect 4400 14110 4440 14170
rect 4400 14090 4410 14110
rect 4430 14090 4440 14110
rect 4400 14035 4440 14090
rect 4400 14005 4405 14035
rect 4435 14005 4440 14035
rect 4400 13955 4440 14005
rect 4400 13925 4405 13955
rect 4435 13925 4440 13955
rect 4400 13875 4440 13925
rect 4400 13845 4405 13875
rect 4435 13845 4440 13875
rect 4400 13795 4440 13845
rect 4400 13765 4405 13795
rect 4435 13765 4440 13795
rect 4400 13715 4440 13765
rect 4400 13685 4405 13715
rect 4435 13685 4440 13715
rect 4400 13635 4440 13685
rect 4400 13605 4405 13635
rect 4435 13605 4440 13635
rect 4400 13555 4440 13605
rect 4400 13525 4405 13555
rect 4435 13525 4440 13555
rect 4400 13475 4440 13525
rect 4400 13445 4405 13475
rect 4435 13445 4440 13475
rect 4400 13390 4440 13445
rect 4400 13370 4410 13390
rect 4430 13370 4440 13390
rect 4400 13310 4440 13370
rect 4400 13290 4410 13310
rect 4430 13290 4440 13310
rect 4400 13230 4440 13290
rect 4400 13210 4410 13230
rect 4430 13210 4440 13230
rect 4400 13150 4440 13210
rect 4400 13130 4410 13150
rect 4430 13130 4440 13150
rect 4400 13075 4440 13130
rect 4400 13045 4405 13075
rect 4435 13045 4440 13075
rect 4400 12995 4440 13045
rect 4400 12965 4405 12995
rect 4435 12965 4440 12995
rect 4400 12915 4440 12965
rect 4400 12885 4405 12915
rect 4435 12885 4440 12915
rect 4400 12835 4440 12885
rect 4400 12805 4405 12835
rect 4435 12805 4440 12835
rect 4400 12755 4440 12805
rect 4400 12725 4405 12755
rect 4435 12725 4440 12755
rect 4400 12675 4440 12725
rect 4400 12645 4405 12675
rect 4435 12645 4440 12675
rect 4400 12595 4440 12645
rect 4400 12565 4405 12595
rect 4435 12565 4440 12595
rect 4400 12515 4440 12565
rect 4400 12485 4405 12515
rect 4435 12485 4440 12515
rect 4400 12430 4440 12485
rect 4400 12410 4410 12430
rect 4430 12410 4440 12430
rect 4400 12355 4440 12410
rect 4400 12325 4405 12355
rect 4435 12325 4440 12355
rect 4400 12275 4440 12325
rect 4400 12245 4405 12275
rect 4435 12245 4440 12275
rect 4400 12195 4440 12245
rect 4400 12165 4405 12195
rect 4435 12165 4440 12195
rect 4400 12115 4440 12165
rect 4400 12085 4405 12115
rect 4435 12085 4440 12115
rect 4400 12035 4440 12085
rect 4400 12005 4405 12035
rect 4435 12005 4440 12035
rect 4400 11955 4440 12005
rect 4400 11925 4405 11955
rect 4435 11925 4440 11955
rect 4400 11875 4440 11925
rect 4400 11845 4405 11875
rect 4435 11845 4440 11875
rect 4400 11795 4440 11845
rect 4400 11765 4405 11795
rect 4435 11765 4440 11795
rect 4400 11715 4440 11765
rect 4400 11685 4405 11715
rect 4435 11685 4440 11715
rect 4400 11635 4440 11685
rect 4400 11605 4405 11635
rect 4435 11605 4440 11635
rect 4400 11555 4440 11605
rect 4400 11525 4405 11555
rect 4435 11525 4440 11555
rect 4400 11475 4440 11525
rect 4400 11445 4405 11475
rect 4435 11445 4440 11475
rect 4400 11395 4440 11445
rect 4400 11365 4405 11395
rect 4435 11365 4440 11395
rect 4400 11315 4440 11365
rect 4400 11285 4405 11315
rect 4435 11285 4440 11315
rect 4400 11235 4440 11285
rect 4400 11205 4405 11235
rect 4435 11205 4440 11235
rect 4400 11155 4440 11205
rect 4400 11125 4405 11155
rect 4435 11125 4440 11155
rect 4400 11075 4440 11125
rect 4400 11045 4405 11075
rect 4435 11045 4440 11075
rect 4400 10990 4440 11045
rect 4400 10970 4410 10990
rect 4430 10970 4440 10990
rect 4400 10915 4440 10970
rect 4400 10885 4405 10915
rect 4435 10885 4440 10915
rect 4400 10835 4440 10885
rect 4400 10805 4405 10835
rect 4435 10805 4440 10835
rect 4400 10755 4440 10805
rect 4400 10725 4405 10755
rect 4435 10725 4440 10755
rect 4400 10675 4440 10725
rect 4400 10645 4405 10675
rect 4435 10645 4440 10675
rect 4400 10595 4440 10645
rect 4400 10565 4405 10595
rect 4435 10565 4440 10595
rect 4400 10515 4440 10565
rect 4400 10485 4405 10515
rect 4435 10485 4440 10515
rect 4400 10435 4440 10485
rect 4400 10405 4405 10435
rect 4435 10405 4440 10435
rect 4400 10355 4440 10405
rect 4400 10325 4405 10355
rect 4435 10325 4440 10355
rect 4400 10270 4440 10325
rect 4400 10250 4410 10270
rect 4430 10250 4440 10270
rect 4400 10190 4440 10250
rect 4400 10170 4410 10190
rect 4430 10170 4440 10190
rect 4400 10110 4440 10170
rect 4400 10090 4410 10110
rect 4430 10090 4440 10110
rect 4400 10030 4440 10090
rect 4400 10010 4410 10030
rect 4430 10010 4440 10030
rect 4400 9955 4440 10010
rect 4400 9925 4405 9955
rect 4435 9925 4440 9955
rect 4400 9875 4440 9925
rect 4400 9845 4405 9875
rect 4435 9845 4440 9875
rect 4400 9795 4440 9845
rect 4400 9765 4405 9795
rect 4435 9765 4440 9795
rect 4400 9715 4440 9765
rect 4400 9685 4405 9715
rect 4435 9685 4440 9715
rect 4400 9635 4440 9685
rect 4400 9605 4405 9635
rect 4435 9605 4440 9635
rect 4400 9555 4440 9605
rect 4400 9525 4405 9555
rect 4435 9525 4440 9555
rect 4400 9475 4440 9525
rect 4400 9445 4405 9475
rect 4435 9445 4440 9475
rect 4400 9395 4440 9445
rect 4400 9365 4405 9395
rect 4435 9365 4440 9395
rect 4400 9310 4440 9365
rect 4400 9290 4410 9310
rect 4430 9290 4440 9310
rect 4400 9230 4440 9290
rect 4400 9210 4410 9230
rect 4430 9210 4440 9230
rect 4400 9150 4440 9210
rect 4400 9130 4410 9150
rect 4430 9130 4440 9150
rect 4400 9070 4440 9130
rect 4400 9050 4410 9070
rect 4430 9050 4440 9070
rect 4400 8995 4440 9050
rect 4400 8965 4405 8995
rect 4435 8965 4440 8995
rect 4400 8915 4440 8965
rect 4400 8885 4405 8915
rect 4435 8885 4440 8915
rect 4400 8835 4440 8885
rect 4400 8805 4405 8835
rect 4435 8805 4440 8835
rect 4400 8755 4440 8805
rect 4400 8725 4405 8755
rect 4435 8725 4440 8755
rect 4400 8675 4440 8725
rect 4400 8645 4405 8675
rect 4435 8645 4440 8675
rect 4400 8595 4440 8645
rect 4400 8565 4405 8595
rect 4435 8565 4440 8595
rect 4400 8515 4440 8565
rect 4400 8485 4405 8515
rect 4435 8485 4440 8515
rect 4400 8435 4440 8485
rect 4400 8405 4405 8435
rect 4435 8405 4440 8435
rect 4400 8350 4440 8405
rect 4400 8330 4410 8350
rect 4430 8330 4440 8350
rect 4400 8275 4440 8330
rect 4400 8245 4405 8275
rect 4435 8245 4440 8275
rect 4400 8195 4440 8245
rect 4400 8165 4405 8195
rect 4435 8165 4440 8195
rect 4400 8115 4440 8165
rect 4400 8085 4405 8115
rect 4435 8085 4440 8115
rect 4400 8035 4440 8085
rect 4400 8005 4405 8035
rect 4435 8005 4440 8035
rect 4400 7955 4440 8005
rect 4400 7925 4405 7955
rect 4435 7925 4440 7955
rect 4400 7875 4440 7925
rect 4400 7845 4405 7875
rect 4435 7845 4440 7875
rect 4400 7795 4440 7845
rect 4400 7765 4405 7795
rect 4435 7765 4440 7795
rect 4400 7715 4440 7765
rect 4400 7685 4405 7715
rect 4435 7685 4440 7715
rect 4400 7635 4440 7685
rect 4400 7605 4405 7635
rect 4435 7605 4440 7635
rect 4400 7555 4440 7605
rect 4400 7525 4405 7555
rect 4435 7525 4440 7555
rect 4400 7475 4440 7525
rect 4400 7445 4405 7475
rect 4435 7445 4440 7475
rect 4400 7395 4440 7445
rect 4400 7365 4405 7395
rect 4435 7365 4440 7395
rect 4400 7315 4440 7365
rect 4400 7285 4405 7315
rect 4435 7285 4440 7315
rect 4400 7235 4440 7285
rect 4400 7205 4405 7235
rect 4435 7205 4440 7235
rect 4400 7155 4440 7205
rect 4400 7125 4405 7155
rect 4435 7125 4440 7155
rect 4400 7075 4440 7125
rect 4400 7045 4405 7075
rect 4435 7045 4440 7075
rect 4400 6995 4440 7045
rect 4400 6965 4405 6995
rect 4435 6965 4440 6995
rect 4400 6910 4440 6965
rect 4400 6890 4410 6910
rect 4430 6890 4440 6910
rect 4400 6835 4440 6890
rect 4400 6805 4405 6835
rect 4435 6805 4440 6835
rect 4400 6755 4440 6805
rect 4400 6725 4405 6755
rect 4435 6725 4440 6755
rect 4400 6675 4440 6725
rect 4400 6645 4405 6675
rect 4435 6645 4440 6675
rect 4400 6595 4440 6645
rect 4400 6565 4405 6595
rect 4435 6565 4440 6595
rect 4400 6515 4440 6565
rect 4400 6485 4405 6515
rect 4435 6485 4440 6515
rect 4400 6435 4440 6485
rect 4400 6405 4405 6435
rect 4435 6405 4440 6435
rect 4400 6355 4440 6405
rect 4400 6325 4405 6355
rect 4435 6325 4440 6355
rect 4400 6275 4440 6325
rect 4400 6245 4405 6275
rect 4435 6245 4440 6275
rect 4400 6190 4440 6245
rect 4400 6170 4410 6190
rect 4430 6170 4440 6190
rect 4400 6110 4440 6170
rect 4400 6090 4410 6110
rect 4430 6090 4440 6110
rect 4400 6030 4440 6090
rect 4400 6010 4410 6030
rect 4430 6010 4440 6030
rect 4400 5950 4440 6010
rect 4400 5930 4410 5950
rect 4430 5930 4440 5950
rect 4400 5875 4440 5930
rect 4400 5845 4405 5875
rect 4435 5845 4440 5875
rect 4400 5795 4440 5845
rect 4400 5765 4405 5795
rect 4435 5765 4440 5795
rect 4400 5715 4440 5765
rect 4400 5685 4405 5715
rect 4435 5685 4440 5715
rect 4400 5635 4440 5685
rect 4400 5605 4405 5635
rect 4435 5605 4440 5635
rect 4400 5555 4440 5605
rect 4400 5525 4405 5555
rect 4435 5525 4440 5555
rect 4400 5475 4440 5525
rect 4400 5445 4405 5475
rect 4435 5445 4440 5475
rect 4400 5395 4440 5445
rect 4400 5365 4405 5395
rect 4435 5365 4440 5395
rect 4400 5315 4440 5365
rect 4400 5285 4405 5315
rect 4435 5285 4440 5315
rect 4400 5235 4440 5285
rect 4400 5205 4405 5235
rect 4435 5205 4440 5235
rect 4400 5155 4440 5205
rect 4400 5125 4405 5155
rect 4435 5125 4440 5155
rect 4400 5075 4440 5125
rect 4400 5045 4405 5075
rect 4435 5045 4440 5075
rect 4400 4995 4440 5045
rect 4400 4965 4405 4995
rect 4435 4965 4440 4995
rect 4400 4915 4440 4965
rect 4400 4885 4405 4915
rect 4435 4885 4440 4915
rect 4400 4830 4440 4885
rect 4400 4810 4410 4830
rect 4430 4810 4440 4830
rect 4400 4755 4440 4810
rect 4400 4725 4405 4755
rect 4435 4725 4440 4755
rect 4400 4675 4440 4725
rect 4400 4645 4405 4675
rect 4435 4645 4440 4675
rect 4400 4590 4440 4645
rect 4400 4570 4410 4590
rect 4430 4570 4440 4590
rect 4400 4515 4440 4570
rect 4400 4485 4405 4515
rect 4435 4485 4440 4515
rect 4400 4435 4440 4485
rect 4400 4405 4405 4435
rect 4435 4405 4440 4435
rect 4400 4355 4440 4405
rect 4400 4325 4405 4355
rect 4435 4325 4440 4355
rect 4400 4275 4440 4325
rect 4400 4245 4405 4275
rect 4435 4245 4440 4275
rect 4400 4195 4440 4245
rect 4400 4165 4405 4195
rect 4435 4165 4440 4195
rect 4400 4115 4440 4165
rect 4400 4085 4405 4115
rect 4435 4085 4440 4115
rect 4400 4035 4440 4085
rect 4400 4005 4405 4035
rect 4435 4005 4440 4035
rect 4400 3955 4440 4005
rect 4400 3925 4405 3955
rect 4435 3925 4440 3955
rect 4400 3875 4440 3925
rect 4400 3845 4405 3875
rect 4435 3845 4440 3875
rect 4400 3790 4440 3845
rect 4400 3770 4410 3790
rect 4430 3770 4440 3790
rect 4400 3715 4440 3770
rect 4400 3685 4405 3715
rect 4435 3685 4440 3715
rect 4400 3635 4440 3685
rect 4400 3605 4405 3635
rect 4435 3605 4440 3635
rect 4400 3550 4440 3605
rect 4400 3530 4410 3550
rect 4430 3530 4440 3550
rect 4400 3475 4440 3530
rect 4400 3445 4405 3475
rect 4435 3445 4440 3475
rect 4400 3395 4440 3445
rect 4400 3365 4405 3395
rect 4435 3365 4440 3395
rect 4400 3310 4440 3365
rect 4400 3290 4410 3310
rect 4430 3290 4440 3310
rect 4400 3235 4440 3290
rect 4400 3205 4405 3235
rect 4435 3205 4440 3235
rect 4400 3155 4440 3205
rect 4400 3125 4405 3155
rect 4435 3125 4440 3155
rect 4400 3075 4440 3125
rect 4400 3045 4405 3075
rect 4435 3045 4440 3075
rect 4400 2995 4440 3045
rect 4400 2965 4405 2995
rect 4435 2965 4440 2995
rect 4400 2915 4440 2965
rect 4400 2885 4405 2915
rect 4435 2885 4440 2915
rect 4400 2835 4440 2885
rect 4400 2805 4405 2835
rect 4435 2805 4440 2835
rect 4400 2755 4440 2805
rect 4400 2725 4405 2755
rect 4435 2725 4440 2755
rect 4400 2675 4440 2725
rect 4400 2645 4405 2675
rect 4435 2645 4440 2675
rect 4400 2595 4440 2645
rect 4400 2565 4405 2595
rect 4435 2565 4440 2595
rect 4400 2515 4440 2565
rect 4400 2485 4405 2515
rect 4435 2485 4440 2515
rect 4400 2435 4440 2485
rect 4400 2405 4405 2435
rect 4435 2405 4440 2435
rect 4400 2355 4440 2405
rect 4400 2325 4405 2355
rect 4435 2325 4440 2355
rect 4400 2275 4440 2325
rect 4400 2245 4405 2275
rect 4435 2245 4440 2275
rect 4400 2195 4440 2245
rect 4400 2165 4405 2195
rect 4435 2165 4440 2195
rect 4400 2115 4440 2165
rect 4400 2085 4405 2115
rect 4435 2085 4440 2115
rect 4400 2035 4440 2085
rect 4400 2005 4405 2035
rect 4435 2005 4440 2035
rect 4400 1955 4440 2005
rect 4400 1925 4405 1955
rect 4435 1925 4440 1955
rect 4400 1870 4440 1925
rect 4400 1850 4410 1870
rect 4430 1850 4440 1870
rect 4400 1790 4440 1850
rect 4400 1770 4410 1790
rect 4430 1770 4440 1790
rect 4400 1715 4440 1770
rect 4400 1685 4405 1715
rect 4435 1685 4440 1715
rect 4400 1635 4440 1685
rect 4400 1605 4405 1635
rect 4435 1605 4440 1635
rect 4400 1555 4440 1605
rect 4400 1525 4405 1555
rect 4435 1525 4440 1555
rect 4400 1475 4440 1525
rect 4400 1445 4405 1475
rect 4435 1445 4440 1475
rect 4400 1395 4440 1445
rect 4400 1365 4405 1395
rect 4435 1365 4440 1395
rect 4400 1315 4440 1365
rect 4400 1285 4405 1315
rect 4435 1285 4440 1315
rect 4400 1235 4440 1285
rect 4400 1205 4405 1235
rect 4435 1205 4440 1235
rect 4400 1155 4440 1205
rect 4400 1125 4405 1155
rect 4435 1125 4440 1155
rect 4400 1075 4440 1125
rect 4400 1045 4405 1075
rect 4435 1045 4440 1075
rect 4400 995 4440 1045
rect 4400 965 4405 995
rect 4435 965 4440 995
rect 4400 910 4440 965
rect 4400 890 4410 910
rect 4430 890 4440 910
rect 4400 835 4440 890
rect 4400 805 4405 835
rect 4435 805 4440 835
rect 4400 755 4440 805
rect 4400 725 4405 755
rect 4435 725 4440 755
rect 4400 675 4440 725
rect 4400 645 4405 675
rect 4435 645 4440 675
rect 4400 595 4440 645
rect 4400 565 4405 595
rect 4435 565 4440 595
rect 4400 515 4440 565
rect 4400 485 4405 515
rect 4435 485 4440 515
rect 4400 430 4440 485
rect 4400 410 4410 430
rect 4430 410 4440 430
rect 4400 350 4440 410
rect 4400 330 4410 350
rect 4430 330 4440 350
rect 4400 275 4440 330
rect 4400 245 4405 275
rect 4435 245 4440 275
rect 4400 195 4440 245
rect 4400 165 4405 195
rect 4435 165 4440 195
rect 4400 115 4440 165
rect 4400 85 4405 115
rect 4435 85 4440 115
rect 4400 35 4440 85
rect 4400 5 4405 35
rect 4435 5 4440 35
rect 4400 0 4440 5
rect 4480 15715 4520 15720
rect 4480 15685 4485 15715
rect 4515 15685 4520 15715
rect 4480 15635 4520 15685
rect 4480 15605 4485 15635
rect 4515 15605 4520 15635
rect 4480 15555 4520 15605
rect 4480 15525 4485 15555
rect 4515 15525 4520 15555
rect 4480 15475 4520 15525
rect 4480 15445 4485 15475
rect 4515 15445 4520 15475
rect 4480 15395 4520 15445
rect 4480 15365 4485 15395
rect 4515 15365 4520 15395
rect 4480 15315 4520 15365
rect 4480 15285 4485 15315
rect 4515 15285 4520 15315
rect 4480 15235 4520 15285
rect 4480 15205 4485 15235
rect 4515 15205 4520 15235
rect 4480 15155 4520 15205
rect 4480 15125 4485 15155
rect 4515 15125 4520 15155
rect 4480 15070 4520 15125
rect 4480 15050 4490 15070
rect 4510 15050 4520 15070
rect 4480 14995 4520 15050
rect 4480 14965 4485 14995
rect 4515 14965 4520 14995
rect 4480 14915 4520 14965
rect 4480 14885 4485 14915
rect 4515 14885 4520 14915
rect 4480 14835 4520 14885
rect 4480 14805 4485 14835
rect 4515 14805 4520 14835
rect 4480 14755 4520 14805
rect 4480 14725 4485 14755
rect 4515 14725 4520 14755
rect 4480 14675 4520 14725
rect 4480 14645 4485 14675
rect 4515 14645 4520 14675
rect 4480 14595 4520 14645
rect 4480 14565 4485 14595
rect 4515 14565 4520 14595
rect 4480 14515 4520 14565
rect 4480 14485 4485 14515
rect 4515 14485 4520 14515
rect 4480 14435 4520 14485
rect 4480 14405 4485 14435
rect 4515 14405 4520 14435
rect 4480 14350 4520 14405
rect 4480 14330 4490 14350
rect 4510 14330 4520 14350
rect 4480 14270 4520 14330
rect 4480 14250 4490 14270
rect 4510 14250 4520 14270
rect 4480 14190 4520 14250
rect 4480 14170 4490 14190
rect 4510 14170 4520 14190
rect 4480 14110 4520 14170
rect 4480 14090 4490 14110
rect 4510 14090 4520 14110
rect 4480 14035 4520 14090
rect 4480 14005 4485 14035
rect 4515 14005 4520 14035
rect 4480 13955 4520 14005
rect 4480 13925 4485 13955
rect 4515 13925 4520 13955
rect 4480 13875 4520 13925
rect 4480 13845 4485 13875
rect 4515 13845 4520 13875
rect 4480 13795 4520 13845
rect 4480 13765 4485 13795
rect 4515 13765 4520 13795
rect 4480 13715 4520 13765
rect 4480 13685 4485 13715
rect 4515 13685 4520 13715
rect 4480 13635 4520 13685
rect 4480 13605 4485 13635
rect 4515 13605 4520 13635
rect 4480 13555 4520 13605
rect 4480 13525 4485 13555
rect 4515 13525 4520 13555
rect 4480 13475 4520 13525
rect 4480 13445 4485 13475
rect 4515 13445 4520 13475
rect 4480 13390 4520 13445
rect 4480 13370 4490 13390
rect 4510 13370 4520 13390
rect 4480 13310 4520 13370
rect 4480 13290 4490 13310
rect 4510 13290 4520 13310
rect 4480 13230 4520 13290
rect 4480 13210 4490 13230
rect 4510 13210 4520 13230
rect 4480 13150 4520 13210
rect 4480 13130 4490 13150
rect 4510 13130 4520 13150
rect 4480 13075 4520 13130
rect 4480 13045 4485 13075
rect 4515 13045 4520 13075
rect 4480 12995 4520 13045
rect 4480 12965 4485 12995
rect 4515 12965 4520 12995
rect 4480 12915 4520 12965
rect 4480 12885 4485 12915
rect 4515 12885 4520 12915
rect 4480 12835 4520 12885
rect 4480 12805 4485 12835
rect 4515 12805 4520 12835
rect 4480 12755 4520 12805
rect 4480 12725 4485 12755
rect 4515 12725 4520 12755
rect 4480 12675 4520 12725
rect 4480 12645 4485 12675
rect 4515 12645 4520 12675
rect 4480 12595 4520 12645
rect 4480 12565 4485 12595
rect 4515 12565 4520 12595
rect 4480 12515 4520 12565
rect 4480 12485 4485 12515
rect 4515 12485 4520 12515
rect 4480 12430 4520 12485
rect 4480 12410 4490 12430
rect 4510 12410 4520 12430
rect 4480 12355 4520 12410
rect 4480 12325 4485 12355
rect 4515 12325 4520 12355
rect 4480 12275 4520 12325
rect 4480 12245 4485 12275
rect 4515 12245 4520 12275
rect 4480 12195 4520 12245
rect 4480 12165 4485 12195
rect 4515 12165 4520 12195
rect 4480 12115 4520 12165
rect 4480 12085 4485 12115
rect 4515 12085 4520 12115
rect 4480 12035 4520 12085
rect 4480 12005 4485 12035
rect 4515 12005 4520 12035
rect 4480 11955 4520 12005
rect 4480 11925 4485 11955
rect 4515 11925 4520 11955
rect 4480 11875 4520 11925
rect 4480 11845 4485 11875
rect 4515 11845 4520 11875
rect 4480 11795 4520 11845
rect 4480 11765 4485 11795
rect 4515 11765 4520 11795
rect 4480 11715 4520 11765
rect 4480 11685 4485 11715
rect 4515 11685 4520 11715
rect 4480 11635 4520 11685
rect 4480 11605 4485 11635
rect 4515 11605 4520 11635
rect 4480 11555 4520 11605
rect 4480 11525 4485 11555
rect 4515 11525 4520 11555
rect 4480 11475 4520 11525
rect 4480 11445 4485 11475
rect 4515 11445 4520 11475
rect 4480 11395 4520 11445
rect 4480 11365 4485 11395
rect 4515 11365 4520 11395
rect 4480 11315 4520 11365
rect 4480 11285 4485 11315
rect 4515 11285 4520 11315
rect 4480 11235 4520 11285
rect 4480 11205 4485 11235
rect 4515 11205 4520 11235
rect 4480 11155 4520 11205
rect 4480 11125 4485 11155
rect 4515 11125 4520 11155
rect 4480 11075 4520 11125
rect 4480 11045 4485 11075
rect 4515 11045 4520 11075
rect 4480 10990 4520 11045
rect 4480 10970 4490 10990
rect 4510 10970 4520 10990
rect 4480 10915 4520 10970
rect 4480 10885 4485 10915
rect 4515 10885 4520 10915
rect 4480 10835 4520 10885
rect 4480 10805 4485 10835
rect 4515 10805 4520 10835
rect 4480 10755 4520 10805
rect 4480 10725 4485 10755
rect 4515 10725 4520 10755
rect 4480 10675 4520 10725
rect 4480 10645 4485 10675
rect 4515 10645 4520 10675
rect 4480 10595 4520 10645
rect 4480 10565 4485 10595
rect 4515 10565 4520 10595
rect 4480 10515 4520 10565
rect 4480 10485 4485 10515
rect 4515 10485 4520 10515
rect 4480 10435 4520 10485
rect 4480 10405 4485 10435
rect 4515 10405 4520 10435
rect 4480 10355 4520 10405
rect 4480 10325 4485 10355
rect 4515 10325 4520 10355
rect 4480 10270 4520 10325
rect 4480 10250 4490 10270
rect 4510 10250 4520 10270
rect 4480 10190 4520 10250
rect 4480 10170 4490 10190
rect 4510 10170 4520 10190
rect 4480 10110 4520 10170
rect 4480 10090 4490 10110
rect 4510 10090 4520 10110
rect 4480 10030 4520 10090
rect 4480 10010 4490 10030
rect 4510 10010 4520 10030
rect 4480 9955 4520 10010
rect 4480 9925 4485 9955
rect 4515 9925 4520 9955
rect 4480 9875 4520 9925
rect 4480 9845 4485 9875
rect 4515 9845 4520 9875
rect 4480 9795 4520 9845
rect 4480 9765 4485 9795
rect 4515 9765 4520 9795
rect 4480 9715 4520 9765
rect 4480 9685 4485 9715
rect 4515 9685 4520 9715
rect 4480 9635 4520 9685
rect 4480 9605 4485 9635
rect 4515 9605 4520 9635
rect 4480 9555 4520 9605
rect 4480 9525 4485 9555
rect 4515 9525 4520 9555
rect 4480 9475 4520 9525
rect 4480 9445 4485 9475
rect 4515 9445 4520 9475
rect 4480 9395 4520 9445
rect 4480 9365 4485 9395
rect 4515 9365 4520 9395
rect 4480 9310 4520 9365
rect 4480 9290 4490 9310
rect 4510 9290 4520 9310
rect 4480 9230 4520 9290
rect 4480 9210 4490 9230
rect 4510 9210 4520 9230
rect 4480 9150 4520 9210
rect 4480 9130 4490 9150
rect 4510 9130 4520 9150
rect 4480 9070 4520 9130
rect 4480 9050 4490 9070
rect 4510 9050 4520 9070
rect 4480 8995 4520 9050
rect 4480 8965 4485 8995
rect 4515 8965 4520 8995
rect 4480 8915 4520 8965
rect 4480 8885 4485 8915
rect 4515 8885 4520 8915
rect 4480 8835 4520 8885
rect 4480 8805 4485 8835
rect 4515 8805 4520 8835
rect 4480 8755 4520 8805
rect 4480 8725 4485 8755
rect 4515 8725 4520 8755
rect 4480 8675 4520 8725
rect 4480 8645 4485 8675
rect 4515 8645 4520 8675
rect 4480 8595 4520 8645
rect 4480 8565 4485 8595
rect 4515 8565 4520 8595
rect 4480 8515 4520 8565
rect 4480 8485 4485 8515
rect 4515 8485 4520 8515
rect 4480 8435 4520 8485
rect 4480 8405 4485 8435
rect 4515 8405 4520 8435
rect 4480 8350 4520 8405
rect 4480 8330 4490 8350
rect 4510 8330 4520 8350
rect 4480 8275 4520 8330
rect 4480 8245 4485 8275
rect 4515 8245 4520 8275
rect 4480 8195 4520 8245
rect 4480 8165 4485 8195
rect 4515 8165 4520 8195
rect 4480 8115 4520 8165
rect 4480 8085 4485 8115
rect 4515 8085 4520 8115
rect 4480 8035 4520 8085
rect 4480 8005 4485 8035
rect 4515 8005 4520 8035
rect 4480 7955 4520 8005
rect 4480 7925 4485 7955
rect 4515 7925 4520 7955
rect 4480 7875 4520 7925
rect 4480 7845 4485 7875
rect 4515 7845 4520 7875
rect 4480 7795 4520 7845
rect 4480 7765 4485 7795
rect 4515 7765 4520 7795
rect 4480 7715 4520 7765
rect 4480 7685 4485 7715
rect 4515 7685 4520 7715
rect 4480 7635 4520 7685
rect 4480 7605 4485 7635
rect 4515 7605 4520 7635
rect 4480 7555 4520 7605
rect 4480 7525 4485 7555
rect 4515 7525 4520 7555
rect 4480 7475 4520 7525
rect 4480 7445 4485 7475
rect 4515 7445 4520 7475
rect 4480 7395 4520 7445
rect 4480 7365 4485 7395
rect 4515 7365 4520 7395
rect 4480 7315 4520 7365
rect 4480 7285 4485 7315
rect 4515 7285 4520 7315
rect 4480 7235 4520 7285
rect 4480 7205 4485 7235
rect 4515 7205 4520 7235
rect 4480 7155 4520 7205
rect 4480 7125 4485 7155
rect 4515 7125 4520 7155
rect 4480 7075 4520 7125
rect 4480 7045 4485 7075
rect 4515 7045 4520 7075
rect 4480 6995 4520 7045
rect 4480 6965 4485 6995
rect 4515 6965 4520 6995
rect 4480 6910 4520 6965
rect 4480 6890 4490 6910
rect 4510 6890 4520 6910
rect 4480 6835 4520 6890
rect 4480 6805 4485 6835
rect 4515 6805 4520 6835
rect 4480 6755 4520 6805
rect 4480 6725 4485 6755
rect 4515 6725 4520 6755
rect 4480 6675 4520 6725
rect 4480 6645 4485 6675
rect 4515 6645 4520 6675
rect 4480 6595 4520 6645
rect 4480 6565 4485 6595
rect 4515 6565 4520 6595
rect 4480 6515 4520 6565
rect 4480 6485 4485 6515
rect 4515 6485 4520 6515
rect 4480 6435 4520 6485
rect 4480 6405 4485 6435
rect 4515 6405 4520 6435
rect 4480 6355 4520 6405
rect 4480 6325 4485 6355
rect 4515 6325 4520 6355
rect 4480 6275 4520 6325
rect 4480 6245 4485 6275
rect 4515 6245 4520 6275
rect 4480 6190 4520 6245
rect 4480 6170 4490 6190
rect 4510 6170 4520 6190
rect 4480 6110 4520 6170
rect 4480 6090 4490 6110
rect 4510 6090 4520 6110
rect 4480 6030 4520 6090
rect 4480 6010 4490 6030
rect 4510 6010 4520 6030
rect 4480 5950 4520 6010
rect 4480 5930 4490 5950
rect 4510 5930 4520 5950
rect 4480 5875 4520 5930
rect 4480 5845 4485 5875
rect 4515 5845 4520 5875
rect 4480 5795 4520 5845
rect 4480 5765 4485 5795
rect 4515 5765 4520 5795
rect 4480 5715 4520 5765
rect 4480 5685 4485 5715
rect 4515 5685 4520 5715
rect 4480 5635 4520 5685
rect 4480 5605 4485 5635
rect 4515 5605 4520 5635
rect 4480 5555 4520 5605
rect 4480 5525 4485 5555
rect 4515 5525 4520 5555
rect 4480 5475 4520 5525
rect 4480 5445 4485 5475
rect 4515 5445 4520 5475
rect 4480 5395 4520 5445
rect 4480 5365 4485 5395
rect 4515 5365 4520 5395
rect 4480 5315 4520 5365
rect 4480 5285 4485 5315
rect 4515 5285 4520 5315
rect 4480 5235 4520 5285
rect 4480 5205 4485 5235
rect 4515 5205 4520 5235
rect 4480 5155 4520 5205
rect 4480 5125 4485 5155
rect 4515 5125 4520 5155
rect 4480 5075 4520 5125
rect 4480 5045 4485 5075
rect 4515 5045 4520 5075
rect 4480 4995 4520 5045
rect 4480 4965 4485 4995
rect 4515 4965 4520 4995
rect 4480 4915 4520 4965
rect 4480 4885 4485 4915
rect 4515 4885 4520 4915
rect 4480 4830 4520 4885
rect 4480 4810 4490 4830
rect 4510 4810 4520 4830
rect 4480 4755 4520 4810
rect 4480 4725 4485 4755
rect 4515 4725 4520 4755
rect 4480 4675 4520 4725
rect 4480 4645 4485 4675
rect 4515 4645 4520 4675
rect 4480 4590 4520 4645
rect 4480 4570 4490 4590
rect 4510 4570 4520 4590
rect 4480 4515 4520 4570
rect 4480 4485 4485 4515
rect 4515 4485 4520 4515
rect 4480 4435 4520 4485
rect 4480 4405 4485 4435
rect 4515 4405 4520 4435
rect 4480 4355 4520 4405
rect 4480 4325 4485 4355
rect 4515 4325 4520 4355
rect 4480 4275 4520 4325
rect 4480 4245 4485 4275
rect 4515 4245 4520 4275
rect 4480 4195 4520 4245
rect 4480 4165 4485 4195
rect 4515 4165 4520 4195
rect 4480 4115 4520 4165
rect 4480 4085 4485 4115
rect 4515 4085 4520 4115
rect 4480 4035 4520 4085
rect 4480 4005 4485 4035
rect 4515 4005 4520 4035
rect 4480 3955 4520 4005
rect 4480 3925 4485 3955
rect 4515 3925 4520 3955
rect 4480 3875 4520 3925
rect 4480 3845 4485 3875
rect 4515 3845 4520 3875
rect 4480 3790 4520 3845
rect 4480 3770 4490 3790
rect 4510 3770 4520 3790
rect 4480 3715 4520 3770
rect 4480 3685 4485 3715
rect 4515 3685 4520 3715
rect 4480 3635 4520 3685
rect 4480 3605 4485 3635
rect 4515 3605 4520 3635
rect 4480 3550 4520 3605
rect 4480 3530 4490 3550
rect 4510 3530 4520 3550
rect 4480 3475 4520 3530
rect 4480 3445 4485 3475
rect 4515 3445 4520 3475
rect 4480 3395 4520 3445
rect 4480 3365 4485 3395
rect 4515 3365 4520 3395
rect 4480 3310 4520 3365
rect 4480 3290 4490 3310
rect 4510 3290 4520 3310
rect 4480 3235 4520 3290
rect 4480 3205 4485 3235
rect 4515 3205 4520 3235
rect 4480 3155 4520 3205
rect 4480 3125 4485 3155
rect 4515 3125 4520 3155
rect 4480 3075 4520 3125
rect 4480 3045 4485 3075
rect 4515 3045 4520 3075
rect 4480 2995 4520 3045
rect 4480 2965 4485 2995
rect 4515 2965 4520 2995
rect 4480 2915 4520 2965
rect 4480 2885 4485 2915
rect 4515 2885 4520 2915
rect 4480 2835 4520 2885
rect 4480 2805 4485 2835
rect 4515 2805 4520 2835
rect 4480 2755 4520 2805
rect 4480 2725 4485 2755
rect 4515 2725 4520 2755
rect 4480 2675 4520 2725
rect 4480 2645 4485 2675
rect 4515 2645 4520 2675
rect 4480 2595 4520 2645
rect 4480 2565 4485 2595
rect 4515 2565 4520 2595
rect 4480 2515 4520 2565
rect 4480 2485 4485 2515
rect 4515 2485 4520 2515
rect 4480 2435 4520 2485
rect 4480 2405 4485 2435
rect 4515 2405 4520 2435
rect 4480 2355 4520 2405
rect 4480 2325 4485 2355
rect 4515 2325 4520 2355
rect 4480 2275 4520 2325
rect 4480 2245 4485 2275
rect 4515 2245 4520 2275
rect 4480 2195 4520 2245
rect 4480 2165 4485 2195
rect 4515 2165 4520 2195
rect 4480 2115 4520 2165
rect 4480 2085 4485 2115
rect 4515 2085 4520 2115
rect 4480 2035 4520 2085
rect 4480 2005 4485 2035
rect 4515 2005 4520 2035
rect 4480 1955 4520 2005
rect 4480 1925 4485 1955
rect 4515 1925 4520 1955
rect 4480 1870 4520 1925
rect 4480 1850 4490 1870
rect 4510 1850 4520 1870
rect 4480 1790 4520 1850
rect 4480 1770 4490 1790
rect 4510 1770 4520 1790
rect 4480 1715 4520 1770
rect 4480 1685 4485 1715
rect 4515 1685 4520 1715
rect 4480 1635 4520 1685
rect 4480 1605 4485 1635
rect 4515 1605 4520 1635
rect 4480 1555 4520 1605
rect 4480 1525 4485 1555
rect 4515 1525 4520 1555
rect 4480 1475 4520 1525
rect 4480 1445 4485 1475
rect 4515 1445 4520 1475
rect 4480 1395 4520 1445
rect 4480 1365 4485 1395
rect 4515 1365 4520 1395
rect 4480 1315 4520 1365
rect 4480 1285 4485 1315
rect 4515 1285 4520 1315
rect 4480 1235 4520 1285
rect 4480 1205 4485 1235
rect 4515 1205 4520 1235
rect 4480 1155 4520 1205
rect 4480 1125 4485 1155
rect 4515 1125 4520 1155
rect 4480 1075 4520 1125
rect 4480 1045 4485 1075
rect 4515 1045 4520 1075
rect 4480 995 4520 1045
rect 4480 965 4485 995
rect 4515 965 4520 995
rect 4480 910 4520 965
rect 4480 890 4490 910
rect 4510 890 4520 910
rect 4480 835 4520 890
rect 4480 805 4485 835
rect 4515 805 4520 835
rect 4480 755 4520 805
rect 4480 725 4485 755
rect 4515 725 4520 755
rect 4480 675 4520 725
rect 4480 645 4485 675
rect 4515 645 4520 675
rect 4480 595 4520 645
rect 4480 565 4485 595
rect 4515 565 4520 595
rect 4480 515 4520 565
rect 4480 485 4485 515
rect 4515 485 4520 515
rect 4480 430 4520 485
rect 4480 410 4490 430
rect 4510 410 4520 430
rect 4480 350 4520 410
rect 4480 330 4490 350
rect 4510 330 4520 350
rect 4480 275 4520 330
rect 4480 245 4485 275
rect 4515 245 4520 275
rect 4480 195 4520 245
rect 4480 165 4485 195
rect 4515 165 4520 195
rect 4480 115 4520 165
rect 4480 85 4485 115
rect 4515 85 4520 115
rect 4480 35 4520 85
rect 4480 5 4485 35
rect 4515 5 4520 35
rect 4480 0 4520 5
rect 4560 15710 4600 15720
rect 4560 15690 4570 15710
rect 4590 15690 4600 15710
rect 4560 15630 4600 15690
rect 4560 15610 4570 15630
rect 4590 15610 4600 15630
rect 4560 15550 4600 15610
rect 4560 15530 4570 15550
rect 4590 15530 4600 15550
rect 4560 15470 4600 15530
rect 4560 15450 4570 15470
rect 4590 15450 4600 15470
rect 4560 15390 4600 15450
rect 4560 15370 4570 15390
rect 4590 15370 4600 15390
rect 4560 15310 4600 15370
rect 4560 15290 4570 15310
rect 4590 15290 4600 15310
rect 4560 15230 4600 15290
rect 4560 15210 4570 15230
rect 4590 15210 4600 15230
rect 4560 15150 4600 15210
rect 4560 15130 4570 15150
rect 4590 15130 4600 15150
rect 4560 15070 4600 15130
rect 4560 15050 4570 15070
rect 4590 15050 4600 15070
rect 4560 14990 4600 15050
rect 4560 14970 4570 14990
rect 4590 14970 4600 14990
rect 4560 14910 4600 14970
rect 4560 14890 4570 14910
rect 4590 14890 4600 14910
rect 4560 14830 4600 14890
rect 4560 14810 4570 14830
rect 4590 14810 4600 14830
rect 4560 14750 4600 14810
rect 4560 14730 4570 14750
rect 4590 14730 4600 14750
rect 4560 14670 4600 14730
rect 4560 14650 4570 14670
rect 4590 14650 4600 14670
rect 4560 14590 4600 14650
rect 4560 14570 4570 14590
rect 4590 14570 4600 14590
rect 4560 14510 4600 14570
rect 4560 14490 4570 14510
rect 4590 14490 4600 14510
rect 4560 14430 4600 14490
rect 4560 14410 4570 14430
rect 4590 14410 4600 14430
rect 4560 14350 4600 14410
rect 4560 14330 4570 14350
rect 4590 14330 4600 14350
rect 4560 14270 4600 14330
rect 4560 14250 4570 14270
rect 4590 14250 4600 14270
rect 4560 14190 4600 14250
rect 4560 14170 4570 14190
rect 4590 14170 4600 14190
rect 4560 14110 4600 14170
rect 4560 14090 4570 14110
rect 4590 14090 4600 14110
rect 4560 14030 4600 14090
rect 4560 14010 4570 14030
rect 4590 14010 4600 14030
rect 4560 13950 4600 14010
rect 4560 13930 4570 13950
rect 4590 13930 4600 13950
rect 4560 13870 4600 13930
rect 4560 13850 4570 13870
rect 4590 13850 4600 13870
rect 4560 13790 4600 13850
rect 4560 13770 4570 13790
rect 4590 13770 4600 13790
rect 4560 13710 4600 13770
rect 4560 13690 4570 13710
rect 4590 13690 4600 13710
rect 4560 13630 4600 13690
rect 4560 13610 4570 13630
rect 4590 13610 4600 13630
rect 4560 13550 4600 13610
rect 4560 13530 4570 13550
rect 4590 13530 4600 13550
rect 4560 13470 4600 13530
rect 4560 13450 4570 13470
rect 4590 13450 4600 13470
rect 4560 13390 4600 13450
rect 4560 13370 4570 13390
rect 4590 13370 4600 13390
rect 4560 13310 4600 13370
rect 4560 13290 4570 13310
rect 4590 13290 4600 13310
rect 4560 13230 4600 13290
rect 4560 13210 4570 13230
rect 4590 13210 4600 13230
rect 4560 13150 4600 13210
rect 4560 13130 4570 13150
rect 4590 13130 4600 13150
rect 4560 13070 4600 13130
rect 4560 13050 4570 13070
rect 4590 13050 4600 13070
rect 4560 12990 4600 13050
rect 4560 12970 4570 12990
rect 4590 12970 4600 12990
rect 4560 12910 4600 12970
rect 4560 12890 4570 12910
rect 4590 12890 4600 12910
rect 4560 12830 4600 12890
rect 4560 12810 4570 12830
rect 4590 12810 4600 12830
rect 4560 12750 4600 12810
rect 4560 12730 4570 12750
rect 4590 12730 4600 12750
rect 4560 12670 4600 12730
rect 4560 12650 4570 12670
rect 4590 12650 4600 12670
rect 4560 12590 4600 12650
rect 4560 12570 4570 12590
rect 4590 12570 4600 12590
rect 4560 12510 4600 12570
rect 4560 12490 4570 12510
rect 4590 12490 4600 12510
rect 4560 12430 4600 12490
rect 4560 12410 4570 12430
rect 4590 12410 4600 12430
rect 4560 12350 4600 12410
rect 4560 12330 4570 12350
rect 4590 12330 4600 12350
rect 4560 12270 4600 12330
rect 4560 12250 4570 12270
rect 4590 12250 4600 12270
rect 4560 12190 4600 12250
rect 4560 12170 4570 12190
rect 4590 12170 4600 12190
rect 4560 12110 4600 12170
rect 4560 12090 4570 12110
rect 4590 12090 4600 12110
rect 4560 12030 4600 12090
rect 4560 12010 4570 12030
rect 4590 12010 4600 12030
rect 4560 11950 4600 12010
rect 4560 11930 4570 11950
rect 4590 11930 4600 11950
rect 4560 11870 4600 11930
rect 4560 11850 4570 11870
rect 4590 11850 4600 11870
rect 4560 11790 4600 11850
rect 4560 11770 4570 11790
rect 4590 11770 4600 11790
rect 4560 11710 4600 11770
rect 4560 11690 4570 11710
rect 4590 11690 4600 11710
rect 4560 11630 4600 11690
rect 4560 11610 4570 11630
rect 4590 11610 4600 11630
rect 4560 11550 4600 11610
rect 4560 11530 4570 11550
rect 4590 11530 4600 11550
rect 4560 11470 4600 11530
rect 4560 11450 4570 11470
rect 4590 11450 4600 11470
rect 4560 11390 4600 11450
rect 4560 11370 4570 11390
rect 4590 11370 4600 11390
rect 4560 11310 4600 11370
rect 4560 11290 4570 11310
rect 4590 11290 4600 11310
rect 4560 11230 4600 11290
rect 4560 11210 4570 11230
rect 4590 11210 4600 11230
rect 4560 11150 4600 11210
rect 4560 11130 4570 11150
rect 4590 11130 4600 11150
rect 4560 11070 4600 11130
rect 4560 11050 4570 11070
rect 4590 11050 4600 11070
rect 4560 10990 4600 11050
rect 4560 10970 4570 10990
rect 4590 10970 4600 10990
rect 4560 10910 4600 10970
rect 4560 10890 4570 10910
rect 4590 10890 4600 10910
rect 4560 10830 4600 10890
rect 4560 10810 4570 10830
rect 4590 10810 4600 10830
rect 4560 10750 4600 10810
rect 4560 10730 4570 10750
rect 4590 10730 4600 10750
rect 4560 10670 4600 10730
rect 4560 10650 4570 10670
rect 4590 10650 4600 10670
rect 4560 10590 4600 10650
rect 4560 10570 4570 10590
rect 4590 10570 4600 10590
rect 4560 10510 4600 10570
rect 4560 10490 4570 10510
rect 4590 10490 4600 10510
rect 4560 10430 4600 10490
rect 4560 10410 4570 10430
rect 4590 10410 4600 10430
rect 4560 10350 4600 10410
rect 4560 10330 4570 10350
rect 4590 10330 4600 10350
rect 4560 10270 4600 10330
rect 4560 10250 4570 10270
rect 4590 10250 4600 10270
rect 4560 10190 4600 10250
rect 4560 10170 4570 10190
rect 4590 10170 4600 10190
rect 4560 10110 4600 10170
rect 4560 10090 4570 10110
rect 4590 10090 4600 10110
rect 4560 10030 4600 10090
rect 4560 10010 4570 10030
rect 4590 10010 4600 10030
rect 4560 9950 4600 10010
rect 4560 9930 4570 9950
rect 4590 9930 4600 9950
rect 4560 9870 4600 9930
rect 4560 9850 4570 9870
rect 4590 9850 4600 9870
rect 4560 9790 4600 9850
rect 4560 9770 4570 9790
rect 4590 9770 4600 9790
rect 4560 9710 4600 9770
rect 4560 9690 4570 9710
rect 4590 9690 4600 9710
rect 4560 9630 4600 9690
rect 4560 9610 4570 9630
rect 4590 9610 4600 9630
rect 4560 9550 4600 9610
rect 4560 9530 4570 9550
rect 4590 9530 4600 9550
rect 4560 9470 4600 9530
rect 4560 9450 4570 9470
rect 4590 9450 4600 9470
rect 4560 9390 4600 9450
rect 4560 9370 4570 9390
rect 4590 9370 4600 9390
rect 4560 9310 4600 9370
rect 4560 9290 4570 9310
rect 4590 9290 4600 9310
rect 4560 9230 4600 9290
rect 4560 9210 4570 9230
rect 4590 9210 4600 9230
rect 4560 9150 4600 9210
rect 4560 9130 4570 9150
rect 4590 9130 4600 9150
rect 4560 9070 4600 9130
rect 4560 9050 4570 9070
rect 4590 9050 4600 9070
rect 4560 8990 4600 9050
rect 4560 8970 4570 8990
rect 4590 8970 4600 8990
rect 4560 8910 4600 8970
rect 4560 8890 4570 8910
rect 4590 8890 4600 8910
rect 4560 8830 4600 8890
rect 4560 8810 4570 8830
rect 4590 8810 4600 8830
rect 4560 8750 4600 8810
rect 4560 8730 4570 8750
rect 4590 8730 4600 8750
rect 4560 8670 4600 8730
rect 4560 8650 4570 8670
rect 4590 8650 4600 8670
rect 4560 8590 4600 8650
rect 4560 8570 4570 8590
rect 4590 8570 4600 8590
rect 4560 8510 4600 8570
rect 4560 8490 4570 8510
rect 4590 8490 4600 8510
rect 4560 8430 4600 8490
rect 4560 8410 4570 8430
rect 4590 8410 4600 8430
rect 4560 8350 4600 8410
rect 4560 8330 4570 8350
rect 4590 8330 4600 8350
rect 4560 8270 4600 8330
rect 4560 8250 4570 8270
rect 4590 8250 4600 8270
rect 4560 8190 4600 8250
rect 4560 8170 4570 8190
rect 4590 8170 4600 8190
rect 4560 8110 4600 8170
rect 4560 8090 4570 8110
rect 4590 8090 4600 8110
rect 4560 8030 4600 8090
rect 4560 8010 4570 8030
rect 4590 8010 4600 8030
rect 4560 7950 4600 8010
rect 4560 7930 4570 7950
rect 4590 7930 4600 7950
rect 4560 7870 4600 7930
rect 4560 7850 4570 7870
rect 4590 7850 4600 7870
rect 4560 7790 4600 7850
rect 4560 7770 4570 7790
rect 4590 7770 4600 7790
rect 4560 7710 4600 7770
rect 4560 7690 4570 7710
rect 4590 7690 4600 7710
rect 4560 7630 4600 7690
rect 4560 7610 4570 7630
rect 4590 7610 4600 7630
rect 4560 7550 4600 7610
rect 4560 7530 4570 7550
rect 4590 7530 4600 7550
rect 4560 7470 4600 7530
rect 4560 7450 4570 7470
rect 4590 7450 4600 7470
rect 4560 7390 4600 7450
rect 4560 7370 4570 7390
rect 4590 7370 4600 7390
rect 4560 7310 4600 7370
rect 4560 7290 4570 7310
rect 4590 7290 4600 7310
rect 4560 7230 4600 7290
rect 4560 7210 4570 7230
rect 4590 7210 4600 7230
rect 4560 7150 4600 7210
rect 4560 7130 4570 7150
rect 4590 7130 4600 7150
rect 4560 7070 4600 7130
rect 4560 7050 4570 7070
rect 4590 7050 4600 7070
rect 4560 6990 4600 7050
rect 4560 6970 4570 6990
rect 4590 6970 4600 6990
rect 4560 6910 4600 6970
rect 4560 6890 4570 6910
rect 4590 6890 4600 6910
rect 4560 6830 4600 6890
rect 4560 6810 4570 6830
rect 4590 6810 4600 6830
rect 4560 6750 4600 6810
rect 4560 6730 4570 6750
rect 4590 6730 4600 6750
rect 4560 6670 4600 6730
rect 4560 6650 4570 6670
rect 4590 6650 4600 6670
rect 4560 6590 4600 6650
rect 4560 6570 4570 6590
rect 4590 6570 4600 6590
rect 4560 6510 4600 6570
rect 4560 6490 4570 6510
rect 4590 6490 4600 6510
rect 4560 6430 4600 6490
rect 4560 6410 4570 6430
rect 4590 6410 4600 6430
rect 4560 6350 4600 6410
rect 4560 6330 4570 6350
rect 4590 6330 4600 6350
rect 4560 6270 4600 6330
rect 4560 6250 4570 6270
rect 4590 6250 4600 6270
rect 4560 6190 4600 6250
rect 4560 6170 4570 6190
rect 4590 6170 4600 6190
rect 4560 6110 4600 6170
rect 4560 6090 4570 6110
rect 4590 6090 4600 6110
rect 4560 6030 4600 6090
rect 4560 6010 4570 6030
rect 4590 6010 4600 6030
rect 4560 5950 4600 6010
rect 4560 5930 4570 5950
rect 4590 5930 4600 5950
rect 4560 5870 4600 5930
rect 4560 5850 4570 5870
rect 4590 5850 4600 5870
rect 4560 5790 4600 5850
rect 4560 5770 4570 5790
rect 4590 5770 4600 5790
rect 4560 5710 4600 5770
rect 4560 5690 4570 5710
rect 4590 5690 4600 5710
rect 4560 5630 4600 5690
rect 4560 5610 4570 5630
rect 4590 5610 4600 5630
rect 4560 5550 4600 5610
rect 4560 5530 4570 5550
rect 4590 5530 4600 5550
rect 4560 5470 4600 5530
rect 4560 5450 4570 5470
rect 4590 5450 4600 5470
rect 4560 5390 4600 5450
rect 4560 5370 4570 5390
rect 4590 5370 4600 5390
rect 4560 5310 4600 5370
rect 4560 5290 4570 5310
rect 4590 5290 4600 5310
rect 4560 5230 4600 5290
rect 4560 5210 4570 5230
rect 4590 5210 4600 5230
rect 4560 5150 4600 5210
rect 4560 5130 4570 5150
rect 4590 5130 4600 5150
rect 4560 5070 4600 5130
rect 4560 5050 4570 5070
rect 4590 5050 4600 5070
rect 4560 4990 4600 5050
rect 4560 4970 4570 4990
rect 4590 4970 4600 4990
rect 4560 4910 4600 4970
rect 4560 4890 4570 4910
rect 4590 4890 4600 4910
rect 4560 4830 4600 4890
rect 4560 4810 4570 4830
rect 4590 4810 4600 4830
rect 4560 4750 4600 4810
rect 4560 4730 4570 4750
rect 4590 4730 4600 4750
rect 4560 4670 4600 4730
rect 4560 4650 4570 4670
rect 4590 4650 4600 4670
rect 4560 4590 4600 4650
rect 4560 4570 4570 4590
rect 4590 4570 4600 4590
rect 4560 4510 4600 4570
rect 4560 4490 4570 4510
rect 4590 4490 4600 4510
rect 4560 4430 4600 4490
rect 4560 4410 4570 4430
rect 4590 4410 4600 4430
rect 4560 4350 4600 4410
rect 4560 4330 4570 4350
rect 4590 4330 4600 4350
rect 4560 4270 4600 4330
rect 4560 4250 4570 4270
rect 4590 4250 4600 4270
rect 4560 4190 4600 4250
rect 4560 4170 4570 4190
rect 4590 4170 4600 4190
rect 4560 4110 4600 4170
rect 4560 4090 4570 4110
rect 4590 4090 4600 4110
rect 4560 4030 4600 4090
rect 4560 4010 4570 4030
rect 4590 4010 4600 4030
rect 4560 3950 4600 4010
rect 4560 3930 4570 3950
rect 4590 3930 4600 3950
rect 4560 3870 4600 3930
rect 4560 3850 4570 3870
rect 4590 3850 4600 3870
rect 4560 3790 4600 3850
rect 4560 3770 4570 3790
rect 4590 3770 4600 3790
rect 4560 3710 4600 3770
rect 4560 3690 4570 3710
rect 4590 3690 4600 3710
rect 4560 3630 4600 3690
rect 4560 3610 4570 3630
rect 4590 3610 4600 3630
rect 4560 3550 4600 3610
rect 4560 3530 4570 3550
rect 4590 3530 4600 3550
rect 4560 3470 4600 3530
rect 4560 3450 4570 3470
rect 4590 3450 4600 3470
rect 4560 3390 4600 3450
rect 4560 3370 4570 3390
rect 4590 3370 4600 3390
rect 4560 3310 4600 3370
rect 4560 3290 4570 3310
rect 4590 3290 4600 3310
rect 4560 3230 4600 3290
rect 4560 3210 4570 3230
rect 4590 3210 4600 3230
rect 4560 3150 4600 3210
rect 4560 3130 4570 3150
rect 4590 3130 4600 3150
rect 4560 3070 4600 3130
rect 4560 3050 4570 3070
rect 4590 3050 4600 3070
rect 4560 2990 4600 3050
rect 4560 2970 4570 2990
rect 4590 2970 4600 2990
rect 4560 2910 4600 2970
rect 4560 2890 4570 2910
rect 4590 2890 4600 2910
rect 4560 2830 4600 2890
rect 4560 2810 4570 2830
rect 4590 2810 4600 2830
rect 4560 2750 4600 2810
rect 4560 2730 4570 2750
rect 4590 2730 4600 2750
rect 4560 2670 4600 2730
rect 4560 2650 4570 2670
rect 4590 2650 4600 2670
rect 4560 2590 4600 2650
rect 4560 2570 4570 2590
rect 4590 2570 4600 2590
rect 4560 2510 4600 2570
rect 4560 2490 4570 2510
rect 4590 2490 4600 2510
rect 4560 2430 4600 2490
rect 4560 2410 4570 2430
rect 4590 2410 4600 2430
rect 4560 2350 4600 2410
rect 4560 2330 4570 2350
rect 4590 2330 4600 2350
rect 4560 2270 4600 2330
rect 4560 2250 4570 2270
rect 4590 2250 4600 2270
rect 4560 2190 4600 2250
rect 4560 2170 4570 2190
rect 4590 2170 4600 2190
rect 4560 2110 4600 2170
rect 4560 2090 4570 2110
rect 4590 2090 4600 2110
rect 4560 2030 4600 2090
rect 4560 2010 4570 2030
rect 4590 2010 4600 2030
rect 4560 1950 4600 2010
rect 4560 1930 4570 1950
rect 4590 1930 4600 1950
rect 4560 1870 4600 1930
rect 4560 1850 4570 1870
rect 4590 1850 4600 1870
rect 4560 1790 4600 1850
rect 4560 1770 4570 1790
rect 4590 1770 4600 1790
rect 4560 1710 4600 1770
rect 4560 1690 4570 1710
rect 4590 1690 4600 1710
rect 4560 1630 4600 1690
rect 4560 1610 4570 1630
rect 4590 1610 4600 1630
rect 4560 1550 4600 1610
rect 4560 1530 4570 1550
rect 4590 1530 4600 1550
rect 4560 1470 4600 1530
rect 4560 1450 4570 1470
rect 4590 1450 4600 1470
rect 4560 1390 4600 1450
rect 4560 1370 4570 1390
rect 4590 1370 4600 1390
rect 4560 1310 4600 1370
rect 4560 1290 4570 1310
rect 4590 1290 4600 1310
rect 4560 1230 4600 1290
rect 4560 1210 4570 1230
rect 4590 1210 4600 1230
rect 4560 1150 4600 1210
rect 4560 1130 4570 1150
rect 4590 1130 4600 1150
rect 4560 1070 4600 1130
rect 4560 1050 4570 1070
rect 4590 1050 4600 1070
rect 4560 990 4600 1050
rect 4560 970 4570 990
rect 4590 970 4600 990
rect 4560 910 4600 970
rect 4560 890 4570 910
rect 4590 890 4600 910
rect 4560 830 4600 890
rect 4560 810 4570 830
rect 4590 810 4600 830
rect 4560 750 4600 810
rect 4560 730 4570 750
rect 4590 730 4600 750
rect 4560 670 4600 730
rect 4560 650 4570 670
rect 4590 650 4600 670
rect 4560 590 4600 650
rect 4560 570 4570 590
rect 4590 570 4600 590
rect 4560 510 4600 570
rect 4560 490 4570 510
rect 4590 490 4600 510
rect 4560 430 4600 490
rect 4560 410 4570 430
rect 4590 410 4600 430
rect 4560 350 4600 410
rect 4560 330 4570 350
rect 4590 330 4600 350
rect 4560 270 4600 330
rect 4560 250 4570 270
rect 4590 250 4600 270
rect 4560 190 4600 250
rect 4560 170 4570 190
rect 4590 170 4600 190
rect 4560 110 4600 170
rect 4560 90 4570 110
rect 4590 90 4600 110
rect 4560 30 4600 90
rect 4560 10 4570 30
rect 4590 10 4600 30
rect 4560 0 4600 10
rect 4640 15715 4680 15720
rect 4640 15685 4645 15715
rect 4675 15685 4680 15715
rect 4640 15635 4680 15685
rect 4640 15605 4645 15635
rect 4675 15605 4680 15635
rect 4640 15555 4680 15605
rect 4640 15525 4645 15555
rect 4675 15525 4680 15555
rect 4640 15475 4680 15525
rect 4640 15445 4645 15475
rect 4675 15445 4680 15475
rect 4640 15395 4680 15445
rect 4640 15365 4645 15395
rect 4675 15365 4680 15395
rect 4640 15315 4680 15365
rect 4640 15285 4645 15315
rect 4675 15285 4680 15315
rect 4640 15235 4680 15285
rect 4640 15205 4645 15235
rect 4675 15205 4680 15235
rect 4640 15155 4680 15205
rect 4640 15125 4645 15155
rect 4675 15125 4680 15155
rect 4640 15070 4680 15125
rect 4640 15050 4650 15070
rect 4670 15050 4680 15070
rect 4640 14995 4680 15050
rect 4640 14965 4645 14995
rect 4675 14965 4680 14995
rect 4640 14915 4680 14965
rect 4640 14885 4645 14915
rect 4675 14885 4680 14915
rect 4640 14835 4680 14885
rect 4640 14805 4645 14835
rect 4675 14805 4680 14835
rect 4640 14755 4680 14805
rect 4640 14725 4645 14755
rect 4675 14725 4680 14755
rect 4640 14675 4680 14725
rect 4640 14645 4645 14675
rect 4675 14645 4680 14675
rect 4640 14595 4680 14645
rect 4640 14565 4645 14595
rect 4675 14565 4680 14595
rect 4640 14515 4680 14565
rect 4640 14485 4645 14515
rect 4675 14485 4680 14515
rect 4640 14435 4680 14485
rect 4640 14405 4645 14435
rect 4675 14405 4680 14435
rect 4640 14350 4680 14405
rect 4640 14330 4650 14350
rect 4670 14330 4680 14350
rect 4640 14270 4680 14330
rect 4640 14250 4650 14270
rect 4670 14250 4680 14270
rect 4640 14190 4680 14250
rect 4640 14170 4650 14190
rect 4670 14170 4680 14190
rect 4640 14110 4680 14170
rect 4640 14090 4650 14110
rect 4670 14090 4680 14110
rect 4640 14035 4680 14090
rect 4640 14005 4645 14035
rect 4675 14005 4680 14035
rect 4640 13955 4680 14005
rect 4640 13925 4645 13955
rect 4675 13925 4680 13955
rect 4640 13875 4680 13925
rect 4640 13845 4645 13875
rect 4675 13845 4680 13875
rect 4640 13795 4680 13845
rect 4640 13765 4645 13795
rect 4675 13765 4680 13795
rect 4640 13715 4680 13765
rect 4640 13685 4645 13715
rect 4675 13685 4680 13715
rect 4640 13635 4680 13685
rect 4640 13605 4645 13635
rect 4675 13605 4680 13635
rect 4640 13555 4680 13605
rect 4640 13525 4645 13555
rect 4675 13525 4680 13555
rect 4640 13475 4680 13525
rect 4640 13445 4645 13475
rect 4675 13445 4680 13475
rect 4640 13390 4680 13445
rect 4640 13370 4650 13390
rect 4670 13370 4680 13390
rect 4640 13310 4680 13370
rect 4640 13290 4650 13310
rect 4670 13290 4680 13310
rect 4640 13230 4680 13290
rect 4640 13210 4650 13230
rect 4670 13210 4680 13230
rect 4640 13150 4680 13210
rect 4640 13130 4650 13150
rect 4670 13130 4680 13150
rect 4640 13075 4680 13130
rect 4640 13045 4645 13075
rect 4675 13045 4680 13075
rect 4640 12995 4680 13045
rect 4640 12965 4645 12995
rect 4675 12965 4680 12995
rect 4640 12915 4680 12965
rect 4640 12885 4645 12915
rect 4675 12885 4680 12915
rect 4640 12835 4680 12885
rect 4640 12805 4645 12835
rect 4675 12805 4680 12835
rect 4640 12755 4680 12805
rect 4640 12725 4645 12755
rect 4675 12725 4680 12755
rect 4640 12675 4680 12725
rect 4640 12645 4645 12675
rect 4675 12645 4680 12675
rect 4640 12595 4680 12645
rect 4640 12565 4645 12595
rect 4675 12565 4680 12595
rect 4640 12515 4680 12565
rect 4640 12485 4645 12515
rect 4675 12485 4680 12515
rect 4640 12430 4680 12485
rect 4640 12410 4650 12430
rect 4670 12410 4680 12430
rect 4640 12355 4680 12410
rect 4640 12325 4645 12355
rect 4675 12325 4680 12355
rect 4640 12275 4680 12325
rect 4640 12245 4645 12275
rect 4675 12245 4680 12275
rect 4640 12195 4680 12245
rect 4640 12165 4645 12195
rect 4675 12165 4680 12195
rect 4640 12115 4680 12165
rect 4640 12085 4645 12115
rect 4675 12085 4680 12115
rect 4640 12035 4680 12085
rect 4640 12005 4645 12035
rect 4675 12005 4680 12035
rect 4640 11955 4680 12005
rect 4640 11925 4645 11955
rect 4675 11925 4680 11955
rect 4640 11875 4680 11925
rect 4640 11845 4645 11875
rect 4675 11845 4680 11875
rect 4640 11795 4680 11845
rect 4640 11765 4645 11795
rect 4675 11765 4680 11795
rect 4640 11715 4680 11765
rect 4640 11685 4645 11715
rect 4675 11685 4680 11715
rect 4640 11635 4680 11685
rect 4640 11605 4645 11635
rect 4675 11605 4680 11635
rect 4640 11555 4680 11605
rect 4640 11525 4645 11555
rect 4675 11525 4680 11555
rect 4640 11475 4680 11525
rect 4640 11445 4645 11475
rect 4675 11445 4680 11475
rect 4640 11395 4680 11445
rect 4640 11365 4645 11395
rect 4675 11365 4680 11395
rect 4640 11315 4680 11365
rect 4640 11285 4645 11315
rect 4675 11285 4680 11315
rect 4640 11235 4680 11285
rect 4640 11205 4645 11235
rect 4675 11205 4680 11235
rect 4640 11155 4680 11205
rect 4640 11125 4645 11155
rect 4675 11125 4680 11155
rect 4640 11075 4680 11125
rect 4640 11045 4645 11075
rect 4675 11045 4680 11075
rect 4640 10990 4680 11045
rect 4640 10970 4650 10990
rect 4670 10970 4680 10990
rect 4640 10915 4680 10970
rect 4640 10885 4645 10915
rect 4675 10885 4680 10915
rect 4640 10835 4680 10885
rect 4640 10805 4645 10835
rect 4675 10805 4680 10835
rect 4640 10755 4680 10805
rect 4640 10725 4645 10755
rect 4675 10725 4680 10755
rect 4640 10675 4680 10725
rect 4640 10645 4645 10675
rect 4675 10645 4680 10675
rect 4640 10595 4680 10645
rect 4640 10565 4645 10595
rect 4675 10565 4680 10595
rect 4640 10515 4680 10565
rect 4640 10485 4645 10515
rect 4675 10485 4680 10515
rect 4640 10435 4680 10485
rect 4640 10405 4645 10435
rect 4675 10405 4680 10435
rect 4640 10355 4680 10405
rect 4640 10325 4645 10355
rect 4675 10325 4680 10355
rect 4640 10270 4680 10325
rect 4640 10250 4650 10270
rect 4670 10250 4680 10270
rect 4640 10190 4680 10250
rect 4640 10170 4650 10190
rect 4670 10170 4680 10190
rect 4640 10110 4680 10170
rect 4640 10090 4650 10110
rect 4670 10090 4680 10110
rect 4640 10030 4680 10090
rect 4640 10010 4650 10030
rect 4670 10010 4680 10030
rect 4640 9955 4680 10010
rect 4640 9925 4645 9955
rect 4675 9925 4680 9955
rect 4640 9875 4680 9925
rect 4640 9845 4645 9875
rect 4675 9845 4680 9875
rect 4640 9795 4680 9845
rect 4640 9765 4645 9795
rect 4675 9765 4680 9795
rect 4640 9715 4680 9765
rect 4640 9685 4645 9715
rect 4675 9685 4680 9715
rect 4640 9635 4680 9685
rect 4640 9605 4645 9635
rect 4675 9605 4680 9635
rect 4640 9555 4680 9605
rect 4640 9525 4645 9555
rect 4675 9525 4680 9555
rect 4640 9475 4680 9525
rect 4640 9445 4645 9475
rect 4675 9445 4680 9475
rect 4640 9395 4680 9445
rect 4640 9365 4645 9395
rect 4675 9365 4680 9395
rect 4640 9310 4680 9365
rect 4640 9290 4650 9310
rect 4670 9290 4680 9310
rect 4640 9230 4680 9290
rect 4640 9210 4650 9230
rect 4670 9210 4680 9230
rect 4640 9150 4680 9210
rect 4640 9130 4650 9150
rect 4670 9130 4680 9150
rect 4640 9070 4680 9130
rect 4640 9050 4650 9070
rect 4670 9050 4680 9070
rect 4640 8995 4680 9050
rect 4640 8965 4645 8995
rect 4675 8965 4680 8995
rect 4640 8915 4680 8965
rect 4640 8885 4645 8915
rect 4675 8885 4680 8915
rect 4640 8835 4680 8885
rect 4640 8805 4645 8835
rect 4675 8805 4680 8835
rect 4640 8755 4680 8805
rect 4640 8725 4645 8755
rect 4675 8725 4680 8755
rect 4640 8675 4680 8725
rect 4640 8645 4645 8675
rect 4675 8645 4680 8675
rect 4640 8595 4680 8645
rect 4640 8565 4645 8595
rect 4675 8565 4680 8595
rect 4640 8515 4680 8565
rect 4640 8485 4645 8515
rect 4675 8485 4680 8515
rect 4640 8435 4680 8485
rect 4640 8405 4645 8435
rect 4675 8405 4680 8435
rect 4640 8350 4680 8405
rect 4640 8330 4650 8350
rect 4670 8330 4680 8350
rect 4640 8275 4680 8330
rect 4640 8245 4645 8275
rect 4675 8245 4680 8275
rect 4640 8195 4680 8245
rect 4640 8165 4645 8195
rect 4675 8165 4680 8195
rect 4640 8115 4680 8165
rect 4640 8085 4645 8115
rect 4675 8085 4680 8115
rect 4640 8035 4680 8085
rect 4640 8005 4645 8035
rect 4675 8005 4680 8035
rect 4640 7955 4680 8005
rect 4640 7925 4645 7955
rect 4675 7925 4680 7955
rect 4640 7875 4680 7925
rect 4640 7845 4645 7875
rect 4675 7845 4680 7875
rect 4640 7795 4680 7845
rect 4640 7765 4645 7795
rect 4675 7765 4680 7795
rect 4640 7715 4680 7765
rect 4640 7685 4645 7715
rect 4675 7685 4680 7715
rect 4640 7635 4680 7685
rect 4640 7605 4645 7635
rect 4675 7605 4680 7635
rect 4640 7555 4680 7605
rect 4640 7525 4645 7555
rect 4675 7525 4680 7555
rect 4640 7475 4680 7525
rect 4640 7445 4645 7475
rect 4675 7445 4680 7475
rect 4640 7395 4680 7445
rect 4640 7365 4645 7395
rect 4675 7365 4680 7395
rect 4640 7315 4680 7365
rect 4640 7285 4645 7315
rect 4675 7285 4680 7315
rect 4640 7235 4680 7285
rect 4640 7205 4645 7235
rect 4675 7205 4680 7235
rect 4640 7155 4680 7205
rect 4640 7125 4645 7155
rect 4675 7125 4680 7155
rect 4640 7075 4680 7125
rect 4640 7045 4645 7075
rect 4675 7045 4680 7075
rect 4640 6995 4680 7045
rect 4640 6965 4645 6995
rect 4675 6965 4680 6995
rect 4640 6910 4680 6965
rect 4640 6890 4650 6910
rect 4670 6890 4680 6910
rect 4640 6835 4680 6890
rect 4640 6805 4645 6835
rect 4675 6805 4680 6835
rect 4640 6755 4680 6805
rect 4640 6725 4645 6755
rect 4675 6725 4680 6755
rect 4640 6675 4680 6725
rect 4640 6645 4645 6675
rect 4675 6645 4680 6675
rect 4640 6595 4680 6645
rect 4640 6565 4645 6595
rect 4675 6565 4680 6595
rect 4640 6515 4680 6565
rect 4640 6485 4645 6515
rect 4675 6485 4680 6515
rect 4640 6435 4680 6485
rect 4640 6405 4645 6435
rect 4675 6405 4680 6435
rect 4640 6355 4680 6405
rect 4640 6325 4645 6355
rect 4675 6325 4680 6355
rect 4640 6275 4680 6325
rect 4640 6245 4645 6275
rect 4675 6245 4680 6275
rect 4640 6190 4680 6245
rect 4640 6170 4650 6190
rect 4670 6170 4680 6190
rect 4640 6110 4680 6170
rect 4640 6090 4650 6110
rect 4670 6090 4680 6110
rect 4640 6030 4680 6090
rect 4640 6010 4650 6030
rect 4670 6010 4680 6030
rect 4640 5950 4680 6010
rect 4640 5930 4650 5950
rect 4670 5930 4680 5950
rect 4640 5875 4680 5930
rect 4640 5845 4645 5875
rect 4675 5845 4680 5875
rect 4640 5795 4680 5845
rect 4640 5765 4645 5795
rect 4675 5765 4680 5795
rect 4640 5715 4680 5765
rect 4640 5685 4645 5715
rect 4675 5685 4680 5715
rect 4640 5635 4680 5685
rect 4640 5605 4645 5635
rect 4675 5605 4680 5635
rect 4640 5555 4680 5605
rect 4640 5525 4645 5555
rect 4675 5525 4680 5555
rect 4640 5475 4680 5525
rect 4640 5445 4645 5475
rect 4675 5445 4680 5475
rect 4640 5395 4680 5445
rect 4640 5365 4645 5395
rect 4675 5365 4680 5395
rect 4640 5315 4680 5365
rect 4640 5285 4645 5315
rect 4675 5285 4680 5315
rect 4640 5235 4680 5285
rect 4640 5205 4645 5235
rect 4675 5205 4680 5235
rect 4640 5155 4680 5205
rect 4640 5125 4645 5155
rect 4675 5125 4680 5155
rect 4640 5075 4680 5125
rect 4640 5045 4645 5075
rect 4675 5045 4680 5075
rect 4640 4995 4680 5045
rect 4640 4965 4645 4995
rect 4675 4965 4680 4995
rect 4640 4915 4680 4965
rect 4640 4885 4645 4915
rect 4675 4885 4680 4915
rect 4640 4830 4680 4885
rect 4640 4810 4650 4830
rect 4670 4810 4680 4830
rect 4640 4755 4680 4810
rect 4640 4725 4645 4755
rect 4675 4725 4680 4755
rect 4640 4675 4680 4725
rect 4640 4645 4645 4675
rect 4675 4645 4680 4675
rect 4640 4590 4680 4645
rect 4640 4570 4650 4590
rect 4670 4570 4680 4590
rect 4640 4515 4680 4570
rect 4640 4485 4645 4515
rect 4675 4485 4680 4515
rect 4640 4435 4680 4485
rect 4640 4405 4645 4435
rect 4675 4405 4680 4435
rect 4640 4355 4680 4405
rect 4640 4325 4645 4355
rect 4675 4325 4680 4355
rect 4640 4275 4680 4325
rect 4640 4245 4645 4275
rect 4675 4245 4680 4275
rect 4640 4195 4680 4245
rect 4640 4165 4645 4195
rect 4675 4165 4680 4195
rect 4640 4115 4680 4165
rect 4640 4085 4645 4115
rect 4675 4085 4680 4115
rect 4640 4035 4680 4085
rect 4640 4005 4645 4035
rect 4675 4005 4680 4035
rect 4640 3955 4680 4005
rect 4640 3925 4645 3955
rect 4675 3925 4680 3955
rect 4640 3875 4680 3925
rect 4640 3845 4645 3875
rect 4675 3845 4680 3875
rect 4640 3790 4680 3845
rect 4640 3770 4650 3790
rect 4670 3770 4680 3790
rect 4640 3715 4680 3770
rect 4640 3685 4645 3715
rect 4675 3685 4680 3715
rect 4640 3635 4680 3685
rect 4640 3605 4645 3635
rect 4675 3605 4680 3635
rect 4640 3550 4680 3605
rect 4640 3530 4650 3550
rect 4670 3530 4680 3550
rect 4640 3475 4680 3530
rect 4640 3445 4645 3475
rect 4675 3445 4680 3475
rect 4640 3395 4680 3445
rect 4640 3365 4645 3395
rect 4675 3365 4680 3395
rect 4640 3310 4680 3365
rect 4640 3290 4650 3310
rect 4670 3290 4680 3310
rect 4640 3235 4680 3290
rect 4640 3205 4645 3235
rect 4675 3205 4680 3235
rect 4640 3155 4680 3205
rect 4640 3125 4645 3155
rect 4675 3125 4680 3155
rect 4640 3075 4680 3125
rect 4640 3045 4645 3075
rect 4675 3045 4680 3075
rect 4640 2995 4680 3045
rect 4640 2965 4645 2995
rect 4675 2965 4680 2995
rect 4640 2915 4680 2965
rect 4640 2885 4645 2915
rect 4675 2885 4680 2915
rect 4640 2835 4680 2885
rect 4640 2805 4645 2835
rect 4675 2805 4680 2835
rect 4640 2755 4680 2805
rect 4640 2725 4645 2755
rect 4675 2725 4680 2755
rect 4640 2675 4680 2725
rect 4640 2645 4645 2675
rect 4675 2645 4680 2675
rect 4640 2595 4680 2645
rect 4640 2565 4645 2595
rect 4675 2565 4680 2595
rect 4640 2515 4680 2565
rect 4640 2485 4645 2515
rect 4675 2485 4680 2515
rect 4640 2435 4680 2485
rect 4640 2405 4645 2435
rect 4675 2405 4680 2435
rect 4640 2355 4680 2405
rect 4640 2325 4645 2355
rect 4675 2325 4680 2355
rect 4640 2275 4680 2325
rect 4640 2245 4645 2275
rect 4675 2245 4680 2275
rect 4640 2195 4680 2245
rect 4640 2165 4645 2195
rect 4675 2165 4680 2195
rect 4640 2115 4680 2165
rect 4640 2085 4645 2115
rect 4675 2085 4680 2115
rect 4640 2035 4680 2085
rect 4640 2005 4645 2035
rect 4675 2005 4680 2035
rect 4640 1955 4680 2005
rect 4640 1925 4645 1955
rect 4675 1925 4680 1955
rect 4640 1870 4680 1925
rect 4640 1850 4650 1870
rect 4670 1850 4680 1870
rect 4640 1790 4680 1850
rect 4640 1770 4650 1790
rect 4670 1770 4680 1790
rect 4640 1715 4680 1770
rect 4640 1685 4645 1715
rect 4675 1685 4680 1715
rect 4640 1635 4680 1685
rect 4640 1605 4645 1635
rect 4675 1605 4680 1635
rect 4640 1555 4680 1605
rect 4640 1525 4645 1555
rect 4675 1525 4680 1555
rect 4640 1475 4680 1525
rect 4640 1445 4645 1475
rect 4675 1445 4680 1475
rect 4640 1395 4680 1445
rect 4640 1365 4645 1395
rect 4675 1365 4680 1395
rect 4640 1315 4680 1365
rect 4640 1285 4645 1315
rect 4675 1285 4680 1315
rect 4640 1235 4680 1285
rect 4640 1205 4645 1235
rect 4675 1205 4680 1235
rect 4640 1155 4680 1205
rect 4640 1125 4645 1155
rect 4675 1125 4680 1155
rect 4640 1075 4680 1125
rect 4640 1045 4645 1075
rect 4675 1045 4680 1075
rect 4640 995 4680 1045
rect 4640 965 4645 995
rect 4675 965 4680 995
rect 4640 910 4680 965
rect 4640 890 4650 910
rect 4670 890 4680 910
rect 4640 835 4680 890
rect 4640 805 4645 835
rect 4675 805 4680 835
rect 4640 755 4680 805
rect 4640 725 4645 755
rect 4675 725 4680 755
rect 4640 675 4680 725
rect 4640 645 4645 675
rect 4675 645 4680 675
rect 4640 595 4680 645
rect 4640 565 4645 595
rect 4675 565 4680 595
rect 4640 515 4680 565
rect 4640 485 4645 515
rect 4675 485 4680 515
rect 4640 430 4680 485
rect 4640 410 4650 430
rect 4670 410 4680 430
rect 4640 350 4680 410
rect 4640 330 4650 350
rect 4670 330 4680 350
rect 4640 275 4680 330
rect 4640 245 4645 275
rect 4675 245 4680 275
rect 4640 195 4680 245
rect 4640 165 4645 195
rect 4675 165 4680 195
rect 4640 115 4680 165
rect 4640 85 4645 115
rect 4675 85 4680 115
rect 4640 35 4680 85
rect 4640 5 4645 35
rect 4675 5 4680 35
rect 4640 0 4680 5
rect 4720 15715 4760 15720
rect 4720 15685 4725 15715
rect 4755 15685 4760 15715
rect 4720 15635 4760 15685
rect 4720 15605 4725 15635
rect 4755 15605 4760 15635
rect 4720 15555 4760 15605
rect 4720 15525 4725 15555
rect 4755 15525 4760 15555
rect 4720 15475 4760 15525
rect 4720 15445 4725 15475
rect 4755 15445 4760 15475
rect 4720 15395 4760 15445
rect 4720 15365 4725 15395
rect 4755 15365 4760 15395
rect 4720 15315 4760 15365
rect 4720 15285 4725 15315
rect 4755 15285 4760 15315
rect 4720 15235 4760 15285
rect 4720 15205 4725 15235
rect 4755 15205 4760 15235
rect 4720 15155 4760 15205
rect 4720 15125 4725 15155
rect 4755 15125 4760 15155
rect 4720 15070 4760 15125
rect 4720 15050 4730 15070
rect 4750 15050 4760 15070
rect 4720 14995 4760 15050
rect 4720 14965 4725 14995
rect 4755 14965 4760 14995
rect 4720 14915 4760 14965
rect 4720 14885 4725 14915
rect 4755 14885 4760 14915
rect 4720 14835 4760 14885
rect 4720 14805 4725 14835
rect 4755 14805 4760 14835
rect 4720 14755 4760 14805
rect 4720 14725 4725 14755
rect 4755 14725 4760 14755
rect 4720 14675 4760 14725
rect 4720 14645 4725 14675
rect 4755 14645 4760 14675
rect 4720 14595 4760 14645
rect 4720 14565 4725 14595
rect 4755 14565 4760 14595
rect 4720 14515 4760 14565
rect 4720 14485 4725 14515
rect 4755 14485 4760 14515
rect 4720 14435 4760 14485
rect 4720 14405 4725 14435
rect 4755 14405 4760 14435
rect 4720 14350 4760 14405
rect 4720 14330 4730 14350
rect 4750 14330 4760 14350
rect 4720 14270 4760 14330
rect 4720 14250 4730 14270
rect 4750 14250 4760 14270
rect 4720 14190 4760 14250
rect 4720 14170 4730 14190
rect 4750 14170 4760 14190
rect 4720 14110 4760 14170
rect 4720 14090 4730 14110
rect 4750 14090 4760 14110
rect 4720 14035 4760 14090
rect 4720 14005 4725 14035
rect 4755 14005 4760 14035
rect 4720 13955 4760 14005
rect 4720 13925 4725 13955
rect 4755 13925 4760 13955
rect 4720 13875 4760 13925
rect 4720 13845 4725 13875
rect 4755 13845 4760 13875
rect 4720 13795 4760 13845
rect 4720 13765 4725 13795
rect 4755 13765 4760 13795
rect 4720 13715 4760 13765
rect 4720 13685 4725 13715
rect 4755 13685 4760 13715
rect 4720 13635 4760 13685
rect 4720 13605 4725 13635
rect 4755 13605 4760 13635
rect 4720 13555 4760 13605
rect 4720 13525 4725 13555
rect 4755 13525 4760 13555
rect 4720 13475 4760 13525
rect 4720 13445 4725 13475
rect 4755 13445 4760 13475
rect 4720 13390 4760 13445
rect 4720 13370 4730 13390
rect 4750 13370 4760 13390
rect 4720 13310 4760 13370
rect 4720 13290 4730 13310
rect 4750 13290 4760 13310
rect 4720 13230 4760 13290
rect 4720 13210 4730 13230
rect 4750 13210 4760 13230
rect 4720 13150 4760 13210
rect 4720 13130 4730 13150
rect 4750 13130 4760 13150
rect 4720 13075 4760 13130
rect 4720 13045 4725 13075
rect 4755 13045 4760 13075
rect 4720 12995 4760 13045
rect 4720 12965 4725 12995
rect 4755 12965 4760 12995
rect 4720 12915 4760 12965
rect 4720 12885 4725 12915
rect 4755 12885 4760 12915
rect 4720 12835 4760 12885
rect 4720 12805 4725 12835
rect 4755 12805 4760 12835
rect 4720 12755 4760 12805
rect 4720 12725 4725 12755
rect 4755 12725 4760 12755
rect 4720 12675 4760 12725
rect 4720 12645 4725 12675
rect 4755 12645 4760 12675
rect 4720 12595 4760 12645
rect 4720 12565 4725 12595
rect 4755 12565 4760 12595
rect 4720 12515 4760 12565
rect 4720 12485 4725 12515
rect 4755 12485 4760 12515
rect 4720 12430 4760 12485
rect 4720 12410 4730 12430
rect 4750 12410 4760 12430
rect 4720 12355 4760 12410
rect 4720 12325 4725 12355
rect 4755 12325 4760 12355
rect 4720 12275 4760 12325
rect 4720 12245 4725 12275
rect 4755 12245 4760 12275
rect 4720 12195 4760 12245
rect 4720 12165 4725 12195
rect 4755 12165 4760 12195
rect 4720 12115 4760 12165
rect 4720 12085 4725 12115
rect 4755 12085 4760 12115
rect 4720 12035 4760 12085
rect 4720 12005 4725 12035
rect 4755 12005 4760 12035
rect 4720 11955 4760 12005
rect 4720 11925 4725 11955
rect 4755 11925 4760 11955
rect 4720 11875 4760 11925
rect 4720 11845 4725 11875
rect 4755 11845 4760 11875
rect 4720 11795 4760 11845
rect 4720 11765 4725 11795
rect 4755 11765 4760 11795
rect 4720 11715 4760 11765
rect 4720 11685 4725 11715
rect 4755 11685 4760 11715
rect 4720 11635 4760 11685
rect 4720 11605 4725 11635
rect 4755 11605 4760 11635
rect 4720 11555 4760 11605
rect 4720 11525 4725 11555
rect 4755 11525 4760 11555
rect 4720 11475 4760 11525
rect 4720 11445 4725 11475
rect 4755 11445 4760 11475
rect 4720 11395 4760 11445
rect 4720 11365 4725 11395
rect 4755 11365 4760 11395
rect 4720 11315 4760 11365
rect 4720 11285 4725 11315
rect 4755 11285 4760 11315
rect 4720 11235 4760 11285
rect 4720 11205 4725 11235
rect 4755 11205 4760 11235
rect 4720 11155 4760 11205
rect 4720 11125 4725 11155
rect 4755 11125 4760 11155
rect 4720 11075 4760 11125
rect 4720 11045 4725 11075
rect 4755 11045 4760 11075
rect 4720 10990 4760 11045
rect 4720 10970 4730 10990
rect 4750 10970 4760 10990
rect 4720 10915 4760 10970
rect 4720 10885 4725 10915
rect 4755 10885 4760 10915
rect 4720 10835 4760 10885
rect 4720 10805 4725 10835
rect 4755 10805 4760 10835
rect 4720 10755 4760 10805
rect 4720 10725 4725 10755
rect 4755 10725 4760 10755
rect 4720 10675 4760 10725
rect 4720 10645 4725 10675
rect 4755 10645 4760 10675
rect 4720 10595 4760 10645
rect 4720 10565 4725 10595
rect 4755 10565 4760 10595
rect 4720 10515 4760 10565
rect 4720 10485 4725 10515
rect 4755 10485 4760 10515
rect 4720 10435 4760 10485
rect 4720 10405 4725 10435
rect 4755 10405 4760 10435
rect 4720 10355 4760 10405
rect 4720 10325 4725 10355
rect 4755 10325 4760 10355
rect 4720 10270 4760 10325
rect 4720 10250 4730 10270
rect 4750 10250 4760 10270
rect 4720 10190 4760 10250
rect 4720 10170 4730 10190
rect 4750 10170 4760 10190
rect 4720 10110 4760 10170
rect 4720 10090 4730 10110
rect 4750 10090 4760 10110
rect 4720 10030 4760 10090
rect 4720 10010 4730 10030
rect 4750 10010 4760 10030
rect 4720 9955 4760 10010
rect 4720 9925 4725 9955
rect 4755 9925 4760 9955
rect 4720 9875 4760 9925
rect 4720 9845 4725 9875
rect 4755 9845 4760 9875
rect 4720 9795 4760 9845
rect 4720 9765 4725 9795
rect 4755 9765 4760 9795
rect 4720 9715 4760 9765
rect 4720 9685 4725 9715
rect 4755 9685 4760 9715
rect 4720 9635 4760 9685
rect 4720 9605 4725 9635
rect 4755 9605 4760 9635
rect 4720 9555 4760 9605
rect 4720 9525 4725 9555
rect 4755 9525 4760 9555
rect 4720 9475 4760 9525
rect 4720 9445 4725 9475
rect 4755 9445 4760 9475
rect 4720 9395 4760 9445
rect 4720 9365 4725 9395
rect 4755 9365 4760 9395
rect 4720 9310 4760 9365
rect 4720 9290 4730 9310
rect 4750 9290 4760 9310
rect 4720 9230 4760 9290
rect 4720 9210 4730 9230
rect 4750 9210 4760 9230
rect 4720 9150 4760 9210
rect 4720 9130 4730 9150
rect 4750 9130 4760 9150
rect 4720 9070 4760 9130
rect 4720 9050 4730 9070
rect 4750 9050 4760 9070
rect 4720 8995 4760 9050
rect 4720 8965 4725 8995
rect 4755 8965 4760 8995
rect 4720 8915 4760 8965
rect 4720 8885 4725 8915
rect 4755 8885 4760 8915
rect 4720 8835 4760 8885
rect 4720 8805 4725 8835
rect 4755 8805 4760 8835
rect 4720 8755 4760 8805
rect 4720 8725 4725 8755
rect 4755 8725 4760 8755
rect 4720 8675 4760 8725
rect 4720 8645 4725 8675
rect 4755 8645 4760 8675
rect 4720 8595 4760 8645
rect 4720 8565 4725 8595
rect 4755 8565 4760 8595
rect 4720 8515 4760 8565
rect 4720 8485 4725 8515
rect 4755 8485 4760 8515
rect 4720 8435 4760 8485
rect 4720 8405 4725 8435
rect 4755 8405 4760 8435
rect 4720 8350 4760 8405
rect 4720 8330 4730 8350
rect 4750 8330 4760 8350
rect 4720 8275 4760 8330
rect 4720 8245 4725 8275
rect 4755 8245 4760 8275
rect 4720 8195 4760 8245
rect 4720 8165 4725 8195
rect 4755 8165 4760 8195
rect 4720 8115 4760 8165
rect 4720 8085 4725 8115
rect 4755 8085 4760 8115
rect 4720 8035 4760 8085
rect 4720 8005 4725 8035
rect 4755 8005 4760 8035
rect 4720 7955 4760 8005
rect 4720 7925 4725 7955
rect 4755 7925 4760 7955
rect 4720 7875 4760 7925
rect 4720 7845 4725 7875
rect 4755 7845 4760 7875
rect 4720 7795 4760 7845
rect 4720 7765 4725 7795
rect 4755 7765 4760 7795
rect 4720 7715 4760 7765
rect 4720 7685 4725 7715
rect 4755 7685 4760 7715
rect 4720 7635 4760 7685
rect 4720 7605 4725 7635
rect 4755 7605 4760 7635
rect 4720 7555 4760 7605
rect 4720 7525 4725 7555
rect 4755 7525 4760 7555
rect 4720 7475 4760 7525
rect 4720 7445 4725 7475
rect 4755 7445 4760 7475
rect 4720 7395 4760 7445
rect 4720 7365 4725 7395
rect 4755 7365 4760 7395
rect 4720 7315 4760 7365
rect 4720 7285 4725 7315
rect 4755 7285 4760 7315
rect 4720 7235 4760 7285
rect 4720 7205 4725 7235
rect 4755 7205 4760 7235
rect 4720 7155 4760 7205
rect 4720 7125 4725 7155
rect 4755 7125 4760 7155
rect 4720 7075 4760 7125
rect 4720 7045 4725 7075
rect 4755 7045 4760 7075
rect 4720 6995 4760 7045
rect 4720 6965 4725 6995
rect 4755 6965 4760 6995
rect 4720 6910 4760 6965
rect 4720 6890 4730 6910
rect 4750 6890 4760 6910
rect 4720 6835 4760 6890
rect 4720 6805 4725 6835
rect 4755 6805 4760 6835
rect 4720 6755 4760 6805
rect 4720 6725 4725 6755
rect 4755 6725 4760 6755
rect 4720 6675 4760 6725
rect 4720 6645 4725 6675
rect 4755 6645 4760 6675
rect 4720 6595 4760 6645
rect 4720 6565 4725 6595
rect 4755 6565 4760 6595
rect 4720 6515 4760 6565
rect 4720 6485 4725 6515
rect 4755 6485 4760 6515
rect 4720 6435 4760 6485
rect 4720 6405 4725 6435
rect 4755 6405 4760 6435
rect 4720 6355 4760 6405
rect 4720 6325 4725 6355
rect 4755 6325 4760 6355
rect 4720 6275 4760 6325
rect 4720 6245 4725 6275
rect 4755 6245 4760 6275
rect 4720 6190 4760 6245
rect 4720 6170 4730 6190
rect 4750 6170 4760 6190
rect 4720 6110 4760 6170
rect 4720 6090 4730 6110
rect 4750 6090 4760 6110
rect 4720 6030 4760 6090
rect 4720 6010 4730 6030
rect 4750 6010 4760 6030
rect 4720 5950 4760 6010
rect 4720 5930 4730 5950
rect 4750 5930 4760 5950
rect 4720 5875 4760 5930
rect 4720 5845 4725 5875
rect 4755 5845 4760 5875
rect 4720 5795 4760 5845
rect 4720 5765 4725 5795
rect 4755 5765 4760 5795
rect 4720 5715 4760 5765
rect 4720 5685 4725 5715
rect 4755 5685 4760 5715
rect 4720 5635 4760 5685
rect 4720 5605 4725 5635
rect 4755 5605 4760 5635
rect 4720 5555 4760 5605
rect 4720 5525 4725 5555
rect 4755 5525 4760 5555
rect 4720 5475 4760 5525
rect 4720 5445 4725 5475
rect 4755 5445 4760 5475
rect 4720 5395 4760 5445
rect 4720 5365 4725 5395
rect 4755 5365 4760 5395
rect 4720 5315 4760 5365
rect 4720 5285 4725 5315
rect 4755 5285 4760 5315
rect 4720 5235 4760 5285
rect 4720 5205 4725 5235
rect 4755 5205 4760 5235
rect 4720 5155 4760 5205
rect 4720 5125 4725 5155
rect 4755 5125 4760 5155
rect 4720 5075 4760 5125
rect 4720 5045 4725 5075
rect 4755 5045 4760 5075
rect 4720 4995 4760 5045
rect 4720 4965 4725 4995
rect 4755 4965 4760 4995
rect 4720 4915 4760 4965
rect 4720 4885 4725 4915
rect 4755 4885 4760 4915
rect 4720 4830 4760 4885
rect 4720 4810 4730 4830
rect 4750 4810 4760 4830
rect 4720 4755 4760 4810
rect 4720 4725 4725 4755
rect 4755 4725 4760 4755
rect 4720 4675 4760 4725
rect 4720 4645 4725 4675
rect 4755 4645 4760 4675
rect 4720 4590 4760 4645
rect 4720 4570 4730 4590
rect 4750 4570 4760 4590
rect 4720 4515 4760 4570
rect 4720 4485 4725 4515
rect 4755 4485 4760 4515
rect 4720 4435 4760 4485
rect 4720 4405 4725 4435
rect 4755 4405 4760 4435
rect 4720 4355 4760 4405
rect 4720 4325 4725 4355
rect 4755 4325 4760 4355
rect 4720 4275 4760 4325
rect 4720 4245 4725 4275
rect 4755 4245 4760 4275
rect 4720 4195 4760 4245
rect 4720 4165 4725 4195
rect 4755 4165 4760 4195
rect 4720 4115 4760 4165
rect 4720 4085 4725 4115
rect 4755 4085 4760 4115
rect 4720 4035 4760 4085
rect 4720 4005 4725 4035
rect 4755 4005 4760 4035
rect 4720 3955 4760 4005
rect 4720 3925 4725 3955
rect 4755 3925 4760 3955
rect 4720 3875 4760 3925
rect 4720 3845 4725 3875
rect 4755 3845 4760 3875
rect 4720 3790 4760 3845
rect 4720 3770 4730 3790
rect 4750 3770 4760 3790
rect 4720 3715 4760 3770
rect 4720 3685 4725 3715
rect 4755 3685 4760 3715
rect 4720 3635 4760 3685
rect 4720 3605 4725 3635
rect 4755 3605 4760 3635
rect 4720 3550 4760 3605
rect 4720 3530 4730 3550
rect 4750 3530 4760 3550
rect 4720 3475 4760 3530
rect 4720 3445 4725 3475
rect 4755 3445 4760 3475
rect 4720 3395 4760 3445
rect 4720 3365 4725 3395
rect 4755 3365 4760 3395
rect 4720 3310 4760 3365
rect 4720 3290 4730 3310
rect 4750 3290 4760 3310
rect 4720 3235 4760 3290
rect 4720 3205 4725 3235
rect 4755 3205 4760 3235
rect 4720 3155 4760 3205
rect 4720 3125 4725 3155
rect 4755 3125 4760 3155
rect 4720 3075 4760 3125
rect 4720 3045 4725 3075
rect 4755 3045 4760 3075
rect 4720 2995 4760 3045
rect 4720 2965 4725 2995
rect 4755 2965 4760 2995
rect 4720 2915 4760 2965
rect 4720 2885 4725 2915
rect 4755 2885 4760 2915
rect 4720 2835 4760 2885
rect 4720 2805 4725 2835
rect 4755 2805 4760 2835
rect 4720 2755 4760 2805
rect 4720 2725 4725 2755
rect 4755 2725 4760 2755
rect 4720 2675 4760 2725
rect 4720 2645 4725 2675
rect 4755 2645 4760 2675
rect 4720 2595 4760 2645
rect 4720 2565 4725 2595
rect 4755 2565 4760 2595
rect 4720 2515 4760 2565
rect 4720 2485 4725 2515
rect 4755 2485 4760 2515
rect 4720 2435 4760 2485
rect 4720 2405 4725 2435
rect 4755 2405 4760 2435
rect 4720 2355 4760 2405
rect 4720 2325 4725 2355
rect 4755 2325 4760 2355
rect 4720 2275 4760 2325
rect 4720 2245 4725 2275
rect 4755 2245 4760 2275
rect 4720 2195 4760 2245
rect 4720 2165 4725 2195
rect 4755 2165 4760 2195
rect 4720 2115 4760 2165
rect 4720 2085 4725 2115
rect 4755 2085 4760 2115
rect 4720 2035 4760 2085
rect 4720 2005 4725 2035
rect 4755 2005 4760 2035
rect 4720 1955 4760 2005
rect 4720 1925 4725 1955
rect 4755 1925 4760 1955
rect 4720 1870 4760 1925
rect 4720 1850 4730 1870
rect 4750 1850 4760 1870
rect 4720 1790 4760 1850
rect 4720 1770 4730 1790
rect 4750 1770 4760 1790
rect 4720 1715 4760 1770
rect 4720 1685 4725 1715
rect 4755 1685 4760 1715
rect 4720 1635 4760 1685
rect 4720 1605 4725 1635
rect 4755 1605 4760 1635
rect 4720 1555 4760 1605
rect 4720 1525 4725 1555
rect 4755 1525 4760 1555
rect 4720 1475 4760 1525
rect 4720 1445 4725 1475
rect 4755 1445 4760 1475
rect 4720 1395 4760 1445
rect 4720 1365 4725 1395
rect 4755 1365 4760 1395
rect 4720 1315 4760 1365
rect 4720 1285 4725 1315
rect 4755 1285 4760 1315
rect 4720 1235 4760 1285
rect 4720 1205 4725 1235
rect 4755 1205 4760 1235
rect 4720 1155 4760 1205
rect 4720 1125 4725 1155
rect 4755 1125 4760 1155
rect 4720 1075 4760 1125
rect 4720 1045 4725 1075
rect 4755 1045 4760 1075
rect 4720 995 4760 1045
rect 4720 965 4725 995
rect 4755 965 4760 995
rect 4720 910 4760 965
rect 4720 890 4730 910
rect 4750 890 4760 910
rect 4720 835 4760 890
rect 4720 805 4725 835
rect 4755 805 4760 835
rect 4720 755 4760 805
rect 4720 725 4725 755
rect 4755 725 4760 755
rect 4720 675 4760 725
rect 4720 645 4725 675
rect 4755 645 4760 675
rect 4720 595 4760 645
rect 4720 565 4725 595
rect 4755 565 4760 595
rect 4720 515 4760 565
rect 4720 485 4725 515
rect 4755 485 4760 515
rect 4720 430 4760 485
rect 4720 410 4730 430
rect 4750 410 4760 430
rect 4720 350 4760 410
rect 4720 330 4730 350
rect 4750 330 4760 350
rect 4720 275 4760 330
rect 4720 245 4725 275
rect 4755 245 4760 275
rect 4720 195 4760 245
rect 4720 165 4725 195
rect 4755 165 4760 195
rect 4720 115 4760 165
rect 4720 85 4725 115
rect 4755 85 4760 115
rect 4720 35 4760 85
rect 4720 5 4725 35
rect 4755 5 4760 35
rect 4720 0 4760 5
rect 4800 15710 4840 15720
rect 4800 15690 4810 15710
rect 4830 15690 4840 15710
rect 4800 15630 4840 15690
rect 4800 15610 4810 15630
rect 4830 15610 4840 15630
rect 4800 15550 4840 15610
rect 4800 15530 4810 15550
rect 4830 15530 4840 15550
rect 4800 15470 4840 15530
rect 4800 15450 4810 15470
rect 4830 15450 4840 15470
rect 4800 15390 4840 15450
rect 4800 15370 4810 15390
rect 4830 15370 4840 15390
rect 4800 15310 4840 15370
rect 4800 15290 4810 15310
rect 4830 15290 4840 15310
rect 4800 15230 4840 15290
rect 4800 15210 4810 15230
rect 4830 15210 4840 15230
rect 4800 15150 4840 15210
rect 4800 15130 4810 15150
rect 4830 15130 4840 15150
rect 4800 15070 4840 15130
rect 4800 15050 4810 15070
rect 4830 15050 4840 15070
rect 4800 14990 4840 15050
rect 4800 14970 4810 14990
rect 4830 14970 4840 14990
rect 4800 14910 4840 14970
rect 4800 14890 4810 14910
rect 4830 14890 4840 14910
rect 4800 14830 4840 14890
rect 4800 14810 4810 14830
rect 4830 14810 4840 14830
rect 4800 14750 4840 14810
rect 4800 14730 4810 14750
rect 4830 14730 4840 14750
rect 4800 14670 4840 14730
rect 4800 14650 4810 14670
rect 4830 14650 4840 14670
rect 4800 14590 4840 14650
rect 4800 14570 4810 14590
rect 4830 14570 4840 14590
rect 4800 14510 4840 14570
rect 4800 14490 4810 14510
rect 4830 14490 4840 14510
rect 4800 14430 4840 14490
rect 4800 14410 4810 14430
rect 4830 14410 4840 14430
rect 4800 14350 4840 14410
rect 4800 14330 4810 14350
rect 4830 14330 4840 14350
rect 4800 14270 4840 14330
rect 4800 14250 4810 14270
rect 4830 14250 4840 14270
rect 4800 14190 4840 14250
rect 4800 14170 4810 14190
rect 4830 14170 4840 14190
rect 4800 14110 4840 14170
rect 4800 14090 4810 14110
rect 4830 14090 4840 14110
rect 4800 14030 4840 14090
rect 4800 14010 4810 14030
rect 4830 14010 4840 14030
rect 4800 13950 4840 14010
rect 4800 13930 4810 13950
rect 4830 13930 4840 13950
rect 4800 13870 4840 13930
rect 4800 13850 4810 13870
rect 4830 13850 4840 13870
rect 4800 13790 4840 13850
rect 4800 13770 4810 13790
rect 4830 13770 4840 13790
rect 4800 13710 4840 13770
rect 4800 13690 4810 13710
rect 4830 13690 4840 13710
rect 4800 13630 4840 13690
rect 4800 13610 4810 13630
rect 4830 13610 4840 13630
rect 4800 13550 4840 13610
rect 4800 13530 4810 13550
rect 4830 13530 4840 13550
rect 4800 13470 4840 13530
rect 4800 13450 4810 13470
rect 4830 13450 4840 13470
rect 4800 13390 4840 13450
rect 4800 13370 4810 13390
rect 4830 13370 4840 13390
rect 4800 13310 4840 13370
rect 4800 13290 4810 13310
rect 4830 13290 4840 13310
rect 4800 13230 4840 13290
rect 4800 13210 4810 13230
rect 4830 13210 4840 13230
rect 4800 13150 4840 13210
rect 4800 13130 4810 13150
rect 4830 13130 4840 13150
rect 4800 13070 4840 13130
rect 4800 13050 4810 13070
rect 4830 13050 4840 13070
rect 4800 12990 4840 13050
rect 4800 12970 4810 12990
rect 4830 12970 4840 12990
rect 4800 12910 4840 12970
rect 4800 12890 4810 12910
rect 4830 12890 4840 12910
rect 4800 12830 4840 12890
rect 4800 12810 4810 12830
rect 4830 12810 4840 12830
rect 4800 12750 4840 12810
rect 4800 12730 4810 12750
rect 4830 12730 4840 12750
rect 4800 12670 4840 12730
rect 4800 12650 4810 12670
rect 4830 12650 4840 12670
rect 4800 12590 4840 12650
rect 4800 12570 4810 12590
rect 4830 12570 4840 12590
rect 4800 12510 4840 12570
rect 4800 12490 4810 12510
rect 4830 12490 4840 12510
rect 4800 12430 4840 12490
rect 4800 12410 4810 12430
rect 4830 12410 4840 12430
rect 4800 12350 4840 12410
rect 4800 12330 4810 12350
rect 4830 12330 4840 12350
rect 4800 12270 4840 12330
rect 4800 12250 4810 12270
rect 4830 12250 4840 12270
rect 4800 12190 4840 12250
rect 4800 12170 4810 12190
rect 4830 12170 4840 12190
rect 4800 12110 4840 12170
rect 4800 12090 4810 12110
rect 4830 12090 4840 12110
rect 4800 12030 4840 12090
rect 4800 12010 4810 12030
rect 4830 12010 4840 12030
rect 4800 11950 4840 12010
rect 4800 11930 4810 11950
rect 4830 11930 4840 11950
rect 4800 11870 4840 11930
rect 4800 11850 4810 11870
rect 4830 11850 4840 11870
rect 4800 11790 4840 11850
rect 4800 11770 4810 11790
rect 4830 11770 4840 11790
rect 4800 11710 4840 11770
rect 4800 11690 4810 11710
rect 4830 11690 4840 11710
rect 4800 11630 4840 11690
rect 4800 11610 4810 11630
rect 4830 11610 4840 11630
rect 4800 11550 4840 11610
rect 4800 11530 4810 11550
rect 4830 11530 4840 11550
rect 4800 11470 4840 11530
rect 4800 11450 4810 11470
rect 4830 11450 4840 11470
rect 4800 11390 4840 11450
rect 4800 11370 4810 11390
rect 4830 11370 4840 11390
rect 4800 11310 4840 11370
rect 4800 11290 4810 11310
rect 4830 11290 4840 11310
rect 4800 11230 4840 11290
rect 4800 11210 4810 11230
rect 4830 11210 4840 11230
rect 4800 11150 4840 11210
rect 4800 11130 4810 11150
rect 4830 11130 4840 11150
rect 4800 11070 4840 11130
rect 4800 11050 4810 11070
rect 4830 11050 4840 11070
rect 4800 10990 4840 11050
rect 4800 10970 4810 10990
rect 4830 10970 4840 10990
rect 4800 10910 4840 10970
rect 4800 10890 4810 10910
rect 4830 10890 4840 10910
rect 4800 10830 4840 10890
rect 4800 10810 4810 10830
rect 4830 10810 4840 10830
rect 4800 10750 4840 10810
rect 4800 10730 4810 10750
rect 4830 10730 4840 10750
rect 4800 10670 4840 10730
rect 4800 10650 4810 10670
rect 4830 10650 4840 10670
rect 4800 10590 4840 10650
rect 4800 10570 4810 10590
rect 4830 10570 4840 10590
rect 4800 10510 4840 10570
rect 4800 10490 4810 10510
rect 4830 10490 4840 10510
rect 4800 10430 4840 10490
rect 4800 10410 4810 10430
rect 4830 10410 4840 10430
rect 4800 10350 4840 10410
rect 4800 10330 4810 10350
rect 4830 10330 4840 10350
rect 4800 10270 4840 10330
rect 4800 10250 4810 10270
rect 4830 10250 4840 10270
rect 4800 10190 4840 10250
rect 4800 10170 4810 10190
rect 4830 10170 4840 10190
rect 4800 10110 4840 10170
rect 4800 10090 4810 10110
rect 4830 10090 4840 10110
rect 4800 10030 4840 10090
rect 4800 10010 4810 10030
rect 4830 10010 4840 10030
rect 4800 9950 4840 10010
rect 4800 9930 4810 9950
rect 4830 9930 4840 9950
rect 4800 9870 4840 9930
rect 4800 9850 4810 9870
rect 4830 9850 4840 9870
rect 4800 9790 4840 9850
rect 4800 9770 4810 9790
rect 4830 9770 4840 9790
rect 4800 9710 4840 9770
rect 4800 9690 4810 9710
rect 4830 9690 4840 9710
rect 4800 9630 4840 9690
rect 4800 9610 4810 9630
rect 4830 9610 4840 9630
rect 4800 9550 4840 9610
rect 4800 9530 4810 9550
rect 4830 9530 4840 9550
rect 4800 9470 4840 9530
rect 4800 9450 4810 9470
rect 4830 9450 4840 9470
rect 4800 9390 4840 9450
rect 4800 9370 4810 9390
rect 4830 9370 4840 9390
rect 4800 9310 4840 9370
rect 4800 9290 4810 9310
rect 4830 9290 4840 9310
rect 4800 9230 4840 9290
rect 4800 9210 4810 9230
rect 4830 9210 4840 9230
rect 4800 9150 4840 9210
rect 4800 9130 4810 9150
rect 4830 9130 4840 9150
rect 4800 9070 4840 9130
rect 4800 9050 4810 9070
rect 4830 9050 4840 9070
rect 4800 8990 4840 9050
rect 4800 8970 4810 8990
rect 4830 8970 4840 8990
rect 4800 8910 4840 8970
rect 4800 8890 4810 8910
rect 4830 8890 4840 8910
rect 4800 8830 4840 8890
rect 4800 8810 4810 8830
rect 4830 8810 4840 8830
rect 4800 8750 4840 8810
rect 4800 8730 4810 8750
rect 4830 8730 4840 8750
rect 4800 8670 4840 8730
rect 4800 8650 4810 8670
rect 4830 8650 4840 8670
rect 4800 8590 4840 8650
rect 4800 8570 4810 8590
rect 4830 8570 4840 8590
rect 4800 8510 4840 8570
rect 4800 8490 4810 8510
rect 4830 8490 4840 8510
rect 4800 8430 4840 8490
rect 4800 8410 4810 8430
rect 4830 8410 4840 8430
rect 4800 8350 4840 8410
rect 4800 8330 4810 8350
rect 4830 8330 4840 8350
rect 4800 8270 4840 8330
rect 4800 8250 4810 8270
rect 4830 8250 4840 8270
rect 4800 8190 4840 8250
rect 4800 8170 4810 8190
rect 4830 8170 4840 8190
rect 4800 8110 4840 8170
rect 4800 8090 4810 8110
rect 4830 8090 4840 8110
rect 4800 8030 4840 8090
rect 4800 8010 4810 8030
rect 4830 8010 4840 8030
rect 4800 7950 4840 8010
rect 4800 7930 4810 7950
rect 4830 7930 4840 7950
rect 4800 7870 4840 7930
rect 4800 7850 4810 7870
rect 4830 7850 4840 7870
rect 4800 7790 4840 7850
rect 4800 7770 4810 7790
rect 4830 7770 4840 7790
rect 4800 7710 4840 7770
rect 4800 7690 4810 7710
rect 4830 7690 4840 7710
rect 4800 7630 4840 7690
rect 4800 7610 4810 7630
rect 4830 7610 4840 7630
rect 4800 7550 4840 7610
rect 4800 7530 4810 7550
rect 4830 7530 4840 7550
rect 4800 7470 4840 7530
rect 4800 7450 4810 7470
rect 4830 7450 4840 7470
rect 4800 7390 4840 7450
rect 4800 7370 4810 7390
rect 4830 7370 4840 7390
rect 4800 7310 4840 7370
rect 4800 7290 4810 7310
rect 4830 7290 4840 7310
rect 4800 7230 4840 7290
rect 4800 7210 4810 7230
rect 4830 7210 4840 7230
rect 4800 7150 4840 7210
rect 4800 7130 4810 7150
rect 4830 7130 4840 7150
rect 4800 7070 4840 7130
rect 4800 7050 4810 7070
rect 4830 7050 4840 7070
rect 4800 6990 4840 7050
rect 4800 6970 4810 6990
rect 4830 6970 4840 6990
rect 4800 6910 4840 6970
rect 4800 6890 4810 6910
rect 4830 6890 4840 6910
rect 4800 6830 4840 6890
rect 4800 6810 4810 6830
rect 4830 6810 4840 6830
rect 4800 6750 4840 6810
rect 4800 6730 4810 6750
rect 4830 6730 4840 6750
rect 4800 6670 4840 6730
rect 4800 6650 4810 6670
rect 4830 6650 4840 6670
rect 4800 6590 4840 6650
rect 4800 6570 4810 6590
rect 4830 6570 4840 6590
rect 4800 6510 4840 6570
rect 4800 6490 4810 6510
rect 4830 6490 4840 6510
rect 4800 6430 4840 6490
rect 4800 6410 4810 6430
rect 4830 6410 4840 6430
rect 4800 6350 4840 6410
rect 4800 6330 4810 6350
rect 4830 6330 4840 6350
rect 4800 6270 4840 6330
rect 4800 6250 4810 6270
rect 4830 6250 4840 6270
rect 4800 6190 4840 6250
rect 4800 6170 4810 6190
rect 4830 6170 4840 6190
rect 4800 6110 4840 6170
rect 4800 6090 4810 6110
rect 4830 6090 4840 6110
rect 4800 6030 4840 6090
rect 4800 6010 4810 6030
rect 4830 6010 4840 6030
rect 4800 5950 4840 6010
rect 4800 5930 4810 5950
rect 4830 5930 4840 5950
rect 4800 5870 4840 5930
rect 4800 5850 4810 5870
rect 4830 5850 4840 5870
rect 4800 5790 4840 5850
rect 4800 5770 4810 5790
rect 4830 5770 4840 5790
rect 4800 5710 4840 5770
rect 4800 5690 4810 5710
rect 4830 5690 4840 5710
rect 4800 5630 4840 5690
rect 4800 5610 4810 5630
rect 4830 5610 4840 5630
rect 4800 5550 4840 5610
rect 4800 5530 4810 5550
rect 4830 5530 4840 5550
rect 4800 5470 4840 5530
rect 4800 5450 4810 5470
rect 4830 5450 4840 5470
rect 4800 5390 4840 5450
rect 4800 5370 4810 5390
rect 4830 5370 4840 5390
rect 4800 5310 4840 5370
rect 4800 5290 4810 5310
rect 4830 5290 4840 5310
rect 4800 5230 4840 5290
rect 4800 5210 4810 5230
rect 4830 5210 4840 5230
rect 4800 5150 4840 5210
rect 4800 5130 4810 5150
rect 4830 5130 4840 5150
rect 4800 5070 4840 5130
rect 4800 5050 4810 5070
rect 4830 5050 4840 5070
rect 4800 4990 4840 5050
rect 4800 4970 4810 4990
rect 4830 4970 4840 4990
rect 4800 4910 4840 4970
rect 4800 4890 4810 4910
rect 4830 4890 4840 4910
rect 4800 4830 4840 4890
rect 4800 4810 4810 4830
rect 4830 4810 4840 4830
rect 4800 4750 4840 4810
rect 4800 4730 4810 4750
rect 4830 4730 4840 4750
rect 4800 4670 4840 4730
rect 4800 4650 4810 4670
rect 4830 4650 4840 4670
rect 4800 4590 4840 4650
rect 4800 4570 4810 4590
rect 4830 4570 4840 4590
rect 4800 4510 4840 4570
rect 4800 4490 4810 4510
rect 4830 4490 4840 4510
rect 4800 4430 4840 4490
rect 4800 4410 4810 4430
rect 4830 4410 4840 4430
rect 4800 4350 4840 4410
rect 4800 4330 4810 4350
rect 4830 4330 4840 4350
rect 4800 4270 4840 4330
rect 4800 4250 4810 4270
rect 4830 4250 4840 4270
rect 4800 4190 4840 4250
rect 4800 4170 4810 4190
rect 4830 4170 4840 4190
rect 4800 4110 4840 4170
rect 4800 4090 4810 4110
rect 4830 4090 4840 4110
rect 4800 4030 4840 4090
rect 4800 4010 4810 4030
rect 4830 4010 4840 4030
rect 4800 3950 4840 4010
rect 4800 3930 4810 3950
rect 4830 3930 4840 3950
rect 4800 3870 4840 3930
rect 4800 3850 4810 3870
rect 4830 3850 4840 3870
rect 4800 3790 4840 3850
rect 4800 3770 4810 3790
rect 4830 3770 4840 3790
rect 4800 3710 4840 3770
rect 4800 3690 4810 3710
rect 4830 3690 4840 3710
rect 4800 3630 4840 3690
rect 4800 3610 4810 3630
rect 4830 3610 4840 3630
rect 4800 3550 4840 3610
rect 4800 3530 4810 3550
rect 4830 3530 4840 3550
rect 4800 3470 4840 3530
rect 4800 3450 4810 3470
rect 4830 3450 4840 3470
rect 4800 3390 4840 3450
rect 4800 3370 4810 3390
rect 4830 3370 4840 3390
rect 4800 3310 4840 3370
rect 4800 3290 4810 3310
rect 4830 3290 4840 3310
rect 4800 3230 4840 3290
rect 4800 3210 4810 3230
rect 4830 3210 4840 3230
rect 4800 3150 4840 3210
rect 4800 3130 4810 3150
rect 4830 3130 4840 3150
rect 4800 3070 4840 3130
rect 4800 3050 4810 3070
rect 4830 3050 4840 3070
rect 4800 2990 4840 3050
rect 4800 2970 4810 2990
rect 4830 2970 4840 2990
rect 4800 2910 4840 2970
rect 4800 2890 4810 2910
rect 4830 2890 4840 2910
rect 4800 2830 4840 2890
rect 4800 2810 4810 2830
rect 4830 2810 4840 2830
rect 4800 2750 4840 2810
rect 4800 2730 4810 2750
rect 4830 2730 4840 2750
rect 4800 2670 4840 2730
rect 4800 2650 4810 2670
rect 4830 2650 4840 2670
rect 4800 2590 4840 2650
rect 4800 2570 4810 2590
rect 4830 2570 4840 2590
rect 4800 2510 4840 2570
rect 4800 2490 4810 2510
rect 4830 2490 4840 2510
rect 4800 2430 4840 2490
rect 4800 2410 4810 2430
rect 4830 2410 4840 2430
rect 4800 2350 4840 2410
rect 4800 2330 4810 2350
rect 4830 2330 4840 2350
rect 4800 2270 4840 2330
rect 4800 2250 4810 2270
rect 4830 2250 4840 2270
rect 4800 2190 4840 2250
rect 4800 2170 4810 2190
rect 4830 2170 4840 2190
rect 4800 2110 4840 2170
rect 4800 2090 4810 2110
rect 4830 2090 4840 2110
rect 4800 2030 4840 2090
rect 4800 2010 4810 2030
rect 4830 2010 4840 2030
rect 4800 1950 4840 2010
rect 4800 1930 4810 1950
rect 4830 1930 4840 1950
rect 4800 1870 4840 1930
rect 4800 1850 4810 1870
rect 4830 1850 4840 1870
rect 4800 1790 4840 1850
rect 4800 1770 4810 1790
rect 4830 1770 4840 1790
rect 4800 1710 4840 1770
rect 4800 1690 4810 1710
rect 4830 1690 4840 1710
rect 4800 1630 4840 1690
rect 4800 1610 4810 1630
rect 4830 1610 4840 1630
rect 4800 1550 4840 1610
rect 4800 1530 4810 1550
rect 4830 1530 4840 1550
rect 4800 1470 4840 1530
rect 4800 1450 4810 1470
rect 4830 1450 4840 1470
rect 4800 1390 4840 1450
rect 4800 1370 4810 1390
rect 4830 1370 4840 1390
rect 4800 1310 4840 1370
rect 4800 1290 4810 1310
rect 4830 1290 4840 1310
rect 4800 1230 4840 1290
rect 4800 1210 4810 1230
rect 4830 1210 4840 1230
rect 4800 1150 4840 1210
rect 4800 1130 4810 1150
rect 4830 1130 4840 1150
rect 4800 1070 4840 1130
rect 4800 1050 4810 1070
rect 4830 1050 4840 1070
rect 4800 990 4840 1050
rect 4800 970 4810 990
rect 4830 970 4840 990
rect 4800 910 4840 970
rect 4800 890 4810 910
rect 4830 890 4840 910
rect 4800 830 4840 890
rect 4800 810 4810 830
rect 4830 810 4840 830
rect 4800 750 4840 810
rect 4800 730 4810 750
rect 4830 730 4840 750
rect 4800 670 4840 730
rect 4800 650 4810 670
rect 4830 650 4840 670
rect 4800 590 4840 650
rect 4800 570 4810 590
rect 4830 570 4840 590
rect 4800 510 4840 570
rect 4800 490 4810 510
rect 4830 490 4840 510
rect 4800 430 4840 490
rect 4800 410 4810 430
rect 4830 410 4840 430
rect 4800 350 4840 410
rect 4800 330 4810 350
rect 4830 330 4840 350
rect 4800 270 4840 330
rect 4800 250 4810 270
rect 4830 250 4840 270
rect 4800 190 4840 250
rect 4800 170 4810 190
rect 4830 170 4840 190
rect 4800 110 4840 170
rect 4800 90 4810 110
rect 4830 90 4840 110
rect 4800 30 4840 90
rect 4800 10 4810 30
rect 4830 10 4840 30
rect 4800 0 4840 10
rect 4880 15715 4920 15720
rect 4880 15685 4885 15715
rect 4915 15685 4920 15715
rect 4880 15635 4920 15685
rect 4880 15605 4885 15635
rect 4915 15605 4920 15635
rect 4880 15555 4920 15605
rect 4880 15525 4885 15555
rect 4915 15525 4920 15555
rect 4880 15475 4920 15525
rect 4880 15445 4885 15475
rect 4915 15445 4920 15475
rect 4880 15395 4920 15445
rect 4880 15365 4885 15395
rect 4915 15365 4920 15395
rect 4880 15315 4920 15365
rect 4880 15285 4885 15315
rect 4915 15285 4920 15315
rect 4880 15235 4920 15285
rect 4880 15205 4885 15235
rect 4915 15205 4920 15235
rect 4880 15155 4920 15205
rect 4880 15125 4885 15155
rect 4915 15125 4920 15155
rect 4880 15070 4920 15125
rect 4880 15050 4890 15070
rect 4910 15050 4920 15070
rect 4880 14995 4920 15050
rect 4880 14965 4885 14995
rect 4915 14965 4920 14995
rect 4880 14915 4920 14965
rect 4880 14885 4885 14915
rect 4915 14885 4920 14915
rect 4880 14835 4920 14885
rect 4880 14805 4885 14835
rect 4915 14805 4920 14835
rect 4880 14755 4920 14805
rect 4880 14725 4885 14755
rect 4915 14725 4920 14755
rect 4880 14675 4920 14725
rect 4880 14645 4885 14675
rect 4915 14645 4920 14675
rect 4880 14595 4920 14645
rect 4880 14565 4885 14595
rect 4915 14565 4920 14595
rect 4880 14515 4920 14565
rect 4880 14485 4885 14515
rect 4915 14485 4920 14515
rect 4880 14435 4920 14485
rect 4880 14405 4885 14435
rect 4915 14405 4920 14435
rect 4880 14350 4920 14405
rect 4880 14330 4890 14350
rect 4910 14330 4920 14350
rect 4880 14270 4920 14330
rect 4880 14250 4890 14270
rect 4910 14250 4920 14270
rect 4880 14190 4920 14250
rect 4880 14170 4890 14190
rect 4910 14170 4920 14190
rect 4880 14110 4920 14170
rect 4880 14090 4890 14110
rect 4910 14090 4920 14110
rect 4880 14035 4920 14090
rect 4880 14005 4885 14035
rect 4915 14005 4920 14035
rect 4880 13955 4920 14005
rect 4880 13925 4885 13955
rect 4915 13925 4920 13955
rect 4880 13875 4920 13925
rect 4880 13845 4885 13875
rect 4915 13845 4920 13875
rect 4880 13795 4920 13845
rect 4880 13765 4885 13795
rect 4915 13765 4920 13795
rect 4880 13715 4920 13765
rect 4880 13685 4885 13715
rect 4915 13685 4920 13715
rect 4880 13635 4920 13685
rect 4880 13605 4885 13635
rect 4915 13605 4920 13635
rect 4880 13555 4920 13605
rect 4880 13525 4885 13555
rect 4915 13525 4920 13555
rect 4880 13475 4920 13525
rect 4880 13445 4885 13475
rect 4915 13445 4920 13475
rect 4880 13390 4920 13445
rect 4880 13370 4890 13390
rect 4910 13370 4920 13390
rect 4880 13310 4920 13370
rect 4880 13290 4890 13310
rect 4910 13290 4920 13310
rect 4880 13230 4920 13290
rect 4880 13210 4890 13230
rect 4910 13210 4920 13230
rect 4880 13150 4920 13210
rect 4880 13130 4890 13150
rect 4910 13130 4920 13150
rect 4880 13075 4920 13130
rect 4880 13045 4885 13075
rect 4915 13045 4920 13075
rect 4880 12995 4920 13045
rect 4880 12965 4885 12995
rect 4915 12965 4920 12995
rect 4880 12915 4920 12965
rect 4880 12885 4885 12915
rect 4915 12885 4920 12915
rect 4880 12835 4920 12885
rect 4880 12805 4885 12835
rect 4915 12805 4920 12835
rect 4880 12755 4920 12805
rect 4880 12725 4885 12755
rect 4915 12725 4920 12755
rect 4880 12675 4920 12725
rect 4880 12645 4885 12675
rect 4915 12645 4920 12675
rect 4880 12595 4920 12645
rect 4880 12565 4885 12595
rect 4915 12565 4920 12595
rect 4880 12515 4920 12565
rect 4880 12485 4885 12515
rect 4915 12485 4920 12515
rect 4880 12430 4920 12485
rect 4880 12410 4890 12430
rect 4910 12410 4920 12430
rect 4880 12355 4920 12410
rect 4880 12325 4885 12355
rect 4915 12325 4920 12355
rect 4880 12275 4920 12325
rect 4880 12245 4885 12275
rect 4915 12245 4920 12275
rect 4880 12195 4920 12245
rect 4880 12165 4885 12195
rect 4915 12165 4920 12195
rect 4880 12115 4920 12165
rect 4880 12085 4885 12115
rect 4915 12085 4920 12115
rect 4880 12035 4920 12085
rect 4880 12005 4885 12035
rect 4915 12005 4920 12035
rect 4880 11955 4920 12005
rect 4880 11925 4885 11955
rect 4915 11925 4920 11955
rect 4880 11875 4920 11925
rect 4880 11845 4885 11875
rect 4915 11845 4920 11875
rect 4880 11795 4920 11845
rect 4880 11765 4885 11795
rect 4915 11765 4920 11795
rect 4880 11715 4920 11765
rect 4880 11685 4885 11715
rect 4915 11685 4920 11715
rect 4880 11635 4920 11685
rect 4880 11605 4885 11635
rect 4915 11605 4920 11635
rect 4880 11555 4920 11605
rect 4880 11525 4885 11555
rect 4915 11525 4920 11555
rect 4880 11475 4920 11525
rect 4880 11445 4885 11475
rect 4915 11445 4920 11475
rect 4880 11395 4920 11445
rect 4880 11365 4885 11395
rect 4915 11365 4920 11395
rect 4880 11315 4920 11365
rect 4880 11285 4885 11315
rect 4915 11285 4920 11315
rect 4880 11235 4920 11285
rect 4880 11205 4885 11235
rect 4915 11205 4920 11235
rect 4880 11155 4920 11205
rect 4880 11125 4885 11155
rect 4915 11125 4920 11155
rect 4880 11075 4920 11125
rect 4880 11045 4885 11075
rect 4915 11045 4920 11075
rect 4880 10990 4920 11045
rect 4880 10970 4890 10990
rect 4910 10970 4920 10990
rect 4880 10915 4920 10970
rect 4880 10885 4885 10915
rect 4915 10885 4920 10915
rect 4880 10835 4920 10885
rect 4880 10805 4885 10835
rect 4915 10805 4920 10835
rect 4880 10755 4920 10805
rect 4880 10725 4885 10755
rect 4915 10725 4920 10755
rect 4880 10675 4920 10725
rect 4880 10645 4885 10675
rect 4915 10645 4920 10675
rect 4880 10595 4920 10645
rect 4880 10565 4885 10595
rect 4915 10565 4920 10595
rect 4880 10515 4920 10565
rect 4880 10485 4885 10515
rect 4915 10485 4920 10515
rect 4880 10435 4920 10485
rect 4880 10405 4885 10435
rect 4915 10405 4920 10435
rect 4880 10355 4920 10405
rect 4880 10325 4885 10355
rect 4915 10325 4920 10355
rect 4880 10270 4920 10325
rect 4880 10250 4890 10270
rect 4910 10250 4920 10270
rect 4880 10190 4920 10250
rect 4880 10170 4890 10190
rect 4910 10170 4920 10190
rect 4880 10110 4920 10170
rect 4880 10090 4890 10110
rect 4910 10090 4920 10110
rect 4880 10030 4920 10090
rect 4880 10010 4890 10030
rect 4910 10010 4920 10030
rect 4880 9955 4920 10010
rect 4880 9925 4885 9955
rect 4915 9925 4920 9955
rect 4880 9875 4920 9925
rect 4880 9845 4885 9875
rect 4915 9845 4920 9875
rect 4880 9795 4920 9845
rect 4880 9765 4885 9795
rect 4915 9765 4920 9795
rect 4880 9715 4920 9765
rect 4880 9685 4885 9715
rect 4915 9685 4920 9715
rect 4880 9635 4920 9685
rect 4880 9605 4885 9635
rect 4915 9605 4920 9635
rect 4880 9555 4920 9605
rect 4880 9525 4885 9555
rect 4915 9525 4920 9555
rect 4880 9475 4920 9525
rect 4880 9445 4885 9475
rect 4915 9445 4920 9475
rect 4880 9395 4920 9445
rect 4880 9365 4885 9395
rect 4915 9365 4920 9395
rect 4880 9310 4920 9365
rect 4880 9290 4890 9310
rect 4910 9290 4920 9310
rect 4880 9230 4920 9290
rect 4880 9210 4890 9230
rect 4910 9210 4920 9230
rect 4880 9150 4920 9210
rect 4880 9130 4890 9150
rect 4910 9130 4920 9150
rect 4880 9070 4920 9130
rect 4880 9050 4890 9070
rect 4910 9050 4920 9070
rect 4880 8995 4920 9050
rect 4880 8965 4885 8995
rect 4915 8965 4920 8995
rect 4880 8915 4920 8965
rect 4880 8885 4885 8915
rect 4915 8885 4920 8915
rect 4880 8835 4920 8885
rect 4880 8805 4885 8835
rect 4915 8805 4920 8835
rect 4880 8755 4920 8805
rect 4880 8725 4885 8755
rect 4915 8725 4920 8755
rect 4880 8675 4920 8725
rect 4880 8645 4885 8675
rect 4915 8645 4920 8675
rect 4880 8595 4920 8645
rect 4880 8565 4885 8595
rect 4915 8565 4920 8595
rect 4880 8515 4920 8565
rect 4880 8485 4885 8515
rect 4915 8485 4920 8515
rect 4880 8435 4920 8485
rect 4880 8405 4885 8435
rect 4915 8405 4920 8435
rect 4880 8350 4920 8405
rect 4880 8330 4890 8350
rect 4910 8330 4920 8350
rect 4880 8275 4920 8330
rect 4880 8245 4885 8275
rect 4915 8245 4920 8275
rect 4880 8195 4920 8245
rect 4880 8165 4885 8195
rect 4915 8165 4920 8195
rect 4880 8115 4920 8165
rect 4880 8085 4885 8115
rect 4915 8085 4920 8115
rect 4880 8035 4920 8085
rect 4880 8005 4885 8035
rect 4915 8005 4920 8035
rect 4880 7955 4920 8005
rect 4880 7925 4885 7955
rect 4915 7925 4920 7955
rect 4880 7875 4920 7925
rect 4880 7845 4885 7875
rect 4915 7845 4920 7875
rect 4880 7795 4920 7845
rect 4880 7765 4885 7795
rect 4915 7765 4920 7795
rect 4880 7715 4920 7765
rect 4880 7685 4885 7715
rect 4915 7685 4920 7715
rect 4880 7635 4920 7685
rect 4880 7605 4885 7635
rect 4915 7605 4920 7635
rect 4880 7555 4920 7605
rect 4880 7525 4885 7555
rect 4915 7525 4920 7555
rect 4880 7475 4920 7525
rect 4880 7445 4885 7475
rect 4915 7445 4920 7475
rect 4880 7395 4920 7445
rect 4880 7365 4885 7395
rect 4915 7365 4920 7395
rect 4880 7315 4920 7365
rect 4880 7285 4885 7315
rect 4915 7285 4920 7315
rect 4880 7235 4920 7285
rect 4880 7205 4885 7235
rect 4915 7205 4920 7235
rect 4880 7155 4920 7205
rect 4880 7125 4885 7155
rect 4915 7125 4920 7155
rect 4880 7075 4920 7125
rect 4880 7045 4885 7075
rect 4915 7045 4920 7075
rect 4880 6995 4920 7045
rect 4880 6965 4885 6995
rect 4915 6965 4920 6995
rect 4880 6910 4920 6965
rect 4880 6890 4890 6910
rect 4910 6890 4920 6910
rect 4880 6835 4920 6890
rect 4880 6805 4885 6835
rect 4915 6805 4920 6835
rect 4880 6755 4920 6805
rect 4880 6725 4885 6755
rect 4915 6725 4920 6755
rect 4880 6675 4920 6725
rect 4880 6645 4885 6675
rect 4915 6645 4920 6675
rect 4880 6595 4920 6645
rect 4880 6565 4885 6595
rect 4915 6565 4920 6595
rect 4880 6515 4920 6565
rect 4880 6485 4885 6515
rect 4915 6485 4920 6515
rect 4880 6435 4920 6485
rect 4880 6405 4885 6435
rect 4915 6405 4920 6435
rect 4880 6355 4920 6405
rect 4880 6325 4885 6355
rect 4915 6325 4920 6355
rect 4880 6275 4920 6325
rect 4880 6245 4885 6275
rect 4915 6245 4920 6275
rect 4880 6190 4920 6245
rect 4880 6170 4890 6190
rect 4910 6170 4920 6190
rect 4880 6110 4920 6170
rect 4880 6090 4890 6110
rect 4910 6090 4920 6110
rect 4880 6030 4920 6090
rect 4880 6010 4890 6030
rect 4910 6010 4920 6030
rect 4880 5950 4920 6010
rect 4880 5930 4890 5950
rect 4910 5930 4920 5950
rect 4880 5875 4920 5930
rect 4880 5845 4885 5875
rect 4915 5845 4920 5875
rect 4880 5795 4920 5845
rect 4880 5765 4885 5795
rect 4915 5765 4920 5795
rect 4880 5715 4920 5765
rect 4880 5685 4885 5715
rect 4915 5685 4920 5715
rect 4880 5635 4920 5685
rect 4880 5605 4885 5635
rect 4915 5605 4920 5635
rect 4880 5555 4920 5605
rect 4880 5525 4885 5555
rect 4915 5525 4920 5555
rect 4880 5475 4920 5525
rect 4880 5445 4885 5475
rect 4915 5445 4920 5475
rect 4880 5395 4920 5445
rect 4880 5365 4885 5395
rect 4915 5365 4920 5395
rect 4880 5315 4920 5365
rect 4880 5285 4885 5315
rect 4915 5285 4920 5315
rect 4880 5235 4920 5285
rect 4880 5205 4885 5235
rect 4915 5205 4920 5235
rect 4880 5155 4920 5205
rect 4880 5125 4885 5155
rect 4915 5125 4920 5155
rect 4880 5075 4920 5125
rect 4880 5045 4885 5075
rect 4915 5045 4920 5075
rect 4880 4995 4920 5045
rect 4880 4965 4885 4995
rect 4915 4965 4920 4995
rect 4880 4915 4920 4965
rect 4880 4885 4885 4915
rect 4915 4885 4920 4915
rect 4880 4830 4920 4885
rect 4880 4810 4890 4830
rect 4910 4810 4920 4830
rect 4880 4755 4920 4810
rect 4880 4725 4885 4755
rect 4915 4725 4920 4755
rect 4880 4675 4920 4725
rect 4880 4645 4885 4675
rect 4915 4645 4920 4675
rect 4880 4590 4920 4645
rect 4880 4570 4890 4590
rect 4910 4570 4920 4590
rect 4880 4515 4920 4570
rect 4880 4485 4885 4515
rect 4915 4485 4920 4515
rect 4880 4435 4920 4485
rect 4880 4405 4885 4435
rect 4915 4405 4920 4435
rect 4880 4355 4920 4405
rect 4880 4325 4885 4355
rect 4915 4325 4920 4355
rect 4880 4275 4920 4325
rect 4880 4245 4885 4275
rect 4915 4245 4920 4275
rect 4880 4195 4920 4245
rect 4880 4165 4885 4195
rect 4915 4165 4920 4195
rect 4880 4115 4920 4165
rect 4880 4085 4885 4115
rect 4915 4085 4920 4115
rect 4880 4035 4920 4085
rect 4880 4005 4885 4035
rect 4915 4005 4920 4035
rect 4880 3955 4920 4005
rect 4880 3925 4885 3955
rect 4915 3925 4920 3955
rect 4880 3875 4920 3925
rect 4880 3845 4885 3875
rect 4915 3845 4920 3875
rect 4880 3790 4920 3845
rect 4880 3770 4890 3790
rect 4910 3770 4920 3790
rect 4880 3715 4920 3770
rect 4880 3685 4885 3715
rect 4915 3685 4920 3715
rect 4880 3635 4920 3685
rect 4880 3605 4885 3635
rect 4915 3605 4920 3635
rect 4880 3550 4920 3605
rect 4880 3530 4890 3550
rect 4910 3530 4920 3550
rect 4880 3475 4920 3530
rect 4880 3445 4885 3475
rect 4915 3445 4920 3475
rect 4880 3395 4920 3445
rect 4880 3365 4885 3395
rect 4915 3365 4920 3395
rect 4880 3310 4920 3365
rect 4880 3290 4890 3310
rect 4910 3290 4920 3310
rect 4880 3235 4920 3290
rect 4880 3205 4885 3235
rect 4915 3205 4920 3235
rect 4880 3155 4920 3205
rect 4880 3125 4885 3155
rect 4915 3125 4920 3155
rect 4880 3075 4920 3125
rect 4880 3045 4885 3075
rect 4915 3045 4920 3075
rect 4880 2995 4920 3045
rect 4880 2965 4885 2995
rect 4915 2965 4920 2995
rect 4880 2915 4920 2965
rect 4880 2885 4885 2915
rect 4915 2885 4920 2915
rect 4880 2835 4920 2885
rect 4880 2805 4885 2835
rect 4915 2805 4920 2835
rect 4880 2755 4920 2805
rect 4880 2725 4885 2755
rect 4915 2725 4920 2755
rect 4880 2675 4920 2725
rect 4880 2645 4885 2675
rect 4915 2645 4920 2675
rect 4880 2595 4920 2645
rect 4880 2565 4885 2595
rect 4915 2565 4920 2595
rect 4880 2515 4920 2565
rect 4880 2485 4885 2515
rect 4915 2485 4920 2515
rect 4880 2435 4920 2485
rect 4880 2405 4885 2435
rect 4915 2405 4920 2435
rect 4880 2355 4920 2405
rect 4880 2325 4885 2355
rect 4915 2325 4920 2355
rect 4880 2275 4920 2325
rect 4880 2245 4885 2275
rect 4915 2245 4920 2275
rect 4880 2195 4920 2245
rect 4880 2165 4885 2195
rect 4915 2165 4920 2195
rect 4880 2115 4920 2165
rect 4880 2085 4885 2115
rect 4915 2085 4920 2115
rect 4880 2035 4920 2085
rect 4880 2005 4885 2035
rect 4915 2005 4920 2035
rect 4880 1955 4920 2005
rect 4880 1925 4885 1955
rect 4915 1925 4920 1955
rect 4880 1870 4920 1925
rect 4880 1850 4890 1870
rect 4910 1850 4920 1870
rect 4880 1790 4920 1850
rect 4880 1770 4890 1790
rect 4910 1770 4920 1790
rect 4880 1715 4920 1770
rect 4880 1685 4885 1715
rect 4915 1685 4920 1715
rect 4880 1635 4920 1685
rect 4880 1605 4885 1635
rect 4915 1605 4920 1635
rect 4880 1555 4920 1605
rect 4880 1525 4885 1555
rect 4915 1525 4920 1555
rect 4880 1475 4920 1525
rect 4880 1445 4885 1475
rect 4915 1445 4920 1475
rect 4880 1395 4920 1445
rect 4880 1365 4885 1395
rect 4915 1365 4920 1395
rect 4880 1315 4920 1365
rect 4880 1285 4885 1315
rect 4915 1285 4920 1315
rect 4880 1235 4920 1285
rect 4880 1205 4885 1235
rect 4915 1205 4920 1235
rect 4880 1155 4920 1205
rect 4880 1125 4885 1155
rect 4915 1125 4920 1155
rect 4880 1075 4920 1125
rect 4880 1045 4885 1075
rect 4915 1045 4920 1075
rect 4880 995 4920 1045
rect 4880 965 4885 995
rect 4915 965 4920 995
rect 4880 910 4920 965
rect 4880 890 4890 910
rect 4910 890 4920 910
rect 4880 835 4920 890
rect 4880 805 4885 835
rect 4915 805 4920 835
rect 4880 755 4920 805
rect 4880 725 4885 755
rect 4915 725 4920 755
rect 4880 675 4920 725
rect 4880 645 4885 675
rect 4915 645 4920 675
rect 4880 595 4920 645
rect 4880 565 4885 595
rect 4915 565 4920 595
rect 4880 515 4920 565
rect 4880 485 4885 515
rect 4915 485 4920 515
rect 4880 430 4920 485
rect 4880 410 4890 430
rect 4910 410 4920 430
rect 4880 350 4920 410
rect 4880 330 4890 350
rect 4910 330 4920 350
rect 4880 275 4920 330
rect 4880 245 4885 275
rect 4915 245 4920 275
rect 4880 195 4920 245
rect 4880 165 4885 195
rect 4915 165 4920 195
rect 4880 115 4920 165
rect 4880 85 4885 115
rect 4915 85 4920 115
rect 4880 35 4920 85
rect 4880 5 4885 35
rect 4915 5 4920 35
rect 4880 0 4920 5
rect 4960 15710 5000 15720
rect 4960 15690 4970 15710
rect 4990 15690 5000 15710
rect 4960 15630 5000 15690
rect 4960 15610 4970 15630
rect 4990 15610 5000 15630
rect 4960 15550 5000 15610
rect 4960 15530 4970 15550
rect 4990 15530 5000 15550
rect 4960 15470 5000 15530
rect 4960 15450 4970 15470
rect 4990 15450 5000 15470
rect 4960 15390 5000 15450
rect 4960 15370 4970 15390
rect 4990 15370 5000 15390
rect 4960 15310 5000 15370
rect 4960 15290 4970 15310
rect 4990 15290 5000 15310
rect 4960 15230 5000 15290
rect 4960 15210 4970 15230
rect 4990 15210 5000 15230
rect 4960 15150 5000 15210
rect 4960 15130 4970 15150
rect 4990 15130 5000 15150
rect 4960 15070 5000 15130
rect 4960 15050 4970 15070
rect 4990 15050 5000 15070
rect 4960 14990 5000 15050
rect 4960 14970 4970 14990
rect 4990 14970 5000 14990
rect 4960 14910 5000 14970
rect 4960 14890 4970 14910
rect 4990 14890 5000 14910
rect 4960 14830 5000 14890
rect 4960 14810 4970 14830
rect 4990 14810 5000 14830
rect 4960 14750 5000 14810
rect 4960 14730 4970 14750
rect 4990 14730 5000 14750
rect 4960 14670 5000 14730
rect 4960 14650 4970 14670
rect 4990 14650 5000 14670
rect 4960 14590 5000 14650
rect 4960 14570 4970 14590
rect 4990 14570 5000 14590
rect 4960 14510 5000 14570
rect 4960 14490 4970 14510
rect 4990 14490 5000 14510
rect 4960 14430 5000 14490
rect 4960 14410 4970 14430
rect 4990 14410 5000 14430
rect 4960 14350 5000 14410
rect 4960 14330 4970 14350
rect 4990 14330 5000 14350
rect 4960 14270 5000 14330
rect 4960 14250 4970 14270
rect 4990 14250 5000 14270
rect 4960 14190 5000 14250
rect 4960 14170 4970 14190
rect 4990 14170 5000 14190
rect 4960 14110 5000 14170
rect 4960 14090 4970 14110
rect 4990 14090 5000 14110
rect 4960 14030 5000 14090
rect 4960 14010 4970 14030
rect 4990 14010 5000 14030
rect 4960 13950 5000 14010
rect 4960 13930 4970 13950
rect 4990 13930 5000 13950
rect 4960 13870 5000 13930
rect 4960 13850 4970 13870
rect 4990 13850 5000 13870
rect 4960 13790 5000 13850
rect 4960 13770 4970 13790
rect 4990 13770 5000 13790
rect 4960 13710 5000 13770
rect 4960 13690 4970 13710
rect 4990 13690 5000 13710
rect 4960 13630 5000 13690
rect 4960 13610 4970 13630
rect 4990 13610 5000 13630
rect 4960 13550 5000 13610
rect 4960 13530 4970 13550
rect 4990 13530 5000 13550
rect 4960 13470 5000 13530
rect 4960 13450 4970 13470
rect 4990 13450 5000 13470
rect 4960 13390 5000 13450
rect 4960 13370 4970 13390
rect 4990 13370 5000 13390
rect 4960 13310 5000 13370
rect 4960 13290 4970 13310
rect 4990 13290 5000 13310
rect 4960 13230 5000 13290
rect 4960 13210 4970 13230
rect 4990 13210 5000 13230
rect 4960 13150 5000 13210
rect 4960 13130 4970 13150
rect 4990 13130 5000 13150
rect 4960 13070 5000 13130
rect 4960 13050 4970 13070
rect 4990 13050 5000 13070
rect 4960 12990 5000 13050
rect 4960 12970 4970 12990
rect 4990 12970 5000 12990
rect 4960 12910 5000 12970
rect 4960 12890 4970 12910
rect 4990 12890 5000 12910
rect 4960 12830 5000 12890
rect 4960 12810 4970 12830
rect 4990 12810 5000 12830
rect 4960 12750 5000 12810
rect 4960 12730 4970 12750
rect 4990 12730 5000 12750
rect 4960 12670 5000 12730
rect 4960 12650 4970 12670
rect 4990 12650 5000 12670
rect 4960 12590 5000 12650
rect 4960 12570 4970 12590
rect 4990 12570 5000 12590
rect 4960 12510 5000 12570
rect 4960 12490 4970 12510
rect 4990 12490 5000 12510
rect 4960 12430 5000 12490
rect 4960 12410 4970 12430
rect 4990 12410 5000 12430
rect 4960 12350 5000 12410
rect 4960 12330 4970 12350
rect 4990 12330 5000 12350
rect 4960 12270 5000 12330
rect 4960 12250 4970 12270
rect 4990 12250 5000 12270
rect 4960 12190 5000 12250
rect 4960 12170 4970 12190
rect 4990 12170 5000 12190
rect 4960 12110 5000 12170
rect 4960 12090 4970 12110
rect 4990 12090 5000 12110
rect 4960 12030 5000 12090
rect 4960 12010 4970 12030
rect 4990 12010 5000 12030
rect 4960 11950 5000 12010
rect 4960 11930 4970 11950
rect 4990 11930 5000 11950
rect 4960 11870 5000 11930
rect 4960 11850 4970 11870
rect 4990 11850 5000 11870
rect 4960 11790 5000 11850
rect 4960 11770 4970 11790
rect 4990 11770 5000 11790
rect 4960 11710 5000 11770
rect 4960 11690 4970 11710
rect 4990 11690 5000 11710
rect 4960 11630 5000 11690
rect 4960 11610 4970 11630
rect 4990 11610 5000 11630
rect 4960 11550 5000 11610
rect 4960 11530 4970 11550
rect 4990 11530 5000 11550
rect 4960 11470 5000 11530
rect 4960 11450 4970 11470
rect 4990 11450 5000 11470
rect 4960 11390 5000 11450
rect 4960 11370 4970 11390
rect 4990 11370 5000 11390
rect 4960 11310 5000 11370
rect 4960 11290 4970 11310
rect 4990 11290 5000 11310
rect 4960 11230 5000 11290
rect 4960 11210 4970 11230
rect 4990 11210 5000 11230
rect 4960 11150 5000 11210
rect 4960 11130 4970 11150
rect 4990 11130 5000 11150
rect 4960 11070 5000 11130
rect 4960 11050 4970 11070
rect 4990 11050 5000 11070
rect 4960 10990 5000 11050
rect 4960 10970 4970 10990
rect 4990 10970 5000 10990
rect 4960 10910 5000 10970
rect 4960 10890 4970 10910
rect 4990 10890 5000 10910
rect 4960 10830 5000 10890
rect 4960 10810 4970 10830
rect 4990 10810 5000 10830
rect 4960 10750 5000 10810
rect 4960 10730 4970 10750
rect 4990 10730 5000 10750
rect 4960 10670 5000 10730
rect 4960 10650 4970 10670
rect 4990 10650 5000 10670
rect 4960 10590 5000 10650
rect 4960 10570 4970 10590
rect 4990 10570 5000 10590
rect 4960 10510 5000 10570
rect 4960 10490 4970 10510
rect 4990 10490 5000 10510
rect 4960 10430 5000 10490
rect 4960 10410 4970 10430
rect 4990 10410 5000 10430
rect 4960 10350 5000 10410
rect 4960 10330 4970 10350
rect 4990 10330 5000 10350
rect 4960 10270 5000 10330
rect 4960 10250 4970 10270
rect 4990 10250 5000 10270
rect 4960 10190 5000 10250
rect 4960 10170 4970 10190
rect 4990 10170 5000 10190
rect 4960 10110 5000 10170
rect 4960 10090 4970 10110
rect 4990 10090 5000 10110
rect 4960 10030 5000 10090
rect 4960 10010 4970 10030
rect 4990 10010 5000 10030
rect 4960 9950 5000 10010
rect 4960 9930 4970 9950
rect 4990 9930 5000 9950
rect 4960 9870 5000 9930
rect 4960 9850 4970 9870
rect 4990 9850 5000 9870
rect 4960 9790 5000 9850
rect 4960 9770 4970 9790
rect 4990 9770 5000 9790
rect 4960 9710 5000 9770
rect 4960 9690 4970 9710
rect 4990 9690 5000 9710
rect 4960 9630 5000 9690
rect 4960 9610 4970 9630
rect 4990 9610 5000 9630
rect 4960 9550 5000 9610
rect 4960 9530 4970 9550
rect 4990 9530 5000 9550
rect 4960 9470 5000 9530
rect 4960 9450 4970 9470
rect 4990 9450 5000 9470
rect 4960 9390 5000 9450
rect 4960 9370 4970 9390
rect 4990 9370 5000 9390
rect 4960 9310 5000 9370
rect 4960 9290 4970 9310
rect 4990 9290 5000 9310
rect 4960 9230 5000 9290
rect 4960 9210 4970 9230
rect 4990 9210 5000 9230
rect 4960 9150 5000 9210
rect 4960 9130 4970 9150
rect 4990 9130 5000 9150
rect 4960 9070 5000 9130
rect 4960 9050 4970 9070
rect 4990 9050 5000 9070
rect 4960 8990 5000 9050
rect 4960 8970 4970 8990
rect 4990 8970 5000 8990
rect 4960 8910 5000 8970
rect 4960 8890 4970 8910
rect 4990 8890 5000 8910
rect 4960 8830 5000 8890
rect 4960 8810 4970 8830
rect 4990 8810 5000 8830
rect 4960 8750 5000 8810
rect 4960 8730 4970 8750
rect 4990 8730 5000 8750
rect 4960 8670 5000 8730
rect 4960 8650 4970 8670
rect 4990 8650 5000 8670
rect 4960 8590 5000 8650
rect 4960 8570 4970 8590
rect 4990 8570 5000 8590
rect 4960 8510 5000 8570
rect 4960 8490 4970 8510
rect 4990 8490 5000 8510
rect 4960 8430 5000 8490
rect 4960 8410 4970 8430
rect 4990 8410 5000 8430
rect 4960 8350 5000 8410
rect 4960 8330 4970 8350
rect 4990 8330 5000 8350
rect 4960 8270 5000 8330
rect 4960 8250 4970 8270
rect 4990 8250 5000 8270
rect 4960 8190 5000 8250
rect 4960 8170 4970 8190
rect 4990 8170 5000 8190
rect 4960 8110 5000 8170
rect 4960 8090 4970 8110
rect 4990 8090 5000 8110
rect 4960 8030 5000 8090
rect 4960 8010 4970 8030
rect 4990 8010 5000 8030
rect 4960 7950 5000 8010
rect 4960 7930 4970 7950
rect 4990 7930 5000 7950
rect 4960 7870 5000 7930
rect 4960 7850 4970 7870
rect 4990 7850 5000 7870
rect 4960 7790 5000 7850
rect 4960 7770 4970 7790
rect 4990 7770 5000 7790
rect 4960 7710 5000 7770
rect 4960 7690 4970 7710
rect 4990 7690 5000 7710
rect 4960 7630 5000 7690
rect 4960 7610 4970 7630
rect 4990 7610 5000 7630
rect 4960 7550 5000 7610
rect 4960 7530 4970 7550
rect 4990 7530 5000 7550
rect 4960 7470 5000 7530
rect 4960 7450 4970 7470
rect 4990 7450 5000 7470
rect 4960 7390 5000 7450
rect 4960 7370 4970 7390
rect 4990 7370 5000 7390
rect 4960 7310 5000 7370
rect 4960 7290 4970 7310
rect 4990 7290 5000 7310
rect 4960 7230 5000 7290
rect 4960 7210 4970 7230
rect 4990 7210 5000 7230
rect 4960 7150 5000 7210
rect 4960 7130 4970 7150
rect 4990 7130 5000 7150
rect 4960 7070 5000 7130
rect 4960 7050 4970 7070
rect 4990 7050 5000 7070
rect 4960 6990 5000 7050
rect 4960 6970 4970 6990
rect 4990 6970 5000 6990
rect 4960 6910 5000 6970
rect 4960 6890 4970 6910
rect 4990 6890 5000 6910
rect 4960 6830 5000 6890
rect 4960 6810 4970 6830
rect 4990 6810 5000 6830
rect 4960 6750 5000 6810
rect 4960 6730 4970 6750
rect 4990 6730 5000 6750
rect 4960 6670 5000 6730
rect 4960 6650 4970 6670
rect 4990 6650 5000 6670
rect 4960 6590 5000 6650
rect 4960 6570 4970 6590
rect 4990 6570 5000 6590
rect 4960 6510 5000 6570
rect 4960 6490 4970 6510
rect 4990 6490 5000 6510
rect 4960 6430 5000 6490
rect 4960 6410 4970 6430
rect 4990 6410 5000 6430
rect 4960 6350 5000 6410
rect 4960 6330 4970 6350
rect 4990 6330 5000 6350
rect 4960 6270 5000 6330
rect 4960 6250 4970 6270
rect 4990 6250 5000 6270
rect 4960 6190 5000 6250
rect 4960 6170 4970 6190
rect 4990 6170 5000 6190
rect 4960 6110 5000 6170
rect 4960 6090 4970 6110
rect 4990 6090 5000 6110
rect 4960 6030 5000 6090
rect 4960 6010 4970 6030
rect 4990 6010 5000 6030
rect 4960 5950 5000 6010
rect 4960 5930 4970 5950
rect 4990 5930 5000 5950
rect 4960 5870 5000 5930
rect 4960 5850 4970 5870
rect 4990 5850 5000 5870
rect 4960 5790 5000 5850
rect 4960 5770 4970 5790
rect 4990 5770 5000 5790
rect 4960 5710 5000 5770
rect 4960 5690 4970 5710
rect 4990 5690 5000 5710
rect 4960 5630 5000 5690
rect 4960 5610 4970 5630
rect 4990 5610 5000 5630
rect 4960 5550 5000 5610
rect 4960 5530 4970 5550
rect 4990 5530 5000 5550
rect 4960 5470 5000 5530
rect 4960 5450 4970 5470
rect 4990 5450 5000 5470
rect 4960 5390 5000 5450
rect 4960 5370 4970 5390
rect 4990 5370 5000 5390
rect 4960 5310 5000 5370
rect 4960 5290 4970 5310
rect 4990 5290 5000 5310
rect 4960 5230 5000 5290
rect 4960 5210 4970 5230
rect 4990 5210 5000 5230
rect 4960 5150 5000 5210
rect 4960 5130 4970 5150
rect 4990 5130 5000 5150
rect 4960 5070 5000 5130
rect 4960 5050 4970 5070
rect 4990 5050 5000 5070
rect 4960 4990 5000 5050
rect 4960 4970 4970 4990
rect 4990 4970 5000 4990
rect 4960 4910 5000 4970
rect 4960 4890 4970 4910
rect 4990 4890 5000 4910
rect 4960 4830 5000 4890
rect 4960 4810 4970 4830
rect 4990 4810 5000 4830
rect 4960 4750 5000 4810
rect 4960 4730 4970 4750
rect 4990 4730 5000 4750
rect 4960 4670 5000 4730
rect 4960 4650 4970 4670
rect 4990 4650 5000 4670
rect 4960 4590 5000 4650
rect 4960 4570 4970 4590
rect 4990 4570 5000 4590
rect 4960 4510 5000 4570
rect 4960 4490 4970 4510
rect 4990 4490 5000 4510
rect 4960 4430 5000 4490
rect 4960 4410 4970 4430
rect 4990 4410 5000 4430
rect 4960 4350 5000 4410
rect 4960 4330 4970 4350
rect 4990 4330 5000 4350
rect 4960 4270 5000 4330
rect 4960 4250 4970 4270
rect 4990 4250 5000 4270
rect 4960 4190 5000 4250
rect 4960 4170 4970 4190
rect 4990 4170 5000 4190
rect 4960 4110 5000 4170
rect 4960 4090 4970 4110
rect 4990 4090 5000 4110
rect 4960 4030 5000 4090
rect 4960 4010 4970 4030
rect 4990 4010 5000 4030
rect 4960 3950 5000 4010
rect 4960 3930 4970 3950
rect 4990 3930 5000 3950
rect 4960 3870 5000 3930
rect 4960 3850 4970 3870
rect 4990 3850 5000 3870
rect 4960 3790 5000 3850
rect 4960 3770 4970 3790
rect 4990 3770 5000 3790
rect 4960 3710 5000 3770
rect 4960 3690 4970 3710
rect 4990 3690 5000 3710
rect 4960 3630 5000 3690
rect 4960 3610 4970 3630
rect 4990 3610 5000 3630
rect 4960 3550 5000 3610
rect 4960 3530 4970 3550
rect 4990 3530 5000 3550
rect 4960 3470 5000 3530
rect 4960 3450 4970 3470
rect 4990 3450 5000 3470
rect 4960 3390 5000 3450
rect 4960 3370 4970 3390
rect 4990 3370 5000 3390
rect 4960 3310 5000 3370
rect 4960 3290 4970 3310
rect 4990 3290 5000 3310
rect 4960 3230 5000 3290
rect 4960 3210 4970 3230
rect 4990 3210 5000 3230
rect 4960 3150 5000 3210
rect 4960 3130 4970 3150
rect 4990 3130 5000 3150
rect 4960 3070 5000 3130
rect 4960 3050 4970 3070
rect 4990 3050 5000 3070
rect 4960 2990 5000 3050
rect 4960 2970 4970 2990
rect 4990 2970 5000 2990
rect 4960 2910 5000 2970
rect 4960 2890 4970 2910
rect 4990 2890 5000 2910
rect 4960 2830 5000 2890
rect 4960 2810 4970 2830
rect 4990 2810 5000 2830
rect 4960 2750 5000 2810
rect 4960 2730 4970 2750
rect 4990 2730 5000 2750
rect 4960 2670 5000 2730
rect 4960 2650 4970 2670
rect 4990 2650 5000 2670
rect 4960 2590 5000 2650
rect 4960 2570 4970 2590
rect 4990 2570 5000 2590
rect 4960 2510 5000 2570
rect 4960 2490 4970 2510
rect 4990 2490 5000 2510
rect 4960 2430 5000 2490
rect 4960 2410 4970 2430
rect 4990 2410 5000 2430
rect 4960 2350 5000 2410
rect 4960 2330 4970 2350
rect 4990 2330 5000 2350
rect 4960 2270 5000 2330
rect 4960 2250 4970 2270
rect 4990 2250 5000 2270
rect 4960 2190 5000 2250
rect 4960 2170 4970 2190
rect 4990 2170 5000 2190
rect 4960 2110 5000 2170
rect 4960 2090 4970 2110
rect 4990 2090 5000 2110
rect 4960 2030 5000 2090
rect 4960 2010 4970 2030
rect 4990 2010 5000 2030
rect 4960 1950 5000 2010
rect 4960 1930 4970 1950
rect 4990 1930 5000 1950
rect 4960 1870 5000 1930
rect 4960 1850 4970 1870
rect 4990 1850 5000 1870
rect 4960 1790 5000 1850
rect 4960 1770 4970 1790
rect 4990 1770 5000 1790
rect 4960 1710 5000 1770
rect 4960 1690 4970 1710
rect 4990 1690 5000 1710
rect 4960 1630 5000 1690
rect 4960 1610 4970 1630
rect 4990 1610 5000 1630
rect 4960 1550 5000 1610
rect 4960 1530 4970 1550
rect 4990 1530 5000 1550
rect 4960 1470 5000 1530
rect 4960 1450 4970 1470
rect 4990 1450 5000 1470
rect 4960 1390 5000 1450
rect 4960 1370 4970 1390
rect 4990 1370 5000 1390
rect 4960 1310 5000 1370
rect 4960 1290 4970 1310
rect 4990 1290 5000 1310
rect 4960 1230 5000 1290
rect 4960 1210 4970 1230
rect 4990 1210 5000 1230
rect 4960 1150 5000 1210
rect 4960 1130 4970 1150
rect 4990 1130 5000 1150
rect 4960 1070 5000 1130
rect 4960 1050 4970 1070
rect 4990 1050 5000 1070
rect 4960 990 5000 1050
rect 4960 970 4970 990
rect 4990 970 5000 990
rect 4960 910 5000 970
rect 4960 890 4970 910
rect 4990 890 5000 910
rect 4960 830 5000 890
rect 4960 810 4970 830
rect 4990 810 5000 830
rect 4960 750 5000 810
rect 4960 730 4970 750
rect 4990 730 5000 750
rect 4960 670 5000 730
rect 4960 650 4970 670
rect 4990 650 5000 670
rect 4960 590 5000 650
rect 4960 570 4970 590
rect 4990 570 5000 590
rect 4960 510 5000 570
rect 4960 490 4970 510
rect 4990 490 5000 510
rect 4960 430 5000 490
rect 4960 410 4970 430
rect 4990 410 5000 430
rect 4960 350 5000 410
rect 4960 330 4970 350
rect 4990 330 5000 350
rect 4960 270 5000 330
rect 4960 250 4970 270
rect 4990 250 5000 270
rect 4960 190 5000 250
rect 4960 170 4970 190
rect 4990 170 5000 190
rect 4960 110 5000 170
rect 4960 90 4970 110
rect 4990 90 5000 110
rect 4960 30 5000 90
rect 4960 10 4970 30
rect 4990 10 5000 30
rect 4960 0 5000 10
rect 5040 15715 5080 15720
rect 5040 15685 5045 15715
rect 5075 15685 5080 15715
rect 5040 15635 5080 15685
rect 5040 15605 5045 15635
rect 5075 15605 5080 15635
rect 5040 15555 5080 15605
rect 5040 15525 5045 15555
rect 5075 15525 5080 15555
rect 5040 15475 5080 15525
rect 5040 15445 5045 15475
rect 5075 15445 5080 15475
rect 5040 15395 5080 15445
rect 5040 15365 5045 15395
rect 5075 15365 5080 15395
rect 5040 15315 5080 15365
rect 5040 15285 5045 15315
rect 5075 15285 5080 15315
rect 5040 15235 5080 15285
rect 5040 15205 5045 15235
rect 5075 15205 5080 15235
rect 5040 15155 5080 15205
rect 5040 15125 5045 15155
rect 5075 15125 5080 15155
rect 5040 15070 5080 15125
rect 5040 15050 5050 15070
rect 5070 15050 5080 15070
rect 5040 14995 5080 15050
rect 5040 14965 5045 14995
rect 5075 14965 5080 14995
rect 5040 14915 5080 14965
rect 5040 14885 5045 14915
rect 5075 14885 5080 14915
rect 5040 14835 5080 14885
rect 5040 14805 5045 14835
rect 5075 14805 5080 14835
rect 5040 14755 5080 14805
rect 5040 14725 5045 14755
rect 5075 14725 5080 14755
rect 5040 14675 5080 14725
rect 5040 14645 5045 14675
rect 5075 14645 5080 14675
rect 5040 14595 5080 14645
rect 5040 14565 5045 14595
rect 5075 14565 5080 14595
rect 5040 14515 5080 14565
rect 5040 14485 5045 14515
rect 5075 14485 5080 14515
rect 5040 14435 5080 14485
rect 5040 14405 5045 14435
rect 5075 14405 5080 14435
rect 5040 14350 5080 14405
rect 5040 14330 5050 14350
rect 5070 14330 5080 14350
rect 5040 14270 5080 14330
rect 5040 14250 5050 14270
rect 5070 14250 5080 14270
rect 5040 14190 5080 14250
rect 5040 14170 5050 14190
rect 5070 14170 5080 14190
rect 5040 14110 5080 14170
rect 5040 14090 5050 14110
rect 5070 14090 5080 14110
rect 5040 14035 5080 14090
rect 5040 14005 5045 14035
rect 5075 14005 5080 14035
rect 5040 13955 5080 14005
rect 5040 13925 5045 13955
rect 5075 13925 5080 13955
rect 5040 13875 5080 13925
rect 5040 13845 5045 13875
rect 5075 13845 5080 13875
rect 5040 13795 5080 13845
rect 5040 13765 5045 13795
rect 5075 13765 5080 13795
rect 5040 13715 5080 13765
rect 5040 13685 5045 13715
rect 5075 13685 5080 13715
rect 5040 13635 5080 13685
rect 5040 13605 5045 13635
rect 5075 13605 5080 13635
rect 5040 13555 5080 13605
rect 5040 13525 5045 13555
rect 5075 13525 5080 13555
rect 5040 13475 5080 13525
rect 5040 13445 5045 13475
rect 5075 13445 5080 13475
rect 5040 13390 5080 13445
rect 5040 13370 5050 13390
rect 5070 13370 5080 13390
rect 5040 13310 5080 13370
rect 5040 13290 5050 13310
rect 5070 13290 5080 13310
rect 5040 13230 5080 13290
rect 5040 13210 5050 13230
rect 5070 13210 5080 13230
rect 5040 13150 5080 13210
rect 5040 13130 5050 13150
rect 5070 13130 5080 13150
rect 5040 13075 5080 13130
rect 5040 13045 5045 13075
rect 5075 13045 5080 13075
rect 5040 12995 5080 13045
rect 5040 12965 5045 12995
rect 5075 12965 5080 12995
rect 5040 12915 5080 12965
rect 5040 12885 5045 12915
rect 5075 12885 5080 12915
rect 5040 12835 5080 12885
rect 5040 12805 5045 12835
rect 5075 12805 5080 12835
rect 5040 12755 5080 12805
rect 5040 12725 5045 12755
rect 5075 12725 5080 12755
rect 5040 12675 5080 12725
rect 5040 12645 5045 12675
rect 5075 12645 5080 12675
rect 5040 12595 5080 12645
rect 5040 12565 5045 12595
rect 5075 12565 5080 12595
rect 5040 12515 5080 12565
rect 5040 12485 5045 12515
rect 5075 12485 5080 12515
rect 5040 12430 5080 12485
rect 5040 12410 5050 12430
rect 5070 12410 5080 12430
rect 5040 12355 5080 12410
rect 5040 12325 5045 12355
rect 5075 12325 5080 12355
rect 5040 12275 5080 12325
rect 5040 12245 5045 12275
rect 5075 12245 5080 12275
rect 5040 12195 5080 12245
rect 5040 12165 5045 12195
rect 5075 12165 5080 12195
rect 5040 12115 5080 12165
rect 5040 12085 5045 12115
rect 5075 12085 5080 12115
rect 5040 12035 5080 12085
rect 5040 12005 5045 12035
rect 5075 12005 5080 12035
rect 5040 11955 5080 12005
rect 5040 11925 5045 11955
rect 5075 11925 5080 11955
rect 5040 11875 5080 11925
rect 5040 11845 5045 11875
rect 5075 11845 5080 11875
rect 5040 11795 5080 11845
rect 5040 11765 5045 11795
rect 5075 11765 5080 11795
rect 5040 11715 5080 11765
rect 5040 11685 5045 11715
rect 5075 11685 5080 11715
rect 5040 11635 5080 11685
rect 5040 11605 5045 11635
rect 5075 11605 5080 11635
rect 5040 11555 5080 11605
rect 5040 11525 5045 11555
rect 5075 11525 5080 11555
rect 5040 11475 5080 11525
rect 5040 11445 5045 11475
rect 5075 11445 5080 11475
rect 5040 11395 5080 11445
rect 5040 11365 5045 11395
rect 5075 11365 5080 11395
rect 5040 11315 5080 11365
rect 5040 11285 5045 11315
rect 5075 11285 5080 11315
rect 5040 11235 5080 11285
rect 5040 11205 5045 11235
rect 5075 11205 5080 11235
rect 5040 11155 5080 11205
rect 5040 11125 5045 11155
rect 5075 11125 5080 11155
rect 5040 11075 5080 11125
rect 5040 11045 5045 11075
rect 5075 11045 5080 11075
rect 5040 10990 5080 11045
rect 5040 10970 5050 10990
rect 5070 10970 5080 10990
rect 5040 10915 5080 10970
rect 5040 10885 5045 10915
rect 5075 10885 5080 10915
rect 5040 10835 5080 10885
rect 5040 10805 5045 10835
rect 5075 10805 5080 10835
rect 5040 10755 5080 10805
rect 5040 10725 5045 10755
rect 5075 10725 5080 10755
rect 5040 10675 5080 10725
rect 5040 10645 5045 10675
rect 5075 10645 5080 10675
rect 5040 10595 5080 10645
rect 5040 10565 5045 10595
rect 5075 10565 5080 10595
rect 5040 10515 5080 10565
rect 5040 10485 5045 10515
rect 5075 10485 5080 10515
rect 5040 10435 5080 10485
rect 5040 10405 5045 10435
rect 5075 10405 5080 10435
rect 5040 10355 5080 10405
rect 5040 10325 5045 10355
rect 5075 10325 5080 10355
rect 5040 10270 5080 10325
rect 5040 10250 5050 10270
rect 5070 10250 5080 10270
rect 5040 10190 5080 10250
rect 5040 10170 5050 10190
rect 5070 10170 5080 10190
rect 5040 10110 5080 10170
rect 5040 10090 5050 10110
rect 5070 10090 5080 10110
rect 5040 10030 5080 10090
rect 5040 10010 5050 10030
rect 5070 10010 5080 10030
rect 5040 9955 5080 10010
rect 5040 9925 5045 9955
rect 5075 9925 5080 9955
rect 5040 9875 5080 9925
rect 5040 9845 5045 9875
rect 5075 9845 5080 9875
rect 5040 9795 5080 9845
rect 5040 9765 5045 9795
rect 5075 9765 5080 9795
rect 5040 9715 5080 9765
rect 5040 9685 5045 9715
rect 5075 9685 5080 9715
rect 5040 9635 5080 9685
rect 5040 9605 5045 9635
rect 5075 9605 5080 9635
rect 5040 9555 5080 9605
rect 5040 9525 5045 9555
rect 5075 9525 5080 9555
rect 5040 9475 5080 9525
rect 5040 9445 5045 9475
rect 5075 9445 5080 9475
rect 5040 9395 5080 9445
rect 5040 9365 5045 9395
rect 5075 9365 5080 9395
rect 5040 9310 5080 9365
rect 5040 9290 5050 9310
rect 5070 9290 5080 9310
rect 5040 9230 5080 9290
rect 5040 9210 5050 9230
rect 5070 9210 5080 9230
rect 5040 9150 5080 9210
rect 5040 9130 5050 9150
rect 5070 9130 5080 9150
rect 5040 9070 5080 9130
rect 5040 9050 5050 9070
rect 5070 9050 5080 9070
rect 5040 8995 5080 9050
rect 5040 8965 5045 8995
rect 5075 8965 5080 8995
rect 5040 8915 5080 8965
rect 5040 8885 5045 8915
rect 5075 8885 5080 8915
rect 5040 8835 5080 8885
rect 5040 8805 5045 8835
rect 5075 8805 5080 8835
rect 5040 8755 5080 8805
rect 5040 8725 5045 8755
rect 5075 8725 5080 8755
rect 5040 8675 5080 8725
rect 5040 8645 5045 8675
rect 5075 8645 5080 8675
rect 5040 8595 5080 8645
rect 5040 8565 5045 8595
rect 5075 8565 5080 8595
rect 5040 8515 5080 8565
rect 5040 8485 5045 8515
rect 5075 8485 5080 8515
rect 5040 8435 5080 8485
rect 5040 8405 5045 8435
rect 5075 8405 5080 8435
rect 5040 8350 5080 8405
rect 5040 8330 5050 8350
rect 5070 8330 5080 8350
rect 5040 8275 5080 8330
rect 5040 8245 5045 8275
rect 5075 8245 5080 8275
rect 5040 8195 5080 8245
rect 5040 8165 5045 8195
rect 5075 8165 5080 8195
rect 5040 8115 5080 8165
rect 5040 8085 5045 8115
rect 5075 8085 5080 8115
rect 5040 8035 5080 8085
rect 5040 8005 5045 8035
rect 5075 8005 5080 8035
rect 5040 7955 5080 8005
rect 5040 7925 5045 7955
rect 5075 7925 5080 7955
rect 5040 7875 5080 7925
rect 5040 7845 5045 7875
rect 5075 7845 5080 7875
rect 5040 7795 5080 7845
rect 5040 7765 5045 7795
rect 5075 7765 5080 7795
rect 5040 7715 5080 7765
rect 5040 7685 5045 7715
rect 5075 7685 5080 7715
rect 5040 7635 5080 7685
rect 5040 7605 5045 7635
rect 5075 7605 5080 7635
rect 5040 7555 5080 7605
rect 5040 7525 5045 7555
rect 5075 7525 5080 7555
rect 5040 7475 5080 7525
rect 5040 7445 5045 7475
rect 5075 7445 5080 7475
rect 5040 7395 5080 7445
rect 5040 7365 5045 7395
rect 5075 7365 5080 7395
rect 5040 7315 5080 7365
rect 5040 7285 5045 7315
rect 5075 7285 5080 7315
rect 5040 7235 5080 7285
rect 5040 7205 5045 7235
rect 5075 7205 5080 7235
rect 5040 7155 5080 7205
rect 5040 7125 5045 7155
rect 5075 7125 5080 7155
rect 5040 7075 5080 7125
rect 5040 7045 5045 7075
rect 5075 7045 5080 7075
rect 5040 6995 5080 7045
rect 5040 6965 5045 6995
rect 5075 6965 5080 6995
rect 5040 6910 5080 6965
rect 5040 6890 5050 6910
rect 5070 6890 5080 6910
rect 5040 6835 5080 6890
rect 5040 6805 5045 6835
rect 5075 6805 5080 6835
rect 5040 6755 5080 6805
rect 5040 6725 5045 6755
rect 5075 6725 5080 6755
rect 5040 6675 5080 6725
rect 5040 6645 5045 6675
rect 5075 6645 5080 6675
rect 5040 6595 5080 6645
rect 5040 6565 5045 6595
rect 5075 6565 5080 6595
rect 5040 6515 5080 6565
rect 5040 6485 5045 6515
rect 5075 6485 5080 6515
rect 5040 6435 5080 6485
rect 5040 6405 5045 6435
rect 5075 6405 5080 6435
rect 5040 6355 5080 6405
rect 5040 6325 5045 6355
rect 5075 6325 5080 6355
rect 5040 6275 5080 6325
rect 5040 6245 5045 6275
rect 5075 6245 5080 6275
rect 5040 6190 5080 6245
rect 5040 6170 5050 6190
rect 5070 6170 5080 6190
rect 5040 6110 5080 6170
rect 5040 6090 5050 6110
rect 5070 6090 5080 6110
rect 5040 6030 5080 6090
rect 5040 6010 5050 6030
rect 5070 6010 5080 6030
rect 5040 5950 5080 6010
rect 5040 5930 5050 5950
rect 5070 5930 5080 5950
rect 5040 5875 5080 5930
rect 5040 5845 5045 5875
rect 5075 5845 5080 5875
rect 5040 5795 5080 5845
rect 5040 5765 5045 5795
rect 5075 5765 5080 5795
rect 5040 5715 5080 5765
rect 5040 5685 5045 5715
rect 5075 5685 5080 5715
rect 5040 5635 5080 5685
rect 5040 5605 5045 5635
rect 5075 5605 5080 5635
rect 5040 5555 5080 5605
rect 5040 5525 5045 5555
rect 5075 5525 5080 5555
rect 5040 5475 5080 5525
rect 5040 5445 5045 5475
rect 5075 5445 5080 5475
rect 5040 5395 5080 5445
rect 5040 5365 5045 5395
rect 5075 5365 5080 5395
rect 5040 5315 5080 5365
rect 5040 5285 5045 5315
rect 5075 5285 5080 5315
rect 5040 5235 5080 5285
rect 5040 5205 5045 5235
rect 5075 5205 5080 5235
rect 5040 5155 5080 5205
rect 5040 5125 5045 5155
rect 5075 5125 5080 5155
rect 5040 5075 5080 5125
rect 5040 5045 5045 5075
rect 5075 5045 5080 5075
rect 5040 4995 5080 5045
rect 5040 4965 5045 4995
rect 5075 4965 5080 4995
rect 5040 4915 5080 4965
rect 5040 4885 5045 4915
rect 5075 4885 5080 4915
rect 5040 4830 5080 4885
rect 5040 4810 5050 4830
rect 5070 4810 5080 4830
rect 5040 4755 5080 4810
rect 5040 4725 5045 4755
rect 5075 4725 5080 4755
rect 5040 4675 5080 4725
rect 5040 4645 5045 4675
rect 5075 4645 5080 4675
rect 5040 4590 5080 4645
rect 5040 4570 5050 4590
rect 5070 4570 5080 4590
rect 5040 4515 5080 4570
rect 5040 4485 5045 4515
rect 5075 4485 5080 4515
rect 5040 4435 5080 4485
rect 5040 4405 5045 4435
rect 5075 4405 5080 4435
rect 5040 4355 5080 4405
rect 5040 4325 5045 4355
rect 5075 4325 5080 4355
rect 5040 4275 5080 4325
rect 5040 4245 5045 4275
rect 5075 4245 5080 4275
rect 5040 4195 5080 4245
rect 5040 4165 5045 4195
rect 5075 4165 5080 4195
rect 5040 4115 5080 4165
rect 5040 4085 5045 4115
rect 5075 4085 5080 4115
rect 5040 4035 5080 4085
rect 5040 4005 5045 4035
rect 5075 4005 5080 4035
rect 5040 3955 5080 4005
rect 5040 3925 5045 3955
rect 5075 3925 5080 3955
rect 5040 3875 5080 3925
rect 5040 3845 5045 3875
rect 5075 3845 5080 3875
rect 5040 3790 5080 3845
rect 5040 3770 5050 3790
rect 5070 3770 5080 3790
rect 5040 3715 5080 3770
rect 5040 3685 5045 3715
rect 5075 3685 5080 3715
rect 5040 3635 5080 3685
rect 5040 3605 5045 3635
rect 5075 3605 5080 3635
rect 5040 3550 5080 3605
rect 5040 3530 5050 3550
rect 5070 3530 5080 3550
rect 5040 3475 5080 3530
rect 5040 3445 5045 3475
rect 5075 3445 5080 3475
rect 5040 3395 5080 3445
rect 5040 3365 5045 3395
rect 5075 3365 5080 3395
rect 5040 3310 5080 3365
rect 5040 3290 5050 3310
rect 5070 3290 5080 3310
rect 5040 3235 5080 3290
rect 5040 3205 5045 3235
rect 5075 3205 5080 3235
rect 5040 3155 5080 3205
rect 5040 3125 5045 3155
rect 5075 3125 5080 3155
rect 5040 3075 5080 3125
rect 5040 3045 5045 3075
rect 5075 3045 5080 3075
rect 5040 2995 5080 3045
rect 5040 2965 5045 2995
rect 5075 2965 5080 2995
rect 5040 2915 5080 2965
rect 5040 2885 5045 2915
rect 5075 2885 5080 2915
rect 5040 2835 5080 2885
rect 5040 2805 5045 2835
rect 5075 2805 5080 2835
rect 5040 2755 5080 2805
rect 5040 2725 5045 2755
rect 5075 2725 5080 2755
rect 5040 2675 5080 2725
rect 5040 2645 5045 2675
rect 5075 2645 5080 2675
rect 5040 2595 5080 2645
rect 5040 2565 5045 2595
rect 5075 2565 5080 2595
rect 5040 2515 5080 2565
rect 5040 2485 5045 2515
rect 5075 2485 5080 2515
rect 5040 2435 5080 2485
rect 5040 2405 5045 2435
rect 5075 2405 5080 2435
rect 5040 2355 5080 2405
rect 5040 2325 5045 2355
rect 5075 2325 5080 2355
rect 5040 2275 5080 2325
rect 5040 2245 5045 2275
rect 5075 2245 5080 2275
rect 5040 2195 5080 2245
rect 5040 2165 5045 2195
rect 5075 2165 5080 2195
rect 5040 2115 5080 2165
rect 5040 2085 5045 2115
rect 5075 2085 5080 2115
rect 5040 2035 5080 2085
rect 5040 2005 5045 2035
rect 5075 2005 5080 2035
rect 5040 1955 5080 2005
rect 5040 1925 5045 1955
rect 5075 1925 5080 1955
rect 5040 1870 5080 1925
rect 5040 1850 5050 1870
rect 5070 1850 5080 1870
rect 5040 1790 5080 1850
rect 5040 1770 5050 1790
rect 5070 1770 5080 1790
rect 5040 1715 5080 1770
rect 5040 1685 5045 1715
rect 5075 1685 5080 1715
rect 5040 1635 5080 1685
rect 5040 1605 5045 1635
rect 5075 1605 5080 1635
rect 5040 1555 5080 1605
rect 5040 1525 5045 1555
rect 5075 1525 5080 1555
rect 5040 1475 5080 1525
rect 5040 1445 5045 1475
rect 5075 1445 5080 1475
rect 5040 1395 5080 1445
rect 5040 1365 5045 1395
rect 5075 1365 5080 1395
rect 5040 1315 5080 1365
rect 5040 1285 5045 1315
rect 5075 1285 5080 1315
rect 5040 1235 5080 1285
rect 5040 1205 5045 1235
rect 5075 1205 5080 1235
rect 5040 1155 5080 1205
rect 5040 1125 5045 1155
rect 5075 1125 5080 1155
rect 5040 1075 5080 1125
rect 5040 1045 5045 1075
rect 5075 1045 5080 1075
rect 5040 995 5080 1045
rect 5040 965 5045 995
rect 5075 965 5080 995
rect 5040 910 5080 965
rect 5040 890 5050 910
rect 5070 890 5080 910
rect 5040 835 5080 890
rect 5040 805 5045 835
rect 5075 805 5080 835
rect 5040 755 5080 805
rect 5040 725 5045 755
rect 5075 725 5080 755
rect 5040 675 5080 725
rect 5040 645 5045 675
rect 5075 645 5080 675
rect 5040 595 5080 645
rect 5040 565 5045 595
rect 5075 565 5080 595
rect 5040 515 5080 565
rect 5040 485 5045 515
rect 5075 485 5080 515
rect 5040 430 5080 485
rect 5040 410 5050 430
rect 5070 410 5080 430
rect 5040 350 5080 410
rect 5040 330 5050 350
rect 5070 330 5080 350
rect 5040 275 5080 330
rect 5040 245 5045 275
rect 5075 245 5080 275
rect 5040 195 5080 245
rect 5040 165 5045 195
rect 5075 165 5080 195
rect 5040 115 5080 165
rect 5040 85 5045 115
rect 5075 85 5080 115
rect 5040 35 5080 85
rect 5040 5 5045 35
rect 5075 5 5080 35
rect 5040 0 5080 5
rect 5120 15710 5160 15720
rect 5120 15690 5130 15710
rect 5150 15690 5160 15710
rect 5120 15630 5160 15690
rect 5120 15610 5130 15630
rect 5150 15610 5160 15630
rect 5120 15550 5160 15610
rect 5120 15530 5130 15550
rect 5150 15530 5160 15550
rect 5120 15470 5160 15530
rect 5120 15450 5130 15470
rect 5150 15450 5160 15470
rect 5120 15390 5160 15450
rect 5120 15370 5130 15390
rect 5150 15370 5160 15390
rect 5120 15310 5160 15370
rect 5120 15290 5130 15310
rect 5150 15290 5160 15310
rect 5120 15230 5160 15290
rect 5120 15210 5130 15230
rect 5150 15210 5160 15230
rect 5120 15150 5160 15210
rect 5120 15130 5130 15150
rect 5150 15130 5160 15150
rect 5120 15070 5160 15130
rect 5120 15050 5130 15070
rect 5150 15050 5160 15070
rect 5120 14990 5160 15050
rect 5120 14970 5130 14990
rect 5150 14970 5160 14990
rect 5120 14910 5160 14970
rect 5120 14890 5130 14910
rect 5150 14890 5160 14910
rect 5120 14830 5160 14890
rect 5120 14810 5130 14830
rect 5150 14810 5160 14830
rect 5120 14750 5160 14810
rect 5120 14730 5130 14750
rect 5150 14730 5160 14750
rect 5120 14670 5160 14730
rect 5120 14650 5130 14670
rect 5150 14650 5160 14670
rect 5120 14590 5160 14650
rect 5120 14570 5130 14590
rect 5150 14570 5160 14590
rect 5120 14510 5160 14570
rect 5120 14490 5130 14510
rect 5150 14490 5160 14510
rect 5120 14430 5160 14490
rect 5120 14410 5130 14430
rect 5150 14410 5160 14430
rect 5120 14350 5160 14410
rect 5120 14330 5130 14350
rect 5150 14330 5160 14350
rect 5120 14270 5160 14330
rect 5120 14250 5130 14270
rect 5150 14250 5160 14270
rect 5120 14190 5160 14250
rect 5120 14170 5130 14190
rect 5150 14170 5160 14190
rect 5120 14110 5160 14170
rect 5120 14090 5130 14110
rect 5150 14090 5160 14110
rect 5120 14030 5160 14090
rect 5120 14010 5130 14030
rect 5150 14010 5160 14030
rect 5120 13950 5160 14010
rect 5120 13930 5130 13950
rect 5150 13930 5160 13950
rect 5120 13870 5160 13930
rect 5120 13850 5130 13870
rect 5150 13850 5160 13870
rect 5120 13790 5160 13850
rect 5120 13770 5130 13790
rect 5150 13770 5160 13790
rect 5120 13710 5160 13770
rect 5120 13690 5130 13710
rect 5150 13690 5160 13710
rect 5120 13630 5160 13690
rect 5120 13610 5130 13630
rect 5150 13610 5160 13630
rect 5120 13550 5160 13610
rect 5120 13530 5130 13550
rect 5150 13530 5160 13550
rect 5120 13470 5160 13530
rect 5120 13450 5130 13470
rect 5150 13450 5160 13470
rect 5120 13390 5160 13450
rect 5120 13370 5130 13390
rect 5150 13370 5160 13390
rect 5120 13310 5160 13370
rect 5120 13290 5130 13310
rect 5150 13290 5160 13310
rect 5120 13230 5160 13290
rect 5120 13210 5130 13230
rect 5150 13210 5160 13230
rect 5120 13150 5160 13210
rect 5120 13130 5130 13150
rect 5150 13130 5160 13150
rect 5120 13070 5160 13130
rect 5120 13050 5130 13070
rect 5150 13050 5160 13070
rect 5120 12990 5160 13050
rect 5120 12970 5130 12990
rect 5150 12970 5160 12990
rect 5120 12910 5160 12970
rect 5120 12890 5130 12910
rect 5150 12890 5160 12910
rect 5120 12830 5160 12890
rect 5120 12810 5130 12830
rect 5150 12810 5160 12830
rect 5120 12750 5160 12810
rect 5120 12730 5130 12750
rect 5150 12730 5160 12750
rect 5120 12670 5160 12730
rect 5120 12650 5130 12670
rect 5150 12650 5160 12670
rect 5120 12590 5160 12650
rect 5120 12570 5130 12590
rect 5150 12570 5160 12590
rect 5120 12510 5160 12570
rect 5120 12490 5130 12510
rect 5150 12490 5160 12510
rect 5120 12430 5160 12490
rect 5120 12410 5130 12430
rect 5150 12410 5160 12430
rect 5120 12350 5160 12410
rect 5120 12330 5130 12350
rect 5150 12330 5160 12350
rect 5120 12270 5160 12330
rect 5120 12250 5130 12270
rect 5150 12250 5160 12270
rect 5120 12190 5160 12250
rect 5120 12170 5130 12190
rect 5150 12170 5160 12190
rect 5120 12110 5160 12170
rect 5120 12090 5130 12110
rect 5150 12090 5160 12110
rect 5120 12030 5160 12090
rect 5120 12010 5130 12030
rect 5150 12010 5160 12030
rect 5120 11950 5160 12010
rect 5120 11930 5130 11950
rect 5150 11930 5160 11950
rect 5120 11870 5160 11930
rect 5120 11850 5130 11870
rect 5150 11850 5160 11870
rect 5120 11790 5160 11850
rect 5120 11770 5130 11790
rect 5150 11770 5160 11790
rect 5120 11710 5160 11770
rect 5120 11690 5130 11710
rect 5150 11690 5160 11710
rect 5120 11630 5160 11690
rect 5120 11610 5130 11630
rect 5150 11610 5160 11630
rect 5120 11550 5160 11610
rect 5120 11530 5130 11550
rect 5150 11530 5160 11550
rect 5120 11470 5160 11530
rect 5120 11450 5130 11470
rect 5150 11450 5160 11470
rect 5120 11390 5160 11450
rect 5120 11370 5130 11390
rect 5150 11370 5160 11390
rect 5120 11310 5160 11370
rect 5120 11290 5130 11310
rect 5150 11290 5160 11310
rect 5120 11230 5160 11290
rect 5120 11210 5130 11230
rect 5150 11210 5160 11230
rect 5120 11150 5160 11210
rect 5120 11130 5130 11150
rect 5150 11130 5160 11150
rect 5120 11070 5160 11130
rect 5120 11050 5130 11070
rect 5150 11050 5160 11070
rect 5120 10990 5160 11050
rect 5120 10970 5130 10990
rect 5150 10970 5160 10990
rect 5120 10910 5160 10970
rect 5120 10890 5130 10910
rect 5150 10890 5160 10910
rect 5120 10830 5160 10890
rect 5120 10810 5130 10830
rect 5150 10810 5160 10830
rect 5120 10750 5160 10810
rect 5120 10730 5130 10750
rect 5150 10730 5160 10750
rect 5120 10670 5160 10730
rect 5120 10650 5130 10670
rect 5150 10650 5160 10670
rect 5120 10590 5160 10650
rect 5120 10570 5130 10590
rect 5150 10570 5160 10590
rect 5120 10510 5160 10570
rect 5120 10490 5130 10510
rect 5150 10490 5160 10510
rect 5120 10430 5160 10490
rect 5120 10410 5130 10430
rect 5150 10410 5160 10430
rect 5120 10350 5160 10410
rect 5120 10330 5130 10350
rect 5150 10330 5160 10350
rect 5120 10270 5160 10330
rect 5120 10250 5130 10270
rect 5150 10250 5160 10270
rect 5120 10190 5160 10250
rect 5120 10170 5130 10190
rect 5150 10170 5160 10190
rect 5120 10110 5160 10170
rect 5120 10090 5130 10110
rect 5150 10090 5160 10110
rect 5120 10030 5160 10090
rect 5120 10010 5130 10030
rect 5150 10010 5160 10030
rect 5120 9950 5160 10010
rect 5120 9930 5130 9950
rect 5150 9930 5160 9950
rect 5120 9870 5160 9930
rect 5120 9850 5130 9870
rect 5150 9850 5160 9870
rect 5120 9790 5160 9850
rect 5120 9770 5130 9790
rect 5150 9770 5160 9790
rect 5120 9710 5160 9770
rect 5120 9690 5130 9710
rect 5150 9690 5160 9710
rect 5120 9630 5160 9690
rect 5120 9610 5130 9630
rect 5150 9610 5160 9630
rect 5120 9550 5160 9610
rect 5120 9530 5130 9550
rect 5150 9530 5160 9550
rect 5120 9470 5160 9530
rect 5120 9450 5130 9470
rect 5150 9450 5160 9470
rect 5120 9390 5160 9450
rect 5120 9370 5130 9390
rect 5150 9370 5160 9390
rect 5120 9310 5160 9370
rect 5120 9290 5130 9310
rect 5150 9290 5160 9310
rect 5120 9230 5160 9290
rect 5120 9210 5130 9230
rect 5150 9210 5160 9230
rect 5120 9150 5160 9210
rect 5120 9130 5130 9150
rect 5150 9130 5160 9150
rect 5120 9070 5160 9130
rect 5120 9050 5130 9070
rect 5150 9050 5160 9070
rect 5120 8990 5160 9050
rect 5120 8970 5130 8990
rect 5150 8970 5160 8990
rect 5120 8910 5160 8970
rect 5120 8890 5130 8910
rect 5150 8890 5160 8910
rect 5120 8830 5160 8890
rect 5120 8810 5130 8830
rect 5150 8810 5160 8830
rect 5120 8750 5160 8810
rect 5120 8730 5130 8750
rect 5150 8730 5160 8750
rect 5120 8670 5160 8730
rect 5120 8650 5130 8670
rect 5150 8650 5160 8670
rect 5120 8590 5160 8650
rect 5120 8570 5130 8590
rect 5150 8570 5160 8590
rect 5120 8510 5160 8570
rect 5120 8490 5130 8510
rect 5150 8490 5160 8510
rect 5120 8430 5160 8490
rect 5120 8410 5130 8430
rect 5150 8410 5160 8430
rect 5120 8350 5160 8410
rect 5120 8330 5130 8350
rect 5150 8330 5160 8350
rect 5120 8270 5160 8330
rect 5120 8250 5130 8270
rect 5150 8250 5160 8270
rect 5120 8190 5160 8250
rect 5120 8170 5130 8190
rect 5150 8170 5160 8190
rect 5120 8110 5160 8170
rect 5120 8090 5130 8110
rect 5150 8090 5160 8110
rect 5120 8030 5160 8090
rect 5120 8010 5130 8030
rect 5150 8010 5160 8030
rect 5120 7950 5160 8010
rect 5120 7930 5130 7950
rect 5150 7930 5160 7950
rect 5120 7870 5160 7930
rect 5120 7850 5130 7870
rect 5150 7850 5160 7870
rect 5120 7790 5160 7850
rect 5120 7770 5130 7790
rect 5150 7770 5160 7790
rect 5120 7710 5160 7770
rect 5120 7690 5130 7710
rect 5150 7690 5160 7710
rect 5120 7630 5160 7690
rect 5120 7610 5130 7630
rect 5150 7610 5160 7630
rect 5120 7550 5160 7610
rect 5120 7530 5130 7550
rect 5150 7530 5160 7550
rect 5120 7470 5160 7530
rect 5120 7450 5130 7470
rect 5150 7450 5160 7470
rect 5120 7390 5160 7450
rect 5120 7370 5130 7390
rect 5150 7370 5160 7390
rect 5120 7310 5160 7370
rect 5120 7290 5130 7310
rect 5150 7290 5160 7310
rect 5120 7230 5160 7290
rect 5120 7210 5130 7230
rect 5150 7210 5160 7230
rect 5120 7150 5160 7210
rect 5120 7130 5130 7150
rect 5150 7130 5160 7150
rect 5120 7070 5160 7130
rect 5120 7050 5130 7070
rect 5150 7050 5160 7070
rect 5120 6990 5160 7050
rect 5120 6970 5130 6990
rect 5150 6970 5160 6990
rect 5120 6910 5160 6970
rect 5120 6890 5130 6910
rect 5150 6890 5160 6910
rect 5120 6830 5160 6890
rect 5120 6810 5130 6830
rect 5150 6810 5160 6830
rect 5120 6750 5160 6810
rect 5120 6730 5130 6750
rect 5150 6730 5160 6750
rect 5120 6670 5160 6730
rect 5120 6650 5130 6670
rect 5150 6650 5160 6670
rect 5120 6590 5160 6650
rect 5120 6570 5130 6590
rect 5150 6570 5160 6590
rect 5120 6510 5160 6570
rect 5120 6490 5130 6510
rect 5150 6490 5160 6510
rect 5120 6430 5160 6490
rect 5120 6410 5130 6430
rect 5150 6410 5160 6430
rect 5120 6350 5160 6410
rect 5120 6330 5130 6350
rect 5150 6330 5160 6350
rect 5120 6270 5160 6330
rect 5120 6250 5130 6270
rect 5150 6250 5160 6270
rect 5120 6190 5160 6250
rect 5120 6170 5130 6190
rect 5150 6170 5160 6190
rect 5120 6110 5160 6170
rect 5120 6090 5130 6110
rect 5150 6090 5160 6110
rect 5120 6030 5160 6090
rect 5120 6010 5130 6030
rect 5150 6010 5160 6030
rect 5120 5950 5160 6010
rect 5120 5930 5130 5950
rect 5150 5930 5160 5950
rect 5120 5870 5160 5930
rect 5120 5850 5130 5870
rect 5150 5850 5160 5870
rect 5120 5790 5160 5850
rect 5120 5770 5130 5790
rect 5150 5770 5160 5790
rect 5120 5710 5160 5770
rect 5120 5690 5130 5710
rect 5150 5690 5160 5710
rect 5120 5630 5160 5690
rect 5120 5610 5130 5630
rect 5150 5610 5160 5630
rect 5120 5550 5160 5610
rect 5120 5530 5130 5550
rect 5150 5530 5160 5550
rect 5120 5470 5160 5530
rect 5120 5450 5130 5470
rect 5150 5450 5160 5470
rect 5120 5390 5160 5450
rect 5120 5370 5130 5390
rect 5150 5370 5160 5390
rect 5120 5310 5160 5370
rect 5120 5290 5130 5310
rect 5150 5290 5160 5310
rect 5120 5230 5160 5290
rect 5120 5210 5130 5230
rect 5150 5210 5160 5230
rect 5120 5150 5160 5210
rect 5120 5130 5130 5150
rect 5150 5130 5160 5150
rect 5120 5070 5160 5130
rect 5120 5050 5130 5070
rect 5150 5050 5160 5070
rect 5120 4990 5160 5050
rect 5120 4970 5130 4990
rect 5150 4970 5160 4990
rect 5120 4910 5160 4970
rect 5120 4890 5130 4910
rect 5150 4890 5160 4910
rect 5120 4830 5160 4890
rect 5120 4810 5130 4830
rect 5150 4810 5160 4830
rect 5120 4750 5160 4810
rect 5120 4730 5130 4750
rect 5150 4730 5160 4750
rect 5120 4670 5160 4730
rect 5120 4650 5130 4670
rect 5150 4650 5160 4670
rect 5120 4590 5160 4650
rect 5120 4570 5130 4590
rect 5150 4570 5160 4590
rect 5120 4510 5160 4570
rect 5120 4490 5130 4510
rect 5150 4490 5160 4510
rect 5120 4430 5160 4490
rect 5120 4410 5130 4430
rect 5150 4410 5160 4430
rect 5120 4350 5160 4410
rect 5120 4330 5130 4350
rect 5150 4330 5160 4350
rect 5120 4270 5160 4330
rect 5120 4250 5130 4270
rect 5150 4250 5160 4270
rect 5120 4190 5160 4250
rect 5120 4170 5130 4190
rect 5150 4170 5160 4190
rect 5120 4110 5160 4170
rect 5120 4090 5130 4110
rect 5150 4090 5160 4110
rect 5120 4030 5160 4090
rect 5120 4010 5130 4030
rect 5150 4010 5160 4030
rect 5120 3950 5160 4010
rect 5120 3930 5130 3950
rect 5150 3930 5160 3950
rect 5120 3870 5160 3930
rect 5120 3850 5130 3870
rect 5150 3850 5160 3870
rect 5120 3790 5160 3850
rect 5120 3770 5130 3790
rect 5150 3770 5160 3790
rect 5120 3710 5160 3770
rect 5120 3690 5130 3710
rect 5150 3690 5160 3710
rect 5120 3630 5160 3690
rect 5120 3610 5130 3630
rect 5150 3610 5160 3630
rect 5120 3550 5160 3610
rect 5120 3530 5130 3550
rect 5150 3530 5160 3550
rect 5120 3470 5160 3530
rect 5120 3450 5130 3470
rect 5150 3450 5160 3470
rect 5120 3390 5160 3450
rect 5120 3370 5130 3390
rect 5150 3370 5160 3390
rect 5120 3310 5160 3370
rect 5120 3290 5130 3310
rect 5150 3290 5160 3310
rect 5120 3230 5160 3290
rect 5120 3210 5130 3230
rect 5150 3210 5160 3230
rect 5120 3150 5160 3210
rect 5120 3130 5130 3150
rect 5150 3130 5160 3150
rect 5120 3070 5160 3130
rect 5120 3050 5130 3070
rect 5150 3050 5160 3070
rect 5120 2990 5160 3050
rect 5120 2970 5130 2990
rect 5150 2970 5160 2990
rect 5120 2910 5160 2970
rect 5120 2890 5130 2910
rect 5150 2890 5160 2910
rect 5120 2830 5160 2890
rect 5120 2810 5130 2830
rect 5150 2810 5160 2830
rect 5120 2750 5160 2810
rect 5120 2730 5130 2750
rect 5150 2730 5160 2750
rect 5120 2670 5160 2730
rect 5120 2650 5130 2670
rect 5150 2650 5160 2670
rect 5120 2590 5160 2650
rect 5120 2570 5130 2590
rect 5150 2570 5160 2590
rect 5120 2510 5160 2570
rect 5120 2490 5130 2510
rect 5150 2490 5160 2510
rect 5120 2430 5160 2490
rect 5120 2410 5130 2430
rect 5150 2410 5160 2430
rect 5120 2350 5160 2410
rect 5120 2330 5130 2350
rect 5150 2330 5160 2350
rect 5120 2270 5160 2330
rect 5120 2250 5130 2270
rect 5150 2250 5160 2270
rect 5120 2190 5160 2250
rect 5120 2170 5130 2190
rect 5150 2170 5160 2190
rect 5120 2110 5160 2170
rect 5120 2090 5130 2110
rect 5150 2090 5160 2110
rect 5120 2030 5160 2090
rect 5120 2010 5130 2030
rect 5150 2010 5160 2030
rect 5120 1950 5160 2010
rect 5120 1930 5130 1950
rect 5150 1930 5160 1950
rect 5120 1870 5160 1930
rect 5120 1850 5130 1870
rect 5150 1850 5160 1870
rect 5120 1790 5160 1850
rect 5120 1770 5130 1790
rect 5150 1770 5160 1790
rect 5120 1710 5160 1770
rect 5120 1690 5130 1710
rect 5150 1690 5160 1710
rect 5120 1630 5160 1690
rect 5120 1610 5130 1630
rect 5150 1610 5160 1630
rect 5120 1550 5160 1610
rect 5120 1530 5130 1550
rect 5150 1530 5160 1550
rect 5120 1470 5160 1530
rect 5120 1450 5130 1470
rect 5150 1450 5160 1470
rect 5120 1390 5160 1450
rect 5120 1370 5130 1390
rect 5150 1370 5160 1390
rect 5120 1310 5160 1370
rect 5120 1290 5130 1310
rect 5150 1290 5160 1310
rect 5120 1230 5160 1290
rect 5120 1210 5130 1230
rect 5150 1210 5160 1230
rect 5120 1150 5160 1210
rect 5120 1130 5130 1150
rect 5150 1130 5160 1150
rect 5120 1070 5160 1130
rect 5120 1050 5130 1070
rect 5150 1050 5160 1070
rect 5120 990 5160 1050
rect 5120 970 5130 990
rect 5150 970 5160 990
rect 5120 910 5160 970
rect 5120 890 5130 910
rect 5150 890 5160 910
rect 5120 830 5160 890
rect 5120 810 5130 830
rect 5150 810 5160 830
rect 5120 750 5160 810
rect 5120 730 5130 750
rect 5150 730 5160 750
rect 5120 670 5160 730
rect 5120 650 5130 670
rect 5150 650 5160 670
rect 5120 590 5160 650
rect 5120 570 5130 590
rect 5150 570 5160 590
rect 5120 510 5160 570
rect 5120 490 5130 510
rect 5150 490 5160 510
rect 5120 430 5160 490
rect 5120 410 5130 430
rect 5150 410 5160 430
rect 5120 350 5160 410
rect 5120 330 5130 350
rect 5150 330 5160 350
rect 5120 270 5160 330
rect 5120 250 5130 270
rect 5150 250 5160 270
rect 5120 190 5160 250
rect 5120 170 5130 190
rect 5150 170 5160 190
rect 5120 110 5160 170
rect 5120 90 5130 110
rect 5150 90 5160 110
rect 5120 30 5160 90
rect 5120 10 5130 30
rect 5150 10 5160 30
rect 5120 0 5160 10
rect 5200 15715 5240 15720
rect 5200 15685 5205 15715
rect 5235 15685 5240 15715
rect 5200 15635 5240 15685
rect 5200 15605 5205 15635
rect 5235 15605 5240 15635
rect 5200 15555 5240 15605
rect 5200 15525 5205 15555
rect 5235 15525 5240 15555
rect 5200 15475 5240 15525
rect 5200 15445 5205 15475
rect 5235 15445 5240 15475
rect 5200 15395 5240 15445
rect 5200 15365 5205 15395
rect 5235 15365 5240 15395
rect 5200 15315 5240 15365
rect 5200 15285 5205 15315
rect 5235 15285 5240 15315
rect 5200 15235 5240 15285
rect 5200 15205 5205 15235
rect 5235 15205 5240 15235
rect 5200 15155 5240 15205
rect 5200 15125 5205 15155
rect 5235 15125 5240 15155
rect 5200 15070 5240 15125
rect 5200 15050 5210 15070
rect 5230 15050 5240 15070
rect 5200 14995 5240 15050
rect 5200 14965 5205 14995
rect 5235 14965 5240 14995
rect 5200 14915 5240 14965
rect 5200 14885 5205 14915
rect 5235 14885 5240 14915
rect 5200 14835 5240 14885
rect 5200 14805 5205 14835
rect 5235 14805 5240 14835
rect 5200 14755 5240 14805
rect 5200 14725 5205 14755
rect 5235 14725 5240 14755
rect 5200 14675 5240 14725
rect 5200 14645 5205 14675
rect 5235 14645 5240 14675
rect 5200 14595 5240 14645
rect 5200 14565 5205 14595
rect 5235 14565 5240 14595
rect 5200 14515 5240 14565
rect 5200 14485 5205 14515
rect 5235 14485 5240 14515
rect 5200 14435 5240 14485
rect 5200 14405 5205 14435
rect 5235 14405 5240 14435
rect 5200 14350 5240 14405
rect 5200 14330 5210 14350
rect 5230 14330 5240 14350
rect 5200 14270 5240 14330
rect 5200 14250 5210 14270
rect 5230 14250 5240 14270
rect 5200 14190 5240 14250
rect 5200 14170 5210 14190
rect 5230 14170 5240 14190
rect 5200 14110 5240 14170
rect 5200 14090 5210 14110
rect 5230 14090 5240 14110
rect 5200 14035 5240 14090
rect 5200 14005 5205 14035
rect 5235 14005 5240 14035
rect 5200 13955 5240 14005
rect 5200 13925 5205 13955
rect 5235 13925 5240 13955
rect 5200 13875 5240 13925
rect 5200 13845 5205 13875
rect 5235 13845 5240 13875
rect 5200 13795 5240 13845
rect 5200 13765 5205 13795
rect 5235 13765 5240 13795
rect 5200 13715 5240 13765
rect 5200 13685 5205 13715
rect 5235 13685 5240 13715
rect 5200 13635 5240 13685
rect 5200 13605 5205 13635
rect 5235 13605 5240 13635
rect 5200 13555 5240 13605
rect 5200 13525 5205 13555
rect 5235 13525 5240 13555
rect 5200 13475 5240 13525
rect 5200 13445 5205 13475
rect 5235 13445 5240 13475
rect 5200 13390 5240 13445
rect 5200 13370 5210 13390
rect 5230 13370 5240 13390
rect 5200 13310 5240 13370
rect 5200 13290 5210 13310
rect 5230 13290 5240 13310
rect 5200 13230 5240 13290
rect 5200 13210 5210 13230
rect 5230 13210 5240 13230
rect 5200 13150 5240 13210
rect 5200 13130 5210 13150
rect 5230 13130 5240 13150
rect 5200 13075 5240 13130
rect 5200 13045 5205 13075
rect 5235 13045 5240 13075
rect 5200 12995 5240 13045
rect 5200 12965 5205 12995
rect 5235 12965 5240 12995
rect 5200 12915 5240 12965
rect 5200 12885 5205 12915
rect 5235 12885 5240 12915
rect 5200 12835 5240 12885
rect 5200 12805 5205 12835
rect 5235 12805 5240 12835
rect 5200 12755 5240 12805
rect 5200 12725 5205 12755
rect 5235 12725 5240 12755
rect 5200 12675 5240 12725
rect 5200 12645 5205 12675
rect 5235 12645 5240 12675
rect 5200 12595 5240 12645
rect 5200 12565 5205 12595
rect 5235 12565 5240 12595
rect 5200 12515 5240 12565
rect 5200 12485 5205 12515
rect 5235 12485 5240 12515
rect 5200 12430 5240 12485
rect 5200 12410 5210 12430
rect 5230 12410 5240 12430
rect 5200 12355 5240 12410
rect 5200 12325 5205 12355
rect 5235 12325 5240 12355
rect 5200 12275 5240 12325
rect 5200 12245 5205 12275
rect 5235 12245 5240 12275
rect 5200 12195 5240 12245
rect 5200 12165 5205 12195
rect 5235 12165 5240 12195
rect 5200 12115 5240 12165
rect 5200 12085 5205 12115
rect 5235 12085 5240 12115
rect 5200 12035 5240 12085
rect 5200 12005 5205 12035
rect 5235 12005 5240 12035
rect 5200 11955 5240 12005
rect 5200 11925 5205 11955
rect 5235 11925 5240 11955
rect 5200 11875 5240 11925
rect 5200 11845 5205 11875
rect 5235 11845 5240 11875
rect 5200 11795 5240 11845
rect 5200 11765 5205 11795
rect 5235 11765 5240 11795
rect 5200 11715 5240 11765
rect 5200 11685 5205 11715
rect 5235 11685 5240 11715
rect 5200 11635 5240 11685
rect 5200 11605 5205 11635
rect 5235 11605 5240 11635
rect 5200 11555 5240 11605
rect 5200 11525 5205 11555
rect 5235 11525 5240 11555
rect 5200 11475 5240 11525
rect 5200 11445 5205 11475
rect 5235 11445 5240 11475
rect 5200 11395 5240 11445
rect 5200 11365 5205 11395
rect 5235 11365 5240 11395
rect 5200 11315 5240 11365
rect 5200 11285 5205 11315
rect 5235 11285 5240 11315
rect 5200 11235 5240 11285
rect 5200 11205 5205 11235
rect 5235 11205 5240 11235
rect 5200 11155 5240 11205
rect 5200 11125 5205 11155
rect 5235 11125 5240 11155
rect 5200 11075 5240 11125
rect 5200 11045 5205 11075
rect 5235 11045 5240 11075
rect 5200 10990 5240 11045
rect 5200 10970 5210 10990
rect 5230 10970 5240 10990
rect 5200 10915 5240 10970
rect 5200 10885 5205 10915
rect 5235 10885 5240 10915
rect 5200 10835 5240 10885
rect 5200 10805 5205 10835
rect 5235 10805 5240 10835
rect 5200 10755 5240 10805
rect 5200 10725 5205 10755
rect 5235 10725 5240 10755
rect 5200 10675 5240 10725
rect 5200 10645 5205 10675
rect 5235 10645 5240 10675
rect 5200 10595 5240 10645
rect 5200 10565 5205 10595
rect 5235 10565 5240 10595
rect 5200 10515 5240 10565
rect 5200 10485 5205 10515
rect 5235 10485 5240 10515
rect 5200 10435 5240 10485
rect 5200 10405 5205 10435
rect 5235 10405 5240 10435
rect 5200 10355 5240 10405
rect 5200 10325 5205 10355
rect 5235 10325 5240 10355
rect 5200 10270 5240 10325
rect 5200 10250 5210 10270
rect 5230 10250 5240 10270
rect 5200 10190 5240 10250
rect 5200 10170 5210 10190
rect 5230 10170 5240 10190
rect 5200 10110 5240 10170
rect 5200 10090 5210 10110
rect 5230 10090 5240 10110
rect 5200 10030 5240 10090
rect 5200 10010 5210 10030
rect 5230 10010 5240 10030
rect 5200 9955 5240 10010
rect 5200 9925 5205 9955
rect 5235 9925 5240 9955
rect 5200 9875 5240 9925
rect 5200 9845 5205 9875
rect 5235 9845 5240 9875
rect 5200 9795 5240 9845
rect 5200 9765 5205 9795
rect 5235 9765 5240 9795
rect 5200 9715 5240 9765
rect 5200 9685 5205 9715
rect 5235 9685 5240 9715
rect 5200 9635 5240 9685
rect 5200 9605 5205 9635
rect 5235 9605 5240 9635
rect 5200 9555 5240 9605
rect 5200 9525 5205 9555
rect 5235 9525 5240 9555
rect 5200 9475 5240 9525
rect 5200 9445 5205 9475
rect 5235 9445 5240 9475
rect 5200 9395 5240 9445
rect 5200 9365 5205 9395
rect 5235 9365 5240 9395
rect 5200 9310 5240 9365
rect 5200 9290 5210 9310
rect 5230 9290 5240 9310
rect 5200 9230 5240 9290
rect 5200 9210 5210 9230
rect 5230 9210 5240 9230
rect 5200 9150 5240 9210
rect 5200 9130 5210 9150
rect 5230 9130 5240 9150
rect 5200 9070 5240 9130
rect 5200 9050 5210 9070
rect 5230 9050 5240 9070
rect 5200 8995 5240 9050
rect 5200 8965 5205 8995
rect 5235 8965 5240 8995
rect 5200 8915 5240 8965
rect 5200 8885 5205 8915
rect 5235 8885 5240 8915
rect 5200 8835 5240 8885
rect 5200 8805 5205 8835
rect 5235 8805 5240 8835
rect 5200 8755 5240 8805
rect 5200 8725 5205 8755
rect 5235 8725 5240 8755
rect 5200 8675 5240 8725
rect 5200 8645 5205 8675
rect 5235 8645 5240 8675
rect 5200 8595 5240 8645
rect 5200 8565 5205 8595
rect 5235 8565 5240 8595
rect 5200 8515 5240 8565
rect 5200 8485 5205 8515
rect 5235 8485 5240 8515
rect 5200 8435 5240 8485
rect 5200 8405 5205 8435
rect 5235 8405 5240 8435
rect 5200 8350 5240 8405
rect 5200 8330 5210 8350
rect 5230 8330 5240 8350
rect 5200 8275 5240 8330
rect 5200 8245 5205 8275
rect 5235 8245 5240 8275
rect 5200 8195 5240 8245
rect 5200 8165 5205 8195
rect 5235 8165 5240 8195
rect 5200 8115 5240 8165
rect 5200 8085 5205 8115
rect 5235 8085 5240 8115
rect 5200 8035 5240 8085
rect 5200 8005 5205 8035
rect 5235 8005 5240 8035
rect 5200 7955 5240 8005
rect 5200 7925 5205 7955
rect 5235 7925 5240 7955
rect 5200 7875 5240 7925
rect 5200 7845 5205 7875
rect 5235 7845 5240 7875
rect 5200 7795 5240 7845
rect 5200 7765 5205 7795
rect 5235 7765 5240 7795
rect 5200 7715 5240 7765
rect 5200 7685 5205 7715
rect 5235 7685 5240 7715
rect 5200 7635 5240 7685
rect 5200 7605 5205 7635
rect 5235 7605 5240 7635
rect 5200 7555 5240 7605
rect 5200 7525 5205 7555
rect 5235 7525 5240 7555
rect 5200 7475 5240 7525
rect 5200 7445 5205 7475
rect 5235 7445 5240 7475
rect 5200 7395 5240 7445
rect 5200 7365 5205 7395
rect 5235 7365 5240 7395
rect 5200 7315 5240 7365
rect 5200 7285 5205 7315
rect 5235 7285 5240 7315
rect 5200 7235 5240 7285
rect 5200 7205 5205 7235
rect 5235 7205 5240 7235
rect 5200 7155 5240 7205
rect 5200 7125 5205 7155
rect 5235 7125 5240 7155
rect 5200 7075 5240 7125
rect 5200 7045 5205 7075
rect 5235 7045 5240 7075
rect 5200 6995 5240 7045
rect 5200 6965 5205 6995
rect 5235 6965 5240 6995
rect 5200 6910 5240 6965
rect 5200 6890 5210 6910
rect 5230 6890 5240 6910
rect 5200 6835 5240 6890
rect 5200 6805 5205 6835
rect 5235 6805 5240 6835
rect 5200 6755 5240 6805
rect 5200 6725 5205 6755
rect 5235 6725 5240 6755
rect 5200 6675 5240 6725
rect 5200 6645 5205 6675
rect 5235 6645 5240 6675
rect 5200 6595 5240 6645
rect 5200 6565 5205 6595
rect 5235 6565 5240 6595
rect 5200 6515 5240 6565
rect 5200 6485 5205 6515
rect 5235 6485 5240 6515
rect 5200 6435 5240 6485
rect 5200 6405 5205 6435
rect 5235 6405 5240 6435
rect 5200 6355 5240 6405
rect 5200 6325 5205 6355
rect 5235 6325 5240 6355
rect 5200 6275 5240 6325
rect 5200 6245 5205 6275
rect 5235 6245 5240 6275
rect 5200 6190 5240 6245
rect 5200 6170 5210 6190
rect 5230 6170 5240 6190
rect 5200 6110 5240 6170
rect 5200 6090 5210 6110
rect 5230 6090 5240 6110
rect 5200 6030 5240 6090
rect 5200 6010 5210 6030
rect 5230 6010 5240 6030
rect 5200 5950 5240 6010
rect 5200 5930 5210 5950
rect 5230 5930 5240 5950
rect 5200 5875 5240 5930
rect 5200 5845 5205 5875
rect 5235 5845 5240 5875
rect 5200 5795 5240 5845
rect 5200 5765 5205 5795
rect 5235 5765 5240 5795
rect 5200 5715 5240 5765
rect 5200 5685 5205 5715
rect 5235 5685 5240 5715
rect 5200 5635 5240 5685
rect 5200 5605 5205 5635
rect 5235 5605 5240 5635
rect 5200 5555 5240 5605
rect 5200 5525 5205 5555
rect 5235 5525 5240 5555
rect 5200 5475 5240 5525
rect 5200 5445 5205 5475
rect 5235 5445 5240 5475
rect 5200 5395 5240 5445
rect 5200 5365 5205 5395
rect 5235 5365 5240 5395
rect 5200 5315 5240 5365
rect 5200 5285 5205 5315
rect 5235 5285 5240 5315
rect 5200 5235 5240 5285
rect 5200 5205 5205 5235
rect 5235 5205 5240 5235
rect 5200 5155 5240 5205
rect 5200 5125 5205 5155
rect 5235 5125 5240 5155
rect 5200 5075 5240 5125
rect 5200 5045 5205 5075
rect 5235 5045 5240 5075
rect 5200 4995 5240 5045
rect 5200 4965 5205 4995
rect 5235 4965 5240 4995
rect 5200 4915 5240 4965
rect 5200 4885 5205 4915
rect 5235 4885 5240 4915
rect 5200 4830 5240 4885
rect 5200 4810 5210 4830
rect 5230 4810 5240 4830
rect 5200 4755 5240 4810
rect 5200 4725 5205 4755
rect 5235 4725 5240 4755
rect 5200 4675 5240 4725
rect 5200 4645 5205 4675
rect 5235 4645 5240 4675
rect 5200 4590 5240 4645
rect 5200 4570 5210 4590
rect 5230 4570 5240 4590
rect 5200 4515 5240 4570
rect 5200 4485 5205 4515
rect 5235 4485 5240 4515
rect 5200 4435 5240 4485
rect 5200 4405 5205 4435
rect 5235 4405 5240 4435
rect 5200 4355 5240 4405
rect 5200 4325 5205 4355
rect 5235 4325 5240 4355
rect 5200 4275 5240 4325
rect 5200 4245 5205 4275
rect 5235 4245 5240 4275
rect 5200 4195 5240 4245
rect 5200 4165 5205 4195
rect 5235 4165 5240 4195
rect 5200 4115 5240 4165
rect 5200 4085 5205 4115
rect 5235 4085 5240 4115
rect 5200 4035 5240 4085
rect 5200 4005 5205 4035
rect 5235 4005 5240 4035
rect 5200 3955 5240 4005
rect 5200 3925 5205 3955
rect 5235 3925 5240 3955
rect 5200 3875 5240 3925
rect 5200 3845 5205 3875
rect 5235 3845 5240 3875
rect 5200 3790 5240 3845
rect 5200 3770 5210 3790
rect 5230 3770 5240 3790
rect 5200 3715 5240 3770
rect 5200 3685 5205 3715
rect 5235 3685 5240 3715
rect 5200 3635 5240 3685
rect 5200 3605 5205 3635
rect 5235 3605 5240 3635
rect 5200 3550 5240 3605
rect 5200 3530 5210 3550
rect 5230 3530 5240 3550
rect 5200 3475 5240 3530
rect 5200 3445 5205 3475
rect 5235 3445 5240 3475
rect 5200 3395 5240 3445
rect 5200 3365 5205 3395
rect 5235 3365 5240 3395
rect 5200 3310 5240 3365
rect 5200 3290 5210 3310
rect 5230 3290 5240 3310
rect 5200 3235 5240 3290
rect 5200 3205 5205 3235
rect 5235 3205 5240 3235
rect 5200 3155 5240 3205
rect 5200 3125 5205 3155
rect 5235 3125 5240 3155
rect 5200 3075 5240 3125
rect 5200 3045 5205 3075
rect 5235 3045 5240 3075
rect 5200 2995 5240 3045
rect 5200 2965 5205 2995
rect 5235 2965 5240 2995
rect 5200 2915 5240 2965
rect 5200 2885 5205 2915
rect 5235 2885 5240 2915
rect 5200 2835 5240 2885
rect 5200 2805 5205 2835
rect 5235 2805 5240 2835
rect 5200 2755 5240 2805
rect 5200 2725 5205 2755
rect 5235 2725 5240 2755
rect 5200 2675 5240 2725
rect 5200 2645 5205 2675
rect 5235 2645 5240 2675
rect 5200 2595 5240 2645
rect 5200 2565 5205 2595
rect 5235 2565 5240 2595
rect 5200 2515 5240 2565
rect 5200 2485 5205 2515
rect 5235 2485 5240 2515
rect 5200 2435 5240 2485
rect 5200 2405 5205 2435
rect 5235 2405 5240 2435
rect 5200 2355 5240 2405
rect 5200 2325 5205 2355
rect 5235 2325 5240 2355
rect 5200 2275 5240 2325
rect 5200 2245 5205 2275
rect 5235 2245 5240 2275
rect 5200 2195 5240 2245
rect 5200 2165 5205 2195
rect 5235 2165 5240 2195
rect 5200 2115 5240 2165
rect 5200 2085 5205 2115
rect 5235 2085 5240 2115
rect 5200 2035 5240 2085
rect 5200 2005 5205 2035
rect 5235 2005 5240 2035
rect 5200 1955 5240 2005
rect 5200 1925 5205 1955
rect 5235 1925 5240 1955
rect 5200 1870 5240 1925
rect 5200 1850 5210 1870
rect 5230 1850 5240 1870
rect 5200 1790 5240 1850
rect 5200 1770 5210 1790
rect 5230 1770 5240 1790
rect 5200 1715 5240 1770
rect 5200 1685 5205 1715
rect 5235 1685 5240 1715
rect 5200 1635 5240 1685
rect 5200 1605 5205 1635
rect 5235 1605 5240 1635
rect 5200 1555 5240 1605
rect 5200 1525 5205 1555
rect 5235 1525 5240 1555
rect 5200 1475 5240 1525
rect 5200 1445 5205 1475
rect 5235 1445 5240 1475
rect 5200 1395 5240 1445
rect 5200 1365 5205 1395
rect 5235 1365 5240 1395
rect 5200 1315 5240 1365
rect 5200 1285 5205 1315
rect 5235 1285 5240 1315
rect 5200 1235 5240 1285
rect 5200 1205 5205 1235
rect 5235 1205 5240 1235
rect 5200 1155 5240 1205
rect 5200 1125 5205 1155
rect 5235 1125 5240 1155
rect 5200 1075 5240 1125
rect 5200 1045 5205 1075
rect 5235 1045 5240 1075
rect 5200 995 5240 1045
rect 5200 965 5205 995
rect 5235 965 5240 995
rect 5200 910 5240 965
rect 5200 890 5210 910
rect 5230 890 5240 910
rect 5200 835 5240 890
rect 5200 805 5205 835
rect 5235 805 5240 835
rect 5200 755 5240 805
rect 5200 725 5205 755
rect 5235 725 5240 755
rect 5200 675 5240 725
rect 5200 645 5205 675
rect 5235 645 5240 675
rect 5200 595 5240 645
rect 5200 565 5205 595
rect 5235 565 5240 595
rect 5200 515 5240 565
rect 5200 485 5205 515
rect 5235 485 5240 515
rect 5200 430 5240 485
rect 5200 410 5210 430
rect 5230 410 5240 430
rect 5200 350 5240 410
rect 5200 330 5210 350
rect 5230 330 5240 350
rect 5200 275 5240 330
rect 5200 245 5205 275
rect 5235 245 5240 275
rect 5200 195 5240 245
rect 5200 165 5205 195
rect 5235 165 5240 195
rect 5200 115 5240 165
rect 5200 85 5205 115
rect 5235 85 5240 115
rect 5200 35 5240 85
rect 5200 5 5205 35
rect 5235 5 5240 35
rect 5200 0 5240 5
rect 5280 15710 5320 15720
rect 5280 15690 5290 15710
rect 5310 15690 5320 15710
rect 5280 15630 5320 15690
rect 5280 15610 5290 15630
rect 5310 15610 5320 15630
rect 5280 15550 5320 15610
rect 5280 15530 5290 15550
rect 5310 15530 5320 15550
rect 5280 15470 5320 15530
rect 5280 15450 5290 15470
rect 5310 15450 5320 15470
rect 5280 15390 5320 15450
rect 5280 15370 5290 15390
rect 5310 15370 5320 15390
rect 5280 15310 5320 15370
rect 5280 15290 5290 15310
rect 5310 15290 5320 15310
rect 5280 15230 5320 15290
rect 5280 15210 5290 15230
rect 5310 15210 5320 15230
rect 5280 15150 5320 15210
rect 5280 15130 5290 15150
rect 5310 15130 5320 15150
rect 5280 15070 5320 15130
rect 5280 15050 5290 15070
rect 5310 15050 5320 15070
rect 5280 14990 5320 15050
rect 5280 14970 5290 14990
rect 5310 14970 5320 14990
rect 5280 14910 5320 14970
rect 5280 14890 5290 14910
rect 5310 14890 5320 14910
rect 5280 14830 5320 14890
rect 5280 14810 5290 14830
rect 5310 14810 5320 14830
rect 5280 14750 5320 14810
rect 5280 14730 5290 14750
rect 5310 14730 5320 14750
rect 5280 14670 5320 14730
rect 5280 14650 5290 14670
rect 5310 14650 5320 14670
rect 5280 14590 5320 14650
rect 5280 14570 5290 14590
rect 5310 14570 5320 14590
rect 5280 14510 5320 14570
rect 5280 14490 5290 14510
rect 5310 14490 5320 14510
rect 5280 14430 5320 14490
rect 5280 14410 5290 14430
rect 5310 14410 5320 14430
rect 5280 14350 5320 14410
rect 5280 14330 5290 14350
rect 5310 14330 5320 14350
rect 5280 14270 5320 14330
rect 5280 14250 5290 14270
rect 5310 14250 5320 14270
rect 5280 14190 5320 14250
rect 5280 14170 5290 14190
rect 5310 14170 5320 14190
rect 5280 14110 5320 14170
rect 5280 14090 5290 14110
rect 5310 14090 5320 14110
rect 5280 14030 5320 14090
rect 5280 14010 5290 14030
rect 5310 14010 5320 14030
rect 5280 13950 5320 14010
rect 5280 13930 5290 13950
rect 5310 13930 5320 13950
rect 5280 13870 5320 13930
rect 5280 13850 5290 13870
rect 5310 13850 5320 13870
rect 5280 13790 5320 13850
rect 5280 13770 5290 13790
rect 5310 13770 5320 13790
rect 5280 13710 5320 13770
rect 5280 13690 5290 13710
rect 5310 13690 5320 13710
rect 5280 13630 5320 13690
rect 5280 13610 5290 13630
rect 5310 13610 5320 13630
rect 5280 13550 5320 13610
rect 5280 13530 5290 13550
rect 5310 13530 5320 13550
rect 5280 13470 5320 13530
rect 5280 13450 5290 13470
rect 5310 13450 5320 13470
rect 5280 13390 5320 13450
rect 5280 13370 5290 13390
rect 5310 13370 5320 13390
rect 5280 13310 5320 13370
rect 5280 13290 5290 13310
rect 5310 13290 5320 13310
rect 5280 13230 5320 13290
rect 5280 13210 5290 13230
rect 5310 13210 5320 13230
rect 5280 13150 5320 13210
rect 5280 13130 5290 13150
rect 5310 13130 5320 13150
rect 5280 13070 5320 13130
rect 5280 13050 5290 13070
rect 5310 13050 5320 13070
rect 5280 12990 5320 13050
rect 5280 12970 5290 12990
rect 5310 12970 5320 12990
rect 5280 12910 5320 12970
rect 5280 12890 5290 12910
rect 5310 12890 5320 12910
rect 5280 12830 5320 12890
rect 5280 12810 5290 12830
rect 5310 12810 5320 12830
rect 5280 12750 5320 12810
rect 5280 12730 5290 12750
rect 5310 12730 5320 12750
rect 5280 12670 5320 12730
rect 5280 12650 5290 12670
rect 5310 12650 5320 12670
rect 5280 12590 5320 12650
rect 5280 12570 5290 12590
rect 5310 12570 5320 12590
rect 5280 12510 5320 12570
rect 5280 12490 5290 12510
rect 5310 12490 5320 12510
rect 5280 12430 5320 12490
rect 5280 12410 5290 12430
rect 5310 12410 5320 12430
rect 5280 12350 5320 12410
rect 5280 12330 5290 12350
rect 5310 12330 5320 12350
rect 5280 12270 5320 12330
rect 5280 12250 5290 12270
rect 5310 12250 5320 12270
rect 5280 12190 5320 12250
rect 5280 12170 5290 12190
rect 5310 12170 5320 12190
rect 5280 12110 5320 12170
rect 5280 12090 5290 12110
rect 5310 12090 5320 12110
rect 5280 12030 5320 12090
rect 5280 12010 5290 12030
rect 5310 12010 5320 12030
rect 5280 11950 5320 12010
rect 5280 11930 5290 11950
rect 5310 11930 5320 11950
rect 5280 11870 5320 11930
rect 5280 11850 5290 11870
rect 5310 11850 5320 11870
rect 5280 11790 5320 11850
rect 5280 11770 5290 11790
rect 5310 11770 5320 11790
rect 5280 11710 5320 11770
rect 5280 11690 5290 11710
rect 5310 11690 5320 11710
rect 5280 11630 5320 11690
rect 5280 11610 5290 11630
rect 5310 11610 5320 11630
rect 5280 11550 5320 11610
rect 5280 11530 5290 11550
rect 5310 11530 5320 11550
rect 5280 11470 5320 11530
rect 5280 11450 5290 11470
rect 5310 11450 5320 11470
rect 5280 11390 5320 11450
rect 5280 11370 5290 11390
rect 5310 11370 5320 11390
rect 5280 11310 5320 11370
rect 5280 11290 5290 11310
rect 5310 11290 5320 11310
rect 5280 11230 5320 11290
rect 5280 11210 5290 11230
rect 5310 11210 5320 11230
rect 5280 11150 5320 11210
rect 5280 11130 5290 11150
rect 5310 11130 5320 11150
rect 5280 11070 5320 11130
rect 5280 11050 5290 11070
rect 5310 11050 5320 11070
rect 5280 10990 5320 11050
rect 5280 10970 5290 10990
rect 5310 10970 5320 10990
rect 5280 10910 5320 10970
rect 5280 10890 5290 10910
rect 5310 10890 5320 10910
rect 5280 10830 5320 10890
rect 5280 10810 5290 10830
rect 5310 10810 5320 10830
rect 5280 10750 5320 10810
rect 5280 10730 5290 10750
rect 5310 10730 5320 10750
rect 5280 10670 5320 10730
rect 5280 10650 5290 10670
rect 5310 10650 5320 10670
rect 5280 10590 5320 10650
rect 5280 10570 5290 10590
rect 5310 10570 5320 10590
rect 5280 10510 5320 10570
rect 5280 10490 5290 10510
rect 5310 10490 5320 10510
rect 5280 10430 5320 10490
rect 5280 10410 5290 10430
rect 5310 10410 5320 10430
rect 5280 10350 5320 10410
rect 5280 10330 5290 10350
rect 5310 10330 5320 10350
rect 5280 10270 5320 10330
rect 5280 10250 5290 10270
rect 5310 10250 5320 10270
rect 5280 10190 5320 10250
rect 5280 10170 5290 10190
rect 5310 10170 5320 10190
rect 5280 10110 5320 10170
rect 5280 10090 5290 10110
rect 5310 10090 5320 10110
rect 5280 10030 5320 10090
rect 5280 10010 5290 10030
rect 5310 10010 5320 10030
rect 5280 9950 5320 10010
rect 5280 9930 5290 9950
rect 5310 9930 5320 9950
rect 5280 9870 5320 9930
rect 5280 9850 5290 9870
rect 5310 9850 5320 9870
rect 5280 9790 5320 9850
rect 5280 9770 5290 9790
rect 5310 9770 5320 9790
rect 5280 9710 5320 9770
rect 5280 9690 5290 9710
rect 5310 9690 5320 9710
rect 5280 9630 5320 9690
rect 5280 9610 5290 9630
rect 5310 9610 5320 9630
rect 5280 9550 5320 9610
rect 5280 9530 5290 9550
rect 5310 9530 5320 9550
rect 5280 9470 5320 9530
rect 5280 9450 5290 9470
rect 5310 9450 5320 9470
rect 5280 9390 5320 9450
rect 5280 9370 5290 9390
rect 5310 9370 5320 9390
rect 5280 9310 5320 9370
rect 5280 9290 5290 9310
rect 5310 9290 5320 9310
rect 5280 9230 5320 9290
rect 5280 9210 5290 9230
rect 5310 9210 5320 9230
rect 5280 9150 5320 9210
rect 5280 9130 5290 9150
rect 5310 9130 5320 9150
rect 5280 9070 5320 9130
rect 5280 9050 5290 9070
rect 5310 9050 5320 9070
rect 5280 8990 5320 9050
rect 5280 8970 5290 8990
rect 5310 8970 5320 8990
rect 5280 8910 5320 8970
rect 5280 8890 5290 8910
rect 5310 8890 5320 8910
rect 5280 8830 5320 8890
rect 5280 8810 5290 8830
rect 5310 8810 5320 8830
rect 5280 8750 5320 8810
rect 5280 8730 5290 8750
rect 5310 8730 5320 8750
rect 5280 8670 5320 8730
rect 5280 8650 5290 8670
rect 5310 8650 5320 8670
rect 5280 8590 5320 8650
rect 5280 8570 5290 8590
rect 5310 8570 5320 8590
rect 5280 8510 5320 8570
rect 5280 8490 5290 8510
rect 5310 8490 5320 8510
rect 5280 8430 5320 8490
rect 5280 8410 5290 8430
rect 5310 8410 5320 8430
rect 5280 8350 5320 8410
rect 5280 8330 5290 8350
rect 5310 8330 5320 8350
rect 5280 8270 5320 8330
rect 5280 8250 5290 8270
rect 5310 8250 5320 8270
rect 5280 8190 5320 8250
rect 5280 8170 5290 8190
rect 5310 8170 5320 8190
rect 5280 8110 5320 8170
rect 5280 8090 5290 8110
rect 5310 8090 5320 8110
rect 5280 8030 5320 8090
rect 5280 8010 5290 8030
rect 5310 8010 5320 8030
rect 5280 7950 5320 8010
rect 5280 7930 5290 7950
rect 5310 7930 5320 7950
rect 5280 7870 5320 7930
rect 5280 7850 5290 7870
rect 5310 7850 5320 7870
rect 5280 7790 5320 7850
rect 5280 7770 5290 7790
rect 5310 7770 5320 7790
rect 5280 7710 5320 7770
rect 5280 7690 5290 7710
rect 5310 7690 5320 7710
rect 5280 7630 5320 7690
rect 5280 7610 5290 7630
rect 5310 7610 5320 7630
rect 5280 7550 5320 7610
rect 5280 7530 5290 7550
rect 5310 7530 5320 7550
rect 5280 7470 5320 7530
rect 5280 7450 5290 7470
rect 5310 7450 5320 7470
rect 5280 7390 5320 7450
rect 5280 7370 5290 7390
rect 5310 7370 5320 7390
rect 5280 7310 5320 7370
rect 5280 7290 5290 7310
rect 5310 7290 5320 7310
rect 5280 7230 5320 7290
rect 5280 7210 5290 7230
rect 5310 7210 5320 7230
rect 5280 7150 5320 7210
rect 5280 7130 5290 7150
rect 5310 7130 5320 7150
rect 5280 7070 5320 7130
rect 5280 7050 5290 7070
rect 5310 7050 5320 7070
rect 5280 6990 5320 7050
rect 5280 6970 5290 6990
rect 5310 6970 5320 6990
rect 5280 6910 5320 6970
rect 5280 6890 5290 6910
rect 5310 6890 5320 6910
rect 5280 6830 5320 6890
rect 5280 6810 5290 6830
rect 5310 6810 5320 6830
rect 5280 6750 5320 6810
rect 5280 6730 5290 6750
rect 5310 6730 5320 6750
rect 5280 6670 5320 6730
rect 5280 6650 5290 6670
rect 5310 6650 5320 6670
rect 5280 6590 5320 6650
rect 5280 6570 5290 6590
rect 5310 6570 5320 6590
rect 5280 6510 5320 6570
rect 5280 6490 5290 6510
rect 5310 6490 5320 6510
rect 5280 6430 5320 6490
rect 5280 6410 5290 6430
rect 5310 6410 5320 6430
rect 5280 6350 5320 6410
rect 5280 6330 5290 6350
rect 5310 6330 5320 6350
rect 5280 6270 5320 6330
rect 5280 6250 5290 6270
rect 5310 6250 5320 6270
rect 5280 6190 5320 6250
rect 5280 6170 5290 6190
rect 5310 6170 5320 6190
rect 5280 6110 5320 6170
rect 5280 6090 5290 6110
rect 5310 6090 5320 6110
rect 5280 6030 5320 6090
rect 5280 6010 5290 6030
rect 5310 6010 5320 6030
rect 5280 5950 5320 6010
rect 5280 5930 5290 5950
rect 5310 5930 5320 5950
rect 5280 5870 5320 5930
rect 5280 5850 5290 5870
rect 5310 5850 5320 5870
rect 5280 5790 5320 5850
rect 5280 5770 5290 5790
rect 5310 5770 5320 5790
rect 5280 5710 5320 5770
rect 5280 5690 5290 5710
rect 5310 5690 5320 5710
rect 5280 5630 5320 5690
rect 5280 5610 5290 5630
rect 5310 5610 5320 5630
rect 5280 5550 5320 5610
rect 5280 5530 5290 5550
rect 5310 5530 5320 5550
rect 5280 5470 5320 5530
rect 5280 5450 5290 5470
rect 5310 5450 5320 5470
rect 5280 5390 5320 5450
rect 5280 5370 5290 5390
rect 5310 5370 5320 5390
rect 5280 5310 5320 5370
rect 5280 5290 5290 5310
rect 5310 5290 5320 5310
rect 5280 5230 5320 5290
rect 5280 5210 5290 5230
rect 5310 5210 5320 5230
rect 5280 5150 5320 5210
rect 5280 5130 5290 5150
rect 5310 5130 5320 5150
rect 5280 5070 5320 5130
rect 5280 5050 5290 5070
rect 5310 5050 5320 5070
rect 5280 4990 5320 5050
rect 5280 4970 5290 4990
rect 5310 4970 5320 4990
rect 5280 4910 5320 4970
rect 5280 4890 5290 4910
rect 5310 4890 5320 4910
rect 5280 4830 5320 4890
rect 5280 4810 5290 4830
rect 5310 4810 5320 4830
rect 5280 4750 5320 4810
rect 5280 4730 5290 4750
rect 5310 4730 5320 4750
rect 5280 4670 5320 4730
rect 5280 4650 5290 4670
rect 5310 4650 5320 4670
rect 5280 4590 5320 4650
rect 5280 4570 5290 4590
rect 5310 4570 5320 4590
rect 5280 4510 5320 4570
rect 5280 4490 5290 4510
rect 5310 4490 5320 4510
rect 5280 4430 5320 4490
rect 5280 4410 5290 4430
rect 5310 4410 5320 4430
rect 5280 4350 5320 4410
rect 5280 4330 5290 4350
rect 5310 4330 5320 4350
rect 5280 4270 5320 4330
rect 5280 4250 5290 4270
rect 5310 4250 5320 4270
rect 5280 4190 5320 4250
rect 5280 4170 5290 4190
rect 5310 4170 5320 4190
rect 5280 4110 5320 4170
rect 5280 4090 5290 4110
rect 5310 4090 5320 4110
rect 5280 4030 5320 4090
rect 5280 4010 5290 4030
rect 5310 4010 5320 4030
rect 5280 3950 5320 4010
rect 5280 3930 5290 3950
rect 5310 3930 5320 3950
rect 5280 3870 5320 3930
rect 5280 3850 5290 3870
rect 5310 3850 5320 3870
rect 5280 3790 5320 3850
rect 5280 3770 5290 3790
rect 5310 3770 5320 3790
rect 5280 3710 5320 3770
rect 5280 3690 5290 3710
rect 5310 3690 5320 3710
rect 5280 3630 5320 3690
rect 5280 3610 5290 3630
rect 5310 3610 5320 3630
rect 5280 3550 5320 3610
rect 5280 3530 5290 3550
rect 5310 3530 5320 3550
rect 5280 3470 5320 3530
rect 5280 3450 5290 3470
rect 5310 3450 5320 3470
rect 5280 3390 5320 3450
rect 5280 3370 5290 3390
rect 5310 3370 5320 3390
rect 5280 3310 5320 3370
rect 5280 3290 5290 3310
rect 5310 3290 5320 3310
rect 5280 3230 5320 3290
rect 5280 3210 5290 3230
rect 5310 3210 5320 3230
rect 5280 3150 5320 3210
rect 5280 3130 5290 3150
rect 5310 3130 5320 3150
rect 5280 3070 5320 3130
rect 5280 3050 5290 3070
rect 5310 3050 5320 3070
rect 5280 2990 5320 3050
rect 5280 2970 5290 2990
rect 5310 2970 5320 2990
rect 5280 2910 5320 2970
rect 5280 2890 5290 2910
rect 5310 2890 5320 2910
rect 5280 2830 5320 2890
rect 5280 2810 5290 2830
rect 5310 2810 5320 2830
rect 5280 2750 5320 2810
rect 5280 2730 5290 2750
rect 5310 2730 5320 2750
rect 5280 2670 5320 2730
rect 5280 2650 5290 2670
rect 5310 2650 5320 2670
rect 5280 2590 5320 2650
rect 5280 2570 5290 2590
rect 5310 2570 5320 2590
rect 5280 2510 5320 2570
rect 5280 2490 5290 2510
rect 5310 2490 5320 2510
rect 5280 2430 5320 2490
rect 5280 2410 5290 2430
rect 5310 2410 5320 2430
rect 5280 2350 5320 2410
rect 5280 2330 5290 2350
rect 5310 2330 5320 2350
rect 5280 2270 5320 2330
rect 5280 2250 5290 2270
rect 5310 2250 5320 2270
rect 5280 2190 5320 2250
rect 5280 2170 5290 2190
rect 5310 2170 5320 2190
rect 5280 2110 5320 2170
rect 5280 2090 5290 2110
rect 5310 2090 5320 2110
rect 5280 2030 5320 2090
rect 5280 2010 5290 2030
rect 5310 2010 5320 2030
rect 5280 1950 5320 2010
rect 5280 1930 5290 1950
rect 5310 1930 5320 1950
rect 5280 1870 5320 1930
rect 5280 1850 5290 1870
rect 5310 1850 5320 1870
rect 5280 1790 5320 1850
rect 5280 1770 5290 1790
rect 5310 1770 5320 1790
rect 5280 1710 5320 1770
rect 5280 1690 5290 1710
rect 5310 1690 5320 1710
rect 5280 1630 5320 1690
rect 5280 1610 5290 1630
rect 5310 1610 5320 1630
rect 5280 1550 5320 1610
rect 5280 1530 5290 1550
rect 5310 1530 5320 1550
rect 5280 1470 5320 1530
rect 5280 1450 5290 1470
rect 5310 1450 5320 1470
rect 5280 1390 5320 1450
rect 5280 1370 5290 1390
rect 5310 1370 5320 1390
rect 5280 1310 5320 1370
rect 5280 1290 5290 1310
rect 5310 1290 5320 1310
rect 5280 1230 5320 1290
rect 5280 1210 5290 1230
rect 5310 1210 5320 1230
rect 5280 1150 5320 1210
rect 5280 1130 5290 1150
rect 5310 1130 5320 1150
rect 5280 1070 5320 1130
rect 5280 1050 5290 1070
rect 5310 1050 5320 1070
rect 5280 990 5320 1050
rect 5280 970 5290 990
rect 5310 970 5320 990
rect 5280 910 5320 970
rect 5280 890 5290 910
rect 5310 890 5320 910
rect 5280 830 5320 890
rect 5280 810 5290 830
rect 5310 810 5320 830
rect 5280 750 5320 810
rect 5280 730 5290 750
rect 5310 730 5320 750
rect 5280 670 5320 730
rect 5280 650 5290 670
rect 5310 650 5320 670
rect 5280 590 5320 650
rect 5280 570 5290 590
rect 5310 570 5320 590
rect 5280 510 5320 570
rect 5280 490 5290 510
rect 5310 490 5320 510
rect 5280 430 5320 490
rect 5280 410 5290 430
rect 5310 410 5320 430
rect 5280 350 5320 410
rect 5280 330 5290 350
rect 5310 330 5320 350
rect 5280 270 5320 330
rect 5280 250 5290 270
rect 5310 250 5320 270
rect 5280 190 5320 250
rect 5280 170 5290 190
rect 5310 170 5320 190
rect 5280 110 5320 170
rect 5280 90 5290 110
rect 5310 90 5320 110
rect 5280 30 5320 90
rect 5280 10 5290 30
rect 5310 10 5320 30
rect 5280 0 5320 10
rect 5360 15715 5400 15720
rect 5360 15685 5365 15715
rect 5395 15685 5400 15715
rect 5360 15635 5400 15685
rect 5360 15605 5365 15635
rect 5395 15605 5400 15635
rect 5360 15555 5400 15605
rect 5360 15525 5365 15555
rect 5395 15525 5400 15555
rect 5360 15475 5400 15525
rect 5360 15445 5365 15475
rect 5395 15445 5400 15475
rect 5360 15395 5400 15445
rect 5360 15365 5365 15395
rect 5395 15365 5400 15395
rect 5360 15315 5400 15365
rect 5360 15285 5365 15315
rect 5395 15285 5400 15315
rect 5360 15235 5400 15285
rect 5360 15205 5365 15235
rect 5395 15205 5400 15235
rect 5360 15155 5400 15205
rect 5360 15125 5365 15155
rect 5395 15125 5400 15155
rect 5360 15070 5400 15125
rect 5360 15050 5370 15070
rect 5390 15050 5400 15070
rect 5360 14995 5400 15050
rect 5360 14965 5365 14995
rect 5395 14965 5400 14995
rect 5360 14915 5400 14965
rect 5360 14885 5365 14915
rect 5395 14885 5400 14915
rect 5360 14835 5400 14885
rect 5360 14805 5365 14835
rect 5395 14805 5400 14835
rect 5360 14755 5400 14805
rect 5360 14725 5365 14755
rect 5395 14725 5400 14755
rect 5360 14675 5400 14725
rect 5360 14645 5365 14675
rect 5395 14645 5400 14675
rect 5360 14595 5400 14645
rect 5360 14565 5365 14595
rect 5395 14565 5400 14595
rect 5360 14515 5400 14565
rect 5360 14485 5365 14515
rect 5395 14485 5400 14515
rect 5360 14435 5400 14485
rect 5360 14405 5365 14435
rect 5395 14405 5400 14435
rect 5360 14350 5400 14405
rect 5360 14330 5370 14350
rect 5390 14330 5400 14350
rect 5360 14270 5400 14330
rect 5360 14250 5370 14270
rect 5390 14250 5400 14270
rect 5360 14190 5400 14250
rect 5360 14170 5370 14190
rect 5390 14170 5400 14190
rect 5360 14110 5400 14170
rect 5360 14090 5370 14110
rect 5390 14090 5400 14110
rect 5360 14035 5400 14090
rect 5360 14005 5365 14035
rect 5395 14005 5400 14035
rect 5360 13955 5400 14005
rect 5360 13925 5365 13955
rect 5395 13925 5400 13955
rect 5360 13875 5400 13925
rect 5360 13845 5365 13875
rect 5395 13845 5400 13875
rect 5360 13795 5400 13845
rect 5360 13765 5365 13795
rect 5395 13765 5400 13795
rect 5360 13715 5400 13765
rect 5360 13685 5365 13715
rect 5395 13685 5400 13715
rect 5360 13635 5400 13685
rect 5360 13605 5365 13635
rect 5395 13605 5400 13635
rect 5360 13555 5400 13605
rect 5360 13525 5365 13555
rect 5395 13525 5400 13555
rect 5360 13475 5400 13525
rect 5360 13445 5365 13475
rect 5395 13445 5400 13475
rect 5360 13390 5400 13445
rect 5360 13370 5370 13390
rect 5390 13370 5400 13390
rect 5360 13310 5400 13370
rect 5360 13290 5370 13310
rect 5390 13290 5400 13310
rect 5360 13230 5400 13290
rect 5360 13210 5370 13230
rect 5390 13210 5400 13230
rect 5360 13150 5400 13210
rect 5360 13130 5370 13150
rect 5390 13130 5400 13150
rect 5360 13075 5400 13130
rect 5360 13045 5365 13075
rect 5395 13045 5400 13075
rect 5360 12995 5400 13045
rect 5360 12965 5365 12995
rect 5395 12965 5400 12995
rect 5360 12915 5400 12965
rect 5360 12885 5365 12915
rect 5395 12885 5400 12915
rect 5360 12835 5400 12885
rect 5360 12805 5365 12835
rect 5395 12805 5400 12835
rect 5360 12755 5400 12805
rect 5360 12725 5365 12755
rect 5395 12725 5400 12755
rect 5360 12675 5400 12725
rect 5360 12645 5365 12675
rect 5395 12645 5400 12675
rect 5360 12595 5400 12645
rect 5360 12565 5365 12595
rect 5395 12565 5400 12595
rect 5360 12515 5400 12565
rect 5360 12485 5365 12515
rect 5395 12485 5400 12515
rect 5360 12430 5400 12485
rect 5360 12410 5370 12430
rect 5390 12410 5400 12430
rect 5360 12355 5400 12410
rect 5360 12325 5365 12355
rect 5395 12325 5400 12355
rect 5360 12275 5400 12325
rect 5360 12245 5365 12275
rect 5395 12245 5400 12275
rect 5360 12195 5400 12245
rect 5360 12165 5365 12195
rect 5395 12165 5400 12195
rect 5360 12115 5400 12165
rect 5360 12085 5365 12115
rect 5395 12085 5400 12115
rect 5360 12035 5400 12085
rect 5360 12005 5365 12035
rect 5395 12005 5400 12035
rect 5360 11955 5400 12005
rect 5360 11925 5365 11955
rect 5395 11925 5400 11955
rect 5360 11875 5400 11925
rect 5360 11845 5365 11875
rect 5395 11845 5400 11875
rect 5360 11795 5400 11845
rect 5360 11765 5365 11795
rect 5395 11765 5400 11795
rect 5360 11715 5400 11765
rect 5360 11685 5365 11715
rect 5395 11685 5400 11715
rect 5360 11635 5400 11685
rect 5360 11605 5365 11635
rect 5395 11605 5400 11635
rect 5360 11555 5400 11605
rect 5360 11525 5365 11555
rect 5395 11525 5400 11555
rect 5360 11475 5400 11525
rect 5360 11445 5365 11475
rect 5395 11445 5400 11475
rect 5360 11395 5400 11445
rect 5360 11365 5365 11395
rect 5395 11365 5400 11395
rect 5360 11315 5400 11365
rect 5360 11285 5365 11315
rect 5395 11285 5400 11315
rect 5360 11235 5400 11285
rect 5360 11205 5365 11235
rect 5395 11205 5400 11235
rect 5360 11155 5400 11205
rect 5360 11125 5365 11155
rect 5395 11125 5400 11155
rect 5360 11075 5400 11125
rect 5360 11045 5365 11075
rect 5395 11045 5400 11075
rect 5360 10990 5400 11045
rect 5360 10970 5370 10990
rect 5390 10970 5400 10990
rect 5360 10915 5400 10970
rect 5360 10885 5365 10915
rect 5395 10885 5400 10915
rect 5360 10835 5400 10885
rect 5360 10805 5365 10835
rect 5395 10805 5400 10835
rect 5360 10755 5400 10805
rect 5360 10725 5365 10755
rect 5395 10725 5400 10755
rect 5360 10675 5400 10725
rect 5360 10645 5365 10675
rect 5395 10645 5400 10675
rect 5360 10595 5400 10645
rect 5360 10565 5365 10595
rect 5395 10565 5400 10595
rect 5360 10515 5400 10565
rect 5360 10485 5365 10515
rect 5395 10485 5400 10515
rect 5360 10435 5400 10485
rect 5360 10405 5365 10435
rect 5395 10405 5400 10435
rect 5360 10355 5400 10405
rect 5360 10325 5365 10355
rect 5395 10325 5400 10355
rect 5360 10270 5400 10325
rect 5360 10250 5370 10270
rect 5390 10250 5400 10270
rect 5360 10190 5400 10250
rect 5360 10170 5370 10190
rect 5390 10170 5400 10190
rect 5360 10110 5400 10170
rect 5360 10090 5370 10110
rect 5390 10090 5400 10110
rect 5360 10030 5400 10090
rect 5360 10010 5370 10030
rect 5390 10010 5400 10030
rect 5360 9955 5400 10010
rect 5360 9925 5365 9955
rect 5395 9925 5400 9955
rect 5360 9875 5400 9925
rect 5360 9845 5365 9875
rect 5395 9845 5400 9875
rect 5360 9795 5400 9845
rect 5360 9765 5365 9795
rect 5395 9765 5400 9795
rect 5360 9715 5400 9765
rect 5360 9685 5365 9715
rect 5395 9685 5400 9715
rect 5360 9635 5400 9685
rect 5360 9605 5365 9635
rect 5395 9605 5400 9635
rect 5360 9555 5400 9605
rect 5360 9525 5365 9555
rect 5395 9525 5400 9555
rect 5360 9475 5400 9525
rect 5360 9445 5365 9475
rect 5395 9445 5400 9475
rect 5360 9395 5400 9445
rect 5360 9365 5365 9395
rect 5395 9365 5400 9395
rect 5360 9310 5400 9365
rect 5360 9290 5370 9310
rect 5390 9290 5400 9310
rect 5360 9230 5400 9290
rect 5360 9210 5370 9230
rect 5390 9210 5400 9230
rect 5360 9150 5400 9210
rect 5360 9130 5370 9150
rect 5390 9130 5400 9150
rect 5360 9070 5400 9130
rect 5360 9050 5370 9070
rect 5390 9050 5400 9070
rect 5360 8995 5400 9050
rect 5360 8965 5365 8995
rect 5395 8965 5400 8995
rect 5360 8915 5400 8965
rect 5360 8885 5365 8915
rect 5395 8885 5400 8915
rect 5360 8835 5400 8885
rect 5360 8805 5365 8835
rect 5395 8805 5400 8835
rect 5360 8755 5400 8805
rect 5360 8725 5365 8755
rect 5395 8725 5400 8755
rect 5360 8675 5400 8725
rect 5360 8645 5365 8675
rect 5395 8645 5400 8675
rect 5360 8595 5400 8645
rect 5360 8565 5365 8595
rect 5395 8565 5400 8595
rect 5360 8515 5400 8565
rect 5360 8485 5365 8515
rect 5395 8485 5400 8515
rect 5360 8435 5400 8485
rect 5360 8405 5365 8435
rect 5395 8405 5400 8435
rect 5360 8350 5400 8405
rect 5360 8330 5370 8350
rect 5390 8330 5400 8350
rect 5360 8275 5400 8330
rect 5360 8245 5365 8275
rect 5395 8245 5400 8275
rect 5360 8195 5400 8245
rect 5360 8165 5365 8195
rect 5395 8165 5400 8195
rect 5360 8115 5400 8165
rect 5360 8085 5365 8115
rect 5395 8085 5400 8115
rect 5360 8035 5400 8085
rect 5360 8005 5365 8035
rect 5395 8005 5400 8035
rect 5360 7955 5400 8005
rect 5360 7925 5365 7955
rect 5395 7925 5400 7955
rect 5360 7875 5400 7925
rect 5360 7845 5365 7875
rect 5395 7845 5400 7875
rect 5360 7795 5400 7845
rect 5360 7765 5365 7795
rect 5395 7765 5400 7795
rect 5360 7715 5400 7765
rect 5360 7685 5365 7715
rect 5395 7685 5400 7715
rect 5360 7635 5400 7685
rect 5360 7605 5365 7635
rect 5395 7605 5400 7635
rect 5360 7555 5400 7605
rect 5360 7525 5365 7555
rect 5395 7525 5400 7555
rect 5360 7475 5400 7525
rect 5360 7445 5365 7475
rect 5395 7445 5400 7475
rect 5360 7395 5400 7445
rect 5360 7365 5365 7395
rect 5395 7365 5400 7395
rect 5360 7315 5400 7365
rect 5360 7285 5365 7315
rect 5395 7285 5400 7315
rect 5360 7235 5400 7285
rect 5360 7205 5365 7235
rect 5395 7205 5400 7235
rect 5360 7155 5400 7205
rect 5360 7125 5365 7155
rect 5395 7125 5400 7155
rect 5360 7075 5400 7125
rect 5360 7045 5365 7075
rect 5395 7045 5400 7075
rect 5360 6995 5400 7045
rect 5360 6965 5365 6995
rect 5395 6965 5400 6995
rect 5360 6910 5400 6965
rect 5360 6890 5370 6910
rect 5390 6890 5400 6910
rect 5360 6835 5400 6890
rect 5360 6805 5365 6835
rect 5395 6805 5400 6835
rect 5360 6755 5400 6805
rect 5360 6725 5365 6755
rect 5395 6725 5400 6755
rect 5360 6675 5400 6725
rect 5360 6645 5365 6675
rect 5395 6645 5400 6675
rect 5360 6595 5400 6645
rect 5360 6565 5365 6595
rect 5395 6565 5400 6595
rect 5360 6515 5400 6565
rect 5360 6485 5365 6515
rect 5395 6485 5400 6515
rect 5360 6435 5400 6485
rect 5360 6405 5365 6435
rect 5395 6405 5400 6435
rect 5360 6355 5400 6405
rect 5360 6325 5365 6355
rect 5395 6325 5400 6355
rect 5360 6275 5400 6325
rect 5360 6245 5365 6275
rect 5395 6245 5400 6275
rect 5360 6190 5400 6245
rect 5360 6170 5370 6190
rect 5390 6170 5400 6190
rect 5360 6110 5400 6170
rect 5360 6090 5370 6110
rect 5390 6090 5400 6110
rect 5360 6030 5400 6090
rect 5360 6010 5370 6030
rect 5390 6010 5400 6030
rect 5360 5950 5400 6010
rect 5360 5930 5370 5950
rect 5390 5930 5400 5950
rect 5360 5875 5400 5930
rect 5360 5845 5365 5875
rect 5395 5845 5400 5875
rect 5360 5795 5400 5845
rect 5360 5765 5365 5795
rect 5395 5765 5400 5795
rect 5360 5715 5400 5765
rect 5360 5685 5365 5715
rect 5395 5685 5400 5715
rect 5360 5635 5400 5685
rect 5360 5605 5365 5635
rect 5395 5605 5400 5635
rect 5360 5555 5400 5605
rect 5360 5525 5365 5555
rect 5395 5525 5400 5555
rect 5360 5475 5400 5525
rect 5360 5445 5365 5475
rect 5395 5445 5400 5475
rect 5360 5395 5400 5445
rect 5360 5365 5365 5395
rect 5395 5365 5400 5395
rect 5360 5315 5400 5365
rect 5360 5285 5365 5315
rect 5395 5285 5400 5315
rect 5360 5235 5400 5285
rect 5360 5205 5365 5235
rect 5395 5205 5400 5235
rect 5360 5155 5400 5205
rect 5360 5125 5365 5155
rect 5395 5125 5400 5155
rect 5360 5075 5400 5125
rect 5360 5045 5365 5075
rect 5395 5045 5400 5075
rect 5360 4995 5400 5045
rect 5360 4965 5365 4995
rect 5395 4965 5400 4995
rect 5360 4915 5400 4965
rect 5360 4885 5365 4915
rect 5395 4885 5400 4915
rect 5360 4830 5400 4885
rect 5360 4810 5370 4830
rect 5390 4810 5400 4830
rect 5360 4755 5400 4810
rect 5360 4725 5365 4755
rect 5395 4725 5400 4755
rect 5360 4675 5400 4725
rect 5360 4645 5365 4675
rect 5395 4645 5400 4675
rect 5360 4590 5400 4645
rect 5360 4570 5370 4590
rect 5390 4570 5400 4590
rect 5360 4515 5400 4570
rect 5360 4485 5365 4515
rect 5395 4485 5400 4515
rect 5360 4435 5400 4485
rect 5360 4405 5365 4435
rect 5395 4405 5400 4435
rect 5360 4355 5400 4405
rect 5360 4325 5365 4355
rect 5395 4325 5400 4355
rect 5360 4275 5400 4325
rect 5360 4245 5365 4275
rect 5395 4245 5400 4275
rect 5360 4195 5400 4245
rect 5360 4165 5365 4195
rect 5395 4165 5400 4195
rect 5360 4115 5400 4165
rect 5360 4085 5365 4115
rect 5395 4085 5400 4115
rect 5360 4035 5400 4085
rect 5360 4005 5365 4035
rect 5395 4005 5400 4035
rect 5360 3955 5400 4005
rect 5360 3925 5365 3955
rect 5395 3925 5400 3955
rect 5360 3875 5400 3925
rect 5360 3845 5365 3875
rect 5395 3845 5400 3875
rect 5360 3790 5400 3845
rect 5360 3770 5370 3790
rect 5390 3770 5400 3790
rect 5360 3715 5400 3770
rect 5360 3685 5365 3715
rect 5395 3685 5400 3715
rect 5360 3635 5400 3685
rect 5360 3605 5365 3635
rect 5395 3605 5400 3635
rect 5360 3550 5400 3605
rect 5360 3530 5370 3550
rect 5390 3530 5400 3550
rect 5360 3475 5400 3530
rect 5360 3445 5365 3475
rect 5395 3445 5400 3475
rect 5360 3395 5400 3445
rect 5360 3365 5365 3395
rect 5395 3365 5400 3395
rect 5360 3310 5400 3365
rect 5360 3290 5370 3310
rect 5390 3290 5400 3310
rect 5360 3235 5400 3290
rect 5360 3205 5365 3235
rect 5395 3205 5400 3235
rect 5360 3155 5400 3205
rect 5360 3125 5365 3155
rect 5395 3125 5400 3155
rect 5360 3075 5400 3125
rect 5360 3045 5365 3075
rect 5395 3045 5400 3075
rect 5360 2995 5400 3045
rect 5360 2965 5365 2995
rect 5395 2965 5400 2995
rect 5360 2915 5400 2965
rect 5360 2885 5365 2915
rect 5395 2885 5400 2915
rect 5360 2835 5400 2885
rect 5360 2805 5365 2835
rect 5395 2805 5400 2835
rect 5360 2755 5400 2805
rect 5360 2725 5365 2755
rect 5395 2725 5400 2755
rect 5360 2675 5400 2725
rect 5360 2645 5365 2675
rect 5395 2645 5400 2675
rect 5360 2595 5400 2645
rect 5360 2565 5365 2595
rect 5395 2565 5400 2595
rect 5360 2515 5400 2565
rect 5360 2485 5365 2515
rect 5395 2485 5400 2515
rect 5360 2435 5400 2485
rect 5360 2405 5365 2435
rect 5395 2405 5400 2435
rect 5360 2355 5400 2405
rect 5360 2325 5365 2355
rect 5395 2325 5400 2355
rect 5360 2275 5400 2325
rect 5360 2245 5365 2275
rect 5395 2245 5400 2275
rect 5360 2195 5400 2245
rect 5360 2165 5365 2195
rect 5395 2165 5400 2195
rect 5360 2115 5400 2165
rect 5360 2085 5365 2115
rect 5395 2085 5400 2115
rect 5360 2035 5400 2085
rect 5360 2005 5365 2035
rect 5395 2005 5400 2035
rect 5360 1955 5400 2005
rect 5360 1925 5365 1955
rect 5395 1925 5400 1955
rect 5360 1870 5400 1925
rect 5360 1850 5370 1870
rect 5390 1850 5400 1870
rect 5360 1790 5400 1850
rect 5360 1770 5370 1790
rect 5390 1770 5400 1790
rect 5360 1715 5400 1770
rect 5360 1685 5365 1715
rect 5395 1685 5400 1715
rect 5360 1635 5400 1685
rect 5360 1605 5365 1635
rect 5395 1605 5400 1635
rect 5360 1555 5400 1605
rect 5360 1525 5365 1555
rect 5395 1525 5400 1555
rect 5360 1475 5400 1525
rect 5360 1445 5365 1475
rect 5395 1445 5400 1475
rect 5360 1395 5400 1445
rect 5360 1365 5365 1395
rect 5395 1365 5400 1395
rect 5360 1315 5400 1365
rect 5360 1285 5365 1315
rect 5395 1285 5400 1315
rect 5360 1235 5400 1285
rect 5360 1205 5365 1235
rect 5395 1205 5400 1235
rect 5360 1155 5400 1205
rect 5360 1125 5365 1155
rect 5395 1125 5400 1155
rect 5360 1075 5400 1125
rect 5360 1045 5365 1075
rect 5395 1045 5400 1075
rect 5360 995 5400 1045
rect 5360 965 5365 995
rect 5395 965 5400 995
rect 5360 910 5400 965
rect 5360 890 5370 910
rect 5390 890 5400 910
rect 5360 835 5400 890
rect 5360 805 5365 835
rect 5395 805 5400 835
rect 5360 755 5400 805
rect 5360 725 5365 755
rect 5395 725 5400 755
rect 5360 675 5400 725
rect 5360 645 5365 675
rect 5395 645 5400 675
rect 5360 595 5400 645
rect 5360 565 5365 595
rect 5395 565 5400 595
rect 5360 515 5400 565
rect 5360 485 5365 515
rect 5395 485 5400 515
rect 5360 430 5400 485
rect 5360 410 5370 430
rect 5390 410 5400 430
rect 5360 350 5400 410
rect 5360 330 5370 350
rect 5390 330 5400 350
rect 5360 275 5400 330
rect 5360 245 5365 275
rect 5395 245 5400 275
rect 5360 195 5400 245
rect 5360 165 5365 195
rect 5395 165 5400 195
rect 5360 115 5400 165
rect 5360 85 5365 115
rect 5395 85 5400 115
rect 5360 35 5400 85
rect 5360 5 5365 35
rect 5395 5 5400 35
rect 5360 0 5400 5
rect 5440 15710 5480 15720
rect 5440 15690 5450 15710
rect 5470 15690 5480 15710
rect 5440 15630 5480 15690
rect 5440 15610 5450 15630
rect 5470 15610 5480 15630
rect 5440 15550 5480 15610
rect 5440 15530 5450 15550
rect 5470 15530 5480 15550
rect 5440 15470 5480 15530
rect 5440 15450 5450 15470
rect 5470 15450 5480 15470
rect 5440 15390 5480 15450
rect 5440 15370 5450 15390
rect 5470 15370 5480 15390
rect 5440 15310 5480 15370
rect 5440 15290 5450 15310
rect 5470 15290 5480 15310
rect 5440 15230 5480 15290
rect 5440 15210 5450 15230
rect 5470 15210 5480 15230
rect 5440 15150 5480 15210
rect 5440 15130 5450 15150
rect 5470 15130 5480 15150
rect 5440 15070 5480 15130
rect 5440 15050 5450 15070
rect 5470 15050 5480 15070
rect 5440 14990 5480 15050
rect 5440 14970 5450 14990
rect 5470 14970 5480 14990
rect 5440 14910 5480 14970
rect 5440 14890 5450 14910
rect 5470 14890 5480 14910
rect 5440 14830 5480 14890
rect 5440 14810 5450 14830
rect 5470 14810 5480 14830
rect 5440 14750 5480 14810
rect 5440 14730 5450 14750
rect 5470 14730 5480 14750
rect 5440 14670 5480 14730
rect 5440 14650 5450 14670
rect 5470 14650 5480 14670
rect 5440 14590 5480 14650
rect 5440 14570 5450 14590
rect 5470 14570 5480 14590
rect 5440 14510 5480 14570
rect 5440 14490 5450 14510
rect 5470 14490 5480 14510
rect 5440 14430 5480 14490
rect 5440 14410 5450 14430
rect 5470 14410 5480 14430
rect 5440 14350 5480 14410
rect 5440 14330 5450 14350
rect 5470 14330 5480 14350
rect 5440 14270 5480 14330
rect 5440 14250 5450 14270
rect 5470 14250 5480 14270
rect 5440 14190 5480 14250
rect 5440 14170 5450 14190
rect 5470 14170 5480 14190
rect 5440 14110 5480 14170
rect 5440 14090 5450 14110
rect 5470 14090 5480 14110
rect 5440 14030 5480 14090
rect 5440 14010 5450 14030
rect 5470 14010 5480 14030
rect 5440 13950 5480 14010
rect 5440 13930 5450 13950
rect 5470 13930 5480 13950
rect 5440 13870 5480 13930
rect 5440 13850 5450 13870
rect 5470 13850 5480 13870
rect 5440 13790 5480 13850
rect 5440 13770 5450 13790
rect 5470 13770 5480 13790
rect 5440 13710 5480 13770
rect 5440 13690 5450 13710
rect 5470 13690 5480 13710
rect 5440 13630 5480 13690
rect 5440 13610 5450 13630
rect 5470 13610 5480 13630
rect 5440 13550 5480 13610
rect 5440 13530 5450 13550
rect 5470 13530 5480 13550
rect 5440 13470 5480 13530
rect 5440 13450 5450 13470
rect 5470 13450 5480 13470
rect 5440 13390 5480 13450
rect 5440 13370 5450 13390
rect 5470 13370 5480 13390
rect 5440 13310 5480 13370
rect 5440 13290 5450 13310
rect 5470 13290 5480 13310
rect 5440 13230 5480 13290
rect 5440 13210 5450 13230
rect 5470 13210 5480 13230
rect 5440 13150 5480 13210
rect 5440 13130 5450 13150
rect 5470 13130 5480 13150
rect 5440 13070 5480 13130
rect 5440 13050 5450 13070
rect 5470 13050 5480 13070
rect 5440 12990 5480 13050
rect 5440 12970 5450 12990
rect 5470 12970 5480 12990
rect 5440 12910 5480 12970
rect 5440 12890 5450 12910
rect 5470 12890 5480 12910
rect 5440 12830 5480 12890
rect 5440 12810 5450 12830
rect 5470 12810 5480 12830
rect 5440 12750 5480 12810
rect 5440 12730 5450 12750
rect 5470 12730 5480 12750
rect 5440 12670 5480 12730
rect 5440 12650 5450 12670
rect 5470 12650 5480 12670
rect 5440 12590 5480 12650
rect 5440 12570 5450 12590
rect 5470 12570 5480 12590
rect 5440 12510 5480 12570
rect 5440 12490 5450 12510
rect 5470 12490 5480 12510
rect 5440 12430 5480 12490
rect 5440 12410 5450 12430
rect 5470 12410 5480 12430
rect 5440 12350 5480 12410
rect 5440 12330 5450 12350
rect 5470 12330 5480 12350
rect 5440 12270 5480 12330
rect 5440 12250 5450 12270
rect 5470 12250 5480 12270
rect 5440 12190 5480 12250
rect 5440 12170 5450 12190
rect 5470 12170 5480 12190
rect 5440 12110 5480 12170
rect 5440 12090 5450 12110
rect 5470 12090 5480 12110
rect 5440 12030 5480 12090
rect 5440 12010 5450 12030
rect 5470 12010 5480 12030
rect 5440 11950 5480 12010
rect 5440 11930 5450 11950
rect 5470 11930 5480 11950
rect 5440 11870 5480 11930
rect 5440 11850 5450 11870
rect 5470 11850 5480 11870
rect 5440 11790 5480 11850
rect 5440 11770 5450 11790
rect 5470 11770 5480 11790
rect 5440 11710 5480 11770
rect 5440 11690 5450 11710
rect 5470 11690 5480 11710
rect 5440 11630 5480 11690
rect 5440 11610 5450 11630
rect 5470 11610 5480 11630
rect 5440 11550 5480 11610
rect 5440 11530 5450 11550
rect 5470 11530 5480 11550
rect 5440 11470 5480 11530
rect 5440 11450 5450 11470
rect 5470 11450 5480 11470
rect 5440 11390 5480 11450
rect 5440 11370 5450 11390
rect 5470 11370 5480 11390
rect 5440 11310 5480 11370
rect 5440 11290 5450 11310
rect 5470 11290 5480 11310
rect 5440 11230 5480 11290
rect 5440 11210 5450 11230
rect 5470 11210 5480 11230
rect 5440 11150 5480 11210
rect 5440 11130 5450 11150
rect 5470 11130 5480 11150
rect 5440 11070 5480 11130
rect 5440 11050 5450 11070
rect 5470 11050 5480 11070
rect 5440 10990 5480 11050
rect 5440 10970 5450 10990
rect 5470 10970 5480 10990
rect 5440 10910 5480 10970
rect 5440 10890 5450 10910
rect 5470 10890 5480 10910
rect 5440 10830 5480 10890
rect 5440 10810 5450 10830
rect 5470 10810 5480 10830
rect 5440 10750 5480 10810
rect 5440 10730 5450 10750
rect 5470 10730 5480 10750
rect 5440 10670 5480 10730
rect 5440 10650 5450 10670
rect 5470 10650 5480 10670
rect 5440 10590 5480 10650
rect 5440 10570 5450 10590
rect 5470 10570 5480 10590
rect 5440 10510 5480 10570
rect 5440 10490 5450 10510
rect 5470 10490 5480 10510
rect 5440 10430 5480 10490
rect 5440 10410 5450 10430
rect 5470 10410 5480 10430
rect 5440 10350 5480 10410
rect 5440 10330 5450 10350
rect 5470 10330 5480 10350
rect 5440 10270 5480 10330
rect 5440 10250 5450 10270
rect 5470 10250 5480 10270
rect 5440 10190 5480 10250
rect 5440 10170 5450 10190
rect 5470 10170 5480 10190
rect 5440 10110 5480 10170
rect 5440 10090 5450 10110
rect 5470 10090 5480 10110
rect 5440 10030 5480 10090
rect 5440 10010 5450 10030
rect 5470 10010 5480 10030
rect 5440 9950 5480 10010
rect 5440 9930 5450 9950
rect 5470 9930 5480 9950
rect 5440 9870 5480 9930
rect 5440 9850 5450 9870
rect 5470 9850 5480 9870
rect 5440 9790 5480 9850
rect 5440 9770 5450 9790
rect 5470 9770 5480 9790
rect 5440 9710 5480 9770
rect 5440 9690 5450 9710
rect 5470 9690 5480 9710
rect 5440 9630 5480 9690
rect 5440 9610 5450 9630
rect 5470 9610 5480 9630
rect 5440 9550 5480 9610
rect 5440 9530 5450 9550
rect 5470 9530 5480 9550
rect 5440 9470 5480 9530
rect 5440 9450 5450 9470
rect 5470 9450 5480 9470
rect 5440 9390 5480 9450
rect 5440 9370 5450 9390
rect 5470 9370 5480 9390
rect 5440 9310 5480 9370
rect 5440 9290 5450 9310
rect 5470 9290 5480 9310
rect 5440 9230 5480 9290
rect 5440 9210 5450 9230
rect 5470 9210 5480 9230
rect 5440 9150 5480 9210
rect 5440 9130 5450 9150
rect 5470 9130 5480 9150
rect 5440 9070 5480 9130
rect 5440 9050 5450 9070
rect 5470 9050 5480 9070
rect 5440 8990 5480 9050
rect 5440 8970 5450 8990
rect 5470 8970 5480 8990
rect 5440 8910 5480 8970
rect 5440 8890 5450 8910
rect 5470 8890 5480 8910
rect 5440 8830 5480 8890
rect 5440 8810 5450 8830
rect 5470 8810 5480 8830
rect 5440 8750 5480 8810
rect 5440 8730 5450 8750
rect 5470 8730 5480 8750
rect 5440 8670 5480 8730
rect 5440 8650 5450 8670
rect 5470 8650 5480 8670
rect 5440 8590 5480 8650
rect 5440 8570 5450 8590
rect 5470 8570 5480 8590
rect 5440 8510 5480 8570
rect 5440 8490 5450 8510
rect 5470 8490 5480 8510
rect 5440 8430 5480 8490
rect 5440 8410 5450 8430
rect 5470 8410 5480 8430
rect 5440 8350 5480 8410
rect 5440 8330 5450 8350
rect 5470 8330 5480 8350
rect 5440 8270 5480 8330
rect 5440 8250 5450 8270
rect 5470 8250 5480 8270
rect 5440 8190 5480 8250
rect 5440 8170 5450 8190
rect 5470 8170 5480 8190
rect 5440 8110 5480 8170
rect 5440 8090 5450 8110
rect 5470 8090 5480 8110
rect 5440 8030 5480 8090
rect 5440 8010 5450 8030
rect 5470 8010 5480 8030
rect 5440 7950 5480 8010
rect 5440 7930 5450 7950
rect 5470 7930 5480 7950
rect 5440 7870 5480 7930
rect 5440 7850 5450 7870
rect 5470 7850 5480 7870
rect 5440 7790 5480 7850
rect 5440 7770 5450 7790
rect 5470 7770 5480 7790
rect 5440 7710 5480 7770
rect 5440 7690 5450 7710
rect 5470 7690 5480 7710
rect 5440 7630 5480 7690
rect 5440 7610 5450 7630
rect 5470 7610 5480 7630
rect 5440 7550 5480 7610
rect 5440 7530 5450 7550
rect 5470 7530 5480 7550
rect 5440 7470 5480 7530
rect 5440 7450 5450 7470
rect 5470 7450 5480 7470
rect 5440 7390 5480 7450
rect 5440 7370 5450 7390
rect 5470 7370 5480 7390
rect 5440 7310 5480 7370
rect 5440 7290 5450 7310
rect 5470 7290 5480 7310
rect 5440 7230 5480 7290
rect 5440 7210 5450 7230
rect 5470 7210 5480 7230
rect 5440 7150 5480 7210
rect 5440 7130 5450 7150
rect 5470 7130 5480 7150
rect 5440 7070 5480 7130
rect 5440 7050 5450 7070
rect 5470 7050 5480 7070
rect 5440 6990 5480 7050
rect 5440 6970 5450 6990
rect 5470 6970 5480 6990
rect 5440 6910 5480 6970
rect 5440 6890 5450 6910
rect 5470 6890 5480 6910
rect 5440 6830 5480 6890
rect 5440 6810 5450 6830
rect 5470 6810 5480 6830
rect 5440 6750 5480 6810
rect 5440 6730 5450 6750
rect 5470 6730 5480 6750
rect 5440 6670 5480 6730
rect 5440 6650 5450 6670
rect 5470 6650 5480 6670
rect 5440 6590 5480 6650
rect 5440 6570 5450 6590
rect 5470 6570 5480 6590
rect 5440 6510 5480 6570
rect 5440 6490 5450 6510
rect 5470 6490 5480 6510
rect 5440 6430 5480 6490
rect 5440 6410 5450 6430
rect 5470 6410 5480 6430
rect 5440 6350 5480 6410
rect 5440 6330 5450 6350
rect 5470 6330 5480 6350
rect 5440 6270 5480 6330
rect 5440 6250 5450 6270
rect 5470 6250 5480 6270
rect 5440 6190 5480 6250
rect 5440 6170 5450 6190
rect 5470 6170 5480 6190
rect 5440 6110 5480 6170
rect 5440 6090 5450 6110
rect 5470 6090 5480 6110
rect 5440 6030 5480 6090
rect 5440 6010 5450 6030
rect 5470 6010 5480 6030
rect 5440 5950 5480 6010
rect 5440 5930 5450 5950
rect 5470 5930 5480 5950
rect 5440 5870 5480 5930
rect 5440 5850 5450 5870
rect 5470 5850 5480 5870
rect 5440 5790 5480 5850
rect 5440 5770 5450 5790
rect 5470 5770 5480 5790
rect 5440 5710 5480 5770
rect 5440 5690 5450 5710
rect 5470 5690 5480 5710
rect 5440 5630 5480 5690
rect 5440 5610 5450 5630
rect 5470 5610 5480 5630
rect 5440 5550 5480 5610
rect 5440 5530 5450 5550
rect 5470 5530 5480 5550
rect 5440 5470 5480 5530
rect 5440 5450 5450 5470
rect 5470 5450 5480 5470
rect 5440 5390 5480 5450
rect 5440 5370 5450 5390
rect 5470 5370 5480 5390
rect 5440 5310 5480 5370
rect 5440 5290 5450 5310
rect 5470 5290 5480 5310
rect 5440 5230 5480 5290
rect 5440 5210 5450 5230
rect 5470 5210 5480 5230
rect 5440 5150 5480 5210
rect 5440 5130 5450 5150
rect 5470 5130 5480 5150
rect 5440 5070 5480 5130
rect 5440 5050 5450 5070
rect 5470 5050 5480 5070
rect 5440 4990 5480 5050
rect 5440 4970 5450 4990
rect 5470 4970 5480 4990
rect 5440 4910 5480 4970
rect 5440 4890 5450 4910
rect 5470 4890 5480 4910
rect 5440 4830 5480 4890
rect 5440 4810 5450 4830
rect 5470 4810 5480 4830
rect 5440 4750 5480 4810
rect 5440 4730 5450 4750
rect 5470 4730 5480 4750
rect 5440 4670 5480 4730
rect 5440 4650 5450 4670
rect 5470 4650 5480 4670
rect 5440 4590 5480 4650
rect 5440 4570 5450 4590
rect 5470 4570 5480 4590
rect 5440 4510 5480 4570
rect 5440 4490 5450 4510
rect 5470 4490 5480 4510
rect 5440 4430 5480 4490
rect 5440 4410 5450 4430
rect 5470 4410 5480 4430
rect 5440 4350 5480 4410
rect 5440 4330 5450 4350
rect 5470 4330 5480 4350
rect 5440 4270 5480 4330
rect 5440 4250 5450 4270
rect 5470 4250 5480 4270
rect 5440 4190 5480 4250
rect 5440 4170 5450 4190
rect 5470 4170 5480 4190
rect 5440 4110 5480 4170
rect 5440 4090 5450 4110
rect 5470 4090 5480 4110
rect 5440 4030 5480 4090
rect 5440 4010 5450 4030
rect 5470 4010 5480 4030
rect 5440 3950 5480 4010
rect 5440 3930 5450 3950
rect 5470 3930 5480 3950
rect 5440 3870 5480 3930
rect 5440 3850 5450 3870
rect 5470 3850 5480 3870
rect 5440 3790 5480 3850
rect 5440 3770 5450 3790
rect 5470 3770 5480 3790
rect 5440 3710 5480 3770
rect 5440 3690 5450 3710
rect 5470 3690 5480 3710
rect 5440 3630 5480 3690
rect 5440 3610 5450 3630
rect 5470 3610 5480 3630
rect 5440 3550 5480 3610
rect 5440 3530 5450 3550
rect 5470 3530 5480 3550
rect 5440 3470 5480 3530
rect 5440 3450 5450 3470
rect 5470 3450 5480 3470
rect 5440 3390 5480 3450
rect 5440 3370 5450 3390
rect 5470 3370 5480 3390
rect 5440 3310 5480 3370
rect 5440 3290 5450 3310
rect 5470 3290 5480 3310
rect 5440 3230 5480 3290
rect 5440 3210 5450 3230
rect 5470 3210 5480 3230
rect 5440 3150 5480 3210
rect 5440 3130 5450 3150
rect 5470 3130 5480 3150
rect 5440 3070 5480 3130
rect 5440 3050 5450 3070
rect 5470 3050 5480 3070
rect 5440 2990 5480 3050
rect 5440 2970 5450 2990
rect 5470 2970 5480 2990
rect 5440 2910 5480 2970
rect 5440 2890 5450 2910
rect 5470 2890 5480 2910
rect 5440 2830 5480 2890
rect 5440 2810 5450 2830
rect 5470 2810 5480 2830
rect 5440 2750 5480 2810
rect 5440 2730 5450 2750
rect 5470 2730 5480 2750
rect 5440 2670 5480 2730
rect 5440 2650 5450 2670
rect 5470 2650 5480 2670
rect 5440 2590 5480 2650
rect 5440 2570 5450 2590
rect 5470 2570 5480 2590
rect 5440 2510 5480 2570
rect 5440 2490 5450 2510
rect 5470 2490 5480 2510
rect 5440 2430 5480 2490
rect 5440 2410 5450 2430
rect 5470 2410 5480 2430
rect 5440 2350 5480 2410
rect 5440 2330 5450 2350
rect 5470 2330 5480 2350
rect 5440 2270 5480 2330
rect 5440 2250 5450 2270
rect 5470 2250 5480 2270
rect 5440 2190 5480 2250
rect 5440 2170 5450 2190
rect 5470 2170 5480 2190
rect 5440 2110 5480 2170
rect 5440 2090 5450 2110
rect 5470 2090 5480 2110
rect 5440 2030 5480 2090
rect 5440 2010 5450 2030
rect 5470 2010 5480 2030
rect 5440 1950 5480 2010
rect 5440 1930 5450 1950
rect 5470 1930 5480 1950
rect 5440 1870 5480 1930
rect 5440 1850 5450 1870
rect 5470 1850 5480 1870
rect 5440 1790 5480 1850
rect 5440 1770 5450 1790
rect 5470 1770 5480 1790
rect 5440 1710 5480 1770
rect 5440 1690 5450 1710
rect 5470 1690 5480 1710
rect 5440 1630 5480 1690
rect 5440 1610 5450 1630
rect 5470 1610 5480 1630
rect 5440 1550 5480 1610
rect 5440 1530 5450 1550
rect 5470 1530 5480 1550
rect 5440 1470 5480 1530
rect 5440 1450 5450 1470
rect 5470 1450 5480 1470
rect 5440 1390 5480 1450
rect 5440 1370 5450 1390
rect 5470 1370 5480 1390
rect 5440 1310 5480 1370
rect 5440 1290 5450 1310
rect 5470 1290 5480 1310
rect 5440 1230 5480 1290
rect 5440 1210 5450 1230
rect 5470 1210 5480 1230
rect 5440 1150 5480 1210
rect 5440 1130 5450 1150
rect 5470 1130 5480 1150
rect 5440 1070 5480 1130
rect 5440 1050 5450 1070
rect 5470 1050 5480 1070
rect 5440 990 5480 1050
rect 5440 970 5450 990
rect 5470 970 5480 990
rect 5440 910 5480 970
rect 5440 890 5450 910
rect 5470 890 5480 910
rect 5440 830 5480 890
rect 5440 810 5450 830
rect 5470 810 5480 830
rect 5440 750 5480 810
rect 5440 730 5450 750
rect 5470 730 5480 750
rect 5440 670 5480 730
rect 5440 650 5450 670
rect 5470 650 5480 670
rect 5440 590 5480 650
rect 5440 570 5450 590
rect 5470 570 5480 590
rect 5440 510 5480 570
rect 5440 490 5450 510
rect 5470 490 5480 510
rect 5440 430 5480 490
rect 5440 410 5450 430
rect 5470 410 5480 430
rect 5440 350 5480 410
rect 5440 330 5450 350
rect 5470 330 5480 350
rect 5440 270 5480 330
rect 5440 250 5450 270
rect 5470 250 5480 270
rect 5440 190 5480 250
rect 5440 170 5450 190
rect 5470 170 5480 190
rect 5440 110 5480 170
rect 5440 90 5450 110
rect 5470 90 5480 110
rect 5440 30 5480 90
rect 5440 10 5450 30
rect 5470 10 5480 30
rect 5440 0 5480 10
rect 5520 15715 5560 15720
rect 5520 15685 5525 15715
rect 5555 15685 5560 15715
rect 5520 15635 5560 15685
rect 5520 15605 5525 15635
rect 5555 15605 5560 15635
rect 5520 15555 5560 15605
rect 5520 15525 5525 15555
rect 5555 15525 5560 15555
rect 5520 15475 5560 15525
rect 5520 15445 5525 15475
rect 5555 15445 5560 15475
rect 5520 15395 5560 15445
rect 5520 15365 5525 15395
rect 5555 15365 5560 15395
rect 5520 15315 5560 15365
rect 5520 15285 5525 15315
rect 5555 15285 5560 15315
rect 5520 15235 5560 15285
rect 5520 15205 5525 15235
rect 5555 15205 5560 15235
rect 5520 15155 5560 15205
rect 5520 15125 5525 15155
rect 5555 15125 5560 15155
rect 5520 15070 5560 15125
rect 5520 15050 5530 15070
rect 5550 15050 5560 15070
rect 5520 14995 5560 15050
rect 5520 14965 5525 14995
rect 5555 14965 5560 14995
rect 5520 14915 5560 14965
rect 5520 14885 5525 14915
rect 5555 14885 5560 14915
rect 5520 14835 5560 14885
rect 5520 14805 5525 14835
rect 5555 14805 5560 14835
rect 5520 14755 5560 14805
rect 5520 14725 5525 14755
rect 5555 14725 5560 14755
rect 5520 14675 5560 14725
rect 5520 14645 5525 14675
rect 5555 14645 5560 14675
rect 5520 14595 5560 14645
rect 5520 14565 5525 14595
rect 5555 14565 5560 14595
rect 5520 14515 5560 14565
rect 5520 14485 5525 14515
rect 5555 14485 5560 14515
rect 5520 14435 5560 14485
rect 5520 14405 5525 14435
rect 5555 14405 5560 14435
rect 5520 14350 5560 14405
rect 5520 14330 5530 14350
rect 5550 14330 5560 14350
rect 5520 14270 5560 14330
rect 5520 14250 5530 14270
rect 5550 14250 5560 14270
rect 5520 14190 5560 14250
rect 5520 14170 5530 14190
rect 5550 14170 5560 14190
rect 5520 14110 5560 14170
rect 5520 14090 5530 14110
rect 5550 14090 5560 14110
rect 5520 14035 5560 14090
rect 5520 14005 5525 14035
rect 5555 14005 5560 14035
rect 5520 13955 5560 14005
rect 5520 13925 5525 13955
rect 5555 13925 5560 13955
rect 5520 13875 5560 13925
rect 5520 13845 5525 13875
rect 5555 13845 5560 13875
rect 5520 13795 5560 13845
rect 5520 13765 5525 13795
rect 5555 13765 5560 13795
rect 5520 13715 5560 13765
rect 5520 13685 5525 13715
rect 5555 13685 5560 13715
rect 5520 13635 5560 13685
rect 5520 13605 5525 13635
rect 5555 13605 5560 13635
rect 5520 13555 5560 13605
rect 5520 13525 5525 13555
rect 5555 13525 5560 13555
rect 5520 13475 5560 13525
rect 5520 13445 5525 13475
rect 5555 13445 5560 13475
rect 5520 13390 5560 13445
rect 5520 13370 5530 13390
rect 5550 13370 5560 13390
rect 5520 13310 5560 13370
rect 5520 13290 5530 13310
rect 5550 13290 5560 13310
rect 5520 13230 5560 13290
rect 5520 13210 5530 13230
rect 5550 13210 5560 13230
rect 5520 13150 5560 13210
rect 5520 13130 5530 13150
rect 5550 13130 5560 13150
rect 5520 13075 5560 13130
rect 5520 13045 5525 13075
rect 5555 13045 5560 13075
rect 5520 12995 5560 13045
rect 5520 12965 5525 12995
rect 5555 12965 5560 12995
rect 5520 12915 5560 12965
rect 5520 12885 5525 12915
rect 5555 12885 5560 12915
rect 5520 12835 5560 12885
rect 5520 12805 5525 12835
rect 5555 12805 5560 12835
rect 5520 12755 5560 12805
rect 5520 12725 5525 12755
rect 5555 12725 5560 12755
rect 5520 12675 5560 12725
rect 5520 12645 5525 12675
rect 5555 12645 5560 12675
rect 5520 12595 5560 12645
rect 5520 12565 5525 12595
rect 5555 12565 5560 12595
rect 5520 12515 5560 12565
rect 5520 12485 5525 12515
rect 5555 12485 5560 12515
rect 5520 12430 5560 12485
rect 5520 12410 5530 12430
rect 5550 12410 5560 12430
rect 5520 12355 5560 12410
rect 5520 12325 5525 12355
rect 5555 12325 5560 12355
rect 5520 12275 5560 12325
rect 5520 12245 5525 12275
rect 5555 12245 5560 12275
rect 5520 12195 5560 12245
rect 5520 12165 5525 12195
rect 5555 12165 5560 12195
rect 5520 12115 5560 12165
rect 5520 12085 5525 12115
rect 5555 12085 5560 12115
rect 5520 12035 5560 12085
rect 5520 12005 5525 12035
rect 5555 12005 5560 12035
rect 5520 11955 5560 12005
rect 5520 11925 5525 11955
rect 5555 11925 5560 11955
rect 5520 11875 5560 11925
rect 5520 11845 5525 11875
rect 5555 11845 5560 11875
rect 5520 11795 5560 11845
rect 5520 11765 5525 11795
rect 5555 11765 5560 11795
rect 5520 11715 5560 11765
rect 5520 11685 5525 11715
rect 5555 11685 5560 11715
rect 5520 11635 5560 11685
rect 5520 11605 5525 11635
rect 5555 11605 5560 11635
rect 5520 11555 5560 11605
rect 5520 11525 5525 11555
rect 5555 11525 5560 11555
rect 5520 11475 5560 11525
rect 5520 11445 5525 11475
rect 5555 11445 5560 11475
rect 5520 11395 5560 11445
rect 5520 11365 5525 11395
rect 5555 11365 5560 11395
rect 5520 11315 5560 11365
rect 5520 11285 5525 11315
rect 5555 11285 5560 11315
rect 5520 11235 5560 11285
rect 5520 11205 5525 11235
rect 5555 11205 5560 11235
rect 5520 11155 5560 11205
rect 5520 11125 5525 11155
rect 5555 11125 5560 11155
rect 5520 11075 5560 11125
rect 5520 11045 5525 11075
rect 5555 11045 5560 11075
rect 5520 10990 5560 11045
rect 5520 10970 5530 10990
rect 5550 10970 5560 10990
rect 5520 10915 5560 10970
rect 5520 10885 5525 10915
rect 5555 10885 5560 10915
rect 5520 10835 5560 10885
rect 5520 10805 5525 10835
rect 5555 10805 5560 10835
rect 5520 10755 5560 10805
rect 5520 10725 5525 10755
rect 5555 10725 5560 10755
rect 5520 10675 5560 10725
rect 5520 10645 5525 10675
rect 5555 10645 5560 10675
rect 5520 10595 5560 10645
rect 5520 10565 5525 10595
rect 5555 10565 5560 10595
rect 5520 10515 5560 10565
rect 5520 10485 5525 10515
rect 5555 10485 5560 10515
rect 5520 10435 5560 10485
rect 5520 10405 5525 10435
rect 5555 10405 5560 10435
rect 5520 10355 5560 10405
rect 5520 10325 5525 10355
rect 5555 10325 5560 10355
rect 5520 10270 5560 10325
rect 5520 10250 5530 10270
rect 5550 10250 5560 10270
rect 5520 10190 5560 10250
rect 5520 10170 5530 10190
rect 5550 10170 5560 10190
rect 5520 10110 5560 10170
rect 5520 10090 5530 10110
rect 5550 10090 5560 10110
rect 5520 10030 5560 10090
rect 5520 10010 5530 10030
rect 5550 10010 5560 10030
rect 5520 9955 5560 10010
rect 5520 9925 5525 9955
rect 5555 9925 5560 9955
rect 5520 9875 5560 9925
rect 5520 9845 5525 9875
rect 5555 9845 5560 9875
rect 5520 9795 5560 9845
rect 5520 9765 5525 9795
rect 5555 9765 5560 9795
rect 5520 9715 5560 9765
rect 5520 9685 5525 9715
rect 5555 9685 5560 9715
rect 5520 9635 5560 9685
rect 5520 9605 5525 9635
rect 5555 9605 5560 9635
rect 5520 9555 5560 9605
rect 5520 9525 5525 9555
rect 5555 9525 5560 9555
rect 5520 9475 5560 9525
rect 5520 9445 5525 9475
rect 5555 9445 5560 9475
rect 5520 9395 5560 9445
rect 5520 9365 5525 9395
rect 5555 9365 5560 9395
rect 5520 9310 5560 9365
rect 5520 9290 5530 9310
rect 5550 9290 5560 9310
rect 5520 9230 5560 9290
rect 5520 9210 5530 9230
rect 5550 9210 5560 9230
rect 5520 9150 5560 9210
rect 5520 9130 5530 9150
rect 5550 9130 5560 9150
rect 5520 9070 5560 9130
rect 5520 9050 5530 9070
rect 5550 9050 5560 9070
rect 5520 8995 5560 9050
rect 5520 8965 5525 8995
rect 5555 8965 5560 8995
rect 5520 8915 5560 8965
rect 5520 8885 5525 8915
rect 5555 8885 5560 8915
rect 5520 8835 5560 8885
rect 5520 8805 5525 8835
rect 5555 8805 5560 8835
rect 5520 8755 5560 8805
rect 5520 8725 5525 8755
rect 5555 8725 5560 8755
rect 5520 8675 5560 8725
rect 5520 8645 5525 8675
rect 5555 8645 5560 8675
rect 5520 8595 5560 8645
rect 5520 8565 5525 8595
rect 5555 8565 5560 8595
rect 5520 8515 5560 8565
rect 5520 8485 5525 8515
rect 5555 8485 5560 8515
rect 5520 8435 5560 8485
rect 5520 8405 5525 8435
rect 5555 8405 5560 8435
rect 5520 8350 5560 8405
rect 5520 8330 5530 8350
rect 5550 8330 5560 8350
rect 5520 8275 5560 8330
rect 5520 8245 5525 8275
rect 5555 8245 5560 8275
rect 5520 8195 5560 8245
rect 5520 8165 5525 8195
rect 5555 8165 5560 8195
rect 5520 8115 5560 8165
rect 5520 8085 5525 8115
rect 5555 8085 5560 8115
rect 5520 8035 5560 8085
rect 5520 8005 5525 8035
rect 5555 8005 5560 8035
rect 5520 7955 5560 8005
rect 5520 7925 5525 7955
rect 5555 7925 5560 7955
rect 5520 7875 5560 7925
rect 5520 7845 5525 7875
rect 5555 7845 5560 7875
rect 5520 7795 5560 7845
rect 5520 7765 5525 7795
rect 5555 7765 5560 7795
rect 5520 7715 5560 7765
rect 5520 7685 5525 7715
rect 5555 7685 5560 7715
rect 5520 7635 5560 7685
rect 5520 7605 5525 7635
rect 5555 7605 5560 7635
rect 5520 7555 5560 7605
rect 5520 7525 5525 7555
rect 5555 7525 5560 7555
rect 5520 7475 5560 7525
rect 5520 7445 5525 7475
rect 5555 7445 5560 7475
rect 5520 7395 5560 7445
rect 5520 7365 5525 7395
rect 5555 7365 5560 7395
rect 5520 7315 5560 7365
rect 5520 7285 5525 7315
rect 5555 7285 5560 7315
rect 5520 7235 5560 7285
rect 5520 7205 5525 7235
rect 5555 7205 5560 7235
rect 5520 7155 5560 7205
rect 5520 7125 5525 7155
rect 5555 7125 5560 7155
rect 5520 7075 5560 7125
rect 5520 7045 5525 7075
rect 5555 7045 5560 7075
rect 5520 6995 5560 7045
rect 5520 6965 5525 6995
rect 5555 6965 5560 6995
rect 5520 6910 5560 6965
rect 5520 6890 5530 6910
rect 5550 6890 5560 6910
rect 5520 6835 5560 6890
rect 5520 6805 5525 6835
rect 5555 6805 5560 6835
rect 5520 6755 5560 6805
rect 5520 6725 5525 6755
rect 5555 6725 5560 6755
rect 5520 6675 5560 6725
rect 5520 6645 5525 6675
rect 5555 6645 5560 6675
rect 5520 6595 5560 6645
rect 5520 6565 5525 6595
rect 5555 6565 5560 6595
rect 5520 6515 5560 6565
rect 5520 6485 5525 6515
rect 5555 6485 5560 6515
rect 5520 6435 5560 6485
rect 5520 6405 5525 6435
rect 5555 6405 5560 6435
rect 5520 6355 5560 6405
rect 5520 6325 5525 6355
rect 5555 6325 5560 6355
rect 5520 6275 5560 6325
rect 5520 6245 5525 6275
rect 5555 6245 5560 6275
rect 5520 6190 5560 6245
rect 5520 6170 5530 6190
rect 5550 6170 5560 6190
rect 5520 6110 5560 6170
rect 5520 6090 5530 6110
rect 5550 6090 5560 6110
rect 5520 6030 5560 6090
rect 5520 6010 5530 6030
rect 5550 6010 5560 6030
rect 5520 5950 5560 6010
rect 5520 5930 5530 5950
rect 5550 5930 5560 5950
rect 5520 5875 5560 5930
rect 5520 5845 5525 5875
rect 5555 5845 5560 5875
rect 5520 5795 5560 5845
rect 5520 5765 5525 5795
rect 5555 5765 5560 5795
rect 5520 5715 5560 5765
rect 5520 5685 5525 5715
rect 5555 5685 5560 5715
rect 5520 5635 5560 5685
rect 5520 5605 5525 5635
rect 5555 5605 5560 5635
rect 5520 5555 5560 5605
rect 5520 5525 5525 5555
rect 5555 5525 5560 5555
rect 5520 5475 5560 5525
rect 5520 5445 5525 5475
rect 5555 5445 5560 5475
rect 5520 5395 5560 5445
rect 5520 5365 5525 5395
rect 5555 5365 5560 5395
rect 5520 5315 5560 5365
rect 5520 5285 5525 5315
rect 5555 5285 5560 5315
rect 5520 5235 5560 5285
rect 5520 5205 5525 5235
rect 5555 5205 5560 5235
rect 5520 5155 5560 5205
rect 5520 5125 5525 5155
rect 5555 5125 5560 5155
rect 5520 5075 5560 5125
rect 5520 5045 5525 5075
rect 5555 5045 5560 5075
rect 5520 4995 5560 5045
rect 5520 4965 5525 4995
rect 5555 4965 5560 4995
rect 5520 4915 5560 4965
rect 5520 4885 5525 4915
rect 5555 4885 5560 4915
rect 5520 4830 5560 4885
rect 5520 4810 5530 4830
rect 5550 4810 5560 4830
rect 5520 4755 5560 4810
rect 5520 4725 5525 4755
rect 5555 4725 5560 4755
rect 5520 4675 5560 4725
rect 5520 4645 5525 4675
rect 5555 4645 5560 4675
rect 5520 4590 5560 4645
rect 5520 4570 5530 4590
rect 5550 4570 5560 4590
rect 5520 4515 5560 4570
rect 5520 4485 5525 4515
rect 5555 4485 5560 4515
rect 5520 4435 5560 4485
rect 5520 4405 5525 4435
rect 5555 4405 5560 4435
rect 5520 4355 5560 4405
rect 5520 4325 5525 4355
rect 5555 4325 5560 4355
rect 5520 4275 5560 4325
rect 5520 4245 5525 4275
rect 5555 4245 5560 4275
rect 5520 4195 5560 4245
rect 5520 4165 5525 4195
rect 5555 4165 5560 4195
rect 5520 4115 5560 4165
rect 5520 4085 5525 4115
rect 5555 4085 5560 4115
rect 5520 4035 5560 4085
rect 5520 4005 5525 4035
rect 5555 4005 5560 4035
rect 5520 3955 5560 4005
rect 5520 3925 5525 3955
rect 5555 3925 5560 3955
rect 5520 3875 5560 3925
rect 5520 3845 5525 3875
rect 5555 3845 5560 3875
rect 5520 3790 5560 3845
rect 5520 3770 5530 3790
rect 5550 3770 5560 3790
rect 5520 3715 5560 3770
rect 5520 3685 5525 3715
rect 5555 3685 5560 3715
rect 5520 3635 5560 3685
rect 5520 3605 5525 3635
rect 5555 3605 5560 3635
rect 5520 3550 5560 3605
rect 5520 3530 5530 3550
rect 5550 3530 5560 3550
rect 5520 3475 5560 3530
rect 5520 3445 5525 3475
rect 5555 3445 5560 3475
rect 5520 3395 5560 3445
rect 5520 3365 5525 3395
rect 5555 3365 5560 3395
rect 5520 3310 5560 3365
rect 5520 3290 5530 3310
rect 5550 3290 5560 3310
rect 5520 3235 5560 3290
rect 5520 3205 5525 3235
rect 5555 3205 5560 3235
rect 5520 3155 5560 3205
rect 5520 3125 5525 3155
rect 5555 3125 5560 3155
rect 5520 3075 5560 3125
rect 5520 3045 5525 3075
rect 5555 3045 5560 3075
rect 5520 2995 5560 3045
rect 5520 2965 5525 2995
rect 5555 2965 5560 2995
rect 5520 2915 5560 2965
rect 5520 2885 5525 2915
rect 5555 2885 5560 2915
rect 5520 2835 5560 2885
rect 5520 2805 5525 2835
rect 5555 2805 5560 2835
rect 5520 2755 5560 2805
rect 5520 2725 5525 2755
rect 5555 2725 5560 2755
rect 5520 2675 5560 2725
rect 5520 2645 5525 2675
rect 5555 2645 5560 2675
rect 5520 2595 5560 2645
rect 5520 2565 5525 2595
rect 5555 2565 5560 2595
rect 5520 2515 5560 2565
rect 5520 2485 5525 2515
rect 5555 2485 5560 2515
rect 5520 2435 5560 2485
rect 5520 2405 5525 2435
rect 5555 2405 5560 2435
rect 5520 2355 5560 2405
rect 5520 2325 5525 2355
rect 5555 2325 5560 2355
rect 5520 2275 5560 2325
rect 5520 2245 5525 2275
rect 5555 2245 5560 2275
rect 5520 2195 5560 2245
rect 5520 2165 5525 2195
rect 5555 2165 5560 2195
rect 5520 2115 5560 2165
rect 5520 2085 5525 2115
rect 5555 2085 5560 2115
rect 5520 2035 5560 2085
rect 5520 2005 5525 2035
rect 5555 2005 5560 2035
rect 5520 1955 5560 2005
rect 5520 1925 5525 1955
rect 5555 1925 5560 1955
rect 5520 1870 5560 1925
rect 5520 1850 5530 1870
rect 5550 1850 5560 1870
rect 5520 1790 5560 1850
rect 5520 1770 5530 1790
rect 5550 1770 5560 1790
rect 5520 1715 5560 1770
rect 5520 1685 5525 1715
rect 5555 1685 5560 1715
rect 5520 1635 5560 1685
rect 5520 1605 5525 1635
rect 5555 1605 5560 1635
rect 5520 1555 5560 1605
rect 5520 1525 5525 1555
rect 5555 1525 5560 1555
rect 5520 1475 5560 1525
rect 5520 1445 5525 1475
rect 5555 1445 5560 1475
rect 5520 1395 5560 1445
rect 5520 1365 5525 1395
rect 5555 1365 5560 1395
rect 5520 1315 5560 1365
rect 5520 1285 5525 1315
rect 5555 1285 5560 1315
rect 5520 1235 5560 1285
rect 5520 1205 5525 1235
rect 5555 1205 5560 1235
rect 5520 1155 5560 1205
rect 5520 1125 5525 1155
rect 5555 1125 5560 1155
rect 5520 1075 5560 1125
rect 5520 1045 5525 1075
rect 5555 1045 5560 1075
rect 5520 995 5560 1045
rect 5520 965 5525 995
rect 5555 965 5560 995
rect 5520 910 5560 965
rect 5520 890 5530 910
rect 5550 890 5560 910
rect 5520 835 5560 890
rect 5520 805 5525 835
rect 5555 805 5560 835
rect 5520 755 5560 805
rect 5520 725 5525 755
rect 5555 725 5560 755
rect 5520 675 5560 725
rect 5520 645 5525 675
rect 5555 645 5560 675
rect 5520 595 5560 645
rect 5520 565 5525 595
rect 5555 565 5560 595
rect 5520 515 5560 565
rect 5520 485 5525 515
rect 5555 485 5560 515
rect 5520 430 5560 485
rect 5520 410 5530 430
rect 5550 410 5560 430
rect 5520 350 5560 410
rect 5520 330 5530 350
rect 5550 330 5560 350
rect 5520 275 5560 330
rect 5520 245 5525 275
rect 5555 245 5560 275
rect 5520 195 5560 245
rect 5520 165 5525 195
rect 5555 165 5560 195
rect 5520 115 5560 165
rect 5520 85 5525 115
rect 5555 85 5560 115
rect 5520 35 5560 85
rect 5520 5 5525 35
rect 5555 5 5560 35
rect 5520 0 5560 5
rect 5600 15710 5640 15720
rect 5600 15690 5610 15710
rect 5630 15690 5640 15710
rect 5600 15630 5640 15690
rect 5600 15610 5610 15630
rect 5630 15610 5640 15630
rect 5600 15550 5640 15610
rect 5600 15530 5610 15550
rect 5630 15530 5640 15550
rect 5600 15470 5640 15530
rect 5600 15450 5610 15470
rect 5630 15450 5640 15470
rect 5600 15390 5640 15450
rect 5600 15370 5610 15390
rect 5630 15370 5640 15390
rect 5600 15310 5640 15370
rect 5600 15290 5610 15310
rect 5630 15290 5640 15310
rect 5600 15230 5640 15290
rect 5600 15210 5610 15230
rect 5630 15210 5640 15230
rect 5600 15150 5640 15210
rect 5600 15130 5610 15150
rect 5630 15130 5640 15150
rect 5600 15070 5640 15130
rect 5600 15050 5610 15070
rect 5630 15050 5640 15070
rect 5600 14990 5640 15050
rect 5600 14970 5610 14990
rect 5630 14970 5640 14990
rect 5600 14910 5640 14970
rect 5600 14890 5610 14910
rect 5630 14890 5640 14910
rect 5600 14830 5640 14890
rect 5600 14810 5610 14830
rect 5630 14810 5640 14830
rect 5600 14750 5640 14810
rect 5600 14730 5610 14750
rect 5630 14730 5640 14750
rect 5600 14670 5640 14730
rect 5600 14650 5610 14670
rect 5630 14650 5640 14670
rect 5600 14590 5640 14650
rect 5600 14570 5610 14590
rect 5630 14570 5640 14590
rect 5600 14510 5640 14570
rect 5600 14490 5610 14510
rect 5630 14490 5640 14510
rect 5600 14430 5640 14490
rect 5600 14410 5610 14430
rect 5630 14410 5640 14430
rect 5600 14350 5640 14410
rect 5600 14330 5610 14350
rect 5630 14330 5640 14350
rect 5600 14270 5640 14330
rect 5600 14250 5610 14270
rect 5630 14250 5640 14270
rect 5600 14190 5640 14250
rect 5600 14170 5610 14190
rect 5630 14170 5640 14190
rect 5600 14110 5640 14170
rect 5600 14090 5610 14110
rect 5630 14090 5640 14110
rect 5600 14030 5640 14090
rect 5600 14010 5610 14030
rect 5630 14010 5640 14030
rect 5600 13950 5640 14010
rect 5600 13930 5610 13950
rect 5630 13930 5640 13950
rect 5600 13870 5640 13930
rect 5600 13850 5610 13870
rect 5630 13850 5640 13870
rect 5600 13790 5640 13850
rect 5600 13770 5610 13790
rect 5630 13770 5640 13790
rect 5600 13710 5640 13770
rect 5600 13690 5610 13710
rect 5630 13690 5640 13710
rect 5600 13630 5640 13690
rect 5600 13610 5610 13630
rect 5630 13610 5640 13630
rect 5600 13550 5640 13610
rect 5600 13530 5610 13550
rect 5630 13530 5640 13550
rect 5600 13470 5640 13530
rect 5600 13450 5610 13470
rect 5630 13450 5640 13470
rect 5600 13390 5640 13450
rect 5600 13370 5610 13390
rect 5630 13370 5640 13390
rect 5600 13310 5640 13370
rect 5600 13290 5610 13310
rect 5630 13290 5640 13310
rect 5600 13230 5640 13290
rect 5600 13210 5610 13230
rect 5630 13210 5640 13230
rect 5600 13150 5640 13210
rect 5600 13130 5610 13150
rect 5630 13130 5640 13150
rect 5600 13070 5640 13130
rect 5600 13050 5610 13070
rect 5630 13050 5640 13070
rect 5600 12990 5640 13050
rect 5600 12970 5610 12990
rect 5630 12970 5640 12990
rect 5600 12910 5640 12970
rect 5600 12890 5610 12910
rect 5630 12890 5640 12910
rect 5600 12830 5640 12890
rect 5600 12810 5610 12830
rect 5630 12810 5640 12830
rect 5600 12750 5640 12810
rect 5600 12730 5610 12750
rect 5630 12730 5640 12750
rect 5600 12670 5640 12730
rect 5600 12650 5610 12670
rect 5630 12650 5640 12670
rect 5600 12590 5640 12650
rect 5600 12570 5610 12590
rect 5630 12570 5640 12590
rect 5600 12510 5640 12570
rect 5600 12490 5610 12510
rect 5630 12490 5640 12510
rect 5600 12430 5640 12490
rect 5600 12410 5610 12430
rect 5630 12410 5640 12430
rect 5600 12350 5640 12410
rect 5600 12330 5610 12350
rect 5630 12330 5640 12350
rect 5600 12270 5640 12330
rect 5600 12250 5610 12270
rect 5630 12250 5640 12270
rect 5600 12190 5640 12250
rect 5600 12170 5610 12190
rect 5630 12170 5640 12190
rect 5600 12110 5640 12170
rect 5600 12090 5610 12110
rect 5630 12090 5640 12110
rect 5600 12030 5640 12090
rect 5600 12010 5610 12030
rect 5630 12010 5640 12030
rect 5600 11950 5640 12010
rect 5600 11930 5610 11950
rect 5630 11930 5640 11950
rect 5600 11870 5640 11930
rect 5600 11850 5610 11870
rect 5630 11850 5640 11870
rect 5600 11790 5640 11850
rect 5600 11770 5610 11790
rect 5630 11770 5640 11790
rect 5600 11710 5640 11770
rect 5600 11690 5610 11710
rect 5630 11690 5640 11710
rect 5600 11630 5640 11690
rect 5600 11610 5610 11630
rect 5630 11610 5640 11630
rect 5600 11550 5640 11610
rect 5600 11530 5610 11550
rect 5630 11530 5640 11550
rect 5600 11470 5640 11530
rect 5600 11450 5610 11470
rect 5630 11450 5640 11470
rect 5600 11390 5640 11450
rect 5600 11370 5610 11390
rect 5630 11370 5640 11390
rect 5600 11310 5640 11370
rect 5600 11290 5610 11310
rect 5630 11290 5640 11310
rect 5600 11230 5640 11290
rect 5600 11210 5610 11230
rect 5630 11210 5640 11230
rect 5600 11150 5640 11210
rect 5600 11130 5610 11150
rect 5630 11130 5640 11150
rect 5600 11070 5640 11130
rect 5600 11050 5610 11070
rect 5630 11050 5640 11070
rect 5600 10990 5640 11050
rect 5600 10970 5610 10990
rect 5630 10970 5640 10990
rect 5600 10910 5640 10970
rect 5600 10890 5610 10910
rect 5630 10890 5640 10910
rect 5600 10830 5640 10890
rect 5600 10810 5610 10830
rect 5630 10810 5640 10830
rect 5600 10750 5640 10810
rect 5600 10730 5610 10750
rect 5630 10730 5640 10750
rect 5600 10670 5640 10730
rect 5600 10650 5610 10670
rect 5630 10650 5640 10670
rect 5600 10590 5640 10650
rect 5600 10570 5610 10590
rect 5630 10570 5640 10590
rect 5600 10510 5640 10570
rect 5600 10490 5610 10510
rect 5630 10490 5640 10510
rect 5600 10430 5640 10490
rect 5600 10410 5610 10430
rect 5630 10410 5640 10430
rect 5600 10350 5640 10410
rect 5600 10330 5610 10350
rect 5630 10330 5640 10350
rect 5600 10270 5640 10330
rect 5600 10250 5610 10270
rect 5630 10250 5640 10270
rect 5600 10190 5640 10250
rect 5600 10170 5610 10190
rect 5630 10170 5640 10190
rect 5600 10110 5640 10170
rect 5600 10090 5610 10110
rect 5630 10090 5640 10110
rect 5600 10030 5640 10090
rect 5600 10010 5610 10030
rect 5630 10010 5640 10030
rect 5600 9950 5640 10010
rect 5600 9930 5610 9950
rect 5630 9930 5640 9950
rect 5600 9870 5640 9930
rect 5600 9850 5610 9870
rect 5630 9850 5640 9870
rect 5600 9790 5640 9850
rect 5600 9770 5610 9790
rect 5630 9770 5640 9790
rect 5600 9710 5640 9770
rect 5600 9690 5610 9710
rect 5630 9690 5640 9710
rect 5600 9630 5640 9690
rect 5600 9610 5610 9630
rect 5630 9610 5640 9630
rect 5600 9550 5640 9610
rect 5600 9530 5610 9550
rect 5630 9530 5640 9550
rect 5600 9470 5640 9530
rect 5600 9450 5610 9470
rect 5630 9450 5640 9470
rect 5600 9390 5640 9450
rect 5600 9370 5610 9390
rect 5630 9370 5640 9390
rect 5600 9310 5640 9370
rect 5600 9290 5610 9310
rect 5630 9290 5640 9310
rect 5600 9230 5640 9290
rect 5600 9210 5610 9230
rect 5630 9210 5640 9230
rect 5600 9150 5640 9210
rect 5600 9130 5610 9150
rect 5630 9130 5640 9150
rect 5600 9070 5640 9130
rect 5600 9050 5610 9070
rect 5630 9050 5640 9070
rect 5600 8990 5640 9050
rect 5600 8970 5610 8990
rect 5630 8970 5640 8990
rect 5600 8910 5640 8970
rect 5600 8890 5610 8910
rect 5630 8890 5640 8910
rect 5600 8830 5640 8890
rect 5600 8810 5610 8830
rect 5630 8810 5640 8830
rect 5600 8750 5640 8810
rect 5600 8730 5610 8750
rect 5630 8730 5640 8750
rect 5600 8670 5640 8730
rect 5600 8650 5610 8670
rect 5630 8650 5640 8670
rect 5600 8590 5640 8650
rect 5600 8570 5610 8590
rect 5630 8570 5640 8590
rect 5600 8510 5640 8570
rect 5600 8490 5610 8510
rect 5630 8490 5640 8510
rect 5600 8430 5640 8490
rect 5600 8410 5610 8430
rect 5630 8410 5640 8430
rect 5600 8350 5640 8410
rect 5600 8330 5610 8350
rect 5630 8330 5640 8350
rect 5600 8270 5640 8330
rect 5600 8250 5610 8270
rect 5630 8250 5640 8270
rect 5600 8190 5640 8250
rect 5600 8170 5610 8190
rect 5630 8170 5640 8190
rect 5600 8110 5640 8170
rect 5600 8090 5610 8110
rect 5630 8090 5640 8110
rect 5600 8030 5640 8090
rect 5600 8010 5610 8030
rect 5630 8010 5640 8030
rect 5600 7950 5640 8010
rect 5600 7930 5610 7950
rect 5630 7930 5640 7950
rect 5600 7870 5640 7930
rect 5600 7850 5610 7870
rect 5630 7850 5640 7870
rect 5600 7790 5640 7850
rect 5600 7770 5610 7790
rect 5630 7770 5640 7790
rect 5600 7710 5640 7770
rect 5600 7690 5610 7710
rect 5630 7690 5640 7710
rect 5600 7630 5640 7690
rect 5600 7610 5610 7630
rect 5630 7610 5640 7630
rect 5600 7550 5640 7610
rect 5600 7530 5610 7550
rect 5630 7530 5640 7550
rect 5600 7470 5640 7530
rect 5600 7450 5610 7470
rect 5630 7450 5640 7470
rect 5600 7390 5640 7450
rect 5600 7370 5610 7390
rect 5630 7370 5640 7390
rect 5600 7310 5640 7370
rect 5600 7290 5610 7310
rect 5630 7290 5640 7310
rect 5600 7230 5640 7290
rect 5600 7210 5610 7230
rect 5630 7210 5640 7230
rect 5600 7150 5640 7210
rect 5600 7130 5610 7150
rect 5630 7130 5640 7150
rect 5600 7070 5640 7130
rect 5600 7050 5610 7070
rect 5630 7050 5640 7070
rect 5600 6990 5640 7050
rect 5600 6970 5610 6990
rect 5630 6970 5640 6990
rect 5600 6910 5640 6970
rect 5600 6890 5610 6910
rect 5630 6890 5640 6910
rect 5600 6830 5640 6890
rect 5600 6810 5610 6830
rect 5630 6810 5640 6830
rect 5600 6750 5640 6810
rect 5600 6730 5610 6750
rect 5630 6730 5640 6750
rect 5600 6670 5640 6730
rect 5600 6650 5610 6670
rect 5630 6650 5640 6670
rect 5600 6590 5640 6650
rect 5600 6570 5610 6590
rect 5630 6570 5640 6590
rect 5600 6510 5640 6570
rect 5600 6490 5610 6510
rect 5630 6490 5640 6510
rect 5600 6430 5640 6490
rect 5600 6410 5610 6430
rect 5630 6410 5640 6430
rect 5600 6350 5640 6410
rect 5600 6330 5610 6350
rect 5630 6330 5640 6350
rect 5600 6270 5640 6330
rect 5600 6250 5610 6270
rect 5630 6250 5640 6270
rect 5600 6190 5640 6250
rect 5600 6170 5610 6190
rect 5630 6170 5640 6190
rect 5600 6110 5640 6170
rect 5600 6090 5610 6110
rect 5630 6090 5640 6110
rect 5600 6030 5640 6090
rect 5600 6010 5610 6030
rect 5630 6010 5640 6030
rect 5600 5950 5640 6010
rect 5600 5930 5610 5950
rect 5630 5930 5640 5950
rect 5600 5870 5640 5930
rect 5600 5850 5610 5870
rect 5630 5850 5640 5870
rect 5600 5790 5640 5850
rect 5600 5770 5610 5790
rect 5630 5770 5640 5790
rect 5600 5710 5640 5770
rect 5600 5690 5610 5710
rect 5630 5690 5640 5710
rect 5600 5630 5640 5690
rect 5600 5610 5610 5630
rect 5630 5610 5640 5630
rect 5600 5550 5640 5610
rect 5600 5530 5610 5550
rect 5630 5530 5640 5550
rect 5600 5470 5640 5530
rect 5600 5450 5610 5470
rect 5630 5450 5640 5470
rect 5600 5390 5640 5450
rect 5600 5370 5610 5390
rect 5630 5370 5640 5390
rect 5600 5310 5640 5370
rect 5600 5290 5610 5310
rect 5630 5290 5640 5310
rect 5600 5230 5640 5290
rect 5600 5210 5610 5230
rect 5630 5210 5640 5230
rect 5600 5150 5640 5210
rect 5600 5130 5610 5150
rect 5630 5130 5640 5150
rect 5600 5070 5640 5130
rect 5600 5050 5610 5070
rect 5630 5050 5640 5070
rect 5600 4990 5640 5050
rect 5600 4970 5610 4990
rect 5630 4970 5640 4990
rect 5600 4910 5640 4970
rect 5600 4890 5610 4910
rect 5630 4890 5640 4910
rect 5600 4830 5640 4890
rect 5600 4810 5610 4830
rect 5630 4810 5640 4830
rect 5600 4750 5640 4810
rect 5600 4730 5610 4750
rect 5630 4730 5640 4750
rect 5600 4670 5640 4730
rect 5600 4650 5610 4670
rect 5630 4650 5640 4670
rect 5600 4590 5640 4650
rect 5600 4570 5610 4590
rect 5630 4570 5640 4590
rect 5600 4510 5640 4570
rect 5600 4490 5610 4510
rect 5630 4490 5640 4510
rect 5600 4430 5640 4490
rect 5600 4410 5610 4430
rect 5630 4410 5640 4430
rect 5600 4350 5640 4410
rect 5600 4330 5610 4350
rect 5630 4330 5640 4350
rect 5600 4270 5640 4330
rect 5600 4250 5610 4270
rect 5630 4250 5640 4270
rect 5600 4190 5640 4250
rect 5600 4170 5610 4190
rect 5630 4170 5640 4190
rect 5600 4110 5640 4170
rect 5600 4090 5610 4110
rect 5630 4090 5640 4110
rect 5600 4030 5640 4090
rect 5600 4010 5610 4030
rect 5630 4010 5640 4030
rect 5600 3950 5640 4010
rect 5600 3930 5610 3950
rect 5630 3930 5640 3950
rect 5600 3870 5640 3930
rect 5600 3850 5610 3870
rect 5630 3850 5640 3870
rect 5600 3790 5640 3850
rect 5600 3770 5610 3790
rect 5630 3770 5640 3790
rect 5600 3710 5640 3770
rect 5600 3690 5610 3710
rect 5630 3690 5640 3710
rect 5600 3630 5640 3690
rect 5600 3610 5610 3630
rect 5630 3610 5640 3630
rect 5600 3550 5640 3610
rect 5600 3530 5610 3550
rect 5630 3530 5640 3550
rect 5600 3470 5640 3530
rect 5600 3450 5610 3470
rect 5630 3450 5640 3470
rect 5600 3390 5640 3450
rect 5600 3370 5610 3390
rect 5630 3370 5640 3390
rect 5600 3310 5640 3370
rect 5600 3290 5610 3310
rect 5630 3290 5640 3310
rect 5600 3230 5640 3290
rect 5600 3210 5610 3230
rect 5630 3210 5640 3230
rect 5600 3150 5640 3210
rect 5600 3130 5610 3150
rect 5630 3130 5640 3150
rect 5600 3070 5640 3130
rect 5600 3050 5610 3070
rect 5630 3050 5640 3070
rect 5600 2990 5640 3050
rect 5600 2970 5610 2990
rect 5630 2970 5640 2990
rect 5600 2910 5640 2970
rect 5600 2890 5610 2910
rect 5630 2890 5640 2910
rect 5600 2830 5640 2890
rect 5600 2810 5610 2830
rect 5630 2810 5640 2830
rect 5600 2750 5640 2810
rect 5600 2730 5610 2750
rect 5630 2730 5640 2750
rect 5600 2670 5640 2730
rect 5600 2650 5610 2670
rect 5630 2650 5640 2670
rect 5600 2590 5640 2650
rect 5600 2570 5610 2590
rect 5630 2570 5640 2590
rect 5600 2510 5640 2570
rect 5600 2490 5610 2510
rect 5630 2490 5640 2510
rect 5600 2430 5640 2490
rect 5600 2410 5610 2430
rect 5630 2410 5640 2430
rect 5600 2350 5640 2410
rect 5600 2330 5610 2350
rect 5630 2330 5640 2350
rect 5600 2270 5640 2330
rect 5600 2250 5610 2270
rect 5630 2250 5640 2270
rect 5600 2190 5640 2250
rect 5600 2170 5610 2190
rect 5630 2170 5640 2190
rect 5600 2110 5640 2170
rect 5600 2090 5610 2110
rect 5630 2090 5640 2110
rect 5600 2030 5640 2090
rect 5600 2010 5610 2030
rect 5630 2010 5640 2030
rect 5600 1950 5640 2010
rect 5600 1930 5610 1950
rect 5630 1930 5640 1950
rect 5600 1870 5640 1930
rect 5600 1850 5610 1870
rect 5630 1850 5640 1870
rect 5600 1790 5640 1850
rect 5600 1770 5610 1790
rect 5630 1770 5640 1790
rect 5600 1710 5640 1770
rect 5600 1690 5610 1710
rect 5630 1690 5640 1710
rect 5600 1630 5640 1690
rect 5600 1610 5610 1630
rect 5630 1610 5640 1630
rect 5600 1550 5640 1610
rect 5600 1530 5610 1550
rect 5630 1530 5640 1550
rect 5600 1470 5640 1530
rect 5600 1450 5610 1470
rect 5630 1450 5640 1470
rect 5600 1390 5640 1450
rect 5600 1370 5610 1390
rect 5630 1370 5640 1390
rect 5600 1310 5640 1370
rect 5600 1290 5610 1310
rect 5630 1290 5640 1310
rect 5600 1230 5640 1290
rect 5600 1210 5610 1230
rect 5630 1210 5640 1230
rect 5600 1150 5640 1210
rect 5600 1130 5610 1150
rect 5630 1130 5640 1150
rect 5600 1070 5640 1130
rect 5600 1050 5610 1070
rect 5630 1050 5640 1070
rect 5600 990 5640 1050
rect 5600 970 5610 990
rect 5630 970 5640 990
rect 5600 910 5640 970
rect 5600 890 5610 910
rect 5630 890 5640 910
rect 5600 830 5640 890
rect 5600 810 5610 830
rect 5630 810 5640 830
rect 5600 750 5640 810
rect 5600 730 5610 750
rect 5630 730 5640 750
rect 5600 670 5640 730
rect 5600 650 5610 670
rect 5630 650 5640 670
rect 5600 590 5640 650
rect 5600 570 5610 590
rect 5630 570 5640 590
rect 5600 510 5640 570
rect 5600 490 5610 510
rect 5630 490 5640 510
rect 5600 430 5640 490
rect 5600 410 5610 430
rect 5630 410 5640 430
rect 5600 350 5640 410
rect 5600 330 5610 350
rect 5630 330 5640 350
rect 5600 270 5640 330
rect 5600 250 5610 270
rect 5630 250 5640 270
rect 5600 190 5640 250
rect 5600 170 5610 190
rect 5630 170 5640 190
rect 5600 110 5640 170
rect 5600 90 5610 110
rect 5630 90 5640 110
rect 5600 30 5640 90
rect 5600 10 5610 30
rect 5630 10 5640 30
rect 5600 0 5640 10
rect 5680 15715 5720 15720
rect 5680 15685 5685 15715
rect 5715 15685 5720 15715
rect 5680 15635 5720 15685
rect 5680 15605 5685 15635
rect 5715 15605 5720 15635
rect 5680 15555 5720 15605
rect 5680 15525 5685 15555
rect 5715 15525 5720 15555
rect 5680 15475 5720 15525
rect 5680 15445 5685 15475
rect 5715 15445 5720 15475
rect 5680 15395 5720 15445
rect 5680 15365 5685 15395
rect 5715 15365 5720 15395
rect 5680 15315 5720 15365
rect 5680 15285 5685 15315
rect 5715 15285 5720 15315
rect 5680 15235 5720 15285
rect 5680 15205 5685 15235
rect 5715 15205 5720 15235
rect 5680 15155 5720 15205
rect 5680 15125 5685 15155
rect 5715 15125 5720 15155
rect 5680 15070 5720 15125
rect 5680 15050 5690 15070
rect 5710 15050 5720 15070
rect 5680 14995 5720 15050
rect 5680 14965 5685 14995
rect 5715 14965 5720 14995
rect 5680 14915 5720 14965
rect 5680 14885 5685 14915
rect 5715 14885 5720 14915
rect 5680 14835 5720 14885
rect 5680 14805 5685 14835
rect 5715 14805 5720 14835
rect 5680 14755 5720 14805
rect 5680 14725 5685 14755
rect 5715 14725 5720 14755
rect 5680 14675 5720 14725
rect 5680 14645 5685 14675
rect 5715 14645 5720 14675
rect 5680 14595 5720 14645
rect 5680 14565 5685 14595
rect 5715 14565 5720 14595
rect 5680 14515 5720 14565
rect 5680 14485 5685 14515
rect 5715 14485 5720 14515
rect 5680 14435 5720 14485
rect 5680 14405 5685 14435
rect 5715 14405 5720 14435
rect 5680 14350 5720 14405
rect 5680 14330 5690 14350
rect 5710 14330 5720 14350
rect 5680 14270 5720 14330
rect 5680 14250 5690 14270
rect 5710 14250 5720 14270
rect 5680 14190 5720 14250
rect 5680 14170 5690 14190
rect 5710 14170 5720 14190
rect 5680 14110 5720 14170
rect 5680 14090 5690 14110
rect 5710 14090 5720 14110
rect 5680 14035 5720 14090
rect 5680 14005 5685 14035
rect 5715 14005 5720 14035
rect 5680 13955 5720 14005
rect 5680 13925 5685 13955
rect 5715 13925 5720 13955
rect 5680 13875 5720 13925
rect 5680 13845 5685 13875
rect 5715 13845 5720 13875
rect 5680 13795 5720 13845
rect 5680 13765 5685 13795
rect 5715 13765 5720 13795
rect 5680 13715 5720 13765
rect 5680 13685 5685 13715
rect 5715 13685 5720 13715
rect 5680 13635 5720 13685
rect 5680 13605 5685 13635
rect 5715 13605 5720 13635
rect 5680 13555 5720 13605
rect 5680 13525 5685 13555
rect 5715 13525 5720 13555
rect 5680 13475 5720 13525
rect 5680 13445 5685 13475
rect 5715 13445 5720 13475
rect 5680 13390 5720 13445
rect 5680 13370 5690 13390
rect 5710 13370 5720 13390
rect 5680 13310 5720 13370
rect 5680 13290 5690 13310
rect 5710 13290 5720 13310
rect 5680 13230 5720 13290
rect 5680 13210 5690 13230
rect 5710 13210 5720 13230
rect 5680 13150 5720 13210
rect 5680 13130 5690 13150
rect 5710 13130 5720 13150
rect 5680 13075 5720 13130
rect 5680 13045 5685 13075
rect 5715 13045 5720 13075
rect 5680 12995 5720 13045
rect 5680 12965 5685 12995
rect 5715 12965 5720 12995
rect 5680 12915 5720 12965
rect 5680 12885 5685 12915
rect 5715 12885 5720 12915
rect 5680 12835 5720 12885
rect 5680 12805 5685 12835
rect 5715 12805 5720 12835
rect 5680 12755 5720 12805
rect 5680 12725 5685 12755
rect 5715 12725 5720 12755
rect 5680 12675 5720 12725
rect 5680 12645 5685 12675
rect 5715 12645 5720 12675
rect 5680 12595 5720 12645
rect 5680 12565 5685 12595
rect 5715 12565 5720 12595
rect 5680 12515 5720 12565
rect 5680 12485 5685 12515
rect 5715 12485 5720 12515
rect 5680 12430 5720 12485
rect 5680 12410 5690 12430
rect 5710 12410 5720 12430
rect 5680 12355 5720 12410
rect 5680 12325 5685 12355
rect 5715 12325 5720 12355
rect 5680 12275 5720 12325
rect 5680 12245 5685 12275
rect 5715 12245 5720 12275
rect 5680 12195 5720 12245
rect 5680 12165 5685 12195
rect 5715 12165 5720 12195
rect 5680 12115 5720 12165
rect 5680 12085 5685 12115
rect 5715 12085 5720 12115
rect 5680 12035 5720 12085
rect 5680 12005 5685 12035
rect 5715 12005 5720 12035
rect 5680 11955 5720 12005
rect 5680 11925 5685 11955
rect 5715 11925 5720 11955
rect 5680 11875 5720 11925
rect 5680 11845 5685 11875
rect 5715 11845 5720 11875
rect 5680 11795 5720 11845
rect 5680 11765 5685 11795
rect 5715 11765 5720 11795
rect 5680 11715 5720 11765
rect 5680 11685 5685 11715
rect 5715 11685 5720 11715
rect 5680 11635 5720 11685
rect 5680 11605 5685 11635
rect 5715 11605 5720 11635
rect 5680 11555 5720 11605
rect 5680 11525 5685 11555
rect 5715 11525 5720 11555
rect 5680 11475 5720 11525
rect 5680 11445 5685 11475
rect 5715 11445 5720 11475
rect 5680 11395 5720 11445
rect 5680 11365 5685 11395
rect 5715 11365 5720 11395
rect 5680 11315 5720 11365
rect 5680 11285 5685 11315
rect 5715 11285 5720 11315
rect 5680 11235 5720 11285
rect 5680 11205 5685 11235
rect 5715 11205 5720 11235
rect 5680 11155 5720 11205
rect 5680 11125 5685 11155
rect 5715 11125 5720 11155
rect 5680 11075 5720 11125
rect 5680 11045 5685 11075
rect 5715 11045 5720 11075
rect 5680 10990 5720 11045
rect 5680 10970 5690 10990
rect 5710 10970 5720 10990
rect 5680 10915 5720 10970
rect 5680 10885 5685 10915
rect 5715 10885 5720 10915
rect 5680 10835 5720 10885
rect 5680 10805 5685 10835
rect 5715 10805 5720 10835
rect 5680 10755 5720 10805
rect 5680 10725 5685 10755
rect 5715 10725 5720 10755
rect 5680 10675 5720 10725
rect 5680 10645 5685 10675
rect 5715 10645 5720 10675
rect 5680 10595 5720 10645
rect 5680 10565 5685 10595
rect 5715 10565 5720 10595
rect 5680 10515 5720 10565
rect 5680 10485 5685 10515
rect 5715 10485 5720 10515
rect 5680 10435 5720 10485
rect 5680 10405 5685 10435
rect 5715 10405 5720 10435
rect 5680 10355 5720 10405
rect 5680 10325 5685 10355
rect 5715 10325 5720 10355
rect 5680 10270 5720 10325
rect 5680 10250 5690 10270
rect 5710 10250 5720 10270
rect 5680 10190 5720 10250
rect 5680 10170 5690 10190
rect 5710 10170 5720 10190
rect 5680 10110 5720 10170
rect 5680 10090 5690 10110
rect 5710 10090 5720 10110
rect 5680 10030 5720 10090
rect 5680 10010 5690 10030
rect 5710 10010 5720 10030
rect 5680 9955 5720 10010
rect 5680 9925 5685 9955
rect 5715 9925 5720 9955
rect 5680 9875 5720 9925
rect 5680 9845 5685 9875
rect 5715 9845 5720 9875
rect 5680 9795 5720 9845
rect 5680 9765 5685 9795
rect 5715 9765 5720 9795
rect 5680 9715 5720 9765
rect 5680 9685 5685 9715
rect 5715 9685 5720 9715
rect 5680 9635 5720 9685
rect 5680 9605 5685 9635
rect 5715 9605 5720 9635
rect 5680 9555 5720 9605
rect 5680 9525 5685 9555
rect 5715 9525 5720 9555
rect 5680 9475 5720 9525
rect 5680 9445 5685 9475
rect 5715 9445 5720 9475
rect 5680 9395 5720 9445
rect 5680 9365 5685 9395
rect 5715 9365 5720 9395
rect 5680 9310 5720 9365
rect 5680 9290 5690 9310
rect 5710 9290 5720 9310
rect 5680 9230 5720 9290
rect 5680 9210 5690 9230
rect 5710 9210 5720 9230
rect 5680 9150 5720 9210
rect 5680 9130 5690 9150
rect 5710 9130 5720 9150
rect 5680 9070 5720 9130
rect 5680 9050 5690 9070
rect 5710 9050 5720 9070
rect 5680 8995 5720 9050
rect 5680 8965 5685 8995
rect 5715 8965 5720 8995
rect 5680 8915 5720 8965
rect 5680 8885 5685 8915
rect 5715 8885 5720 8915
rect 5680 8835 5720 8885
rect 5680 8805 5685 8835
rect 5715 8805 5720 8835
rect 5680 8755 5720 8805
rect 5680 8725 5685 8755
rect 5715 8725 5720 8755
rect 5680 8675 5720 8725
rect 5680 8645 5685 8675
rect 5715 8645 5720 8675
rect 5680 8595 5720 8645
rect 5680 8565 5685 8595
rect 5715 8565 5720 8595
rect 5680 8515 5720 8565
rect 5680 8485 5685 8515
rect 5715 8485 5720 8515
rect 5680 8435 5720 8485
rect 5680 8405 5685 8435
rect 5715 8405 5720 8435
rect 5680 8350 5720 8405
rect 5680 8330 5690 8350
rect 5710 8330 5720 8350
rect 5680 8275 5720 8330
rect 5680 8245 5685 8275
rect 5715 8245 5720 8275
rect 5680 8195 5720 8245
rect 5680 8165 5685 8195
rect 5715 8165 5720 8195
rect 5680 8115 5720 8165
rect 5680 8085 5685 8115
rect 5715 8085 5720 8115
rect 5680 8035 5720 8085
rect 5680 8005 5685 8035
rect 5715 8005 5720 8035
rect 5680 7955 5720 8005
rect 5680 7925 5685 7955
rect 5715 7925 5720 7955
rect 5680 7875 5720 7925
rect 5680 7845 5685 7875
rect 5715 7845 5720 7875
rect 5680 7795 5720 7845
rect 5680 7765 5685 7795
rect 5715 7765 5720 7795
rect 5680 7715 5720 7765
rect 5680 7685 5685 7715
rect 5715 7685 5720 7715
rect 5680 7635 5720 7685
rect 5680 7605 5685 7635
rect 5715 7605 5720 7635
rect 5680 7555 5720 7605
rect 5680 7525 5685 7555
rect 5715 7525 5720 7555
rect 5680 7475 5720 7525
rect 5680 7445 5685 7475
rect 5715 7445 5720 7475
rect 5680 7395 5720 7445
rect 5680 7365 5685 7395
rect 5715 7365 5720 7395
rect 5680 7315 5720 7365
rect 5680 7285 5685 7315
rect 5715 7285 5720 7315
rect 5680 7235 5720 7285
rect 5680 7205 5685 7235
rect 5715 7205 5720 7235
rect 5680 7155 5720 7205
rect 5680 7125 5685 7155
rect 5715 7125 5720 7155
rect 5680 7075 5720 7125
rect 5680 7045 5685 7075
rect 5715 7045 5720 7075
rect 5680 6995 5720 7045
rect 5680 6965 5685 6995
rect 5715 6965 5720 6995
rect 5680 6910 5720 6965
rect 5680 6890 5690 6910
rect 5710 6890 5720 6910
rect 5680 6835 5720 6890
rect 5680 6805 5685 6835
rect 5715 6805 5720 6835
rect 5680 6755 5720 6805
rect 5680 6725 5685 6755
rect 5715 6725 5720 6755
rect 5680 6675 5720 6725
rect 5680 6645 5685 6675
rect 5715 6645 5720 6675
rect 5680 6595 5720 6645
rect 5680 6565 5685 6595
rect 5715 6565 5720 6595
rect 5680 6515 5720 6565
rect 5680 6485 5685 6515
rect 5715 6485 5720 6515
rect 5680 6435 5720 6485
rect 5680 6405 5685 6435
rect 5715 6405 5720 6435
rect 5680 6355 5720 6405
rect 5680 6325 5685 6355
rect 5715 6325 5720 6355
rect 5680 6275 5720 6325
rect 5680 6245 5685 6275
rect 5715 6245 5720 6275
rect 5680 6190 5720 6245
rect 5680 6170 5690 6190
rect 5710 6170 5720 6190
rect 5680 6110 5720 6170
rect 5680 6090 5690 6110
rect 5710 6090 5720 6110
rect 5680 6030 5720 6090
rect 5680 6010 5690 6030
rect 5710 6010 5720 6030
rect 5680 5950 5720 6010
rect 5680 5930 5690 5950
rect 5710 5930 5720 5950
rect 5680 5875 5720 5930
rect 5680 5845 5685 5875
rect 5715 5845 5720 5875
rect 5680 5795 5720 5845
rect 5680 5765 5685 5795
rect 5715 5765 5720 5795
rect 5680 5715 5720 5765
rect 5680 5685 5685 5715
rect 5715 5685 5720 5715
rect 5680 5635 5720 5685
rect 5680 5605 5685 5635
rect 5715 5605 5720 5635
rect 5680 5555 5720 5605
rect 5680 5525 5685 5555
rect 5715 5525 5720 5555
rect 5680 5475 5720 5525
rect 5680 5445 5685 5475
rect 5715 5445 5720 5475
rect 5680 5395 5720 5445
rect 5680 5365 5685 5395
rect 5715 5365 5720 5395
rect 5680 5315 5720 5365
rect 5680 5285 5685 5315
rect 5715 5285 5720 5315
rect 5680 5235 5720 5285
rect 5680 5205 5685 5235
rect 5715 5205 5720 5235
rect 5680 5155 5720 5205
rect 5680 5125 5685 5155
rect 5715 5125 5720 5155
rect 5680 5075 5720 5125
rect 5680 5045 5685 5075
rect 5715 5045 5720 5075
rect 5680 4995 5720 5045
rect 5680 4965 5685 4995
rect 5715 4965 5720 4995
rect 5680 4915 5720 4965
rect 5680 4885 5685 4915
rect 5715 4885 5720 4915
rect 5680 4830 5720 4885
rect 5680 4810 5690 4830
rect 5710 4810 5720 4830
rect 5680 4755 5720 4810
rect 5680 4725 5685 4755
rect 5715 4725 5720 4755
rect 5680 4675 5720 4725
rect 5680 4645 5685 4675
rect 5715 4645 5720 4675
rect 5680 4590 5720 4645
rect 5680 4570 5690 4590
rect 5710 4570 5720 4590
rect 5680 4515 5720 4570
rect 5680 4485 5685 4515
rect 5715 4485 5720 4515
rect 5680 4435 5720 4485
rect 5680 4405 5685 4435
rect 5715 4405 5720 4435
rect 5680 4355 5720 4405
rect 5680 4325 5685 4355
rect 5715 4325 5720 4355
rect 5680 4275 5720 4325
rect 5680 4245 5685 4275
rect 5715 4245 5720 4275
rect 5680 4195 5720 4245
rect 5680 4165 5685 4195
rect 5715 4165 5720 4195
rect 5680 4115 5720 4165
rect 5680 4085 5685 4115
rect 5715 4085 5720 4115
rect 5680 4035 5720 4085
rect 5680 4005 5685 4035
rect 5715 4005 5720 4035
rect 5680 3955 5720 4005
rect 5680 3925 5685 3955
rect 5715 3925 5720 3955
rect 5680 3875 5720 3925
rect 5680 3845 5685 3875
rect 5715 3845 5720 3875
rect 5680 3790 5720 3845
rect 5680 3770 5690 3790
rect 5710 3770 5720 3790
rect 5680 3715 5720 3770
rect 5680 3685 5685 3715
rect 5715 3685 5720 3715
rect 5680 3635 5720 3685
rect 5680 3605 5685 3635
rect 5715 3605 5720 3635
rect 5680 3550 5720 3605
rect 5680 3530 5690 3550
rect 5710 3530 5720 3550
rect 5680 3475 5720 3530
rect 5680 3445 5685 3475
rect 5715 3445 5720 3475
rect 5680 3395 5720 3445
rect 5680 3365 5685 3395
rect 5715 3365 5720 3395
rect 5680 3310 5720 3365
rect 5680 3290 5690 3310
rect 5710 3290 5720 3310
rect 5680 3235 5720 3290
rect 5680 3205 5685 3235
rect 5715 3205 5720 3235
rect 5680 3155 5720 3205
rect 5680 3125 5685 3155
rect 5715 3125 5720 3155
rect 5680 3075 5720 3125
rect 5680 3045 5685 3075
rect 5715 3045 5720 3075
rect 5680 2995 5720 3045
rect 5680 2965 5685 2995
rect 5715 2965 5720 2995
rect 5680 2915 5720 2965
rect 5680 2885 5685 2915
rect 5715 2885 5720 2915
rect 5680 2835 5720 2885
rect 5680 2805 5685 2835
rect 5715 2805 5720 2835
rect 5680 2755 5720 2805
rect 5680 2725 5685 2755
rect 5715 2725 5720 2755
rect 5680 2675 5720 2725
rect 5680 2645 5685 2675
rect 5715 2645 5720 2675
rect 5680 2595 5720 2645
rect 5680 2565 5685 2595
rect 5715 2565 5720 2595
rect 5680 2515 5720 2565
rect 5680 2485 5685 2515
rect 5715 2485 5720 2515
rect 5680 2435 5720 2485
rect 5680 2405 5685 2435
rect 5715 2405 5720 2435
rect 5680 2355 5720 2405
rect 5680 2325 5685 2355
rect 5715 2325 5720 2355
rect 5680 2275 5720 2325
rect 5680 2245 5685 2275
rect 5715 2245 5720 2275
rect 5680 2195 5720 2245
rect 5680 2165 5685 2195
rect 5715 2165 5720 2195
rect 5680 2115 5720 2165
rect 5680 2085 5685 2115
rect 5715 2085 5720 2115
rect 5680 2035 5720 2085
rect 5680 2005 5685 2035
rect 5715 2005 5720 2035
rect 5680 1955 5720 2005
rect 5680 1925 5685 1955
rect 5715 1925 5720 1955
rect 5680 1870 5720 1925
rect 5680 1850 5690 1870
rect 5710 1850 5720 1870
rect 5680 1790 5720 1850
rect 5680 1770 5690 1790
rect 5710 1770 5720 1790
rect 5680 1715 5720 1770
rect 5680 1685 5685 1715
rect 5715 1685 5720 1715
rect 5680 1635 5720 1685
rect 5680 1605 5685 1635
rect 5715 1605 5720 1635
rect 5680 1555 5720 1605
rect 5680 1525 5685 1555
rect 5715 1525 5720 1555
rect 5680 1475 5720 1525
rect 5680 1445 5685 1475
rect 5715 1445 5720 1475
rect 5680 1395 5720 1445
rect 5680 1365 5685 1395
rect 5715 1365 5720 1395
rect 5680 1315 5720 1365
rect 5680 1285 5685 1315
rect 5715 1285 5720 1315
rect 5680 1235 5720 1285
rect 5680 1205 5685 1235
rect 5715 1205 5720 1235
rect 5680 1155 5720 1205
rect 5680 1125 5685 1155
rect 5715 1125 5720 1155
rect 5680 1075 5720 1125
rect 5680 1045 5685 1075
rect 5715 1045 5720 1075
rect 5680 995 5720 1045
rect 5680 965 5685 995
rect 5715 965 5720 995
rect 5680 910 5720 965
rect 5680 890 5690 910
rect 5710 890 5720 910
rect 5680 835 5720 890
rect 5680 805 5685 835
rect 5715 805 5720 835
rect 5680 755 5720 805
rect 5680 725 5685 755
rect 5715 725 5720 755
rect 5680 675 5720 725
rect 5680 645 5685 675
rect 5715 645 5720 675
rect 5680 595 5720 645
rect 5680 565 5685 595
rect 5715 565 5720 595
rect 5680 515 5720 565
rect 5680 485 5685 515
rect 5715 485 5720 515
rect 5680 430 5720 485
rect 5680 410 5690 430
rect 5710 410 5720 430
rect 5680 350 5720 410
rect 5680 330 5690 350
rect 5710 330 5720 350
rect 5680 275 5720 330
rect 5680 245 5685 275
rect 5715 245 5720 275
rect 5680 195 5720 245
rect 5680 165 5685 195
rect 5715 165 5720 195
rect 5680 115 5720 165
rect 5680 85 5685 115
rect 5715 85 5720 115
rect 5680 35 5720 85
rect 5680 5 5685 35
rect 5715 5 5720 35
rect 5680 0 5720 5
rect 5760 15715 5800 15720
rect 5760 15685 5765 15715
rect 5795 15685 5800 15715
rect 5760 15635 5800 15685
rect 5760 15605 5765 15635
rect 5795 15605 5800 15635
rect 5760 15555 5800 15605
rect 5760 15525 5765 15555
rect 5795 15525 5800 15555
rect 5760 15475 5800 15525
rect 5760 15445 5765 15475
rect 5795 15445 5800 15475
rect 5760 15395 5800 15445
rect 5760 15365 5765 15395
rect 5795 15365 5800 15395
rect 5760 15315 5800 15365
rect 5760 15285 5765 15315
rect 5795 15285 5800 15315
rect 5760 15235 5800 15285
rect 5760 15205 5765 15235
rect 5795 15205 5800 15235
rect 5760 15155 5800 15205
rect 5760 15125 5765 15155
rect 5795 15125 5800 15155
rect 5760 15070 5800 15125
rect 5760 15050 5770 15070
rect 5790 15050 5800 15070
rect 5760 14995 5800 15050
rect 5760 14965 5765 14995
rect 5795 14965 5800 14995
rect 5760 14915 5800 14965
rect 5760 14885 5765 14915
rect 5795 14885 5800 14915
rect 5760 14835 5800 14885
rect 5760 14805 5765 14835
rect 5795 14805 5800 14835
rect 5760 14755 5800 14805
rect 5760 14725 5765 14755
rect 5795 14725 5800 14755
rect 5760 14675 5800 14725
rect 5760 14645 5765 14675
rect 5795 14645 5800 14675
rect 5760 14595 5800 14645
rect 5760 14565 5765 14595
rect 5795 14565 5800 14595
rect 5760 14515 5800 14565
rect 5760 14485 5765 14515
rect 5795 14485 5800 14515
rect 5760 14435 5800 14485
rect 5760 14405 5765 14435
rect 5795 14405 5800 14435
rect 5760 14350 5800 14405
rect 5760 14330 5770 14350
rect 5790 14330 5800 14350
rect 5760 14270 5800 14330
rect 5760 14250 5770 14270
rect 5790 14250 5800 14270
rect 5760 14190 5800 14250
rect 5760 14170 5770 14190
rect 5790 14170 5800 14190
rect 5760 14110 5800 14170
rect 5760 14090 5770 14110
rect 5790 14090 5800 14110
rect 5760 14035 5800 14090
rect 5760 14005 5765 14035
rect 5795 14005 5800 14035
rect 5760 13955 5800 14005
rect 5760 13925 5765 13955
rect 5795 13925 5800 13955
rect 5760 13875 5800 13925
rect 5760 13845 5765 13875
rect 5795 13845 5800 13875
rect 5760 13795 5800 13845
rect 5760 13765 5765 13795
rect 5795 13765 5800 13795
rect 5760 13715 5800 13765
rect 5760 13685 5765 13715
rect 5795 13685 5800 13715
rect 5760 13635 5800 13685
rect 5760 13605 5765 13635
rect 5795 13605 5800 13635
rect 5760 13555 5800 13605
rect 5760 13525 5765 13555
rect 5795 13525 5800 13555
rect 5760 13475 5800 13525
rect 5760 13445 5765 13475
rect 5795 13445 5800 13475
rect 5760 13390 5800 13445
rect 5760 13370 5770 13390
rect 5790 13370 5800 13390
rect 5760 13310 5800 13370
rect 5760 13290 5770 13310
rect 5790 13290 5800 13310
rect 5760 13230 5800 13290
rect 5760 13210 5770 13230
rect 5790 13210 5800 13230
rect 5760 13150 5800 13210
rect 5760 13130 5770 13150
rect 5790 13130 5800 13150
rect 5760 13075 5800 13130
rect 5760 13045 5765 13075
rect 5795 13045 5800 13075
rect 5760 12995 5800 13045
rect 5760 12965 5765 12995
rect 5795 12965 5800 12995
rect 5760 12915 5800 12965
rect 5760 12885 5765 12915
rect 5795 12885 5800 12915
rect 5760 12835 5800 12885
rect 5760 12805 5765 12835
rect 5795 12805 5800 12835
rect 5760 12755 5800 12805
rect 5760 12725 5765 12755
rect 5795 12725 5800 12755
rect 5760 12675 5800 12725
rect 5760 12645 5765 12675
rect 5795 12645 5800 12675
rect 5760 12595 5800 12645
rect 5760 12565 5765 12595
rect 5795 12565 5800 12595
rect 5760 12515 5800 12565
rect 5760 12485 5765 12515
rect 5795 12485 5800 12515
rect 5760 12430 5800 12485
rect 5760 12410 5770 12430
rect 5790 12410 5800 12430
rect 5760 12355 5800 12410
rect 5760 12325 5765 12355
rect 5795 12325 5800 12355
rect 5760 12275 5800 12325
rect 5760 12245 5765 12275
rect 5795 12245 5800 12275
rect 5760 12195 5800 12245
rect 5760 12165 5765 12195
rect 5795 12165 5800 12195
rect 5760 12115 5800 12165
rect 5760 12085 5765 12115
rect 5795 12085 5800 12115
rect 5760 12035 5800 12085
rect 5760 12005 5765 12035
rect 5795 12005 5800 12035
rect 5760 11955 5800 12005
rect 5760 11925 5765 11955
rect 5795 11925 5800 11955
rect 5760 11875 5800 11925
rect 5760 11845 5765 11875
rect 5795 11845 5800 11875
rect 5760 11795 5800 11845
rect 5760 11765 5765 11795
rect 5795 11765 5800 11795
rect 5760 11715 5800 11765
rect 5760 11685 5765 11715
rect 5795 11685 5800 11715
rect 5760 11635 5800 11685
rect 5760 11605 5765 11635
rect 5795 11605 5800 11635
rect 5760 11555 5800 11605
rect 5760 11525 5765 11555
rect 5795 11525 5800 11555
rect 5760 11475 5800 11525
rect 5760 11445 5765 11475
rect 5795 11445 5800 11475
rect 5760 11395 5800 11445
rect 5760 11365 5765 11395
rect 5795 11365 5800 11395
rect 5760 11315 5800 11365
rect 5760 11285 5765 11315
rect 5795 11285 5800 11315
rect 5760 11235 5800 11285
rect 5760 11205 5765 11235
rect 5795 11205 5800 11235
rect 5760 11155 5800 11205
rect 5760 11125 5765 11155
rect 5795 11125 5800 11155
rect 5760 11075 5800 11125
rect 5760 11045 5765 11075
rect 5795 11045 5800 11075
rect 5760 10990 5800 11045
rect 5760 10970 5770 10990
rect 5790 10970 5800 10990
rect 5760 10915 5800 10970
rect 5760 10885 5765 10915
rect 5795 10885 5800 10915
rect 5760 10835 5800 10885
rect 5760 10805 5765 10835
rect 5795 10805 5800 10835
rect 5760 10755 5800 10805
rect 5760 10725 5765 10755
rect 5795 10725 5800 10755
rect 5760 10675 5800 10725
rect 5760 10645 5765 10675
rect 5795 10645 5800 10675
rect 5760 10595 5800 10645
rect 5760 10565 5765 10595
rect 5795 10565 5800 10595
rect 5760 10515 5800 10565
rect 5760 10485 5765 10515
rect 5795 10485 5800 10515
rect 5760 10435 5800 10485
rect 5760 10405 5765 10435
rect 5795 10405 5800 10435
rect 5760 10355 5800 10405
rect 5760 10325 5765 10355
rect 5795 10325 5800 10355
rect 5760 10270 5800 10325
rect 5760 10250 5770 10270
rect 5790 10250 5800 10270
rect 5760 10190 5800 10250
rect 5760 10170 5770 10190
rect 5790 10170 5800 10190
rect 5760 10110 5800 10170
rect 5760 10090 5770 10110
rect 5790 10090 5800 10110
rect 5760 10030 5800 10090
rect 5760 10010 5770 10030
rect 5790 10010 5800 10030
rect 5760 9955 5800 10010
rect 5760 9925 5765 9955
rect 5795 9925 5800 9955
rect 5760 9875 5800 9925
rect 5760 9845 5765 9875
rect 5795 9845 5800 9875
rect 5760 9795 5800 9845
rect 5760 9765 5765 9795
rect 5795 9765 5800 9795
rect 5760 9715 5800 9765
rect 5760 9685 5765 9715
rect 5795 9685 5800 9715
rect 5760 9635 5800 9685
rect 5760 9605 5765 9635
rect 5795 9605 5800 9635
rect 5760 9555 5800 9605
rect 5760 9525 5765 9555
rect 5795 9525 5800 9555
rect 5760 9475 5800 9525
rect 5760 9445 5765 9475
rect 5795 9445 5800 9475
rect 5760 9395 5800 9445
rect 5760 9365 5765 9395
rect 5795 9365 5800 9395
rect 5760 9310 5800 9365
rect 5760 9290 5770 9310
rect 5790 9290 5800 9310
rect 5760 9230 5800 9290
rect 5760 9210 5770 9230
rect 5790 9210 5800 9230
rect 5760 9150 5800 9210
rect 5760 9130 5770 9150
rect 5790 9130 5800 9150
rect 5760 9070 5800 9130
rect 5760 9050 5770 9070
rect 5790 9050 5800 9070
rect 5760 8995 5800 9050
rect 5760 8965 5765 8995
rect 5795 8965 5800 8995
rect 5760 8915 5800 8965
rect 5760 8885 5765 8915
rect 5795 8885 5800 8915
rect 5760 8835 5800 8885
rect 5760 8805 5765 8835
rect 5795 8805 5800 8835
rect 5760 8755 5800 8805
rect 5760 8725 5765 8755
rect 5795 8725 5800 8755
rect 5760 8675 5800 8725
rect 5760 8645 5765 8675
rect 5795 8645 5800 8675
rect 5760 8595 5800 8645
rect 5760 8565 5765 8595
rect 5795 8565 5800 8595
rect 5760 8515 5800 8565
rect 5760 8485 5765 8515
rect 5795 8485 5800 8515
rect 5760 8435 5800 8485
rect 5760 8405 5765 8435
rect 5795 8405 5800 8435
rect 5760 8350 5800 8405
rect 5760 8330 5770 8350
rect 5790 8330 5800 8350
rect 5760 8275 5800 8330
rect 5760 8245 5765 8275
rect 5795 8245 5800 8275
rect 5760 8195 5800 8245
rect 5760 8165 5765 8195
rect 5795 8165 5800 8195
rect 5760 8115 5800 8165
rect 5760 8085 5765 8115
rect 5795 8085 5800 8115
rect 5760 8035 5800 8085
rect 5760 8005 5765 8035
rect 5795 8005 5800 8035
rect 5760 7955 5800 8005
rect 5760 7925 5765 7955
rect 5795 7925 5800 7955
rect 5760 7875 5800 7925
rect 5760 7845 5765 7875
rect 5795 7845 5800 7875
rect 5760 7795 5800 7845
rect 5760 7765 5765 7795
rect 5795 7765 5800 7795
rect 5760 7715 5800 7765
rect 5760 7685 5765 7715
rect 5795 7685 5800 7715
rect 5760 7635 5800 7685
rect 5760 7605 5765 7635
rect 5795 7605 5800 7635
rect 5760 7555 5800 7605
rect 5760 7525 5765 7555
rect 5795 7525 5800 7555
rect 5760 7475 5800 7525
rect 5760 7445 5765 7475
rect 5795 7445 5800 7475
rect 5760 7395 5800 7445
rect 5760 7365 5765 7395
rect 5795 7365 5800 7395
rect 5760 7315 5800 7365
rect 5760 7285 5765 7315
rect 5795 7285 5800 7315
rect 5760 7235 5800 7285
rect 5760 7205 5765 7235
rect 5795 7205 5800 7235
rect 5760 7155 5800 7205
rect 5760 7125 5765 7155
rect 5795 7125 5800 7155
rect 5760 7075 5800 7125
rect 5760 7045 5765 7075
rect 5795 7045 5800 7075
rect 5760 6995 5800 7045
rect 5760 6965 5765 6995
rect 5795 6965 5800 6995
rect 5760 6910 5800 6965
rect 5760 6890 5770 6910
rect 5790 6890 5800 6910
rect 5760 6835 5800 6890
rect 5760 6805 5765 6835
rect 5795 6805 5800 6835
rect 5760 6755 5800 6805
rect 5760 6725 5765 6755
rect 5795 6725 5800 6755
rect 5760 6675 5800 6725
rect 5760 6645 5765 6675
rect 5795 6645 5800 6675
rect 5760 6595 5800 6645
rect 5760 6565 5765 6595
rect 5795 6565 5800 6595
rect 5760 6515 5800 6565
rect 5760 6485 5765 6515
rect 5795 6485 5800 6515
rect 5760 6435 5800 6485
rect 5760 6405 5765 6435
rect 5795 6405 5800 6435
rect 5760 6355 5800 6405
rect 5760 6325 5765 6355
rect 5795 6325 5800 6355
rect 5760 6275 5800 6325
rect 5760 6245 5765 6275
rect 5795 6245 5800 6275
rect 5760 6190 5800 6245
rect 5760 6170 5770 6190
rect 5790 6170 5800 6190
rect 5760 6110 5800 6170
rect 5760 6090 5770 6110
rect 5790 6090 5800 6110
rect 5760 6030 5800 6090
rect 5760 6010 5770 6030
rect 5790 6010 5800 6030
rect 5760 5950 5800 6010
rect 5760 5930 5770 5950
rect 5790 5930 5800 5950
rect 5760 5875 5800 5930
rect 5760 5845 5765 5875
rect 5795 5845 5800 5875
rect 5760 5795 5800 5845
rect 5760 5765 5765 5795
rect 5795 5765 5800 5795
rect 5760 5715 5800 5765
rect 5760 5685 5765 5715
rect 5795 5685 5800 5715
rect 5760 5635 5800 5685
rect 5760 5605 5765 5635
rect 5795 5605 5800 5635
rect 5760 5555 5800 5605
rect 5760 5525 5765 5555
rect 5795 5525 5800 5555
rect 5760 5475 5800 5525
rect 5760 5445 5765 5475
rect 5795 5445 5800 5475
rect 5760 5395 5800 5445
rect 5760 5365 5765 5395
rect 5795 5365 5800 5395
rect 5760 5315 5800 5365
rect 5760 5285 5765 5315
rect 5795 5285 5800 5315
rect 5760 5235 5800 5285
rect 5760 5205 5765 5235
rect 5795 5205 5800 5235
rect 5760 5155 5800 5205
rect 5760 5125 5765 5155
rect 5795 5125 5800 5155
rect 5760 5075 5800 5125
rect 5760 5045 5765 5075
rect 5795 5045 5800 5075
rect 5760 4995 5800 5045
rect 5760 4965 5765 4995
rect 5795 4965 5800 4995
rect 5760 4915 5800 4965
rect 5760 4885 5765 4915
rect 5795 4885 5800 4915
rect 5760 4830 5800 4885
rect 5760 4810 5770 4830
rect 5790 4810 5800 4830
rect 5760 4755 5800 4810
rect 5760 4725 5765 4755
rect 5795 4725 5800 4755
rect 5760 4675 5800 4725
rect 5760 4645 5765 4675
rect 5795 4645 5800 4675
rect 5760 4590 5800 4645
rect 5760 4570 5770 4590
rect 5790 4570 5800 4590
rect 5760 4515 5800 4570
rect 5760 4485 5765 4515
rect 5795 4485 5800 4515
rect 5760 4435 5800 4485
rect 5760 4405 5765 4435
rect 5795 4405 5800 4435
rect 5760 4355 5800 4405
rect 5760 4325 5765 4355
rect 5795 4325 5800 4355
rect 5760 4275 5800 4325
rect 5760 4245 5765 4275
rect 5795 4245 5800 4275
rect 5760 4195 5800 4245
rect 5760 4165 5765 4195
rect 5795 4165 5800 4195
rect 5760 4115 5800 4165
rect 5760 4085 5765 4115
rect 5795 4085 5800 4115
rect 5760 4035 5800 4085
rect 5760 4005 5765 4035
rect 5795 4005 5800 4035
rect 5760 3955 5800 4005
rect 5760 3925 5765 3955
rect 5795 3925 5800 3955
rect 5760 3875 5800 3925
rect 5760 3845 5765 3875
rect 5795 3845 5800 3875
rect 5760 3790 5800 3845
rect 5760 3770 5770 3790
rect 5790 3770 5800 3790
rect 5760 3715 5800 3770
rect 5760 3685 5765 3715
rect 5795 3685 5800 3715
rect 5760 3635 5800 3685
rect 5760 3605 5765 3635
rect 5795 3605 5800 3635
rect 5760 3550 5800 3605
rect 5760 3530 5770 3550
rect 5790 3530 5800 3550
rect 5760 3475 5800 3530
rect 5760 3445 5765 3475
rect 5795 3445 5800 3475
rect 5760 3395 5800 3445
rect 5760 3365 5765 3395
rect 5795 3365 5800 3395
rect 5760 3310 5800 3365
rect 5760 3290 5770 3310
rect 5790 3290 5800 3310
rect 5760 3235 5800 3290
rect 5760 3205 5765 3235
rect 5795 3205 5800 3235
rect 5760 3155 5800 3205
rect 5760 3125 5765 3155
rect 5795 3125 5800 3155
rect 5760 3075 5800 3125
rect 5760 3045 5765 3075
rect 5795 3045 5800 3075
rect 5760 2995 5800 3045
rect 5760 2965 5765 2995
rect 5795 2965 5800 2995
rect 5760 2915 5800 2965
rect 5760 2885 5765 2915
rect 5795 2885 5800 2915
rect 5760 2835 5800 2885
rect 5760 2805 5765 2835
rect 5795 2805 5800 2835
rect 5760 2755 5800 2805
rect 5760 2725 5765 2755
rect 5795 2725 5800 2755
rect 5760 2675 5800 2725
rect 5760 2645 5765 2675
rect 5795 2645 5800 2675
rect 5760 2595 5800 2645
rect 5760 2565 5765 2595
rect 5795 2565 5800 2595
rect 5760 2515 5800 2565
rect 5760 2485 5765 2515
rect 5795 2485 5800 2515
rect 5760 2435 5800 2485
rect 5760 2405 5765 2435
rect 5795 2405 5800 2435
rect 5760 2355 5800 2405
rect 5760 2325 5765 2355
rect 5795 2325 5800 2355
rect 5760 2275 5800 2325
rect 5760 2245 5765 2275
rect 5795 2245 5800 2275
rect 5760 2195 5800 2245
rect 5760 2165 5765 2195
rect 5795 2165 5800 2195
rect 5760 2115 5800 2165
rect 5760 2085 5765 2115
rect 5795 2085 5800 2115
rect 5760 2035 5800 2085
rect 5760 2005 5765 2035
rect 5795 2005 5800 2035
rect 5760 1955 5800 2005
rect 5760 1925 5765 1955
rect 5795 1925 5800 1955
rect 5760 1870 5800 1925
rect 5760 1850 5770 1870
rect 5790 1850 5800 1870
rect 5760 1790 5800 1850
rect 5760 1770 5770 1790
rect 5790 1770 5800 1790
rect 5760 1715 5800 1770
rect 5760 1685 5765 1715
rect 5795 1685 5800 1715
rect 5760 1635 5800 1685
rect 5760 1605 5765 1635
rect 5795 1605 5800 1635
rect 5760 1555 5800 1605
rect 5760 1525 5765 1555
rect 5795 1525 5800 1555
rect 5760 1475 5800 1525
rect 5760 1445 5765 1475
rect 5795 1445 5800 1475
rect 5760 1395 5800 1445
rect 5760 1365 5765 1395
rect 5795 1365 5800 1395
rect 5760 1315 5800 1365
rect 5760 1285 5765 1315
rect 5795 1285 5800 1315
rect 5760 1235 5800 1285
rect 5760 1205 5765 1235
rect 5795 1205 5800 1235
rect 5760 1155 5800 1205
rect 5760 1125 5765 1155
rect 5795 1125 5800 1155
rect 5760 1075 5800 1125
rect 5760 1045 5765 1075
rect 5795 1045 5800 1075
rect 5760 995 5800 1045
rect 5760 965 5765 995
rect 5795 965 5800 995
rect 5760 910 5800 965
rect 5760 890 5770 910
rect 5790 890 5800 910
rect 5760 835 5800 890
rect 5760 805 5765 835
rect 5795 805 5800 835
rect 5760 755 5800 805
rect 5760 725 5765 755
rect 5795 725 5800 755
rect 5760 675 5800 725
rect 5760 645 5765 675
rect 5795 645 5800 675
rect 5760 595 5800 645
rect 5760 565 5765 595
rect 5795 565 5800 595
rect 5760 515 5800 565
rect 5760 485 5765 515
rect 5795 485 5800 515
rect 5760 430 5800 485
rect 5760 410 5770 430
rect 5790 410 5800 430
rect 5760 350 5800 410
rect 5760 330 5770 350
rect 5790 330 5800 350
rect 5760 275 5800 330
rect 5760 245 5765 275
rect 5795 245 5800 275
rect 5760 195 5800 245
rect 5760 165 5765 195
rect 5795 165 5800 195
rect 5760 115 5800 165
rect 5760 85 5765 115
rect 5795 85 5800 115
rect 5760 35 5800 85
rect 5760 5 5765 35
rect 5795 5 5800 35
rect 5760 0 5800 5
rect 5840 15710 5880 15720
rect 5840 15690 5850 15710
rect 5870 15690 5880 15710
rect 5840 15630 5880 15690
rect 5840 15610 5850 15630
rect 5870 15610 5880 15630
rect 5840 15550 5880 15610
rect 5840 15530 5850 15550
rect 5870 15530 5880 15550
rect 5840 15470 5880 15530
rect 5840 15450 5850 15470
rect 5870 15450 5880 15470
rect 5840 15390 5880 15450
rect 5840 15370 5850 15390
rect 5870 15370 5880 15390
rect 5840 15310 5880 15370
rect 5840 15290 5850 15310
rect 5870 15290 5880 15310
rect 5840 15230 5880 15290
rect 5840 15210 5850 15230
rect 5870 15210 5880 15230
rect 5840 15150 5880 15210
rect 5840 15130 5850 15150
rect 5870 15130 5880 15150
rect 5840 15070 5880 15130
rect 5840 15050 5850 15070
rect 5870 15050 5880 15070
rect 5840 14990 5880 15050
rect 5840 14970 5850 14990
rect 5870 14970 5880 14990
rect 5840 14910 5880 14970
rect 5840 14890 5850 14910
rect 5870 14890 5880 14910
rect 5840 14830 5880 14890
rect 5840 14810 5850 14830
rect 5870 14810 5880 14830
rect 5840 14750 5880 14810
rect 5840 14730 5850 14750
rect 5870 14730 5880 14750
rect 5840 14670 5880 14730
rect 5840 14650 5850 14670
rect 5870 14650 5880 14670
rect 5840 14590 5880 14650
rect 5840 14570 5850 14590
rect 5870 14570 5880 14590
rect 5840 14510 5880 14570
rect 5840 14490 5850 14510
rect 5870 14490 5880 14510
rect 5840 14430 5880 14490
rect 5840 14410 5850 14430
rect 5870 14410 5880 14430
rect 5840 14350 5880 14410
rect 5840 14330 5850 14350
rect 5870 14330 5880 14350
rect 5840 14270 5880 14330
rect 5840 14250 5850 14270
rect 5870 14250 5880 14270
rect 5840 14190 5880 14250
rect 5840 14170 5850 14190
rect 5870 14170 5880 14190
rect 5840 14110 5880 14170
rect 5840 14090 5850 14110
rect 5870 14090 5880 14110
rect 5840 14030 5880 14090
rect 5840 14010 5850 14030
rect 5870 14010 5880 14030
rect 5840 13950 5880 14010
rect 5840 13930 5850 13950
rect 5870 13930 5880 13950
rect 5840 13870 5880 13930
rect 5840 13850 5850 13870
rect 5870 13850 5880 13870
rect 5840 13790 5880 13850
rect 5840 13770 5850 13790
rect 5870 13770 5880 13790
rect 5840 13710 5880 13770
rect 5840 13690 5850 13710
rect 5870 13690 5880 13710
rect 5840 13630 5880 13690
rect 5840 13610 5850 13630
rect 5870 13610 5880 13630
rect 5840 13550 5880 13610
rect 5840 13530 5850 13550
rect 5870 13530 5880 13550
rect 5840 13470 5880 13530
rect 5840 13450 5850 13470
rect 5870 13450 5880 13470
rect 5840 13390 5880 13450
rect 5840 13370 5850 13390
rect 5870 13370 5880 13390
rect 5840 13310 5880 13370
rect 5840 13290 5850 13310
rect 5870 13290 5880 13310
rect 5840 13230 5880 13290
rect 5840 13210 5850 13230
rect 5870 13210 5880 13230
rect 5840 13150 5880 13210
rect 5840 13130 5850 13150
rect 5870 13130 5880 13150
rect 5840 13070 5880 13130
rect 5840 13050 5850 13070
rect 5870 13050 5880 13070
rect 5840 12990 5880 13050
rect 5840 12970 5850 12990
rect 5870 12970 5880 12990
rect 5840 12910 5880 12970
rect 5840 12890 5850 12910
rect 5870 12890 5880 12910
rect 5840 12830 5880 12890
rect 5840 12810 5850 12830
rect 5870 12810 5880 12830
rect 5840 12750 5880 12810
rect 5840 12730 5850 12750
rect 5870 12730 5880 12750
rect 5840 12670 5880 12730
rect 5840 12650 5850 12670
rect 5870 12650 5880 12670
rect 5840 12590 5880 12650
rect 5840 12570 5850 12590
rect 5870 12570 5880 12590
rect 5840 12510 5880 12570
rect 5840 12490 5850 12510
rect 5870 12490 5880 12510
rect 5840 12430 5880 12490
rect 5840 12410 5850 12430
rect 5870 12410 5880 12430
rect 5840 12350 5880 12410
rect 5840 12330 5850 12350
rect 5870 12330 5880 12350
rect 5840 12270 5880 12330
rect 5840 12250 5850 12270
rect 5870 12250 5880 12270
rect 5840 12190 5880 12250
rect 5840 12170 5850 12190
rect 5870 12170 5880 12190
rect 5840 12110 5880 12170
rect 5840 12090 5850 12110
rect 5870 12090 5880 12110
rect 5840 12030 5880 12090
rect 5840 12010 5850 12030
rect 5870 12010 5880 12030
rect 5840 11950 5880 12010
rect 5840 11930 5850 11950
rect 5870 11930 5880 11950
rect 5840 11870 5880 11930
rect 5840 11850 5850 11870
rect 5870 11850 5880 11870
rect 5840 11790 5880 11850
rect 5840 11770 5850 11790
rect 5870 11770 5880 11790
rect 5840 11710 5880 11770
rect 5840 11690 5850 11710
rect 5870 11690 5880 11710
rect 5840 11630 5880 11690
rect 5840 11610 5850 11630
rect 5870 11610 5880 11630
rect 5840 11550 5880 11610
rect 5840 11530 5850 11550
rect 5870 11530 5880 11550
rect 5840 11470 5880 11530
rect 5840 11450 5850 11470
rect 5870 11450 5880 11470
rect 5840 11390 5880 11450
rect 5840 11370 5850 11390
rect 5870 11370 5880 11390
rect 5840 11310 5880 11370
rect 5840 11290 5850 11310
rect 5870 11290 5880 11310
rect 5840 11230 5880 11290
rect 5840 11210 5850 11230
rect 5870 11210 5880 11230
rect 5840 11150 5880 11210
rect 5840 11130 5850 11150
rect 5870 11130 5880 11150
rect 5840 11070 5880 11130
rect 5840 11050 5850 11070
rect 5870 11050 5880 11070
rect 5840 10990 5880 11050
rect 5840 10970 5850 10990
rect 5870 10970 5880 10990
rect 5840 10910 5880 10970
rect 5840 10890 5850 10910
rect 5870 10890 5880 10910
rect 5840 10830 5880 10890
rect 5840 10810 5850 10830
rect 5870 10810 5880 10830
rect 5840 10750 5880 10810
rect 5840 10730 5850 10750
rect 5870 10730 5880 10750
rect 5840 10670 5880 10730
rect 5840 10650 5850 10670
rect 5870 10650 5880 10670
rect 5840 10590 5880 10650
rect 5840 10570 5850 10590
rect 5870 10570 5880 10590
rect 5840 10510 5880 10570
rect 5840 10490 5850 10510
rect 5870 10490 5880 10510
rect 5840 10430 5880 10490
rect 5840 10410 5850 10430
rect 5870 10410 5880 10430
rect 5840 10350 5880 10410
rect 5840 10330 5850 10350
rect 5870 10330 5880 10350
rect 5840 10270 5880 10330
rect 5840 10250 5850 10270
rect 5870 10250 5880 10270
rect 5840 10190 5880 10250
rect 5840 10170 5850 10190
rect 5870 10170 5880 10190
rect 5840 10110 5880 10170
rect 5840 10090 5850 10110
rect 5870 10090 5880 10110
rect 5840 10030 5880 10090
rect 5840 10010 5850 10030
rect 5870 10010 5880 10030
rect 5840 9950 5880 10010
rect 5840 9930 5850 9950
rect 5870 9930 5880 9950
rect 5840 9870 5880 9930
rect 5840 9850 5850 9870
rect 5870 9850 5880 9870
rect 5840 9790 5880 9850
rect 5840 9770 5850 9790
rect 5870 9770 5880 9790
rect 5840 9710 5880 9770
rect 5840 9690 5850 9710
rect 5870 9690 5880 9710
rect 5840 9630 5880 9690
rect 5840 9610 5850 9630
rect 5870 9610 5880 9630
rect 5840 9550 5880 9610
rect 5840 9530 5850 9550
rect 5870 9530 5880 9550
rect 5840 9470 5880 9530
rect 5840 9450 5850 9470
rect 5870 9450 5880 9470
rect 5840 9390 5880 9450
rect 5840 9370 5850 9390
rect 5870 9370 5880 9390
rect 5840 9310 5880 9370
rect 5840 9290 5850 9310
rect 5870 9290 5880 9310
rect 5840 9230 5880 9290
rect 5840 9210 5850 9230
rect 5870 9210 5880 9230
rect 5840 9150 5880 9210
rect 5840 9130 5850 9150
rect 5870 9130 5880 9150
rect 5840 9070 5880 9130
rect 5840 9050 5850 9070
rect 5870 9050 5880 9070
rect 5840 8990 5880 9050
rect 5840 8970 5850 8990
rect 5870 8970 5880 8990
rect 5840 8910 5880 8970
rect 5840 8890 5850 8910
rect 5870 8890 5880 8910
rect 5840 8830 5880 8890
rect 5840 8810 5850 8830
rect 5870 8810 5880 8830
rect 5840 8750 5880 8810
rect 5840 8730 5850 8750
rect 5870 8730 5880 8750
rect 5840 8670 5880 8730
rect 5840 8650 5850 8670
rect 5870 8650 5880 8670
rect 5840 8590 5880 8650
rect 5840 8570 5850 8590
rect 5870 8570 5880 8590
rect 5840 8510 5880 8570
rect 5840 8490 5850 8510
rect 5870 8490 5880 8510
rect 5840 8430 5880 8490
rect 5840 8410 5850 8430
rect 5870 8410 5880 8430
rect 5840 8350 5880 8410
rect 5840 8330 5850 8350
rect 5870 8330 5880 8350
rect 5840 8270 5880 8330
rect 5840 8250 5850 8270
rect 5870 8250 5880 8270
rect 5840 8190 5880 8250
rect 5840 8170 5850 8190
rect 5870 8170 5880 8190
rect 5840 8110 5880 8170
rect 5840 8090 5850 8110
rect 5870 8090 5880 8110
rect 5840 8030 5880 8090
rect 5840 8010 5850 8030
rect 5870 8010 5880 8030
rect 5840 7950 5880 8010
rect 5840 7930 5850 7950
rect 5870 7930 5880 7950
rect 5840 7870 5880 7930
rect 5840 7850 5850 7870
rect 5870 7850 5880 7870
rect 5840 7790 5880 7850
rect 5840 7770 5850 7790
rect 5870 7770 5880 7790
rect 5840 7710 5880 7770
rect 5840 7690 5850 7710
rect 5870 7690 5880 7710
rect 5840 7630 5880 7690
rect 5840 7610 5850 7630
rect 5870 7610 5880 7630
rect 5840 7550 5880 7610
rect 5840 7530 5850 7550
rect 5870 7530 5880 7550
rect 5840 7470 5880 7530
rect 5840 7450 5850 7470
rect 5870 7450 5880 7470
rect 5840 7390 5880 7450
rect 5840 7370 5850 7390
rect 5870 7370 5880 7390
rect 5840 7310 5880 7370
rect 5840 7290 5850 7310
rect 5870 7290 5880 7310
rect 5840 7230 5880 7290
rect 5840 7210 5850 7230
rect 5870 7210 5880 7230
rect 5840 7150 5880 7210
rect 5840 7130 5850 7150
rect 5870 7130 5880 7150
rect 5840 7070 5880 7130
rect 5840 7050 5850 7070
rect 5870 7050 5880 7070
rect 5840 6990 5880 7050
rect 5840 6970 5850 6990
rect 5870 6970 5880 6990
rect 5840 6910 5880 6970
rect 5840 6890 5850 6910
rect 5870 6890 5880 6910
rect 5840 6830 5880 6890
rect 5840 6810 5850 6830
rect 5870 6810 5880 6830
rect 5840 6750 5880 6810
rect 5840 6730 5850 6750
rect 5870 6730 5880 6750
rect 5840 6670 5880 6730
rect 5840 6650 5850 6670
rect 5870 6650 5880 6670
rect 5840 6590 5880 6650
rect 5840 6570 5850 6590
rect 5870 6570 5880 6590
rect 5840 6510 5880 6570
rect 5840 6490 5850 6510
rect 5870 6490 5880 6510
rect 5840 6430 5880 6490
rect 5840 6410 5850 6430
rect 5870 6410 5880 6430
rect 5840 6350 5880 6410
rect 5840 6330 5850 6350
rect 5870 6330 5880 6350
rect 5840 6270 5880 6330
rect 5840 6250 5850 6270
rect 5870 6250 5880 6270
rect 5840 6190 5880 6250
rect 5840 6170 5850 6190
rect 5870 6170 5880 6190
rect 5840 6110 5880 6170
rect 5840 6090 5850 6110
rect 5870 6090 5880 6110
rect 5840 6030 5880 6090
rect 5840 6010 5850 6030
rect 5870 6010 5880 6030
rect 5840 5950 5880 6010
rect 5840 5930 5850 5950
rect 5870 5930 5880 5950
rect 5840 5870 5880 5930
rect 5840 5850 5850 5870
rect 5870 5850 5880 5870
rect 5840 5790 5880 5850
rect 5840 5770 5850 5790
rect 5870 5770 5880 5790
rect 5840 5710 5880 5770
rect 5840 5690 5850 5710
rect 5870 5690 5880 5710
rect 5840 5630 5880 5690
rect 5840 5610 5850 5630
rect 5870 5610 5880 5630
rect 5840 5550 5880 5610
rect 5840 5530 5850 5550
rect 5870 5530 5880 5550
rect 5840 5470 5880 5530
rect 5840 5450 5850 5470
rect 5870 5450 5880 5470
rect 5840 5390 5880 5450
rect 5840 5370 5850 5390
rect 5870 5370 5880 5390
rect 5840 5310 5880 5370
rect 5840 5290 5850 5310
rect 5870 5290 5880 5310
rect 5840 5230 5880 5290
rect 5840 5210 5850 5230
rect 5870 5210 5880 5230
rect 5840 5150 5880 5210
rect 5840 5130 5850 5150
rect 5870 5130 5880 5150
rect 5840 5070 5880 5130
rect 5840 5050 5850 5070
rect 5870 5050 5880 5070
rect 5840 4990 5880 5050
rect 5840 4970 5850 4990
rect 5870 4970 5880 4990
rect 5840 4910 5880 4970
rect 5840 4890 5850 4910
rect 5870 4890 5880 4910
rect 5840 4830 5880 4890
rect 5840 4810 5850 4830
rect 5870 4810 5880 4830
rect 5840 4750 5880 4810
rect 5840 4730 5850 4750
rect 5870 4730 5880 4750
rect 5840 4670 5880 4730
rect 5840 4650 5850 4670
rect 5870 4650 5880 4670
rect 5840 4590 5880 4650
rect 5840 4570 5850 4590
rect 5870 4570 5880 4590
rect 5840 4510 5880 4570
rect 5840 4490 5850 4510
rect 5870 4490 5880 4510
rect 5840 4430 5880 4490
rect 5840 4410 5850 4430
rect 5870 4410 5880 4430
rect 5840 4350 5880 4410
rect 5840 4330 5850 4350
rect 5870 4330 5880 4350
rect 5840 4270 5880 4330
rect 5840 4250 5850 4270
rect 5870 4250 5880 4270
rect 5840 4190 5880 4250
rect 5840 4170 5850 4190
rect 5870 4170 5880 4190
rect 5840 4110 5880 4170
rect 5840 4090 5850 4110
rect 5870 4090 5880 4110
rect 5840 4030 5880 4090
rect 5840 4010 5850 4030
rect 5870 4010 5880 4030
rect 5840 3950 5880 4010
rect 5840 3930 5850 3950
rect 5870 3930 5880 3950
rect 5840 3870 5880 3930
rect 5840 3850 5850 3870
rect 5870 3850 5880 3870
rect 5840 3790 5880 3850
rect 5840 3770 5850 3790
rect 5870 3770 5880 3790
rect 5840 3710 5880 3770
rect 5840 3690 5850 3710
rect 5870 3690 5880 3710
rect 5840 3630 5880 3690
rect 5840 3610 5850 3630
rect 5870 3610 5880 3630
rect 5840 3550 5880 3610
rect 5840 3530 5850 3550
rect 5870 3530 5880 3550
rect 5840 3470 5880 3530
rect 5840 3450 5850 3470
rect 5870 3450 5880 3470
rect 5840 3390 5880 3450
rect 5840 3370 5850 3390
rect 5870 3370 5880 3390
rect 5840 3310 5880 3370
rect 5840 3290 5850 3310
rect 5870 3290 5880 3310
rect 5840 3230 5880 3290
rect 5840 3210 5850 3230
rect 5870 3210 5880 3230
rect 5840 3150 5880 3210
rect 5840 3130 5850 3150
rect 5870 3130 5880 3150
rect 5840 3070 5880 3130
rect 5840 3050 5850 3070
rect 5870 3050 5880 3070
rect 5840 2990 5880 3050
rect 5840 2970 5850 2990
rect 5870 2970 5880 2990
rect 5840 2910 5880 2970
rect 5840 2890 5850 2910
rect 5870 2890 5880 2910
rect 5840 2830 5880 2890
rect 5840 2810 5850 2830
rect 5870 2810 5880 2830
rect 5840 2750 5880 2810
rect 5840 2730 5850 2750
rect 5870 2730 5880 2750
rect 5840 2670 5880 2730
rect 5840 2650 5850 2670
rect 5870 2650 5880 2670
rect 5840 2590 5880 2650
rect 5840 2570 5850 2590
rect 5870 2570 5880 2590
rect 5840 2510 5880 2570
rect 5840 2490 5850 2510
rect 5870 2490 5880 2510
rect 5840 2430 5880 2490
rect 5840 2410 5850 2430
rect 5870 2410 5880 2430
rect 5840 2350 5880 2410
rect 5840 2330 5850 2350
rect 5870 2330 5880 2350
rect 5840 2270 5880 2330
rect 5840 2250 5850 2270
rect 5870 2250 5880 2270
rect 5840 2190 5880 2250
rect 5840 2170 5850 2190
rect 5870 2170 5880 2190
rect 5840 2110 5880 2170
rect 5840 2090 5850 2110
rect 5870 2090 5880 2110
rect 5840 2030 5880 2090
rect 5840 2010 5850 2030
rect 5870 2010 5880 2030
rect 5840 1950 5880 2010
rect 5840 1930 5850 1950
rect 5870 1930 5880 1950
rect 5840 1870 5880 1930
rect 5840 1850 5850 1870
rect 5870 1850 5880 1870
rect 5840 1790 5880 1850
rect 5840 1770 5850 1790
rect 5870 1770 5880 1790
rect 5840 1710 5880 1770
rect 5840 1690 5850 1710
rect 5870 1690 5880 1710
rect 5840 1630 5880 1690
rect 5840 1610 5850 1630
rect 5870 1610 5880 1630
rect 5840 1550 5880 1610
rect 5840 1530 5850 1550
rect 5870 1530 5880 1550
rect 5840 1470 5880 1530
rect 5840 1450 5850 1470
rect 5870 1450 5880 1470
rect 5840 1390 5880 1450
rect 5840 1370 5850 1390
rect 5870 1370 5880 1390
rect 5840 1310 5880 1370
rect 5840 1290 5850 1310
rect 5870 1290 5880 1310
rect 5840 1230 5880 1290
rect 5840 1210 5850 1230
rect 5870 1210 5880 1230
rect 5840 1150 5880 1210
rect 5840 1130 5850 1150
rect 5870 1130 5880 1150
rect 5840 1070 5880 1130
rect 5840 1050 5850 1070
rect 5870 1050 5880 1070
rect 5840 990 5880 1050
rect 5840 970 5850 990
rect 5870 970 5880 990
rect 5840 910 5880 970
rect 5840 890 5850 910
rect 5870 890 5880 910
rect 5840 830 5880 890
rect 5840 810 5850 830
rect 5870 810 5880 830
rect 5840 750 5880 810
rect 5840 730 5850 750
rect 5870 730 5880 750
rect 5840 670 5880 730
rect 5840 650 5850 670
rect 5870 650 5880 670
rect 5840 590 5880 650
rect 5840 570 5850 590
rect 5870 570 5880 590
rect 5840 510 5880 570
rect 5840 490 5850 510
rect 5870 490 5880 510
rect 5840 430 5880 490
rect 5840 410 5850 430
rect 5870 410 5880 430
rect 5840 350 5880 410
rect 5840 330 5850 350
rect 5870 330 5880 350
rect 5840 270 5880 330
rect 5840 250 5850 270
rect 5870 250 5880 270
rect 5840 190 5880 250
rect 5840 170 5850 190
rect 5870 170 5880 190
rect 5840 110 5880 170
rect 5840 90 5850 110
rect 5870 90 5880 110
rect 5840 30 5880 90
rect 5840 10 5850 30
rect 5870 10 5880 30
rect 5840 0 5880 10
rect 5920 15715 5960 15720
rect 5920 15685 5925 15715
rect 5955 15685 5960 15715
rect 5920 15635 5960 15685
rect 5920 15605 5925 15635
rect 5955 15605 5960 15635
rect 5920 15555 5960 15605
rect 5920 15525 5925 15555
rect 5955 15525 5960 15555
rect 5920 15475 5960 15525
rect 5920 15445 5925 15475
rect 5955 15445 5960 15475
rect 5920 15395 5960 15445
rect 5920 15365 5925 15395
rect 5955 15365 5960 15395
rect 5920 15315 5960 15365
rect 5920 15285 5925 15315
rect 5955 15285 5960 15315
rect 5920 15235 5960 15285
rect 5920 15205 5925 15235
rect 5955 15205 5960 15235
rect 5920 15155 5960 15205
rect 5920 15125 5925 15155
rect 5955 15125 5960 15155
rect 5920 15070 5960 15125
rect 5920 15050 5930 15070
rect 5950 15050 5960 15070
rect 5920 14995 5960 15050
rect 5920 14965 5925 14995
rect 5955 14965 5960 14995
rect 5920 14915 5960 14965
rect 5920 14885 5925 14915
rect 5955 14885 5960 14915
rect 5920 14835 5960 14885
rect 5920 14805 5925 14835
rect 5955 14805 5960 14835
rect 5920 14755 5960 14805
rect 5920 14725 5925 14755
rect 5955 14725 5960 14755
rect 5920 14675 5960 14725
rect 5920 14645 5925 14675
rect 5955 14645 5960 14675
rect 5920 14595 5960 14645
rect 5920 14565 5925 14595
rect 5955 14565 5960 14595
rect 5920 14515 5960 14565
rect 5920 14485 5925 14515
rect 5955 14485 5960 14515
rect 5920 14435 5960 14485
rect 5920 14405 5925 14435
rect 5955 14405 5960 14435
rect 5920 14350 5960 14405
rect 5920 14330 5930 14350
rect 5950 14330 5960 14350
rect 5920 14270 5960 14330
rect 5920 14250 5930 14270
rect 5950 14250 5960 14270
rect 5920 14190 5960 14250
rect 5920 14170 5930 14190
rect 5950 14170 5960 14190
rect 5920 14110 5960 14170
rect 5920 14090 5930 14110
rect 5950 14090 5960 14110
rect 5920 14035 5960 14090
rect 5920 14005 5925 14035
rect 5955 14005 5960 14035
rect 5920 13955 5960 14005
rect 5920 13925 5925 13955
rect 5955 13925 5960 13955
rect 5920 13875 5960 13925
rect 5920 13845 5925 13875
rect 5955 13845 5960 13875
rect 5920 13795 5960 13845
rect 5920 13765 5925 13795
rect 5955 13765 5960 13795
rect 5920 13715 5960 13765
rect 5920 13685 5925 13715
rect 5955 13685 5960 13715
rect 5920 13635 5960 13685
rect 5920 13605 5925 13635
rect 5955 13605 5960 13635
rect 5920 13555 5960 13605
rect 5920 13525 5925 13555
rect 5955 13525 5960 13555
rect 5920 13475 5960 13525
rect 5920 13445 5925 13475
rect 5955 13445 5960 13475
rect 5920 13390 5960 13445
rect 5920 13370 5930 13390
rect 5950 13370 5960 13390
rect 5920 13310 5960 13370
rect 5920 13290 5930 13310
rect 5950 13290 5960 13310
rect 5920 13230 5960 13290
rect 5920 13210 5930 13230
rect 5950 13210 5960 13230
rect 5920 13150 5960 13210
rect 5920 13130 5930 13150
rect 5950 13130 5960 13150
rect 5920 13075 5960 13130
rect 5920 13045 5925 13075
rect 5955 13045 5960 13075
rect 5920 12995 5960 13045
rect 5920 12965 5925 12995
rect 5955 12965 5960 12995
rect 5920 12915 5960 12965
rect 5920 12885 5925 12915
rect 5955 12885 5960 12915
rect 5920 12835 5960 12885
rect 5920 12805 5925 12835
rect 5955 12805 5960 12835
rect 5920 12755 5960 12805
rect 5920 12725 5925 12755
rect 5955 12725 5960 12755
rect 5920 12675 5960 12725
rect 5920 12645 5925 12675
rect 5955 12645 5960 12675
rect 5920 12595 5960 12645
rect 5920 12565 5925 12595
rect 5955 12565 5960 12595
rect 5920 12515 5960 12565
rect 5920 12485 5925 12515
rect 5955 12485 5960 12515
rect 5920 12430 5960 12485
rect 5920 12410 5930 12430
rect 5950 12410 5960 12430
rect 5920 12355 5960 12410
rect 5920 12325 5925 12355
rect 5955 12325 5960 12355
rect 5920 12275 5960 12325
rect 5920 12245 5925 12275
rect 5955 12245 5960 12275
rect 5920 12195 5960 12245
rect 5920 12165 5925 12195
rect 5955 12165 5960 12195
rect 5920 12115 5960 12165
rect 5920 12085 5925 12115
rect 5955 12085 5960 12115
rect 5920 12035 5960 12085
rect 5920 12005 5925 12035
rect 5955 12005 5960 12035
rect 5920 11955 5960 12005
rect 5920 11925 5925 11955
rect 5955 11925 5960 11955
rect 5920 11875 5960 11925
rect 5920 11845 5925 11875
rect 5955 11845 5960 11875
rect 5920 11795 5960 11845
rect 5920 11765 5925 11795
rect 5955 11765 5960 11795
rect 5920 11715 5960 11765
rect 5920 11685 5925 11715
rect 5955 11685 5960 11715
rect 5920 11635 5960 11685
rect 5920 11605 5925 11635
rect 5955 11605 5960 11635
rect 5920 11555 5960 11605
rect 5920 11525 5925 11555
rect 5955 11525 5960 11555
rect 5920 11475 5960 11525
rect 5920 11445 5925 11475
rect 5955 11445 5960 11475
rect 5920 11395 5960 11445
rect 5920 11365 5925 11395
rect 5955 11365 5960 11395
rect 5920 11315 5960 11365
rect 5920 11285 5925 11315
rect 5955 11285 5960 11315
rect 5920 11235 5960 11285
rect 5920 11205 5925 11235
rect 5955 11205 5960 11235
rect 5920 11155 5960 11205
rect 5920 11125 5925 11155
rect 5955 11125 5960 11155
rect 5920 11075 5960 11125
rect 5920 11045 5925 11075
rect 5955 11045 5960 11075
rect 5920 10990 5960 11045
rect 5920 10970 5930 10990
rect 5950 10970 5960 10990
rect 5920 10915 5960 10970
rect 5920 10885 5925 10915
rect 5955 10885 5960 10915
rect 5920 10835 5960 10885
rect 5920 10805 5925 10835
rect 5955 10805 5960 10835
rect 5920 10755 5960 10805
rect 5920 10725 5925 10755
rect 5955 10725 5960 10755
rect 5920 10675 5960 10725
rect 5920 10645 5925 10675
rect 5955 10645 5960 10675
rect 5920 10595 5960 10645
rect 5920 10565 5925 10595
rect 5955 10565 5960 10595
rect 5920 10515 5960 10565
rect 5920 10485 5925 10515
rect 5955 10485 5960 10515
rect 5920 10435 5960 10485
rect 5920 10405 5925 10435
rect 5955 10405 5960 10435
rect 5920 10355 5960 10405
rect 5920 10325 5925 10355
rect 5955 10325 5960 10355
rect 5920 10270 5960 10325
rect 5920 10250 5930 10270
rect 5950 10250 5960 10270
rect 5920 10190 5960 10250
rect 5920 10170 5930 10190
rect 5950 10170 5960 10190
rect 5920 10110 5960 10170
rect 5920 10090 5930 10110
rect 5950 10090 5960 10110
rect 5920 10030 5960 10090
rect 5920 10010 5930 10030
rect 5950 10010 5960 10030
rect 5920 9955 5960 10010
rect 5920 9925 5925 9955
rect 5955 9925 5960 9955
rect 5920 9875 5960 9925
rect 5920 9845 5925 9875
rect 5955 9845 5960 9875
rect 5920 9795 5960 9845
rect 5920 9765 5925 9795
rect 5955 9765 5960 9795
rect 5920 9715 5960 9765
rect 5920 9685 5925 9715
rect 5955 9685 5960 9715
rect 5920 9635 5960 9685
rect 5920 9605 5925 9635
rect 5955 9605 5960 9635
rect 5920 9555 5960 9605
rect 5920 9525 5925 9555
rect 5955 9525 5960 9555
rect 5920 9475 5960 9525
rect 5920 9445 5925 9475
rect 5955 9445 5960 9475
rect 5920 9395 5960 9445
rect 5920 9365 5925 9395
rect 5955 9365 5960 9395
rect 5920 9310 5960 9365
rect 5920 9290 5930 9310
rect 5950 9290 5960 9310
rect 5920 9230 5960 9290
rect 5920 9210 5930 9230
rect 5950 9210 5960 9230
rect 5920 9150 5960 9210
rect 5920 9130 5930 9150
rect 5950 9130 5960 9150
rect 5920 9070 5960 9130
rect 5920 9050 5930 9070
rect 5950 9050 5960 9070
rect 5920 8995 5960 9050
rect 5920 8965 5925 8995
rect 5955 8965 5960 8995
rect 5920 8915 5960 8965
rect 5920 8885 5925 8915
rect 5955 8885 5960 8915
rect 5920 8835 5960 8885
rect 5920 8805 5925 8835
rect 5955 8805 5960 8835
rect 5920 8755 5960 8805
rect 5920 8725 5925 8755
rect 5955 8725 5960 8755
rect 5920 8675 5960 8725
rect 5920 8645 5925 8675
rect 5955 8645 5960 8675
rect 5920 8595 5960 8645
rect 5920 8565 5925 8595
rect 5955 8565 5960 8595
rect 5920 8515 5960 8565
rect 5920 8485 5925 8515
rect 5955 8485 5960 8515
rect 5920 8435 5960 8485
rect 5920 8405 5925 8435
rect 5955 8405 5960 8435
rect 5920 8350 5960 8405
rect 5920 8330 5930 8350
rect 5950 8330 5960 8350
rect 5920 8275 5960 8330
rect 5920 8245 5925 8275
rect 5955 8245 5960 8275
rect 5920 8195 5960 8245
rect 5920 8165 5925 8195
rect 5955 8165 5960 8195
rect 5920 8115 5960 8165
rect 5920 8085 5925 8115
rect 5955 8085 5960 8115
rect 5920 8035 5960 8085
rect 5920 8005 5925 8035
rect 5955 8005 5960 8035
rect 5920 7955 5960 8005
rect 5920 7925 5925 7955
rect 5955 7925 5960 7955
rect 5920 7875 5960 7925
rect 5920 7845 5925 7875
rect 5955 7845 5960 7875
rect 5920 7795 5960 7845
rect 5920 7765 5925 7795
rect 5955 7765 5960 7795
rect 5920 7715 5960 7765
rect 5920 7685 5925 7715
rect 5955 7685 5960 7715
rect 5920 7635 5960 7685
rect 5920 7605 5925 7635
rect 5955 7605 5960 7635
rect 5920 7555 5960 7605
rect 5920 7525 5925 7555
rect 5955 7525 5960 7555
rect 5920 7475 5960 7525
rect 5920 7445 5925 7475
rect 5955 7445 5960 7475
rect 5920 7395 5960 7445
rect 5920 7365 5925 7395
rect 5955 7365 5960 7395
rect 5920 7315 5960 7365
rect 5920 7285 5925 7315
rect 5955 7285 5960 7315
rect 5920 7235 5960 7285
rect 5920 7205 5925 7235
rect 5955 7205 5960 7235
rect 5920 7155 5960 7205
rect 5920 7125 5925 7155
rect 5955 7125 5960 7155
rect 5920 7075 5960 7125
rect 5920 7045 5925 7075
rect 5955 7045 5960 7075
rect 5920 6995 5960 7045
rect 5920 6965 5925 6995
rect 5955 6965 5960 6995
rect 5920 6910 5960 6965
rect 5920 6890 5930 6910
rect 5950 6890 5960 6910
rect 5920 6835 5960 6890
rect 5920 6805 5925 6835
rect 5955 6805 5960 6835
rect 5920 6755 5960 6805
rect 5920 6725 5925 6755
rect 5955 6725 5960 6755
rect 5920 6675 5960 6725
rect 5920 6645 5925 6675
rect 5955 6645 5960 6675
rect 5920 6595 5960 6645
rect 5920 6565 5925 6595
rect 5955 6565 5960 6595
rect 5920 6515 5960 6565
rect 5920 6485 5925 6515
rect 5955 6485 5960 6515
rect 5920 6435 5960 6485
rect 5920 6405 5925 6435
rect 5955 6405 5960 6435
rect 5920 6355 5960 6405
rect 5920 6325 5925 6355
rect 5955 6325 5960 6355
rect 5920 6275 5960 6325
rect 5920 6245 5925 6275
rect 5955 6245 5960 6275
rect 5920 6190 5960 6245
rect 5920 6170 5930 6190
rect 5950 6170 5960 6190
rect 5920 6110 5960 6170
rect 5920 6090 5930 6110
rect 5950 6090 5960 6110
rect 5920 6030 5960 6090
rect 5920 6010 5930 6030
rect 5950 6010 5960 6030
rect 5920 5950 5960 6010
rect 5920 5930 5930 5950
rect 5950 5930 5960 5950
rect 5920 5875 5960 5930
rect 5920 5845 5925 5875
rect 5955 5845 5960 5875
rect 5920 5795 5960 5845
rect 5920 5765 5925 5795
rect 5955 5765 5960 5795
rect 5920 5715 5960 5765
rect 5920 5685 5925 5715
rect 5955 5685 5960 5715
rect 5920 5635 5960 5685
rect 5920 5605 5925 5635
rect 5955 5605 5960 5635
rect 5920 5555 5960 5605
rect 5920 5525 5925 5555
rect 5955 5525 5960 5555
rect 5920 5475 5960 5525
rect 5920 5445 5925 5475
rect 5955 5445 5960 5475
rect 5920 5395 5960 5445
rect 5920 5365 5925 5395
rect 5955 5365 5960 5395
rect 5920 5315 5960 5365
rect 5920 5285 5925 5315
rect 5955 5285 5960 5315
rect 5920 5235 5960 5285
rect 5920 5205 5925 5235
rect 5955 5205 5960 5235
rect 5920 5155 5960 5205
rect 5920 5125 5925 5155
rect 5955 5125 5960 5155
rect 5920 5075 5960 5125
rect 5920 5045 5925 5075
rect 5955 5045 5960 5075
rect 5920 4995 5960 5045
rect 5920 4965 5925 4995
rect 5955 4965 5960 4995
rect 5920 4915 5960 4965
rect 5920 4885 5925 4915
rect 5955 4885 5960 4915
rect 5920 4830 5960 4885
rect 5920 4810 5930 4830
rect 5950 4810 5960 4830
rect 5920 4755 5960 4810
rect 5920 4725 5925 4755
rect 5955 4725 5960 4755
rect 5920 4675 5960 4725
rect 5920 4645 5925 4675
rect 5955 4645 5960 4675
rect 5920 4590 5960 4645
rect 5920 4570 5930 4590
rect 5950 4570 5960 4590
rect 5920 4515 5960 4570
rect 5920 4485 5925 4515
rect 5955 4485 5960 4515
rect 5920 4435 5960 4485
rect 5920 4405 5925 4435
rect 5955 4405 5960 4435
rect 5920 4355 5960 4405
rect 5920 4325 5925 4355
rect 5955 4325 5960 4355
rect 5920 4275 5960 4325
rect 5920 4245 5925 4275
rect 5955 4245 5960 4275
rect 5920 4195 5960 4245
rect 5920 4165 5925 4195
rect 5955 4165 5960 4195
rect 5920 4115 5960 4165
rect 5920 4085 5925 4115
rect 5955 4085 5960 4115
rect 5920 4035 5960 4085
rect 5920 4005 5925 4035
rect 5955 4005 5960 4035
rect 5920 3955 5960 4005
rect 5920 3925 5925 3955
rect 5955 3925 5960 3955
rect 5920 3875 5960 3925
rect 5920 3845 5925 3875
rect 5955 3845 5960 3875
rect 5920 3790 5960 3845
rect 5920 3770 5930 3790
rect 5950 3770 5960 3790
rect 5920 3715 5960 3770
rect 5920 3685 5925 3715
rect 5955 3685 5960 3715
rect 5920 3635 5960 3685
rect 5920 3605 5925 3635
rect 5955 3605 5960 3635
rect 5920 3550 5960 3605
rect 5920 3530 5930 3550
rect 5950 3530 5960 3550
rect 5920 3475 5960 3530
rect 5920 3445 5925 3475
rect 5955 3445 5960 3475
rect 5920 3395 5960 3445
rect 5920 3365 5925 3395
rect 5955 3365 5960 3395
rect 5920 3310 5960 3365
rect 5920 3290 5930 3310
rect 5950 3290 5960 3310
rect 5920 3235 5960 3290
rect 5920 3205 5925 3235
rect 5955 3205 5960 3235
rect 5920 3155 5960 3205
rect 5920 3125 5925 3155
rect 5955 3125 5960 3155
rect 5920 3075 5960 3125
rect 5920 3045 5925 3075
rect 5955 3045 5960 3075
rect 5920 2995 5960 3045
rect 5920 2965 5925 2995
rect 5955 2965 5960 2995
rect 5920 2915 5960 2965
rect 5920 2885 5925 2915
rect 5955 2885 5960 2915
rect 5920 2835 5960 2885
rect 5920 2805 5925 2835
rect 5955 2805 5960 2835
rect 5920 2755 5960 2805
rect 5920 2725 5925 2755
rect 5955 2725 5960 2755
rect 5920 2675 5960 2725
rect 5920 2645 5925 2675
rect 5955 2645 5960 2675
rect 5920 2595 5960 2645
rect 5920 2565 5925 2595
rect 5955 2565 5960 2595
rect 5920 2515 5960 2565
rect 5920 2485 5925 2515
rect 5955 2485 5960 2515
rect 5920 2435 5960 2485
rect 5920 2405 5925 2435
rect 5955 2405 5960 2435
rect 5920 2355 5960 2405
rect 5920 2325 5925 2355
rect 5955 2325 5960 2355
rect 5920 2275 5960 2325
rect 5920 2245 5925 2275
rect 5955 2245 5960 2275
rect 5920 2195 5960 2245
rect 5920 2165 5925 2195
rect 5955 2165 5960 2195
rect 5920 2115 5960 2165
rect 5920 2085 5925 2115
rect 5955 2085 5960 2115
rect 5920 2035 5960 2085
rect 5920 2005 5925 2035
rect 5955 2005 5960 2035
rect 5920 1955 5960 2005
rect 5920 1925 5925 1955
rect 5955 1925 5960 1955
rect 5920 1870 5960 1925
rect 5920 1850 5930 1870
rect 5950 1850 5960 1870
rect 5920 1790 5960 1850
rect 5920 1770 5930 1790
rect 5950 1770 5960 1790
rect 5920 1715 5960 1770
rect 5920 1685 5925 1715
rect 5955 1685 5960 1715
rect 5920 1635 5960 1685
rect 5920 1605 5925 1635
rect 5955 1605 5960 1635
rect 5920 1555 5960 1605
rect 5920 1525 5925 1555
rect 5955 1525 5960 1555
rect 5920 1475 5960 1525
rect 5920 1445 5925 1475
rect 5955 1445 5960 1475
rect 5920 1395 5960 1445
rect 5920 1365 5925 1395
rect 5955 1365 5960 1395
rect 5920 1315 5960 1365
rect 5920 1285 5925 1315
rect 5955 1285 5960 1315
rect 5920 1235 5960 1285
rect 5920 1205 5925 1235
rect 5955 1205 5960 1235
rect 5920 1155 5960 1205
rect 5920 1125 5925 1155
rect 5955 1125 5960 1155
rect 5920 1075 5960 1125
rect 5920 1045 5925 1075
rect 5955 1045 5960 1075
rect 5920 995 5960 1045
rect 5920 965 5925 995
rect 5955 965 5960 995
rect 5920 910 5960 965
rect 5920 890 5930 910
rect 5950 890 5960 910
rect 5920 835 5960 890
rect 5920 805 5925 835
rect 5955 805 5960 835
rect 5920 755 5960 805
rect 5920 725 5925 755
rect 5955 725 5960 755
rect 5920 675 5960 725
rect 5920 645 5925 675
rect 5955 645 5960 675
rect 5920 595 5960 645
rect 5920 565 5925 595
rect 5955 565 5960 595
rect 5920 515 5960 565
rect 5920 485 5925 515
rect 5955 485 5960 515
rect 5920 430 5960 485
rect 5920 410 5930 430
rect 5950 410 5960 430
rect 5920 350 5960 410
rect 5920 330 5930 350
rect 5950 330 5960 350
rect 5920 275 5960 330
rect 5920 245 5925 275
rect 5955 245 5960 275
rect 5920 195 5960 245
rect 5920 165 5925 195
rect 5955 165 5960 195
rect 5920 115 5960 165
rect 5920 85 5925 115
rect 5955 85 5960 115
rect 5920 35 5960 85
rect 5920 5 5925 35
rect 5955 5 5960 35
rect 5920 0 5960 5
rect 6000 15715 6040 15720
rect 6000 15685 6005 15715
rect 6035 15685 6040 15715
rect 6000 15635 6040 15685
rect 6000 15605 6005 15635
rect 6035 15605 6040 15635
rect 6000 15555 6040 15605
rect 6000 15525 6005 15555
rect 6035 15525 6040 15555
rect 6000 15475 6040 15525
rect 6000 15445 6005 15475
rect 6035 15445 6040 15475
rect 6000 15395 6040 15445
rect 6000 15365 6005 15395
rect 6035 15365 6040 15395
rect 6000 15315 6040 15365
rect 6000 15285 6005 15315
rect 6035 15285 6040 15315
rect 6000 15235 6040 15285
rect 6000 15205 6005 15235
rect 6035 15205 6040 15235
rect 6000 15155 6040 15205
rect 6000 15125 6005 15155
rect 6035 15125 6040 15155
rect 6000 15070 6040 15125
rect 6000 15050 6010 15070
rect 6030 15050 6040 15070
rect 6000 14995 6040 15050
rect 6000 14965 6005 14995
rect 6035 14965 6040 14995
rect 6000 14915 6040 14965
rect 6000 14885 6005 14915
rect 6035 14885 6040 14915
rect 6000 14835 6040 14885
rect 6000 14805 6005 14835
rect 6035 14805 6040 14835
rect 6000 14755 6040 14805
rect 6000 14725 6005 14755
rect 6035 14725 6040 14755
rect 6000 14675 6040 14725
rect 6000 14645 6005 14675
rect 6035 14645 6040 14675
rect 6000 14595 6040 14645
rect 6000 14565 6005 14595
rect 6035 14565 6040 14595
rect 6000 14515 6040 14565
rect 6000 14485 6005 14515
rect 6035 14485 6040 14515
rect 6000 14435 6040 14485
rect 6000 14405 6005 14435
rect 6035 14405 6040 14435
rect 6000 14350 6040 14405
rect 6000 14330 6010 14350
rect 6030 14330 6040 14350
rect 6000 14270 6040 14330
rect 6000 14250 6010 14270
rect 6030 14250 6040 14270
rect 6000 14190 6040 14250
rect 6000 14170 6010 14190
rect 6030 14170 6040 14190
rect 6000 14110 6040 14170
rect 6000 14090 6010 14110
rect 6030 14090 6040 14110
rect 6000 14035 6040 14090
rect 6000 14005 6005 14035
rect 6035 14005 6040 14035
rect 6000 13955 6040 14005
rect 6000 13925 6005 13955
rect 6035 13925 6040 13955
rect 6000 13875 6040 13925
rect 6000 13845 6005 13875
rect 6035 13845 6040 13875
rect 6000 13795 6040 13845
rect 6000 13765 6005 13795
rect 6035 13765 6040 13795
rect 6000 13715 6040 13765
rect 6000 13685 6005 13715
rect 6035 13685 6040 13715
rect 6000 13635 6040 13685
rect 6000 13605 6005 13635
rect 6035 13605 6040 13635
rect 6000 13555 6040 13605
rect 6000 13525 6005 13555
rect 6035 13525 6040 13555
rect 6000 13475 6040 13525
rect 6000 13445 6005 13475
rect 6035 13445 6040 13475
rect 6000 13390 6040 13445
rect 6000 13370 6010 13390
rect 6030 13370 6040 13390
rect 6000 13310 6040 13370
rect 6000 13290 6010 13310
rect 6030 13290 6040 13310
rect 6000 13230 6040 13290
rect 6000 13210 6010 13230
rect 6030 13210 6040 13230
rect 6000 13150 6040 13210
rect 6000 13130 6010 13150
rect 6030 13130 6040 13150
rect 6000 13075 6040 13130
rect 6000 13045 6005 13075
rect 6035 13045 6040 13075
rect 6000 12995 6040 13045
rect 6000 12965 6005 12995
rect 6035 12965 6040 12995
rect 6000 12915 6040 12965
rect 6000 12885 6005 12915
rect 6035 12885 6040 12915
rect 6000 12835 6040 12885
rect 6000 12805 6005 12835
rect 6035 12805 6040 12835
rect 6000 12755 6040 12805
rect 6000 12725 6005 12755
rect 6035 12725 6040 12755
rect 6000 12675 6040 12725
rect 6000 12645 6005 12675
rect 6035 12645 6040 12675
rect 6000 12595 6040 12645
rect 6000 12565 6005 12595
rect 6035 12565 6040 12595
rect 6000 12515 6040 12565
rect 6000 12485 6005 12515
rect 6035 12485 6040 12515
rect 6000 12430 6040 12485
rect 6000 12410 6010 12430
rect 6030 12410 6040 12430
rect 6000 12355 6040 12410
rect 6000 12325 6005 12355
rect 6035 12325 6040 12355
rect 6000 12275 6040 12325
rect 6000 12245 6005 12275
rect 6035 12245 6040 12275
rect 6000 12195 6040 12245
rect 6000 12165 6005 12195
rect 6035 12165 6040 12195
rect 6000 12115 6040 12165
rect 6000 12085 6005 12115
rect 6035 12085 6040 12115
rect 6000 12035 6040 12085
rect 6000 12005 6005 12035
rect 6035 12005 6040 12035
rect 6000 11955 6040 12005
rect 6000 11925 6005 11955
rect 6035 11925 6040 11955
rect 6000 11875 6040 11925
rect 6000 11845 6005 11875
rect 6035 11845 6040 11875
rect 6000 11795 6040 11845
rect 6000 11765 6005 11795
rect 6035 11765 6040 11795
rect 6000 11715 6040 11765
rect 6000 11685 6005 11715
rect 6035 11685 6040 11715
rect 6000 11635 6040 11685
rect 6000 11605 6005 11635
rect 6035 11605 6040 11635
rect 6000 11555 6040 11605
rect 6000 11525 6005 11555
rect 6035 11525 6040 11555
rect 6000 11475 6040 11525
rect 6000 11445 6005 11475
rect 6035 11445 6040 11475
rect 6000 11395 6040 11445
rect 6000 11365 6005 11395
rect 6035 11365 6040 11395
rect 6000 11315 6040 11365
rect 6000 11285 6005 11315
rect 6035 11285 6040 11315
rect 6000 11235 6040 11285
rect 6000 11205 6005 11235
rect 6035 11205 6040 11235
rect 6000 11155 6040 11205
rect 6000 11125 6005 11155
rect 6035 11125 6040 11155
rect 6000 11075 6040 11125
rect 6000 11045 6005 11075
rect 6035 11045 6040 11075
rect 6000 10990 6040 11045
rect 6000 10970 6010 10990
rect 6030 10970 6040 10990
rect 6000 10915 6040 10970
rect 6000 10885 6005 10915
rect 6035 10885 6040 10915
rect 6000 10835 6040 10885
rect 6000 10805 6005 10835
rect 6035 10805 6040 10835
rect 6000 10755 6040 10805
rect 6000 10725 6005 10755
rect 6035 10725 6040 10755
rect 6000 10675 6040 10725
rect 6000 10645 6005 10675
rect 6035 10645 6040 10675
rect 6000 10595 6040 10645
rect 6000 10565 6005 10595
rect 6035 10565 6040 10595
rect 6000 10515 6040 10565
rect 6000 10485 6005 10515
rect 6035 10485 6040 10515
rect 6000 10435 6040 10485
rect 6000 10405 6005 10435
rect 6035 10405 6040 10435
rect 6000 10355 6040 10405
rect 6000 10325 6005 10355
rect 6035 10325 6040 10355
rect 6000 10270 6040 10325
rect 6000 10250 6010 10270
rect 6030 10250 6040 10270
rect 6000 10190 6040 10250
rect 6000 10170 6010 10190
rect 6030 10170 6040 10190
rect 6000 10110 6040 10170
rect 6000 10090 6010 10110
rect 6030 10090 6040 10110
rect 6000 10030 6040 10090
rect 6000 10010 6010 10030
rect 6030 10010 6040 10030
rect 6000 9955 6040 10010
rect 6000 9925 6005 9955
rect 6035 9925 6040 9955
rect 6000 9875 6040 9925
rect 6000 9845 6005 9875
rect 6035 9845 6040 9875
rect 6000 9795 6040 9845
rect 6000 9765 6005 9795
rect 6035 9765 6040 9795
rect 6000 9715 6040 9765
rect 6000 9685 6005 9715
rect 6035 9685 6040 9715
rect 6000 9635 6040 9685
rect 6000 9605 6005 9635
rect 6035 9605 6040 9635
rect 6000 9555 6040 9605
rect 6000 9525 6005 9555
rect 6035 9525 6040 9555
rect 6000 9475 6040 9525
rect 6000 9445 6005 9475
rect 6035 9445 6040 9475
rect 6000 9395 6040 9445
rect 6000 9365 6005 9395
rect 6035 9365 6040 9395
rect 6000 9310 6040 9365
rect 6000 9290 6010 9310
rect 6030 9290 6040 9310
rect 6000 9230 6040 9290
rect 6000 9210 6010 9230
rect 6030 9210 6040 9230
rect 6000 9150 6040 9210
rect 6000 9130 6010 9150
rect 6030 9130 6040 9150
rect 6000 9070 6040 9130
rect 6000 9050 6010 9070
rect 6030 9050 6040 9070
rect 6000 8995 6040 9050
rect 6000 8965 6005 8995
rect 6035 8965 6040 8995
rect 6000 8915 6040 8965
rect 6000 8885 6005 8915
rect 6035 8885 6040 8915
rect 6000 8835 6040 8885
rect 6000 8805 6005 8835
rect 6035 8805 6040 8835
rect 6000 8755 6040 8805
rect 6000 8725 6005 8755
rect 6035 8725 6040 8755
rect 6000 8675 6040 8725
rect 6000 8645 6005 8675
rect 6035 8645 6040 8675
rect 6000 8595 6040 8645
rect 6000 8565 6005 8595
rect 6035 8565 6040 8595
rect 6000 8515 6040 8565
rect 6000 8485 6005 8515
rect 6035 8485 6040 8515
rect 6000 8435 6040 8485
rect 6000 8405 6005 8435
rect 6035 8405 6040 8435
rect 6000 8350 6040 8405
rect 6000 8330 6010 8350
rect 6030 8330 6040 8350
rect 6000 8275 6040 8330
rect 6000 8245 6005 8275
rect 6035 8245 6040 8275
rect 6000 8195 6040 8245
rect 6000 8165 6005 8195
rect 6035 8165 6040 8195
rect 6000 8115 6040 8165
rect 6000 8085 6005 8115
rect 6035 8085 6040 8115
rect 6000 8035 6040 8085
rect 6000 8005 6005 8035
rect 6035 8005 6040 8035
rect 6000 7955 6040 8005
rect 6000 7925 6005 7955
rect 6035 7925 6040 7955
rect 6000 7875 6040 7925
rect 6000 7845 6005 7875
rect 6035 7845 6040 7875
rect 6000 7795 6040 7845
rect 6000 7765 6005 7795
rect 6035 7765 6040 7795
rect 6000 7715 6040 7765
rect 6000 7685 6005 7715
rect 6035 7685 6040 7715
rect 6000 7635 6040 7685
rect 6000 7605 6005 7635
rect 6035 7605 6040 7635
rect 6000 7555 6040 7605
rect 6000 7525 6005 7555
rect 6035 7525 6040 7555
rect 6000 7475 6040 7525
rect 6000 7445 6005 7475
rect 6035 7445 6040 7475
rect 6000 7395 6040 7445
rect 6000 7365 6005 7395
rect 6035 7365 6040 7395
rect 6000 7315 6040 7365
rect 6000 7285 6005 7315
rect 6035 7285 6040 7315
rect 6000 7235 6040 7285
rect 6000 7205 6005 7235
rect 6035 7205 6040 7235
rect 6000 7155 6040 7205
rect 6000 7125 6005 7155
rect 6035 7125 6040 7155
rect 6000 7075 6040 7125
rect 6000 7045 6005 7075
rect 6035 7045 6040 7075
rect 6000 6995 6040 7045
rect 6000 6965 6005 6995
rect 6035 6965 6040 6995
rect 6000 6910 6040 6965
rect 6000 6890 6010 6910
rect 6030 6890 6040 6910
rect 6000 6835 6040 6890
rect 6000 6805 6005 6835
rect 6035 6805 6040 6835
rect 6000 6755 6040 6805
rect 6000 6725 6005 6755
rect 6035 6725 6040 6755
rect 6000 6675 6040 6725
rect 6000 6645 6005 6675
rect 6035 6645 6040 6675
rect 6000 6595 6040 6645
rect 6000 6565 6005 6595
rect 6035 6565 6040 6595
rect 6000 6515 6040 6565
rect 6000 6485 6005 6515
rect 6035 6485 6040 6515
rect 6000 6435 6040 6485
rect 6000 6405 6005 6435
rect 6035 6405 6040 6435
rect 6000 6355 6040 6405
rect 6000 6325 6005 6355
rect 6035 6325 6040 6355
rect 6000 6275 6040 6325
rect 6000 6245 6005 6275
rect 6035 6245 6040 6275
rect 6000 6190 6040 6245
rect 6000 6170 6010 6190
rect 6030 6170 6040 6190
rect 6000 6110 6040 6170
rect 6000 6090 6010 6110
rect 6030 6090 6040 6110
rect 6000 6030 6040 6090
rect 6000 6010 6010 6030
rect 6030 6010 6040 6030
rect 6000 5950 6040 6010
rect 6000 5930 6010 5950
rect 6030 5930 6040 5950
rect 6000 5875 6040 5930
rect 6000 5845 6005 5875
rect 6035 5845 6040 5875
rect 6000 5795 6040 5845
rect 6000 5765 6005 5795
rect 6035 5765 6040 5795
rect 6000 5715 6040 5765
rect 6000 5685 6005 5715
rect 6035 5685 6040 5715
rect 6000 5635 6040 5685
rect 6000 5605 6005 5635
rect 6035 5605 6040 5635
rect 6000 5555 6040 5605
rect 6000 5525 6005 5555
rect 6035 5525 6040 5555
rect 6000 5475 6040 5525
rect 6000 5445 6005 5475
rect 6035 5445 6040 5475
rect 6000 5395 6040 5445
rect 6000 5365 6005 5395
rect 6035 5365 6040 5395
rect 6000 5315 6040 5365
rect 6000 5285 6005 5315
rect 6035 5285 6040 5315
rect 6000 5235 6040 5285
rect 6000 5205 6005 5235
rect 6035 5205 6040 5235
rect 6000 5155 6040 5205
rect 6000 5125 6005 5155
rect 6035 5125 6040 5155
rect 6000 5075 6040 5125
rect 6000 5045 6005 5075
rect 6035 5045 6040 5075
rect 6000 4995 6040 5045
rect 6000 4965 6005 4995
rect 6035 4965 6040 4995
rect 6000 4915 6040 4965
rect 6000 4885 6005 4915
rect 6035 4885 6040 4915
rect 6000 4830 6040 4885
rect 6000 4810 6010 4830
rect 6030 4810 6040 4830
rect 6000 4755 6040 4810
rect 6000 4725 6005 4755
rect 6035 4725 6040 4755
rect 6000 4675 6040 4725
rect 6000 4645 6005 4675
rect 6035 4645 6040 4675
rect 6000 4590 6040 4645
rect 6000 4570 6010 4590
rect 6030 4570 6040 4590
rect 6000 4515 6040 4570
rect 6000 4485 6005 4515
rect 6035 4485 6040 4515
rect 6000 4435 6040 4485
rect 6000 4405 6005 4435
rect 6035 4405 6040 4435
rect 6000 4355 6040 4405
rect 6000 4325 6005 4355
rect 6035 4325 6040 4355
rect 6000 4275 6040 4325
rect 6000 4245 6005 4275
rect 6035 4245 6040 4275
rect 6000 4195 6040 4245
rect 6000 4165 6005 4195
rect 6035 4165 6040 4195
rect 6000 4115 6040 4165
rect 6000 4085 6005 4115
rect 6035 4085 6040 4115
rect 6000 4035 6040 4085
rect 6000 4005 6005 4035
rect 6035 4005 6040 4035
rect 6000 3955 6040 4005
rect 6000 3925 6005 3955
rect 6035 3925 6040 3955
rect 6000 3875 6040 3925
rect 6000 3845 6005 3875
rect 6035 3845 6040 3875
rect 6000 3790 6040 3845
rect 6000 3770 6010 3790
rect 6030 3770 6040 3790
rect 6000 3715 6040 3770
rect 6000 3685 6005 3715
rect 6035 3685 6040 3715
rect 6000 3635 6040 3685
rect 6000 3605 6005 3635
rect 6035 3605 6040 3635
rect 6000 3550 6040 3605
rect 6000 3530 6010 3550
rect 6030 3530 6040 3550
rect 6000 3475 6040 3530
rect 6000 3445 6005 3475
rect 6035 3445 6040 3475
rect 6000 3395 6040 3445
rect 6000 3365 6005 3395
rect 6035 3365 6040 3395
rect 6000 3310 6040 3365
rect 6000 3290 6010 3310
rect 6030 3290 6040 3310
rect 6000 3235 6040 3290
rect 6000 3205 6005 3235
rect 6035 3205 6040 3235
rect 6000 3155 6040 3205
rect 6000 3125 6005 3155
rect 6035 3125 6040 3155
rect 6000 3075 6040 3125
rect 6000 3045 6005 3075
rect 6035 3045 6040 3075
rect 6000 2995 6040 3045
rect 6000 2965 6005 2995
rect 6035 2965 6040 2995
rect 6000 2915 6040 2965
rect 6000 2885 6005 2915
rect 6035 2885 6040 2915
rect 6000 2835 6040 2885
rect 6000 2805 6005 2835
rect 6035 2805 6040 2835
rect 6000 2755 6040 2805
rect 6000 2725 6005 2755
rect 6035 2725 6040 2755
rect 6000 2675 6040 2725
rect 6000 2645 6005 2675
rect 6035 2645 6040 2675
rect 6000 2595 6040 2645
rect 6000 2565 6005 2595
rect 6035 2565 6040 2595
rect 6000 2515 6040 2565
rect 6000 2485 6005 2515
rect 6035 2485 6040 2515
rect 6000 2435 6040 2485
rect 6000 2405 6005 2435
rect 6035 2405 6040 2435
rect 6000 2355 6040 2405
rect 6000 2325 6005 2355
rect 6035 2325 6040 2355
rect 6000 2275 6040 2325
rect 6000 2245 6005 2275
rect 6035 2245 6040 2275
rect 6000 2195 6040 2245
rect 6000 2165 6005 2195
rect 6035 2165 6040 2195
rect 6000 2115 6040 2165
rect 6000 2085 6005 2115
rect 6035 2085 6040 2115
rect 6000 2035 6040 2085
rect 6000 2005 6005 2035
rect 6035 2005 6040 2035
rect 6000 1955 6040 2005
rect 6000 1925 6005 1955
rect 6035 1925 6040 1955
rect 6000 1870 6040 1925
rect 6000 1850 6010 1870
rect 6030 1850 6040 1870
rect 6000 1790 6040 1850
rect 6000 1770 6010 1790
rect 6030 1770 6040 1790
rect 6000 1715 6040 1770
rect 6000 1685 6005 1715
rect 6035 1685 6040 1715
rect 6000 1635 6040 1685
rect 6000 1605 6005 1635
rect 6035 1605 6040 1635
rect 6000 1555 6040 1605
rect 6000 1525 6005 1555
rect 6035 1525 6040 1555
rect 6000 1475 6040 1525
rect 6000 1445 6005 1475
rect 6035 1445 6040 1475
rect 6000 1395 6040 1445
rect 6000 1365 6005 1395
rect 6035 1365 6040 1395
rect 6000 1315 6040 1365
rect 6000 1285 6005 1315
rect 6035 1285 6040 1315
rect 6000 1235 6040 1285
rect 6000 1205 6005 1235
rect 6035 1205 6040 1235
rect 6000 1155 6040 1205
rect 6000 1125 6005 1155
rect 6035 1125 6040 1155
rect 6000 1075 6040 1125
rect 6000 1045 6005 1075
rect 6035 1045 6040 1075
rect 6000 995 6040 1045
rect 6000 965 6005 995
rect 6035 965 6040 995
rect 6000 910 6040 965
rect 6000 890 6010 910
rect 6030 890 6040 910
rect 6000 835 6040 890
rect 6000 805 6005 835
rect 6035 805 6040 835
rect 6000 755 6040 805
rect 6000 725 6005 755
rect 6035 725 6040 755
rect 6000 675 6040 725
rect 6000 645 6005 675
rect 6035 645 6040 675
rect 6000 595 6040 645
rect 6000 565 6005 595
rect 6035 565 6040 595
rect 6000 515 6040 565
rect 6000 485 6005 515
rect 6035 485 6040 515
rect 6000 430 6040 485
rect 6000 410 6010 430
rect 6030 410 6040 430
rect 6000 350 6040 410
rect 6000 330 6010 350
rect 6030 330 6040 350
rect 6000 275 6040 330
rect 6000 245 6005 275
rect 6035 245 6040 275
rect 6000 195 6040 245
rect 6000 165 6005 195
rect 6035 165 6040 195
rect 6000 115 6040 165
rect 6000 85 6005 115
rect 6035 85 6040 115
rect 6000 35 6040 85
rect 6000 5 6005 35
rect 6035 5 6040 35
rect 6000 0 6040 5
rect 6080 15710 6120 15720
rect 6080 15690 6090 15710
rect 6110 15690 6120 15710
rect 6080 15630 6120 15690
rect 6080 15610 6090 15630
rect 6110 15610 6120 15630
rect 6080 15550 6120 15610
rect 6080 15530 6090 15550
rect 6110 15530 6120 15550
rect 6080 15470 6120 15530
rect 6080 15450 6090 15470
rect 6110 15450 6120 15470
rect 6080 15390 6120 15450
rect 6080 15370 6090 15390
rect 6110 15370 6120 15390
rect 6080 15310 6120 15370
rect 6080 15290 6090 15310
rect 6110 15290 6120 15310
rect 6080 15230 6120 15290
rect 6080 15210 6090 15230
rect 6110 15210 6120 15230
rect 6080 15150 6120 15210
rect 6080 15130 6090 15150
rect 6110 15130 6120 15150
rect 6080 15070 6120 15130
rect 6080 15050 6090 15070
rect 6110 15050 6120 15070
rect 6080 14990 6120 15050
rect 6080 14970 6090 14990
rect 6110 14970 6120 14990
rect 6080 14910 6120 14970
rect 6080 14890 6090 14910
rect 6110 14890 6120 14910
rect 6080 14830 6120 14890
rect 6080 14810 6090 14830
rect 6110 14810 6120 14830
rect 6080 14750 6120 14810
rect 6080 14730 6090 14750
rect 6110 14730 6120 14750
rect 6080 14670 6120 14730
rect 6080 14650 6090 14670
rect 6110 14650 6120 14670
rect 6080 14590 6120 14650
rect 6080 14570 6090 14590
rect 6110 14570 6120 14590
rect 6080 14510 6120 14570
rect 6080 14490 6090 14510
rect 6110 14490 6120 14510
rect 6080 14430 6120 14490
rect 6080 14410 6090 14430
rect 6110 14410 6120 14430
rect 6080 14350 6120 14410
rect 6080 14330 6090 14350
rect 6110 14330 6120 14350
rect 6080 14270 6120 14330
rect 6080 14250 6090 14270
rect 6110 14250 6120 14270
rect 6080 14190 6120 14250
rect 6080 14170 6090 14190
rect 6110 14170 6120 14190
rect 6080 14110 6120 14170
rect 6080 14090 6090 14110
rect 6110 14090 6120 14110
rect 6080 14030 6120 14090
rect 6080 14010 6090 14030
rect 6110 14010 6120 14030
rect 6080 13950 6120 14010
rect 6080 13930 6090 13950
rect 6110 13930 6120 13950
rect 6080 13870 6120 13930
rect 6080 13850 6090 13870
rect 6110 13850 6120 13870
rect 6080 13790 6120 13850
rect 6080 13770 6090 13790
rect 6110 13770 6120 13790
rect 6080 13710 6120 13770
rect 6080 13690 6090 13710
rect 6110 13690 6120 13710
rect 6080 13630 6120 13690
rect 6080 13610 6090 13630
rect 6110 13610 6120 13630
rect 6080 13550 6120 13610
rect 6080 13530 6090 13550
rect 6110 13530 6120 13550
rect 6080 13470 6120 13530
rect 6080 13450 6090 13470
rect 6110 13450 6120 13470
rect 6080 13390 6120 13450
rect 6080 13370 6090 13390
rect 6110 13370 6120 13390
rect 6080 13310 6120 13370
rect 6080 13290 6090 13310
rect 6110 13290 6120 13310
rect 6080 13230 6120 13290
rect 6080 13210 6090 13230
rect 6110 13210 6120 13230
rect 6080 13150 6120 13210
rect 6080 13130 6090 13150
rect 6110 13130 6120 13150
rect 6080 13070 6120 13130
rect 6080 13050 6090 13070
rect 6110 13050 6120 13070
rect 6080 12990 6120 13050
rect 6080 12970 6090 12990
rect 6110 12970 6120 12990
rect 6080 12910 6120 12970
rect 6080 12890 6090 12910
rect 6110 12890 6120 12910
rect 6080 12830 6120 12890
rect 6080 12810 6090 12830
rect 6110 12810 6120 12830
rect 6080 12750 6120 12810
rect 6080 12730 6090 12750
rect 6110 12730 6120 12750
rect 6080 12670 6120 12730
rect 6080 12650 6090 12670
rect 6110 12650 6120 12670
rect 6080 12590 6120 12650
rect 6080 12570 6090 12590
rect 6110 12570 6120 12590
rect 6080 12510 6120 12570
rect 6080 12490 6090 12510
rect 6110 12490 6120 12510
rect 6080 12430 6120 12490
rect 6080 12410 6090 12430
rect 6110 12410 6120 12430
rect 6080 12350 6120 12410
rect 6080 12330 6090 12350
rect 6110 12330 6120 12350
rect 6080 12270 6120 12330
rect 6080 12250 6090 12270
rect 6110 12250 6120 12270
rect 6080 12190 6120 12250
rect 6080 12170 6090 12190
rect 6110 12170 6120 12190
rect 6080 12110 6120 12170
rect 6080 12090 6090 12110
rect 6110 12090 6120 12110
rect 6080 12030 6120 12090
rect 6080 12010 6090 12030
rect 6110 12010 6120 12030
rect 6080 11950 6120 12010
rect 6080 11930 6090 11950
rect 6110 11930 6120 11950
rect 6080 11870 6120 11930
rect 6080 11850 6090 11870
rect 6110 11850 6120 11870
rect 6080 11790 6120 11850
rect 6080 11770 6090 11790
rect 6110 11770 6120 11790
rect 6080 11710 6120 11770
rect 6080 11690 6090 11710
rect 6110 11690 6120 11710
rect 6080 11630 6120 11690
rect 6080 11610 6090 11630
rect 6110 11610 6120 11630
rect 6080 11550 6120 11610
rect 6080 11530 6090 11550
rect 6110 11530 6120 11550
rect 6080 11470 6120 11530
rect 6080 11450 6090 11470
rect 6110 11450 6120 11470
rect 6080 11390 6120 11450
rect 6080 11370 6090 11390
rect 6110 11370 6120 11390
rect 6080 11310 6120 11370
rect 6080 11290 6090 11310
rect 6110 11290 6120 11310
rect 6080 11230 6120 11290
rect 6080 11210 6090 11230
rect 6110 11210 6120 11230
rect 6080 11150 6120 11210
rect 6080 11130 6090 11150
rect 6110 11130 6120 11150
rect 6080 11070 6120 11130
rect 6080 11050 6090 11070
rect 6110 11050 6120 11070
rect 6080 10990 6120 11050
rect 6080 10970 6090 10990
rect 6110 10970 6120 10990
rect 6080 10910 6120 10970
rect 6080 10890 6090 10910
rect 6110 10890 6120 10910
rect 6080 10830 6120 10890
rect 6080 10810 6090 10830
rect 6110 10810 6120 10830
rect 6080 10750 6120 10810
rect 6080 10730 6090 10750
rect 6110 10730 6120 10750
rect 6080 10670 6120 10730
rect 6080 10650 6090 10670
rect 6110 10650 6120 10670
rect 6080 10590 6120 10650
rect 6080 10570 6090 10590
rect 6110 10570 6120 10590
rect 6080 10510 6120 10570
rect 6080 10490 6090 10510
rect 6110 10490 6120 10510
rect 6080 10430 6120 10490
rect 6080 10410 6090 10430
rect 6110 10410 6120 10430
rect 6080 10350 6120 10410
rect 6080 10330 6090 10350
rect 6110 10330 6120 10350
rect 6080 10270 6120 10330
rect 6080 10250 6090 10270
rect 6110 10250 6120 10270
rect 6080 10190 6120 10250
rect 6080 10170 6090 10190
rect 6110 10170 6120 10190
rect 6080 10110 6120 10170
rect 6080 10090 6090 10110
rect 6110 10090 6120 10110
rect 6080 10030 6120 10090
rect 6080 10010 6090 10030
rect 6110 10010 6120 10030
rect 6080 9950 6120 10010
rect 6080 9930 6090 9950
rect 6110 9930 6120 9950
rect 6080 9870 6120 9930
rect 6080 9850 6090 9870
rect 6110 9850 6120 9870
rect 6080 9790 6120 9850
rect 6080 9770 6090 9790
rect 6110 9770 6120 9790
rect 6080 9710 6120 9770
rect 6080 9690 6090 9710
rect 6110 9690 6120 9710
rect 6080 9630 6120 9690
rect 6080 9610 6090 9630
rect 6110 9610 6120 9630
rect 6080 9550 6120 9610
rect 6080 9530 6090 9550
rect 6110 9530 6120 9550
rect 6080 9470 6120 9530
rect 6080 9450 6090 9470
rect 6110 9450 6120 9470
rect 6080 9390 6120 9450
rect 6080 9370 6090 9390
rect 6110 9370 6120 9390
rect 6080 9310 6120 9370
rect 6080 9290 6090 9310
rect 6110 9290 6120 9310
rect 6080 9230 6120 9290
rect 6080 9210 6090 9230
rect 6110 9210 6120 9230
rect 6080 9150 6120 9210
rect 6080 9130 6090 9150
rect 6110 9130 6120 9150
rect 6080 9070 6120 9130
rect 6080 9050 6090 9070
rect 6110 9050 6120 9070
rect 6080 8990 6120 9050
rect 6080 8970 6090 8990
rect 6110 8970 6120 8990
rect 6080 8910 6120 8970
rect 6080 8890 6090 8910
rect 6110 8890 6120 8910
rect 6080 8830 6120 8890
rect 6080 8810 6090 8830
rect 6110 8810 6120 8830
rect 6080 8750 6120 8810
rect 6080 8730 6090 8750
rect 6110 8730 6120 8750
rect 6080 8670 6120 8730
rect 6080 8650 6090 8670
rect 6110 8650 6120 8670
rect 6080 8590 6120 8650
rect 6080 8570 6090 8590
rect 6110 8570 6120 8590
rect 6080 8510 6120 8570
rect 6080 8490 6090 8510
rect 6110 8490 6120 8510
rect 6080 8430 6120 8490
rect 6080 8410 6090 8430
rect 6110 8410 6120 8430
rect 6080 8350 6120 8410
rect 6080 8330 6090 8350
rect 6110 8330 6120 8350
rect 6080 8270 6120 8330
rect 6080 8250 6090 8270
rect 6110 8250 6120 8270
rect 6080 8190 6120 8250
rect 6080 8170 6090 8190
rect 6110 8170 6120 8190
rect 6080 8110 6120 8170
rect 6080 8090 6090 8110
rect 6110 8090 6120 8110
rect 6080 8030 6120 8090
rect 6080 8010 6090 8030
rect 6110 8010 6120 8030
rect 6080 7950 6120 8010
rect 6080 7930 6090 7950
rect 6110 7930 6120 7950
rect 6080 7870 6120 7930
rect 6080 7850 6090 7870
rect 6110 7850 6120 7870
rect 6080 7790 6120 7850
rect 6080 7770 6090 7790
rect 6110 7770 6120 7790
rect 6080 7710 6120 7770
rect 6080 7690 6090 7710
rect 6110 7690 6120 7710
rect 6080 7630 6120 7690
rect 6080 7610 6090 7630
rect 6110 7610 6120 7630
rect 6080 7550 6120 7610
rect 6080 7530 6090 7550
rect 6110 7530 6120 7550
rect 6080 7470 6120 7530
rect 6080 7450 6090 7470
rect 6110 7450 6120 7470
rect 6080 7390 6120 7450
rect 6080 7370 6090 7390
rect 6110 7370 6120 7390
rect 6080 7310 6120 7370
rect 6080 7290 6090 7310
rect 6110 7290 6120 7310
rect 6080 7230 6120 7290
rect 6080 7210 6090 7230
rect 6110 7210 6120 7230
rect 6080 7150 6120 7210
rect 6080 7130 6090 7150
rect 6110 7130 6120 7150
rect 6080 7070 6120 7130
rect 6080 7050 6090 7070
rect 6110 7050 6120 7070
rect 6080 6990 6120 7050
rect 6080 6970 6090 6990
rect 6110 6970 6120 6990
rect 6080 6910 6120 6970
rect 6080 6890 6090 6910
rect 6110 6890 6120 6910
rect 6080 6830 6120 6890
rect 6080 6810 6090 6830
rect 6110 6810 6120 6830
rect 6080 6750 6120 6810
rect 6080 6730 6090 6750
rect 6110 6730 6120 6750
rect 6080 6670 6120 6730
rect 6080 6650 6090 6670
rect 6110 6650 6120 6670
rect 6080 6590 6120 6650
rect 6080 6570 6090 6590
rect 6110 6570 6120 6590
rect 6080 6510 6120 6570
rect 6080 6490 6090 6510
rect 6110 6490 6120 6510
rect 6080 6430 6120 6490
rect 6080 6410 6090 6430
rect 6110 6410 6120 6430
rect 6080 6350 6120 6410
rect 6080 6330 6090 6350
rect 6110 6330 6120 6350
rect 6080 6270 6120 6330
rect 6080 6250 6090 6270
rect 6110 6250 6120 6270
rect 6080 6190 6120 6250
rect 6080 6170 6090 6190
rect 6110 6170 6120 6190
rect 6080 6110 6120 6170
rect 6080 6090 6090 6110
rect 6110 6090 6120 6110
rect 6080 6030 6120 6090
rect 6080 6010 6090 6030
rect 6110 6010 6120 6030
rect 6080 5950 6120 6010
rect 6080 5930 6090 5950
rect 6110 5930 6120 5950
rect 6080 5870 6120 5930
rect 6080 5850 6090 5870
rect 6110 5850 6120 5870
rect 6080 5790 6120 5850
rect 6080 5770 6090 5790
rect 6110 5770 6120 5790
rect 6080 5710 6120 5770
rect 6080 5690 6090 5710
rect 6110 5690 6120 5710
rect 6080 5630 6120 5690
rect 6080 5610 6090 5630
rect 6110 5610 6120 5630
rect 6080 5550 6120 5610
rect 6080 5530 6090 5550
rect 6110 5530 6120 5550
rect 6080 5470 6120 5530
rect 6080 5450 6090 5470
rect 6110 5450 6120 5470
rect 6080 5390 6120 5450
rect 6080 5370 6090 5390
rect 6110 5370 6120 5390
rect 6080 5310 6120 5370
rect 6080 5290 6090 5310
rect 6110 5290 6120 5310
rect 6080 5230 6120 5290
rect 6080 5210 6090 5230
rect 6110 5210 6120 5230
rect 6080 5150 6120 5210
rect 6080 5130 6090 5150
rect 6110 5130 6120 5150
rect 6080 5070 6120 5130
rect 6080 5050 6090 5070
rect 6110 5050 6120 5070
rect 6080 4990 6120 5050
rect 6080 4970 6090 4990
rect 6110 4970 6120 4990
rect 6080 4910 6120 4970
rect 6080 4890 6090 4910
rect 6110 4890 6120 4910
rect 6080 4830 6120 4890
rect 6080 4810 6090 4830
rect 6110 4810 6120 4830
rect 6080 4750 6120 4810
rect 6080 4730 6090 4750
rect 6110 4730 6120 4750
rect 6080 4670 6120 4730
rect 6080 4650 6090 4670
rect 6110 4650 6120 4670
rect 6080 4590 6120 4650
rect 6080 4570 6090 4590
rect 6110 4570 6120 4590
rect 6080 4510 6120 4570
rect 6080 4490 6090 4510
rect 6110 4490 6120 4510
rect 6080 4430 6120 4490
rect 6080 4410 6090 4430
rect 6110 4410 6120 4430
rect 6080 4350 6120 4410
rect 6080 4330 6090 4350
rect 6110 4330 6120 4350
rect 6080 4270 6120 4330
rect 6080 4250 6090 4270
rect 6110 4250 6120 4270
rect 6080 4190 6120 4250
rect 6080 4170 6090 4190
rect 6110 4170 6120 4190
rect 6080 4110 6120 4170
rect 6080 4090 6090 4110
rect 6110 4090 6120 4110
rect 6080 4030 6120 4090
rect 6080 4010 6090 4030
rect 6110 4010 6120 4030
rect 6080 3950 6120 4010
rect 6080 3930 6090 3950
rect 6110 3930 6120 3950
rect 6080 3870 6120 3930
rect 6080 3850 6090 3870
rect 6110 3850 6120 3870
rect 6080 3790 6120 3850
rect 6080 3770 6090 3790
rect 6110 3770 6120 3790
rect 6080 3710 6120 3770
rect 6080 3690 6090 3710
rect 6110 3690 6120 3710
rect 6080 3630 6120 3690
rect 6080 3610 6090 3630
rect 6110 3610 6120 3630
rect 6080 3550 6120 3610
rect 6080 3530 6090 3550
rect 6110 3530 6120 3550
rect 6080 3470 6120 3530
rect 6080 3450 6090 3470
rect 6110 3450 6120 3470
rect 6080 3390 6120 3450
rect 6080 3370 6090 3390
rect 6110 3370 6120 3390
rect 6080 3310 6120 3370
rect 6080 3290 6090 3310
rect 6110 3290 6120 3310
rect 6080 3230 6120 3290
rect 6080 3210 6090 3230
rect 6110 3210 6120 3230
rect 6080 3150 6120 3210
rect 6080 3130 6090 3150
rect 6110 3130 6120 3150
rect 6080 3070 6120 3130
rect 6080 3050 6090 3070
rect 6110 3050 6120 3070
rect 6080 2990 6120 3050
rect 6080 2970 6090 2990
rect 6110 2970 6120 2990
rect 6080 2910 6120 2970
rect 6080 2890 6090 2910
rect 6110 2890 6120 2910
rect 6080 2830 6120 2890
rect 6080 2810 6090 2830
rect 6110 2810 6120 2830
rect 6080 2750 6120 2810
rect 6080 2730 6090 2750
rect 6110 2730 6120 2750
rect 6080 2670 6120 2730
rect 6080 2650 6090 2670
rect 6110 2650 6120 2670
rect 6080 2590 6120 2650
rect 6080 2570 6090 2590
rect 6110 2570 6120 2590
rect 6080 2510 6120 2570
rect 6080 2490 6090 2510
rect 6110 2490 6120 2510
rect 6080 2430 6120 2490
rect 6080 2410 6090 2430
rect 6110 2410 6120 2430
rect 6080 2350 6120 2410
rect 6080 2330 6090 2350
rect 6110 2330 6120 2350
rect 6080 2270 6120 2330
rect 6080 2250 6090 2270
rect 6110 2250 6120 2270
rect 6080 2190 6120 2250
rect 6080 2170 6090 2190
rect 6110 2170 6120 2190
rect 6080 2110 6120 2170
rect 6080 2090 6090 2110
rect 6110 2090 6120 2110
rect 6080 2030 6120 2090
rect 6080 2010 6090 2030
rect 6110 2010 6120 2030
rect 6080 1950 6120 2010
rect 6080 1930 6090 1950
rect 6110 1930 6120 1950
rect 6080 1870 6120 1930
rect 6080 1850 6090 1870
rect 6110 1850 6120 1870
rect 6080 1790 6120 1850
rect 6080 1770 6090 1790
rect 6110 1770 6120 1790
rect 6080 1710 6120 1770
rect 6080 1690 6090 1710
rect 6110 1690 6120 1710
rect 6080 1630 6120 1690
rect 6080 1610 6090 1630
rect 6110 1610 6120 1630
rect 6080 1550 6120 1610
rect 6080 1530 6090 1550
rect 6110 1530 6120 1550
rect 6080 1470 6120 1530
rect 6080 1450 6090 1470
rect 6110 1450 6120 1470
rect 6080 1390 6120 1450
rect 6080 1370 6090 1390
rect 6110 1370 6120 1390
rect 6080 1310 6120 1370
rect 6080 1290 6090 1310
rect 6110 1290 6120 1310
rect 6080 1230 6120 1290
rect 6080 1210 6090 1230
rect 6110 1210 6120 1230
rect 6080 1150 6120 1210
rect 6080 1130 6090 1150
rect 6110 1130 6120 1150
rect 6080 1070 6120 1130
rect 6080 1050 6090 1070
rect 6110 1050 6120 1070
rect 6080 990 6120 1050
rect 6080 970 6090 990
rect 6110 970 6120 990
rect 6080 910 6120 970
rect 6080 890 6090 910
rect 6110 890 6120 910
rect 6080 830 6120 890
rect 6080 810 6090 830
rect 6110 810 6120 830
rect 6080 750 6120 810
rect 6080 730 6090 750
rect 6110 730 6120 750
rect 6080 670 6120 730
rect 6080 650 6090 670
rect 6110 650 6120 670
rect 6080 590 6120 650
rect 6080 570 6090 590
rect 6110 570 6120 590
rect 6080 510 6120 570
rect 6080 490 6090 510
rect 6110 490 6120 510
rect 6080 430 6120 490
rect 6080 410 6090 430
rect 6110 410 6120 430
rect 6080 350 6120 410
rect 6080 330 6090 350
rect 6110 330 6120 350
rect 6080 270 6120 330
rect 6080 250 6090 270
rect 6110 250 6120 270
rect 6080 190 6120 250
rect 6080 170 6090 190
rect 6110 170 6120 190
rect 6080 110 6120 170
rect 6080 90 6090 110
rect 6110 90 6120 110
rect 6080 30 6120 90
rect 6080 10 6090 30
rect 6110 10 6120 30
rect 6080 0 6120 10
rect 6160 15715 6200 15720
rect 6160 15685 6165 15715
rect 6195 15685 6200 15715
rect 6160 15635 6200 15685
rect 6160 15605 6165 15635
rect 6195 15605 6200 15635
rect 6160 15555 6200 15605
rect 6160 15525 6165 15555
rect 6195 15525 6200 15555
rect 6160 15475 6200 15525
rect 6160 15445 6165 15475
rect 6195 15445 6200 15475
rect 6160 15395 6200 15445
rect 6160 15365 6165 15395
rect 6195 15365 6200 15395
rect 6160 15315 6200 15365
rect 6160 15285 6165 15315
rect 6195 15285 6200 15315
rect 6160 15235 6200 15285
rect 6160 15205 6165 15235
rect 6195 15205 6200 15235
rect 6160 15155 6200 15205
rect 6160 15125 6165 15155
rect 6195 15125 6200 15155
rect 6160 15070 6200 15125
rect 6160 15050 6170 15070
rect 6190 15050 6200 15070
rect 6160 14995 6200 15050
rect 6160 14965 6165 14995
rect 6195 14965 6200 14995
rect 6160 14915 6200 14965
rect 6160 14885 6165 14915
rect 6195 14885 6200 14915
rect 6160 14835 6200 14885
rect 6160 14805 6165 14835
rect 6195 14805 6200 14835
rect 6160 14755 6200 14805
rect 6160 14725 6165 14755
rect 6195 14725 6200 14755
rect 6160 14675 6200 14725
rect 6160 14645 6165 14675
rect 6195 14645 6200 14675
rect 6160 14595 6200 14645
rect 6160 14565 6165 14595
rect 6195 14565 6200 14595
rect 6160 14515 6200 14565
rect 6160 14485 6165 14515
rect 6195 14485 6200 14515
rect 6160 14435 6200 14485
rect 6160 14405 6165 14435
rect 6195 14405 6200 14435
rect 6160 14350 6200 14405
rect 6160 14330 6170 14350
rect 6190 14330 6200 14350
rect 6160 14270 6200 14330
rect 6160 14250 6170 14270
rect 6190 14250 6200 14270
rect 6160 14190 6200 14250
rect 6160 14170 6170 14190
rect 6190 14170 6200 14190
rect 6160 14110 6200 14170
rect 6160 14090 6170 14110
rect 6190 14090 6200 14110
rect 6160 14035 6200 14090
rect 6160 14005 6165 14035
rect 6195 14005 6200 14035
rect 6160 13955 6200 14005
rect 6160 13925 6165 13955
rect 6195 13925 6200 13955
rect 6160 13875 6200 13925
rect 6160 13845 6165 13875
rect 6195 13845 6200 13875
rect 6160 13795 6200 13845
rect 6160 13765 6165 13795
rect 6195 13765 6200 13795
rect 6160 13715 6200 13765
rect 6160 13685 6165 13715
rect 6195 13685 6200 13715
rect 6160 13635 6200 13685
rect 6160 13605 6165 13635
rect 6195 13605 6200 13635
rect 6160 13555 6200 13605
rect 6160 13525 6165 13555
rect 6195 13525 6200 13555
rect 6160 13475 6200 13525
rect 6160 13445 6165 13475
rect 6195 13445 6200 13475
rect 6160 13390 6200 13445
rect 6160 13370 6170 13390
rect 6190 13370 6200 13390
rect 6160 13310 6200 13370
rect 6160 13290 6170 13310
rect 6190 13290 6200 13310
rect 6160 13230 6200 13290
rect 6160 13210 6170 13230
rect 6190 13210 6200 13230
rect 6160 13150 6200 13210
rect 6160 13130 6170 13150
rect 6190 13130 6200 13150
rect 6160 13075 6200 13130
rect 6160 13045 6165 13075
rect 6195 13045 6200 13075
rect 6160 12995 6200 13045
rect 6160 12965 6165 12995
rect 6195 12965 6200 12995
rect 6160 12915 6200 12965
rect 6160 12885 6165 12915
rect 6195 12885 6200 12915
rect 6160 12835 6200 12885
rect 6160 12805 6165 12835
rect 6195 12805 6200 12835
rect 6160 12755 6200 12805
rect 6160 12725 6165 12755
rect 6195 12725 6200 12755
rect 6160 12675 6200 12725
rect 6160 12645 6165 12675
rect 6195 12645 6200 12675
rect 6160 12595 6200 12645
rect 6160 12565 6165 12595
rect 6195 12565 6200 12595
rect 6160 12515 6200 12565
rect 6160 12485 6165 12515
rect 6195 12485 6200 12515
rect 6160 12430 6200 12485
rect 6160 12410 6170 12430
rect 6190 12410 6200 12430
rect 6160 12355 6200 12410
rect 6160 12325 6165 12355
rect 6195 12325 6200 12355
rect 6160 12275 6200 12325
rect 6160 12245 6165 12275
rect 6195 12245 6200 12275
rect 6160 12195 6200 12245
rect 6160 12165 6165 12195
rect 6195 12165 6200 12195
rect 6160 12115 6200 12165
rect 6160 12085 6165 12115
rect 6195 12085 6200 12115
rect 6160 12035 6200 12085
rect 6160 12005 6165 12035
rect 6195 12005 6200 12035
rect 6160 11955 6200 12005
rect 6160 11925 6165 11955
rect 6195 11925 6200 11955
rect 6160 11875 6200 11925
rect 6160 11845 6165 11875
rect 6195 11845 6200 11875
rect 6160 11795 6200 11845
rect 6160 11765 6165 11795
rect 6195 11765 6200 11795
rect 6160 11715 6200 11765
rect 6160 11685 6165 11715
rect 6195 11685 6200 11715
rect 6160 11635 6200 11685
rect 6160 11605 6165 11635
rect 6195 11605 6200 11635
rect 6160 11555 6200 11605
rect 6160 11525 6165 11555
rect 6195 11525 6200 11555
rect 6160 11475 6200 11525
rect 6160 11445 6165 11475
rect 6195 11445 6200 11475
rect 6160 11395 6200 11445
rect 6160 11365 6165 11395
rect 6195 11365 6200 11395
rect 6160 11315 6200 11365
rect 6160 11285 6165 11315
rect 6195 11285 6200 11315
rect 6160 11235 6200 11285
rect 6160 11205 6165 11235
rect 6195 11205 6200 11235
rect 6160 11155 6200 11205
rect 6160 11125 6165 11155
rect 6195 11125 6200 11155
rect 6160 11075 6200 11125
rect 6160 11045 6165 11075
rect 6195 11045 6200 11075
rect 6160 10990 6200 11045
rect 6160 10970 6170 10990
rect 6190 10970 6200 10990
rect 6160 10915 6200 10970
rect 6160 10885 6165 10915
rect 6195 10885 6200 10915
rect 6160 10835 6200 10885
rect 6160 10805 6165 10835
rect 6195 10805 6200 10835
rect 6160 10755 6200 10805
rect 6160 10725 6165 10755
rect 6195 10725 6200 10755
rect 6160 10675 6200 10725
rect 6160 10645 6165 10675
rect 6195 10645 6200 10675
rect 6160 10595 6200 10645
rect 6160 10565 6165 10595
rect 6195 10565 6200 10595
rect 6160 10515 6200 10565
rect 6160 10485 6165 10515
rect 6195 10485 6200 10515
rect 6160 10435 6200 10485
rect 6160 10405 6165 10435
rect 6195 10405 6200 10435
rect 6160 10355 6200 10405
rect 6160 10325 6165 10355
rect 6195 10325 6200 10355
rect 6160 10270 6200 10325
rect 6160 10250 6170 10270
rect 6190 10250 6200 10270
rect 6160 10190 6200 10250
rect 6160 10170 6170 10190
rect 6190 10170 6200 10190
rect 6160 10110 6200 10170
rect 6160 10090 6170 10110
rect 6190 10090 6200 10110
rect 6160 10030 6200 10090
rect 6160 10010 6170 10030
rect 6190 10010 6200 10030
rect 6160 9955 6200 10010
rect 6160 9925 6165 9955
rect 6195 9925 6200 9955
rect 6160 9875 6200 9925
rect 6160 9845 6165 9875
rect 6195 9845 6200 9875
rect 6160 9795 6200 9845
rect 6160 9765 6165 9795
rect 6195 9765 6200 9795
rect 6160 9715 6200 9765
rect 6160 9685 6165 9715
rect 6195 9685 6200 9715
rect 6160 9635 6200 9685
rect 6160 9605 6165 9635
rect 6195 9605 6200 9635
rect 6160 9555 6200 9605
rect 6160 9525 6165 9555
rect 6195 9525 6200 9555
rect 6160 9475 6200 9525
rect 6160 9445 6165 9475
rect 6195 9445 6200 9475
rect 6160 9395 6200 9445
rect 6160 9365 6165 9395
rect 6195 9365 6200 9395
rect 6160 9310 6200 9365
rect 6160 9290 6170 9310
rect 6190 9290 6200 9310
rect 6160 9230 6200 9290
rect 6160 9210 6170 9230
rect 6190 9210 6200 9230
rect 6160 9150 6200 9210
rect 6160 9130 6170 9150
rect 6190 9130 6200 9150
rect 6160 9070 6200 9130
rect 6160 9050 6170 9070
rect 6190 9050 6200 9070
rect 6160 8995 6200 9050
rect 6160 8965 6165 8995
rect 6195 8965 6200 8995
rect 6160 8915 6200 8965
rect 6160 8885 6165 8915
rect 6195 8885 6200 8915
rect 6160 8835 6200 8885
rect 6160 8805 6165 8835
rect 6195 8805 6200 8835
rect 6160 8755 6200 8805
rect 6160 8725 6165 8755
rect 6195 8725 6200 8755
rect 6160 8675 6200 8725
rect 6160 8645 6165 8675
rect 6195 8645 6200 8675
rect 6160 8595 6200 8645
rect 6160 8565 6165 8595
rect 6195 8565 6200 8595
rect 6160 8515 6200 8565
rect 6160 8485 6165 8515
rect 6195 8485 6200 8515
rect 6160 8435 6200 8485
rect 6160 8405 6165 8435
rect 6195 8405 6200 8435
rect 6160 8350 6200 8405
rect 6160 8330 6170 8350
rect 6190 8330 6200 8350
rect 6160 8275 6200 8330
rect 6160 8245 6165 8275
rect 6195 8245 6200 8275
rect 6160 8195 6200 8245
rect 6160 8165 6165 8195
rect 6195 8165 6200 8195
rect 6160 8115 6200 8165
rect 6160 8085 6165 8115
rect 6195 8085 6200 8115
rect 6160 8035 6200 8085
rect 6160 8005 6165 8035
rect 6195 8005 6200 8035
rect 6160 7955 6200 8005
rect 6160 7925 6165 7955
rect 6195 7925 6200 7955
rect 6160 7875 6200 7925
rect 6160 7845 6165 7875
rect 6195 7845 6200 7875
rect 6160 7795 6200 7845
rect 6160 7765 6165 7795
rect 6195 7765 6200 7795
rect 6160 7715 6200 7765
rect 6160 7685 6165 7715
rect 6195 7685 6200 7715
rect 6160 7635 6200 7685
rect 6160 7605 6165 7635
rect 6195 7605 6200 7635
rect 6160 7555 6200 7605
rect 6160 7525 6165 7555
rect 6195 7525 6200 7555
rect 6160 7475 6200 7525
rect 6160 7445 6165 7475
rect 6195 7445 6200 7475
rect 6160 7395 6200 7445
rect 6160 7365 6165 7395
rect 6195 7365 6200 7395
rect 6160 7315 6200 7365
rect 6160 7285 6165 7315
rect 6195 7285 6200 7315
rect 6160 7235 6200 7285
rect 6160 7205 6165 7235
rect 6195 7205 6200 7235
rect 6160 7155 6200 7205
rect 6160 7125 6165 7155
rect 6195 7125 6200 7155
rect 6160 7075 6200 7125
rect 6160 7045 6165 7075
rect 6195 7045 6200 7075
rect 6160 6995 6200 7045
rect 6160 6965 6165 6995
rect 6195 6965 6200 6995
rect 6160 6910 6200 6965
rect 6160 6890 6170 6910
rect 6190 6890 6200 6910
rect 6160 6835 6200 6890
rect 6160 6805 6165 6835
rect 6195 6805 6200 6835
rect 6160 6755 6200 6805
rect 6160 6725 6165 6755
rect 6195 6725 6200 6755
rect 6160 6675 6200 6725
rect 6160 6645 6165 6675
rect 6195 6645 6200 6675
rect 6160 6595 6200 6645
rect 6160 6565 6165 6595
rect 6195 6565 6200 6595
rect 6160 6515 6200 6565
rect 6160 6485 6165 6515
rect 6195 6485 6200 6515
rect 6160 6435 6200 6485
rect 6160 6405 6165 6435
rect 6195 6405 6200 6435
rect 6160 6355 6200 6405
rect 6160 6325 6165 6355
rect 6195 6325 6200 6355
rect 6160 6275 6200 6325
rect 6160 6245 6165 6275
rect 6195 6245 6200 6275
rect 6160 6190 6200 6245
rect 6160 6170 6170 6190
rect 6190 6170 6200 6190
rect 6160 6110 6200 6170
rect 6160 6090 6170 6110
rect 6190 6090 6200 6110
rect 6160 6030 6200 6090
rect 6160 6010 6170 6030
rect 6190 6010 6200 6030
rect 6160 5950 6200 6010
rect 6160 5930 6170 5950
rect 6190 5930 6200 5950
rect 6160 5875 6200 5930
rect 6160 5845 6165 5875
rect 6195 5845 6200 5875
rect 6160 5795 6200 5845
rect 6160 5765 6165 5795
rect 6195 5765 6200 5795
rect 6160 5715 6200 5765
rect 6160 5685 6165 5715
rect 6195 5685 6200 5715
rect 6160 5635 6200 5685
rect 6160 5605 6165 5635
rect 6195 5605 6200 5635
rect 6160 5555 6200 5605
rect 6160 5525 6165 5555
rect 6195 5525 6200 5555
rect 6160 5475 6200 5525
rect 6160 5445 6165 5475
rect 6195 5445 6200 5475
rect 6160 5395 6200 5445
rect 6160 5365 6165 5395
rect 6195 5365 6200 5395
rect 6160 5315 6200 5365
rect 6160 5285 6165 5315
rect 6195 5285 6200 5315
rect 6160 5235 6200 5285
rect 6160 5205 6165 5235
rect 6195 5205 6200 5235
rect 6160 5155 6200 5205
rect 6160 5125 6165 5155
rect 6195 5125 6200 5155
rect 6160 5075 6200 5125
rect 6160 5045 6165 5075
rect 6195 5045 6200 5075
rect 6160 4995 6200 5045
rect 6160 4965 6165 4995
rect 6195 4965 6200 4995
rect 6160 4915 6200 4965
rect 6160 4885 6165 4915
rect 6195 4885 6200 4915
rect 6160 4830 6200 4885
rect 6160 4810 6170 4830
rect 6190 4810 6200 4830
rect 6160 4755 6200 4810
rect 6160 4725 6165 4755
rect 6195 4725 6200 4755
rect 6160 4675 6200 4725
rect 6160 4645 6165 4675
rect 6195 4645 6200 4675
rect 6160 4590 6200 4645
rect 6160 4570 6170 4590
rect 6190 4570 6200 4590
rect 6160 4515 6200 4570
rect 6160 4485 6165 4515
rect 6195 4485 6200 4515
rect 6160 4435 6200 4485
rect 6160 4405 6165 4435
rect 6195 4405 6200 4435
rect 6160 4355 6200 4405
rect 6160 4325 6165 4355
rect 6195 4325 6200 4355
rect 6160 4275 6200 4325
rect 6160 4245 6165 4275
rect 6195 4245 6200 4275
rect 6160 4195 6200 4245
rect 6160 4165 6165 4195
rect 6195 4165 6200 4195
rect 6160 4115 6200 4165
rect 6160 4085 6165 4115
rect 6195 4085 6200 4115
rect 6160 4035 6200 4085
rect 6160 4005 6165 4035
rect 6195 4005 6200 4035
rect 6160 3955 6200 4005
rect 6160 3925 6165 3955
rect 6195 3925 6200 3955
rect 6160 3875 6200 3925
rect 6160 3845 6165 3875
rect 6195 3845 6200 3875
rect 6160 3790 6200 3845
rect 6160 3770 6170 3790
rect 6190 3770 6200 3790
rect 6160 3715 6200 3770
rect 6160 3685 6165 3715
rect 6195 3685 6200 3715
rect 6160 3635 6200 3685
rect 6160 3605 6165 3635
rect 6195 3605 6200 3635
rect 6160 3550 6200 3605
rect 6160 3530 6170 3550
rect 6190 3530 6200 3550
rect 6160 3475 6200 3530
rect 6160 3445 6165 3475
rect 6195 3445 6200 3475
rect 6160 3395 6200 3445
rect 6160 3365 6165 3395
rect 6195 3365 6200 3395
rect 6160 3310 6200 3365
rect 6160 3290 6170 3310
rect 6190 3290 6200 3310
rect 6160 3235 6200 3290
rect 6160 3205 6165 3235
rect 6195 3205 6200 3235
rect 6160 3155 6200 3205
rect 6160 3125 6165 3155
rect 6195 3125 6200 3155
rect 6160 3075 6200 3125
rect 6160 3045 6165 3075
rect 6195 3045 6200 3075
rect 6160 2995 6200 3045
rect 6160 2965 6165 2995
rect 6195 2965 6200 2995
rect 6160 2915 6200 2965
rect 6160 2885 6165 2915
rect 6195 2885 6200 2915
rect 6160 2835 6200 2885
rect 6160 2805 6165 2835
rect 6195 2805 6200 2835
rect 6160 2755 6200 2805
rect 6160 2725 6165 2755
rect 6195 2725 6200 2755
rect 6160 2675 6200 2725
rect 6160 2645 6165 2675
rect 6195 2645 6200 2675
rect 6160 2595 6200 2645
rect 6160 2565 6165 2595
rect 6195 2565 6200 2595
rect 6160 2515 6200 2565
rect 6160 2485 6165 2515
rect 6195 2485 6200 2515
rect 6160 2435 6200 2485
rect 6160 2405 6165 2435
rect 6195 2405 6200 2435
rect 6160 2355 6200 2405
rect 6160 2325 6165 2355
rect 6195 2325 6200 2355
rect 6160 2275 6200 2325
rect 6160 2245 6165 2275
rect 6195 2245 6200 2275
rect 6160 2195 6200 2245
rect 6160 2165 6165 2195
rect 6195 2165 6200 2195
rect 6160 2115 6200 2165
rect 6160 2085 6165 2115
rect 6195 2085 6200 2115
rect 6160 2035 6200 2085
rect 6160 2005 6165 2035
rect 6195 2005 6200 2035
rect 6160 1955 6200 2005
rect 6160 1925 6165 1955
rect 6195 1925 6200 1955
rect 6160 1870 6200 1925
rect 6160 1850 6170 1870
rect 6190 1850 6200 1870
rect 6160 1790 6200 1850
rect 6160 1770 6170 1790
rect 6190 1770 6200 1790
rect 6160 1715 6200 1770
rect 6160 1685 6165 1715
rect 6195 1685 6200 1715
rect 6160 1635 6200 1685
rect 6160 1605 6165 1635
rect 6195 1605 6200 1635
rect 6160 1555 6200 1605
rect 6160 1525 6165 1555
rect 6195 1525 6200 1555
rect 6160 1475 6200 1525
rect 6160 1445 6165 1475
rect 6195 1445 6200 1475
rect 6160 1395 6200 1445
rect 6160 1365 6165 1395
rect 6195 1365 6200 1395
rect 6160 1315 6200 1365
rect 6160 1285 6165 1315
rect 6195 1285 6200 1315
rect 6160 1235 6200 1285
rect 6160 1205 6165 1235
rect 6195 1205 6200 1235
rect 6160 1155 6200 1205
rect 6160 1125 6165 1155
rect 6195 1125 6200 1155
rect 6160 1075 6200 1125
rect 6160 1045 6165 1075
rect 6195 1045 6200 1075
rect 6160 995 6200 1045
rect 6160 965 6165 995
rect 6195 965 6200 995
rect 6160 910 6200 965
rect 6160 890 6170 910
rect 6190 890 6200 910
rect 6160 835 6200 890
rect 6160 805 6165 835
rect 6195 805 6200 835
rect 6160 755 6200 805
rect 6160 725 6165 755
rect 6195 725 6200 755
rect 6160 675 6200 725
rect 6160 645 6165 675
rect 6195 645 6200 675
rect 6160 595 6200 645
rect 6160 565 6165 595
rect 6195 565 6200 595
rect 6160 515 6200 565
rect 6160 485 6165 515
rect 6195 485 6200 515
rect 6160 430 6200 485
rect 6160 410 6170 430
rect 6190 410 6200 430
rect 6160 350 6200 410
rect 6160 330 6170 350
rect 6190 330 6200 350
rect 6160 275 6200 330
rect 6160 245 6165 275
rect 6195 245 6200 275
rect 6160 195 6200 245
rect 6160 165 6165 195
rect 6195 165 6200 195
rect 6160 115 6200 165
rect 6160 85 6165 115
rect 6195 85 6200 115
rect 6160 35 6200 85
rect 6160 5 6165 35
rect 6195 5 6200 35
rect 6160 0 6200 5
<< via1 >>
rect 4245 15710 4275 15715
rect 4245 15690 4250 15710
rect 4250 15690 4270 15710
rect 4270 15690 4275 15710
rect 4245 15685 4275 15690
rect 4245 15630 4275 15635
rect 4245 15610 4250 15630
rect 4250 15610 4270 15630
rect 4270 15610 4275 15630
rect 4245 15605 4275 15610
rect 4245 15550 4275 15555
rect 4245 15530 4250 15550
rect 4250 15530 4270 15550
rect 4270 15530 4275 15550
rect 4245 15525 4275 15530
rect 4245 15470 4275 15475
rect 4245 15450 4250 15470
rect 4250 15450 4270 15470
rect 4270 15450 4275 15470
rect 4245 15445 4275 15450
rect 4245 15390 4275 15395
rect 4245 15370 4250 15390
rect 4250 15370 4270 15390
rect 4270 15370 4275 15390
rect 4245 15365 4275 15370
rect 4245 15310 4275 15315
rect 4245 15290 4250 15310
rect 4250 15290 4270 15310
rect 4270 15290 4275 15310
rect 4245 15285 4275 15290
rect 4245 15230 4275 15235
rect 4245 15210 4250 15230
rect 4250 15210 4270 15230
rect 4270 15210 4275 15230
rect 4245 15205 4275 15210
rect 4245 15150 4275 15155
rect 4245 15130 4250 15150
rect 4250 15130 4270 15150
rect 4270 15130 4275 15150
rect 4245 15125 4275 15130
rect 4245 14990 4275 14995
rect 4245 14970 4250 14990
rect 4250 14970 4270 14990
rect 4270 14970 4275 14990
rect 4245 14965 4275 14970
rect 4245 14910 4275 14915
rect 4245 14890 4250 14910
rect 4250 14890 4270 14910
rect 4270 14890 4275 14910
rect 4245 14885 4275 14890
rect 4245 14830 4275 14835
rect 4245 14810 4250 14830
rect 4250 14810 4270 14830
rect 4270 14810 4275 14830
rect 4245 14805 4275 14810
rect 4245 14750 4275 14755
rect 4245 14730 4250 14750
rect 4250 14730 4270 14750
rect 4270 14730 4275 14750
rect 4245 14725 4275 14730
rect 4245 14670 4275 14675
rect 4245 14650 4250 14670
rect 4250 14650 4270 14670
rect 4270 14650 4275 14670
rect 4245 14645 4275 14650
rect 4245 14590 4275 14595
rect 4245 14570 4250 14590
rect 4250 14570 4270 14590
rect 4270 14570 4275 14590
rect 4245 14565 4275 14570
rect 4245 14510 4275 14515
rect 4245 14490 4250 14510
rect 4250 14490 4270 14510
rect 4270 14490 4275 14510
rect 4245 14485 4275 14490
rect 4245 14430 4275 14435
rect 4245 14410 4250 14430
rect 4250 14410 4270 14430
rect 4270 14410 4275 14430
rect 4245 14405 4275 14410
rect 4245 14030 4275 14035
rect 4245 14010 4250 14030
rect 4250 14010 4270 14030
rect 4270 14010 4275 14030
rect 4245 14005 4275 14010
rect 4245 13950 4275 13955
rect 4245 13930 4250 13950
rect 4250 13930 4270 13950
rect 4270 13930 4275 13950
rect 4245 13925 4275 13930
rect 4245 13870 4275 13875
rect 4245 13850 4250 13870
rect 4250 13850 4270 13870
rect 4270 13850 4275 13870
rect 4245 13845 4275 13850
rect 4245 13790 4275 13795
rect 4245 13770 4250 13790
rect 4250 13770 4270 13790
rect 4270 13770 4275 13790
rect 4245 13765 4275 13770
rect 4245 13710 4275 13715
rect 4245 13690 4250 13710
rect 4250 13690 4270 13710
rect 4270 13690 4275 13710
rect 4245 13685 4275 13690
rect 4245 13630 4275 13635
rect 4245 13610 4250 13630
rect 4250 13610 4270 13630
rect 4270 13610 4275 13630
rect 4245 13605 4275 13610
rect 4245 13550 4275 13555
rect 4245 13530 4250 13550
rect 4250 13530 4270 13550
rect 4270 13530 4275 13550
rect 4245 13525 4275 13530
rect 4245 13470 4275 13475
rect 4245 13450 4250 13470
rect 4250 13450 4270 13470
rect 4270 13450 4275 13470
rect 4245 13445 4275 13450
rect 4245 13070 4275 13075
rect 4245 13050 4250 13070
rect 4250 13050 4270 13070
rect 4270 13050 4275 13070
rect 4245 13045 4275 13050
rect 4245 12990 4275 12995
rect 4245 12970 4250 12990
rect 4250 12970 4270 12990
rect 4270 12970 4275 12990
rect 4245 12965 4275 12970
rect 4245 12910 4275 12915
rect 4245 12890 4250 12910
rect 4250 12890 4270 12910
rect 4270 12890 4275 12910
rect 4245 12885 4275 12890
rect 4245 12830 4275 12835
rect 4245 12810 4250 12830
rect 4250 12810 4270 12830
rect 4270 12810 4275 12830
rect 4245 12805 4275 12810
rect 4245 12750 4275 12755
rect 4245 12730 4250 12750
rect 4250 12730 4270 12750
rect 4270 12730 4275 12750
rect 4245 12725 4275 12730
rect 4245 12670 4275 12675
rect 4245 12650 4250 12670
rect 4250 12650 4270 12670
rect 4270 12650 4275 12670
rect 4245 12645 4275 12650
rect 4245 12590 4275 12595
rect 4245 12570 4250 12590
rect 4250 12570 4270 12590
rect 4270 12570 4275 12590
rect 4245 12565 4275 12570
rect 4245 12510 4275 12515
rect 4245 12490 4250 12510
rect 4250 12490 4270 12510
rect 4270 12490 4275 12510
rect 4245 12485 4275 12490
rect 4245 12350 4275 12355
rect 4245 12330 4250 12350
rect 4250 12330 4270 12350
rect 4270 12330 4275 12350
rect 4245 12325 4275 12330
rect 4245 12270 4275 12275
rect 4245 12250 4250 12270
rect 4250 12250 4270 12270
rect 4270 12250 4275 12270
rect 4245 12245 4275 12250
rect 4245 12190 4275 12195
rect 4245 12170 4250 12190
rect 4250 12170 4270 12190
rect 4270 12170 4275 12190
rect 4245 12165 4275 12170
rect 4245 12110 4275 12115
rect 4245 12090 4250 12110
rect 4250 12090 4270 12110
rect 4270 12090 4275 12110
rect 4245 12085 4275 12090
rect 4245 12030 4275 12035
rect 4245 12010 4250 12030
rect 4250 12010 4270 12030
rect 4270 12010 4275 12030
rect 4245 12005 4275 12010
rect 4245 11950 4275 11955
rect 4245 11930 4250 11950
rect 4250 11930 4270 11950
rect 4270 11930 4275 11950
rect 4245 11925 4275 11930
rect 4245 11870 4275 11875
rect 4245 11850 4250 11870
rect 4250 11850 4270 11870
rect 4270 11850 4275 11870
rect 4245 11845 4275 11850
rect 4245 11790 4275 11795
rect 4245 11770 4250 11790
rect 4250 11770 4270 11790
rect 4270 11770 4275 11790
rect 4245 11765 4275 11770
rect 4245 11710 4275 11715
rect 4245 11690 4250 11710
rect 4250 11690 4270 11710
rect 4270 11690 4275 11710
rect 4245 11685 4275 11690
rect 4245 11630 4275 11635
rect 4245 11610 4250 11630
rect 4250 11610 4270 11630
rect 4270 11610 4275 11630
rect 4245 11605 4275 11610
rect 4245 11550 4275 11555
rect 4245 11530 4250 11550
rect 4250 11530 4270 11550
rect 4270 11530 4275 11550
rect 4245 11525 4275 11530
rect 4245 11470 4275 11475
rect 4245 11450 4250 11470
rect 4250 11450 4270 11470
rect 4270 11450 4275 11470
rect 4245 11445 4275 11450
rect 4245 11390 4275 11395
rect 4245 11370 4250 11390
rect 4250 11370 4270 11390
rect 4270 11370 4275 11390
rect 4245 11365 4275 11370
rect 4245 11310 4275 11315
rect 4245 11290 4250 11310
rect 4250 11290 4270 11310
rect 4270 11290 4275 11310
rect 4245 11285 4275 11290
rect 4245 11230 4275 11235
rect 4245 11210 4250 11230
rect 4250 11210 4270 11230
rect 4270 11210 4275 11230
rect 4245 11205 4275 11210
rect 4245 11150 4275 11155
rect 4245 11130 4250 11150
rect 4250 11130 4270 11150
rect 4270 11130 4275 11150
rect 4245 11125 4275 11130
rect 4245 11070 4275 11075
rect 4245 11050 4250 11070
rect 4250 11050 4270 11070
rect 4270 11050 4275 11070
rect 4245 11045 4275 11050
rect 4245 10910 4275 10915
rect 4245 10890 4250 10910
rect 4250 10890 4270 10910
rect 4270 10890 4275 10910
rect 4245 10885 4275 10890
rect 4245 10830 4275 10835
rect 4245 10810 4250 10830
rect 4250 10810 4270 10830
rect 4270 10810 4275 10830
rect 4245 10805 4275 10810
rect 4245 10750 4275 10755
rect 4245 10730 4250 10750
rect 4250 10730 4270 10750
rect 4270 10730 4275 10750
rect 4245 10725 4275 10730
rect 4245 10670 4275 10675
rect 4245 10650 4250 10670
rect 4250 10650 4270 10670
rect 4270 10650 4275 10670
rect 4245 10645 4275 10650
rect 4245 10590 4275 10595
rect 4245 10570 4250 10590
rect 4250 10570 4270 10590
rect 4270 10570 4275 10590
rect 4245 10565 4275 10570
rect 4245 10510 4275 10515
rect 4245 10490 4250 10510
rect 4250 10490 4270 10510
rect 4270 10490 4275 10510
rect 4245 10485 4275 10490
rect 4245 10430 4275 10435
rect 4245 10410 4250 10430
rect 4250 10410 4270 10430
rect 4270 10410 4275 10430
rect 4245 10405 4275 10410
rect 4245 10350 4275 10355
rect 4245 10330 4250 10350
rect 4250 10330 4270 10350
rect 4270 10330 4275 10350
rect 4245 10325 4275 10330
rect 4245 9950 4275 9955
rect 4245 9930 4250 9950
rect 4250 9930 4270 9950
rect 4270 9930 4275 9950
rect 4245 9925 4275 9930
rect 4245 9870 4275 9875
rect 4245 9850 4250 9870
rect 4250 9850 4270 9870
rect 4270 9850 4275 9870
rect 4245 9845 4275 9850
rect 4245 9790 4275 9795
rect 4245 9770 4250 9790
rect 4250 9770 4270 9790
rect 4270 9770 4275 9790
rect 4245 9765 4275 9770
rect 4245 9710 4275 9715
rect 4245 9690 4250 9710
rect 4250 9690 4270 9710
rect 4270 9690 4275 9710
rect 4245 9685 4275 9690
rect 4245 9630 4275 9635
rect 4245 9610 4250 9630
rect 4250 9610 4270 9630
rect 4270 9610 4275 9630
rect 4245 9605 4275 9610
rect 4245 9550 4275 9555
rect 4245 9530 4250 9550
rect 4250 9530 4270 9550
rect 4270 9530 4275 9550
rect 4245 9525 4275 9530
rect 4245 9470 4275 9475
rect 4245 9450 4250 9470
rect 4250 9450 4270 9470
rect 4270 9450 4275 9470
rect 4245 9445 4275 9450
rect 4245 9390 4275 9395
rect 4245 9370 4250 9390
rect 4250 9370 4270 9390
rect 4270 9370 4275 9390
rect 4245 9365 4275 9370
rect 4245 8990 4275 8995
rect 4245 8970 4250 8990
rect 4250 8970 4270 8990
rect 4270 8970 4275 8990
rect 4245 8965 4275 8970
rect 4245 8910 4275 8915
rect 4245 8890 4250 8910
rect 4250 8890 4270 8910
rect 4270 8890 4275 8910
rect 4245 8885 4275 8890
rect 4245 8830 4275 8835
rect 4245 8810 4250 8830
rect 4250 8810 4270 8830
rect 4270 8810 4275 8830
rect 4245 8805 4275 8810
rect 4245 8750 4275 8755
rect 4245 8730 4250 8750
rect 4250 8730 4270 8750
rect 4270 8730 4275 8750
rect 4245 8725 4275 8730
rect 4245 8670 4275 8675
rect 4245 8650 4250 8670
rect 4250 8650 4270 8670
rect 4270 8650 4275 8670
rect 4245 8645 4275 8650
rect 4245 8590 4275 8595
rect 4245 8570 4250 8590
rect 4250 8570 4270 8590
rect 4270 8570 4275 8590
rect 4245 8565 4275 8570
rect 4245 8510 4275 8515
rect 4245 8490 4250 8510
rect 4250 8490 4270 8510
rect 4270 8490 4275 8510
rect 4245 8485 4275 8490
rect 4245 8430 4275 8435
rect 4245 8410 4250 8430
rect 4250 8410 4270 8430
rect 4270 8410 4275 8430
rect 4245 8405 4275 8410
rect 4245 8270 4275 8275
rect 4245 8250 4250 8270
rect 4250 8250 4270 8270
rect 4270 8250 4275 8270
rect 4245 8245 4275 8250
rect 4245 8190 4275 8195
rect 4245 8170 4250 8190
rect 4250 8170 4270 8190
rect 4270 8170 4275 8190
rect 4245 8165 4275 8170
rect 4245 8110 4275 8115
rect 4245 8090 4250 8110
rect 4250 8090 4270 8110
rect 4270 8090 4275 8110
rect 4245 8085 4275 8090
rect 4245 8030 4275 8035
rect 4245 8010 4250 8030
rect 4250 8010 4270 8030
rect 4270 8010 4275 8030
rect 4245 8005 4275 8010
rect 4245 7950 4275 7955
rect 4245 7930 4250 7950
rect 4250 7930 4270 7950
rect 4270 7930 4275 7950
rect 4245 7925 4275 7930
rect 4245 7870 4275 7875
rect 4245 7850 4250 7870
rect 4250 7850 4270 7870
rect 4270 7850 4275 7870
rect 4245 7845 4275 7850
rect 4245 7790 4275 7795
rect 4245 7770 4250 7790
rect 4250 7770 4270 7790
rect 4270 7770 4275 7790
rect 4245 7765 4275 7770
rect 4245 7710 4275 7715
rect 4245 7690 4250 7710
rect 4250 7690 4270 7710
rect 4270 7690 4275 7710
rect 4245 7685 4275 7690
rect 4245 7630 4275 7635
rect 4245 7610 4250 7630
rect 4250 7610 4270 7630
rect 4270 7610 4275 7630
rect 4245 7605 4275 7610
rect 4245 7550 4275 7555
rect 4245 7530 4250 7550
rect 4250 7530 4270 7550
rect 4270 7530 4275 7550
rect 4245 7525 4275 7530
rect 4245 7470 4275 7475
rect 4245 7450 4250 7470
rect 4250 7450 4270 7470
rect 4270 7450 4275 7470
rect 4245 7445 4275 7450
rect 4245 7390 4275 7395
rect 4245 7370 4250 7390
rect 4250 7370 4270 7390
rect 4270 7370 4275 7390
rect 4245 7365 4275 7370
rect 4245 7310 4275 7315
rect 4245 7290 4250 7310
rect 4250 7290 4270 7310
rect 4270 7290 4275 7310
rect 4245 7285 4275 7290
rect 4245 7230 4275 7235
rect 4245 7210 4250 7230
rect 4250 7210 4270 7230
rect 4270 7210 4275 7230
rect 4245 7205 4275 7210
rect 4245 7150 4275 7155
rect 4245 7130 4250 7150
rect 4250 7130 4270 7150
rect 4270 7130 4275 7150
rect 4245 7125 4275 7130
rect 4245 7070 4275 7075
rect 4245 7050 4250 7070
rect 4250 7050 4270 7070
rect 4270 7050 4275 7070
rect 4245 7045 4275 7050
rect 4245 6990 4275 6995
rect 4245 6970 4250 6990
rect 4250 6970 4270 6990
rect 4270 6970 4275 6990
rect 4245 6965 4275 6970
rect 4245 6830 4275 6835
rect 4245 6810 4250 6830
rect 4250 6810 4270 6830
rect 4270 6810 4275 6830
rect 4245 6805 4275 6810
rect 4245 6750 4275 6755
rect 4245 6730 4250 6750
rect 4250 6730 4270 6750
rect 4270 6730 4275 6750
rect 4245 6725 4275 6730
rect 4245 6670 4275 6675
rect 4245 6650 4250 6670
rect 4250 6650 4270 6670
rect 4270 6650 4275 6670
rect 4245 6645 4275 6650
rect 4245 6590 4275 6595
rect 4245 6570 4250 6590
rect 4250 6570 4270 6590
rect 4270 6570 4275 6590
rect 4245 6565 4275 6570
rect 4245 6510 4275 6515
rect 4245 6490 4250 6510
rect 4250 6490 4270 6510
rect 4270 6490 4275 6510
rect 4245 6485 4275 6490
rect 4245 6430 4275 6435
rect 4245 6410 4250 6430
rect 4250 6410 4270 6430
rect 4270 6410 4275 6430
rect 4245 6405 4275 6410
rect 4245 6350 4275 6355
rect 4245 6330 4250 6350
rect 4250 6330 4270 6350
rect 4270 6330 4275 6350
rect 4245 6325 4275 6330
rect 4245 6270 4275 6275
rect 4245 6250 4250 6270
rect 4250 6250 4270 6270
rect 4270 6250 4275 6270
rect 4245 6245 4275 6250
rect 4245 5870 4275 5875
rect 4245 5850 4250 5870
rect 4250 5850 4270 5870
rect 4270 5850 4275 5870
rect 4245 5845 4275 5850
rect 4245 5790 4275 5795
rect 4245 5770 4250 5790
rect 4250 5770 4270 5790
rect 4270 5770 4275 5790
rect 4245 5765 4275 5770
rect 4245 5710 4275 5715
rect 4245 5690 4250 5710
rect 4250 5690 4270 5710
rect 4270 5690 4275 5710
rect 4245 5685 4275 5690
rect 4245 5630 4275 5635
rect 4245 5610 4250 5630
rect 4250 5610 4270 5630
rect 4270 5610 4275 5630
rect 4245 5605 4275 5610
rect 4245 5550 4275 5555
rect 4245 5530 4250 5550
rect 4250 5530 4270 5550
rect 4270 5530 4275 5550
rect 4245 5525 4275 5530
rect 4245 5470 4275 5475
rect 4245 5450 4250 5470
rect 4250 5450 4270 5470
rect 4270 5450 4275 5470
rect 4245 5445 4275 5450
rect 4245 5390 4275 5395
rect 4245 5370 4250 5390
rect 4250 5370 4270 5390
rect 4270 5370 4275 5390
rect 4245 5365 4275 5370
rect 4245 5310 4275 5315
rect 4245 5290 4250 5310
rect 4250 5290 4270 5310
rect 4270 5290 4275 5310
rect 4245 5285 4275 5290
rect 4245 5230 4275 5235
rect 4245 5210 4250 5230
rect 4250 5210 4270 5230
rect 4270 5210 4275 5230
rect 4245 5205 4275 5210
rect 4245 5150 4275 5155
rect 4245 5130 4250 5150
rect 4250 5130 4270 5150
rect 4270 5130 4275 5150
rect 4245 5125 4275 5130
rect 4245 5070 4275 5075
rect 4245 5050 4250 5070
rect 4250 5050 4270 5070
rect 4270 5050 4275 5070
rect 4245 5045 4275 5050
rect 4245 4990 4275 4995
rect 4245 4970 4250 4990
rect 4250 4970 4270 4990
rect 4270 4970 4275 4990
rect 4245 4965 4275 4970
rect 4245 4910 4275 4915
rect 4245 4890 4250 4910
rect 4250 4890 4270 4910
rect 4270 4890 4275 4910
rect 4245 4885 4275 4890
rect 4245 4750 4275 4755
rect 4245 4730 4250 4750
rect 4250 4730 4270 4750
rect 4270 4730 4275 4750
rect 4245 4725 4275 4730
rect 4245 4670 4275 4675
rect 4245 4650 4250 4670
rect 4250 4650 4270 4670
rect 4270 4650 4275 4670
rect 4245 4645 4275 4650
rect 4245 4510 4275 4515
rect 4245 4490 4250 4510
rect 4250 4490 4270 4510
rect 4270 4490 4275 4510
rect 4245 4485 4275 4490
rect 4245 4430 4275 4435
rect 4245 4410 4250 4430
rect 4250 4410 4270 4430
rect 4270 4410 4275 4430
rect 4245 4405 4275 4410
rect 4245 4350 4275 4355
rect 4245 4330 4250 4350
rect 4250 4330 4270 4350
rect 4270 4330 4275 4350
rect 4245 4325 4275 4330
rect 4245 4270 4275 4275
rect 4245 4250 4250 4270
rect 4250 4250 4270 4270
rect 4270 4250 4275 4270
rect 4245 4245 4275 4250
rect 4245 4190 4275 4195
rect 4245 4170 4250 4190
rect 4250 4170 4270 4190
rect 4270 4170 4275 4190
rect 4245 4165 4275 4170
rect 4245 4110 4275 4115
rect 4245 4090 4250 4110
rect 4250 4090 4270 4110
rect 4270 4090 4275 4110
rect 4245 4085 4275 4090
rect 4245 4030 4275 4035
rect 4245 4010 4250 4030
rect 4250 4010 4270 4030
rect 4270 4010 4275 4030
rect 4245 4005 4275 4010
rect 4245 3950 4275 3955
rect 4245 3930 4250 3950
rect 4250 3930 4270 3950
rect 4270 3930 4275 3950
rect 4245 3925 4275 3930
rect 4245 3870 4275 3875
rect 4245 3850 4250 3870
rect 4250 3850 4270 3870
rect 4270 3850 4275 3870
rect 4245 3845 4275 3850
rect 4245 3710 4275 3715
rect 4245 3690 4250 3710
rect 4250 3690 4270 3710
rect 4270 3690 4275 3710
rect 4245 3685 4275 3690
rect 4245 3630 4275 3635
rect 4245 3610 4250 3630
rect 4250 3610 4270 3630
rect 4270 3610 4275 3630
rect 4245 3605 4275 3610
rect 4245 3470 4275 3475
rect 4245 3450 4250 3470
rect 4250 3450 4270 3470
rect 4270 3450 4275 3470
rect 4245 3445 4275 3450
rect 4245 3390 4275 3395
rect 4245 3370 4250 3390
rect 4250 3370 4270 3390
rect 4270 3370 4275 3390
rect 4245 3365 4275 3370
rect 4245 3230 4275 3235
rect 4245 3210 4250 3230
rect 4250 3210 4270 3230
rect 4270 3210 4275 3230
rect 4245 3205 4275 3210
rect 4245 3150 4275 3155
rect 4245 3130 4250 3150
rect 4250 3130 4270 3150
rect 4270 3130 4275 3150
rect 4245 3125 4275 3130
rect 4245 3070 4275 3075
rect 4245 3050 4250 3070
rect 4250 3050 4270 3070
rect 4270 3050 4275 3070
rect 4245 3045 4275 3050
rect 4245 2990 4275 2995
rect 4245 2970 4250 2990
rect 4250 2970 4270 2990
rect 4270 2970 4275 2990
rect 4245 2965 4275 2970
rect 4245 2910 4275 2915
rect 4245 2890 4250 2910
rect 4250 2890 4270 2910
rect 4270 2890 4275 2910
rect 4245 2885 4275 2890
rect 4245 2830 4275 2835
rect 4245 2810 4250 2830
rect 4250 2810 4270 2830
rect 4270 2810 4275 2830
rect 4245 2805 4275 2810
rect 4245 2750 4275 2755
rect 4245 2730 4250 2750
rect 4250 2730 4270 2750
rect 4270 2730 4275 2750
rect 4245 2725 4275 2730
rect 4245 2670 4275 2675
rect 4245 2650 4250 2670
rect 4250 2650 4270 2670
rect 4270 2650 4275 2670
rect 4245 2645 4275 2650
rect 4245 2590 4275 2595
rect 4245 2570 4250 2590
rect 4250 2570 4270 2590
rect 4270 2570 4275 2590
rect 4245 2565 4275 2570
rect 4245 2510 4275 2515
rect 4245 2490 4250 2510
rect 4250 2490 4270 2510
rect 4270 2490 4275 2510
rect 4245 2485 4275 2490
rect 4245 2430 4275 2435
rect 4245 2410 4250 2430
rect 4250 2410 4270 2430
rect 4270 2410 4275 2430
rect 4245 2405 4275 2410
rect 4245 2350 4275 2355
rect 4245 2330 4250 2350
rect 4250 2330 4270 2350
rect 4270 2330 4275 2350
rect 4245 2325 4275 2330
rect 4245 2270 4275 2275
rect 4245 2250 4250 2270
rect 4250 2250 4270 2270
rect 4270 2250 4275 2270
rect 4245 2245 4275 2250
rect 4245 2190 4275 2195
rect 4245 2170 4250 2190
rect 4250 2170 4270 2190
rect 4270 2170 4275 2190
rect 4245 2165 4275 2170
rect 4245 2110 4275 2115
rect 4245 2090 4250 2110
rect 4250 2090 4270 2110
rect 4270 2090 4275 2110
rect 4245 2085 4275 2090
rect 4245 2030 4275 2035
rect 4245 2010 4250 2030
rect 4250 2010 4270 2030
rect 4270 2010 4275 2030
rect 4245 2005 4275 2010
rect 4245 1950 4275 1955
rect 4245 1930 4250 1950
rect 4250 1930 4270 1950
rect 4270 1930 4275 1950
rect 4245 1925 4275 1930
rect 4245 1710 4275 1715
rect 4245 1690 4250 1710
rect 4250 1690 4270 1710
rect 4270 1690 4275 1710
rect 4245 1685 4275 1690
rect 4245 1630 4275 1635
rect 4245 1610 4250 1630
rect 4250 1610 4270 1630
rect 4270 1610 4275 1630
rect 4245 1605 4275 1610
rect 4245 1550 4275 1555
rect 4245 1530 4250 1550
rect 4250 1530 4270 1550
rect 4270 1530 4275 1550
rect 4245 1525 4275 1530
rect 4245 1470 4275 1475
rect 4245 1450 4250 1470
rect 4250 1450 4270 1470
rect 4270 1450 4275 1470
rect 4245 1445 4275 1450
rect 4245 1390 4275 1395
rect 4245 1370 4250 1390
rect 4250 1370 4270 1390
rect 4270 1370 4275 1390
rect 4245 1365 4275 1370
rect 4245 1310 4275 1315
rect 4245 1290 4250 1310
rect 4250 1290 4270 1310
rect 4270 1290 4275 1310
rect 4245 1285 4275 1290
rect 4245 1230 4275 1235
rect 4245 1210 4250 1230
rect 4250 1210 4270 1230
rect 4270 1210 4275 1230
rect 4245 1205 4275 1210
rect 4245 1150 4275 1155
rect 4245 1130 4250 1150
rect 4250 1130 4270 1150
rect 4270 1130 4275 1150
rect 4245 1125 4275 1130
rect 4245 1070 4275 1075
rect 4245 1050 4250 1070
rect 4250 1050 4270 1070
rect 4270 1050 4275 1070
rect 4245 1045 4275 1050
rect 4245 990 4275 995
rect 4245 970 4250 990
rect 4250 970 4270 990
rect 4270 970 4275 990
rect 4245 965 4275 970
rect 4245 830 4275 835
rect 4245 810 4250 830
rect 4250 810 4270 830
rect 4270 810 4275 830
rect 4245 805 4275 810
rect 4245 750 4275 755
rect 4245 730 4250 750
rect 4250 730 4270 750
rect 4270 730 4275 750
rect 4245 725 4275 730
rect 4245 670 4275 675
rect 4245 650 4250 670
rect 4250 650 4270 670
rect 4270 650 4275 670
rect 4245 645 4275 650
rect 4245 590 4275 595
rect 4245 570 4250 590
rect 4250 570 4270 590
rect 4270 570 4275 590
rect 4245 565 4275 570
rect 4245 510 4275 515
rect 4245 490 4250 510
rect 4250 490 4270 510
rect 4270 490 4275 510
rect 4245 485 4275 490
rect 4245 270 4275 275
rect 4245 250 4250 270
rect 4250 250 4270 270
rect 4270 250 4275 270
rect 4245 245 4275 250
rect 4245 190 4275 195
rect 4245 170 4250 190
rect 4250 170 4270 190
rect 4270 170 4275 190
rect 4245 165 4275 170
rect 4245 110 4275 115
rect 4245 90 4250 110
rect 4250 90 4270 110
rect 4270 90 4275 110
rect 4245 85 4275 90
rect 4245 30 4275 35
rect 4245 10 4250 30
rect 4250 10 4270 30
rect 4270 10 4275 30
rect 4245 5 4275 10
rect 4405 15710 4435 15715
rect 4405 15690 4410 15710
rect 4410 15690 4430 15710
rect 4430 15690 4435 15710
rect 4405 15685 4435 15690
rect 4405 15630 4435 15635
rect 4405 15610 4410 15630
rect 4410 15610 4430 15630
rect 4430 15610 4435 15630
rect 4405 15605 4435 15610
rect 4405 15550 4435 15555
rect 4405 15530 4410 15550
rect 4410 15530 4430 15550
rect 4430 15530 4435 15550
rect 4405 15525 4435 15530
rect 4405 15470 4435 15475
rect 4405 15450 4410 15470
rect 4410 15450 4430 15470
rect 4430 15450 4435 15470
rect 4405 15445 4435 15450
rect 4405 15390 4435 15395
rect 4405 15370 4410 15390
rect 4410 15370 4430 15390
rect 4430 15370 4435 15390
rect 4405 15365 4435 15370
rect 4405 15310 4435 15315
rect 4405 15290 4410 15310
rect 4410 15290 4430 15310
rect 4430 15290 4435 15310
rect 4405 15285 4435 15290
rect 4405 15230 4435 15235
rect 4405 15210 4410 15230
rect 4410 15210 4430 15230
rect 4430 15210 4435 15230
rect 4405 15205 4435 15210
rect 4405 15150 4435 15155
rect 4405 15130 4410 15150
rect 4410 15130 4430 15150
rect 4430 15130 4435 15150
rect 4405 15125 4435 15130
rect 4405 14990 4435 14995
rect 4405 14970 4410 14990
rect 4410 14970 4430 14990
rect 4430 14970 4435 14990
rect 4405 14965 4435 14970
rect 4405 14910 4435 14915
rect 4405 14890 4410 14910
rect 4410 14890 4430 14910
rect 4430 14890 4435 14910
rect 4405 14885 4435 14890
rect 4405 14830 4435 14835
rect 4405 14810 4410 14830
rect 4410 14810 4430 14830
rect 4430 14810 4435 14830
rect 4405 14805 4435 14810
rect 4405 14750 4435 14755
rect 4405 14730 4410 14750
rect 4410 14730 4430 14750
rect 4430 14730 4435 14750
rect 4405 14725 4435 14730
rect 4405 14670 4435 14675
rect 4405 14650 4410 14670
rect 4410 14650 4430 14670
rect 4430 14650 4435 14670
rect 4405 14645 4435 14650
rect 4405 14590 4435 14595
rect 4405 14570 4410 14590
rect 4410 14570 4430 14590
rect 4430 14570 4435 14590
rect 4405 14565 4435 14570
rect 4405 14510 4435 14515
rect 4405 14490 4410 14510
rect 4410 14490 4430 14510
rect 4430 14490 4435 14510
rect 4405 14485 4435 14490
rect 4405 14430 4435 14435
rect 4405 14410 4410 14430
rect 4410 14410 4430 14430
rect 4430 14410 4435 14430
rect 4405 14405 4435 14410
rect 4405 14030 4435 14035
rect 4405 14010 4410 14030
rect 4410 14010 4430 14030
rect 4430 14010 4435 14030
rect 4405 14005 4435 14010
rect 4405 13950 4435 13955
rect 4405 13930 4410 13950
rect 4410 13930 4430 13950
rect 4430 13930 4435 13950
rect 4405 13925 4435 13930
rect 4405 13870 4435 13875
rect 4405 13850 4410 13870
rect 4410 13850 4430 13870
rect 4430 13850 4435 13870
rect 4405 13845 4435 13850
rect 4405 13790 4435 13795
rect 4405 13770 4410 13790
rect 4410 13770 4430 13790
rect 4430 13770 4435 13790
rect 4405 13765 4435 13770
rect 4405 13710 4435 13715
rect 4405 13690 4410 13710
rect 4410 13690 4430 13710
rect 4430 13690 4435 13710
rect 4405 13685 4435 13690
rect 4405 13630 4435 13635
rect 4405 13610 4410 13630
rect 4410 13610 4430 13630
rect 4430 13610 4435 13630
rect 4405 13605 4435 13610
rect 4405 13550 4435 13555
rect 4405 13530 4410 13550
rect 4410 13530 4430 13550
rect 4430 13530 4435 13550
rect 4405 13525 4435 13530
rect 4405 13470 4435 13475
rect 4405 13450 4410 13470
rect 4410 13450 4430 13470
rect 4430 13450 4435 13470
rect 4405 13445 4435 13450
rect 4405 13070 4435 13075
rect 4405 13050 4410 13070
rect 4410 13050 4430 13070
rect 4430 13050 4435 13070
rect 4405 13045 4435 13050
rect 4405 12990 4435 12995
rect 4405 12970 4410 12990
rect 4410 12970 4430 12990
rect 4430 12970 4435 12990
rect 4405 12965 4435 12970
rect 4405 12910 4435 12915
rect 4405 12890 4410 12910
rect 4410 12890 4430 12910
rect 4430 12890 4435 12910
rect 4405 12885 4435 12890
rect 4405 12830 4435 12835
rect 4405 12810 4410 12830
rect 4410 12810 4430 12830
rect 4430 12810 4435 12830
rect 4405 12805 4435 12810
rect 4405 12750 4435 12755
rect 4405 12730 4410 12750
rect 4410 12730 4430 12750
rect 4430 12730 4435 12750
rect 4405 12725 4435 12730
rect 4405 12670 4435 12675
rect 4405 12650 4410 12670
rect 4410 12650 4430 12670
rect 4430 12650 4435 12670
rect 4405 12645 4435 12650
rect 4405 12590 4435 12595
rect 4405 12570 4410 12590
rect 4410 12570 4430 12590
rect 4430 12570 4435 12590
rect 4405 12565 4435 12570
rect 4405 12510 4435 12515
rect 4405 12490 4410 12510
rect 4410 12490 4430 12510
rect 4430 12490 4435 12510
rect 4405 12485 4435 12490
rect 4405 12350 4435 12355
rect 4405 12330 4410 12350
rect 4410 12330 4430 12350
rect 4430 12330 4435 12350
rect 4405 12325 4435 12330
rect 4405 12270 4435 12275
rect 4405 12250 4410 12270
rect 4410 12250 4430 12270
rect 4430 12250 4435 12270
rect 4405 12245 4435 12250
rect 4405 12190 4435 12195
rect 4405 12170 4410 12190
rect 4410 12170 4430 12190
rect 4430 12170 4435 12190
rect 4405 12165 4435 12170
rect 4405 12110 4435 12115
rect 4405 12090 4410 12110
rect 4410 12090 4430 12110
rect 4430 12090 4435 12110
rect 4405 12085 4435 12090
rect 4405 12030 4435 12035
rect 4405 12010 4410 12030
rect 4410 12010 4430 12030
rect 4430 12010 4435 12030
rect 4405 12005 4435 12010
rect 4405 11950 4435 11955
rect 4405 11930 4410 11950
rect 4410 11930 4430 11950
rect 4430 11930 4435 11950
rect 4405 11925 4435 11930
rect 4405 11870 4435 11875
rect 4405 11850 4410 11870
rect 4410 11850 4430 11870
rect 4430 11850 4435 11870
rect 4405 11845 4435 11850
rect 4405 11790 4435 11795
rect 4405 11770 4410 11790
rect 4410 11770 4430 11790
rect 4430 11770 4435 11790
rect 4405 11765 4435 11770
rect 4405 11710 4435 11715
rect 4405 11690 4410 11710
rect 4410 11690 4430 11710
rect 4430 11690 4435 11710
rect 4405 11685 4435 11690
rect 4405 11630 4435 11635
rect 4405 11610 4410 11630
rect 4410 11610 4430 11630
rect 4430 11610 4435 11630
rect 4405 11605 4435 11610
rect 4405 11550 4435 11555
rect 4405 11530 4410 11550
rect 4410 11530 4430 11550
rect 4430 11530 4435 11550
rect 4405 11525 4435 11530
rect 4405 11470 4435 11475
rect 4405 11450 4410 11470
rect 4410 11450 4430 11470
rect 4430 11450 4435 11470
rect 4405 11445 4435 11450
rect 4405 11390 4435 11395
rect 4405 11370 4410 11390
rect 4410 11370 4430 11390
rect 4430 11370 4435 11390
rect 4405 11365 4435 11370
rect 4405 11310 4435 11315
rect 4405 11290 4410 11310
rect 4410 11290 4430 11310
rect 4430 11290 4435 11310
rect 4405 11285 4435 11290
rect 4405 11230 4435 11235
rect 4405 11210 4410 11230
rect 4410 11210 4430 11230
rect 4430 11210 4435 11230
rect 4405 11205 4435 11210
rect 4405 11150 4435 11155
rect 4405 11130 4410 11150
rect 4410 11130 4430 11150
rect 4430 11130 4435 11150
rect 4405 11125 4435 11130
rect 4405 11070 4435 11075
rect 4405 11050 4410 11070
rect 4410 11050 4430 11070
rect 4430 11050 4435 11070
rect 4405 11045 4435 11050
rect 4405 10910 4435 10915
rect 4405 10890 4410 10910
rect 4410 10890 4430 10910
rect 4430 10890 4435 10910
rect 4405 10885 4435 10890
rect 4405 10830 4435 10835
rect 4405 10810 4410 10830
rect 4410 10810 4430 10830
rect 4430 10810 4435 10830
rect 4405 10805 4435 10810
rect 4405 10750 4435 10755
rect 4405 10730 4410 10750
rect 4410 10730 4430 10750
rect 4430 10730 4435 10750
rect 4405 10725 4435 10730
rect 4405 10670 4435 10675
rect 4405 10650 4410 10670
rect 4410 10650 4430 10670
rect 4430 10650 4435 10670
rect 4405 10645 4435 10650
rect 4405 10590 4435 10595
rect 4405 10570 4410 10590
rect 4410 10570 4430 10590
rect 4430 10570 4435 10590
rect 4405 10565 4435 10570
rect 4405 10510 4435 10515
rect 4405 10490 4410 10510
rect 4410 10490 4430 10510
rect 4430 10490 4435 10510
rect 4405 10485 4435 10490
rect 4405 10430 4435 10435
rect 4405 10410 4410 10430
rect 4410 10410 4430 10430
rect 4430 10410 4435 10430
rect 4405 10405 4435 10410
rect 4405 10350 4435 10355
rect 4405 10330 4410 10350
rect 4410 10330 4430 10350
rect 4430 10330 4435 10350
rect 4405 10325 4435 10330
rect 4405 9950 4435 9955
rect 4405 9930 4410 9950
rect 4410 9930 4430 9950
rect 4430 9930 4435 9950
rect 4405 9925 4435 9930
rect 4405 9870 4435 9875
rect 4405 9850 4410 9870
rect 4410 9850 4430 9870
rect 4430 9850 4435 9870
rect 4405 9845 4435 9850
rect 4405 9790 4435 9795
rect 4405 9770 4410 9790
rect 4410 9770 4430 9790
rect 4430 9770 4435 9790
rect 4405 9765 4435 9770
rect 4405 9710 4435 9715
rect 4405 9690 4410 9710
rect 4410 9690 4430 9710
rect 4430 9690 4435 9710
rect 4405 9685 4435 9690
rect 4405 9630 4435 9635
rect 4405 9610 4410 9630
rect 4410 9610 4430 9630
rect 4430 9610 4435 9630
rect 4405 9605 4435 9610
rect 4405 9550 4435 9555
rect 4405 9530 4410 9550
rect 4410 9530 4430 9550
rect 4430 9530 4435 9550
rect 4405 9525 4435 9530
rect 4405 9470 4435 9475
rect 4405 9450 4410 9470
rect 4410 9450 4430 9470
rect 4430 9450 4435 9470
rect 4405 9445 4435 9450
rect 4405 9390 4435 9395
rect 4405 9370 4410 9390
rect 4410 9370 4430 9390
rect 4430 9370 4435 9390
rect 4405 9365 4435 9370
rect 4405 8990 4435 8995
rect 4405 8970 4410 8990
rect 4410 8970 4430 8990
rect 4430 8970 4435 8990
rect 4405 8965 4435 8970
rect 4405 8910 4435 8915
rect 4405 8890 4410 8910
rect 4410 8890 4430 8910
rect 4430 8890 4435 8910
rect 4405 8885 4435 8890
rect 4405 8830 4435 8835
rect 4405 8810 4410 8830
rect 4410 8810 4430 8830
rect 4430 8810 4435 8830
rect 4405 8805 4435 8810
rect 4405 8750 4435 8755
rect 4405 8730 4410 8750
rect 4410 8730 4430 8750
rect 4430 8730 4435 8750
rect 4405 8725 4435 8730
rect 4405 8670 4435 8675
rect 4405 8650 4410 8670
rect 4410 8650 4430 8670
rect 4430 8650 4435 8670
rect 4405 8645 4435 8650
rect 4405 8590 4435 8595
rect 4405 8570 4410 8590
rect 4410 8570 4430 8590
rect 4430 8570 4435 8590
rect 4405 8565 4435 8570
rect 4405 8510 4435 8515
rect 4405 8490 4410 8510
rect 4410 8490 4430 8510
rect 4430 8490 4435 8510
rect 4405 8485 4435 8490
rect 4405 8430 4435 8435
rect 4405 8410 4410 8430
rect 4410 8410 4430 8430
rect 4430 8410 4435 8430
rect 4405 8405 4435 8410
rect 4405 8270 4435 8275
rect 4405 8250 4410 8270
rect 4410 8250 4430 8270
rect 4430 8250 4435 8270
rect 4405 8245 4435 8250
rect 4405 8190 4435 8195
rect 4405 8170 4410 8190
rect 4410 8170 4430 8190
rect 4430 8170 4435 8190
rect 4405 8165 4435 8170
rect 4405 8110 4435 8115
rect 4405 8090 4410 8110
rect 4410 8090 4430 8110
rect 4430 8090 4435 8110
rect 4405 8085 4435 8090
rect 4405 8030 4435 8035
rect 4405 8010 4410 8030
rect 4410 8010 4430 8030
rect 4430 8010 4435 8030
rect 4405 8005 4435 8010
rect 4405 7950 4435 7955
rect 4405 7930 4410 7950
rect 4410 7930 4430 7950
rect 4430 7930 4435 7950
rect 4405 7925 4435 7930
rect 4405 7870 4435 7875
rect 4405 7850 4410 7870
rect 4410 7850 4430 7870
rect 4430 7850 4435 7870
rect 4405 7845 4435 7850
rect 4405 7790 4435 7795
rect 4405 7770 4410 7790
rect 4410 7770 4430 7790
rect 4430 7770 4435 7790
rect 4405 7765 4435 7770
rect 4405 7710 4435 7715
rect 4405 7690 4410 7710
rect 4410 7690 4430 7710
rect 4430 7690 4435 7710
rect 4405 7685 4435 7690
rect 4405 7630 4435 7635
rect 4405 7610 4410 7630
rect 4410 7610 4430 7630
rect 4430 7610 4435 7630
rect 4405 7605 4435 7610
rect 4405 7550 4435 7555
rect 4405 7530 4410 7550
rect 4410 7530 4430 7550
rect 4430 7530 4435 7550
rect 4405 7525 4435 7530
rect 4405 7470 4435 7475
rect 4405 7450 4410 7470
rect 4410 7450 4430 7470
rect 4430 7450 4435 7470
rect 4405 7445 4435 7450
rect 4405 7390 4435 7395
rect 4405 7370 4410 7390
rect 4410 7370 4430 7390
rect 4430 7370 4435 7390
rect 4405 7365 4435 7370
rect 4405 7310 4435 7315
rect 4405 7290 4410 7310
rect 4410 7290 4430 7310
rect 4430 7290 4435 7310
rect 4405 7285 4435 7290
rect 4405 7230 4435 7235
rect 4405 7210 4410 7230
rect 4410 7210 4430 7230
rect 4430 7210 4435 7230
rect 4405 7205 4435 7210
rect 4405 7150 4435 7155
rect 4405 7130 4410 7150
rect 4410 7130 4430 7150
rect 4430 7130 4435 7150
rect 4405 7125 4435 7130
rect 4405 7070 4435 7075
rect 4405 7050 4410 7070
rect 4410 7050 4430 7070
rect 4430 7050 4435 7070
rect 4405 7045 4435 7050
rect 4405 6990 4435 6995
rect 4405 6970 4410 6990
rect 4410 6970 4430 6990
rect 4430 6970 4435 6990
rect 4405 6965 4435 6970
rect 4405 6830 4435 6835
rect 4405 6810 4410 6830
rect 4410 6810 4430 6830
rect 4430 6810 4435 6830
rect 4405 6805 4435 6810
rect 4405 6750 4435 6755
rect 4405 6730 4410 6750
rect 4410 6730 4430 6750
rect 4430 6730 4435 6750
rect 4405 6725 4435 6730
rect 4405 6670 4435 6675
rect 4405 6650 4410 6670
rect 4410 6650 4430 6670
rect 4430 6650 4435 6670
rect 4405 6645 4435 6650
rect 4405 6590 4435 6595
rect 4405 6570 4410 6590
rect 4410 6570 4430 6590
rect 4430 6570 4435 6590
rect 4405 6565 4435 6570
rect 4405 6510 4435 6515
rect 4405 6490 4410 6510
rect 4410 6490 4430 6510
rect 4430 6490 4435 6510
rect 4405 6485 4435 6490
rect 4405 6430 4435 6435
rect 4405 6410 4410 6430
rect 4410 6410 4430 6430
rect 4430 6410 4435 6430
rect 4405 6405 4435 6410
rect 4405 6350 4435 6355
rect 4405 6330 4410 6350
rect 4410 6330 4430 6350
rect 4430 6330 4435 6350
rect 4405 6325 4435 6330
rect 4405 6270 4435 6275
rect 4405 6250 4410 6270
rect 4410 6250 4430 6270
rect 4430 6250 4435 6270
rect 4405 6245 4435 6250
rect 4405 5870 4435 5875
rect 4405 5850 4410 5870
rect 4410 5850 4430 5870
rect 4430 5850 4435 5870
rect 4405 5845 4435 5850
rect 4405 5790 4435 5795
rect 4405 5770 4410 5790
rect 4410 5770 4430 5790
rect 4430 5770 4435 5790
rect 4405 5765 4435 5770
rect 4405 5710 4435 5715
rect 4405 5690 4410 5710
rect 4410 5690 4430 5710
rect 4430 5690 4435 5710
rect 4405 5685 4435 5690
rect 4405 5630 4435 5635
rect 4405 5610 4410 5630
rect 4410 5610 4430 5630
rect 4430 5610 4435 5630
rect 4405 5605 4435 5610
rect 4405 5550 4435 5555
rect 4405 5530 4410 5550
rect 4410 5530 4430 5550
rect 4430 5530 4435 5550
rect 4405 5525 4435 5530
rect 4405 5470 4435 5475
rect 4405 5450 4410 5470
rect 4410 5450 4430 5470
rect 4430 5450 4435 5470
rect 4405 5445 4435 5450
rect 4405 5390 4435 5395
rect 4405 5370 4410 5390
rect 4410 5370 4430 5390
rect 4430 5370 4435 5390
rect 4405 5365 4435 5370
rect 4405 5310 4435 5315
rect 4405 5290 4410 5310
rect 4410 5290 4430 5310
rect 4430 5290 4435 5310
rect 4405 5285 4435 5290
rect 4405 5230 4435 5235
rect 4405 5210 4410 5230
rect 4410 5210 4430 5230
rect 4430 5210 4435 5230
rect 4405 5205 4435 5210
rect 4405 5150 4435 5155
rect 4405 5130 4410 5150
rect 4410 5130 4430 5150
rect 4430 5130 4435 5150
rect 4405 5125 4435 5130
rect 4405 5070 4435 5075
rect 4405 5050 4410 5070
rect 4410 5050 4430 5070
rect 4430 5050 4435 5070
rect 4405 5045 4435 5050
rect 4405 4990 4435 4995
rect 4405 4970 4410 4990
rect 4410 4970 4430 4990
rect 4430 4970 4435 4990
rect 4405 4965 4435 4970
rect 4405 4910 4435 4915
rect 4405 4890 4410 4910
rect 4410 4890 4430 4910
rect 4430 4890 4435 4910
rect 4405 4885 4435 4890
rect 4405 4750 4435 4755
rect 4405 4730 4410 4750
rect 4410 4730 4430 4750
rect 4430 4730 4435 4750
rect 4405 4725 4435 4730
rect 4405 4670 4435 4675
rect 4405 4650 4410 4670
rect 4410 4650 4430 4670
rect 4430 4650 4435 4670
rect 4405 4645 4435 4650
rect 4405 4510 4435 4515
rect 4405 4490 4410 4510
rect 4410 4490 4430 4510
rect 4430 4490 4435 4510
rect 4405 4485 4435 4490
rect 4405 4430 4435 4435
rect 4405 4410 4410 4430
rect 4410 4410 4430 4430
rect 4430 4410 4435 4430
rect 4405 4405 4435 4410
rect 4405 4350 4435 4355
rect 4405 4330 4410 4350
rect 4410 4330 4430 4350
rect 4430 4330 4435 4350
rect 4405 4325 4435 4330
rect 4405 4270 4435 4275
rect 4405 4250 4410 4270
rect 4410 4250 4430 4270
rect 4430 4250 4435 4270
rect 4405 4245 4435 4250
rect 4405 4190 4435 4195
rect 4405 4170 4410 4190
rect 4410 4170 4430 4190
rect 4430 4170 4435 4190
rect 4405 4165 4435 4170
rect 4405 4110 4435 4115
rect 4405 4090 4410 4110
rect 4410 4090 4430 4110
rect 4430 4090 4435 4110
rect 4405 4085 4435 4090
rect 4405 4030 4435 4035
rect 4405 4010 4410 4030
rect 4410 4010 4430 4030
rect 4430 4010 4435 4030
rect 4405 4005 4435 4010
rect 4405 3950 4435 3955
rect 4405 3930 4410 3950
rect 4410 3930 4430 3950
rect 4430 3930 4435 3950
rect 4405 3925 4435 3930
rect 4405 3870 4435 3875
rect 4405 3850 4410 3870
rect 4410 3850 4430 3870
rect 4430 3850 4435 3870
rect 4405 3845 4435 3850
rect 4405 3710 4435 3715
rect 4405 3690 4410 3710
rect 4410 3690 4430 3710
rect 4430 3690 4435 3710
rect 4405 3685 4435 3690
rect 4405 3630 4435 3635
rect 4405 3610 4410 3630
rect 4410 3610 4430 3630
rect 4430 3610 4435 3630
rect 4405 3605 4435 3610
rect 4405 3470 4435 3475
rect 4405 3450 4410 3470
rect 4410 3450 4430 3470
rect 4430 3450 4435 3470
rect 4405 3445 4435 3450
rect 4405 3390 4435 3395
rect 4405 3370 4410 3390
rect 4410 3370 4430 3390
rect 4430 3370 4435 3390
rect 4405 3365 4435 3370
rect 4405 3230 4435 3235
rect 4405 3210 4410 3230
rect 4410 3210 4430 3230
rect 4430 3210 4435 3230
rect 4405 3205 4435 3210
rect 4405 3150 4435 3155
rect 4405 3130 4410 3150
rect 4410 3130 4430 3150
rect 4430 3130 4435 3150
rect 4405 3125 4435 3130
rect 4405 3070 4435 3075
rect 4405 3050 4410 3070
rect 4410 3050 4430 3070
rect 4430 3050 4435 3070
rect 4405 3045 4435 3050
rect 4405 2990 4435 2995
rect 4405 2970 4410 2990
rect 4410 2970 4430 2990
rect 4430 2970 4435 2990
rect 4405 2965 4435 2970
rect 4405 2910 4435 2915
rect 4405 2890 4410 2910
rect 4410 2890 4430 2910
rect 4430 2890 4435 2910
rect 4405 2885 4435 2890
rect 4405 2830 4435 2835
rect 4405 2810 4410 2830
rect 4410 2810 4430 2830
rect 4430 2810 4435 2830
rect 4405 2805 4435 2810
rect 4405 2750 4435 2755
rect 4405 2730 4410 2750
rect 4410 2730 4430 2750
rect 4430 2730 4435 2750
rect 4405 2725 4435 2730
rect 4405 2670 4435 2675
rect 4405 2650 4410 2670
rect 4410 2650 4430 2670
rect 4430 2650 4435 2670
rect 4405 2645 4435 2650
rect 4405 2590 4435 2595
rect 4405 2570 4410 2590
rect 4410 2570 4430 2590
rect 4430 2570 4435 2590
rect 4405 2565 4435 2570
rect 4405 2510 4435 2515
rect 4405 2490 4410 2510
rect 4410 2490 4430 2510
rect 4430 2490 4435 2510
rect 4405 2485 4435 2490
rect 4405 2430 4435 2435
rect 4405 2410 4410 2430
rect 4410 2410 4430 2430
rect 4430 2410 4435 2430
rect 4405 2405 4435 2410
rect 4405 2350 4435 2355
rect 4405 2330 4410 2350
rect 4410 2330 4430 2350
rect 4430 2330 4435 2350
rect 4405 2325 4435 2330
rect 4405 2270 4435 2275
rect 4405 2250 4410 2270
rect 4410 2250 4430 2270
rect 4430 2250 4435 2270
rect 4405 2245 4435 2250
rect 4405 2190 4435 2195
rect 4405 2170 4410 2190
rect 4410 2170 4430 2190
rect 4430 2170 4435 2190
rect 4405 2165 4435 2170
rect 4405 2110 4435 2115
rect 4405 2090 4410 2110
rect 4410 2090 4430 2110
rect 4430 2090 4435 2110
rect 4405 2085 4435 2090
rect 4405 2030 4435 2035
rect 4405 2010 4410 2030
rect 4410 2010 4430 2030
rect 4430 2010 4435 2030
rect 4405 2005 4435 2010
rect 4405 1950 4435 1955
rect 4405 1930 4410 1950
rect 4410 1930 4430 1950
rect 4430 1930 4435 1950
rect 4405 1925 4435 1930
rect 4405 1710 4435 1715
rect 4405 1690 4410 1710
rect 4410 1690 4430 1710
rect 4430 1690 4435 1710
rect 4405 1685 4435 1690
rect 4405 1630 4435 1635
rect 4405 1610 4410 1630
rect 4410 1610 4430 1630
rect 4430 1610 4435 1630
rect 4405 1605 4435 1610
rect 4405 1550 4435 1555
rect 4405 1530 4410 1550
rect 4410 1530 4430 1550
rect 4430 1530 4435 1550
rect 4405 1525 4435 1530
rect 4405 1470 4435 1475
rect 4405 1450 4410 1470
rect 4410 1450 4430 1470
rect 4430 1450 4435 1470
rect 4405 1445 4435 1450
rect 4405 1390 4435 1395
rect 4405 1370 4410 1390
rect 4410 1370 4430 1390
rect 4430 1370 4435 1390
rect 4405 1365 4435 1370
rect 4405 1310 4435 1315
rect 4405 1290 4410 1310
rect 4410 1290 4430 1310
rect 4430 1290 4435 1310
rect 4405 1285 4435 1290
rect 4405 1230 4435 1235
rect 4405 1210 4410 1230
rect 4410 1210 4430 1230
rect 4430 1210 4435 1230
rect 4405 1205 4435 1210
rect 4405 1150 4435 1155
rect 4405 1130 4410 1150
rect 4410 1130 4430 1150
rect 4430 1130 4435 1150
rect 4405 1125 4435 1130
rect 4405 1070 4435 1075
rect 4405 1050 4410 1070
rect 4410 1050 4430 1070
rect 4430 1050 4435 1070
rect 4405 1045 4435 1050
rect 4405 990 4435 995
rect 4405 970 4410 990
rect 4410 970 4430 990
rect 4430 970 4435 990
rect 4405 965 4435 970
rect 4405 830 4435 835
rect 4405 810 4410 830
rect 4410 810 4430 830
rect 4430 810 4435 830
rect 4405 805 4435 810
rect 4405 750 4435 755
rect 4405 730 4410 750
rect 4410 730 4430 750
rect 4430 730 4435 750
rect 4405 725 4435 730
rect 4405 670 4435 675
rect 4405 650 4410 670
rect 4410 650 4430 670
rect 4430 650 4435 670
rect 4405 645 4435 650
rect 4405 590 4435 595
rect 4405 570 4410 590
rect 4410 570 4430 590
rect 4430 570 4435 590
rect 4405 565 4435 570
rect 4405 510 4435 515
rect 4405 490 4410 510
rect 4410 490 4430 510
rect 4430 490 4435 510
rect 4405 485 4435 490
rect 4405 270 4435 275
rect 4405 250 4410 270
rect 4410 250 4430 270
rect 4430 250 4435 270
rect 4405 245 4435 250
rect 4405 190 4435 195
rect 4405 170 4410 190
rect 4410 170 4430 190
rect 4430 170 4435 190
rect 4405 165 4435 170
rect 4405 110 4435 115
rect 4405 90 4410 110
rect 4410 90 4430 110
rect 4430 90 4435 110
rect 4405 85 4435 90
rect 4405 30 4435 35
rect 4405 10 4410 30
rect 4410 10 4430 30
rect 4430 10 4435 30
rect 4405 5 4435 10
rect 4485 15710 4515 15715
rect 4485 15690 4490 15710
rect 4490 15690 4510 15710
rect 4510 15690 4515 15710
rect 4485 15685 4515 15690
rect 4485 15630 4515 15635
rect 4485 15610 4490 15630
rect 4490 15610 4510 15630
rect 4510 15610 4515 15630
rect 4485 15605 4515 15610
rect 4485 15550 4515 15555
rect 4485 15530 4490 15550
rect 4490 15530 4510 15550
rect 4510 15530 4515 15550
rect 4485 15525 4515 15530
rect 4485 15470 4515 15475
rect 4485 15450 4490 15470
rect 4490 15450 4510 15470
rect 4510 15450 4515 15470
rect 4485 15445 4515 15450
rect 4485 15390 4515 15395
rect 4485 15370 4490 15390
rect 4490 15370 4510 15390
rect 4510 15370 4515 15390
rect 4485 15365 4515 15370
rect 4485 15310 4515 15315
rect 4485 15290 4490 15310
rect 4490 15290 4510 15310
rect 4510 15290 4515 15310
rect 4485 15285 4515 15290
rect 4485 15230 4515 15235
rect 4485 15210 4490 15230
rect 4490 15210 4510 15230
rect 4510 15210 4515 15230
rect 4485 15205 4515 15210
rect 4485 15150 4515 15155
rect 4485 15130 4490 15150
rect 4490 15130 4510 15150
rect 4510 15130 4515 15150
rect 4485 15125 4515 15130
rect 4485 14990 4515 14995
rect 4485 14970 4490 14990
rect 4490 14970 4510 14990
rect 4510 14970 4515 14990
rect 4485 14965 4515 14970
rect 4485 14910 4515 14915
rect 4485 14890 4490 14910
rect 4490 14890 4510 14910
rect 4510 14890 4515 14910
rect 4485 14885 4515 14890
rect 4485 14830 4515 14835
rect 4485 14810 4490 14830
rect 4490 14810 4510 14830
rect 4510 14810 4515 14830
rect 4485 14805 4515 14810
rect 4485 14750 4515 14755
rect 4485 14730 4490 14750
rect 4490 14730 4510 14750
rect 4510 14730 4515 14750
rect 4485 14725 4515 14730
rect 4485 14670 4515 14675
rect 4485 14650 4490 14670
rect 4490 14650 4510 14670
rect 4510 14650 4515 14670
rect 4485 14645 4515 14650
rect 4485 14590 4515 14595
rect 4485 14570 4490 14590
rect 4490 14570 4510 14590
rect 4510 14570 4515 14590
rect 4485 14565 4515 14570
rect 4485 14510 4515 14515
rect 4485 14490 4490 14510
rect 4490 14490 4510 14510
rect 4510 14490 4515 14510
rect 4485 14485 4515 14490
rect 4485 14430 4515 14435
rect 4485 14410 4490 14430
rect 4490 14410 4510 14430
rect 4510 14410 4515 14430
rect 4485 14405 4515 14410
rect 4485 14030 4515 14035
rect 4485 14010 4490 14030
rect 4490 14010 4510 14030
rect 4510 14010 4515 14030
rect 4485 14005 4515 14010
rect 4485 13950 4515 13955
rect 4485 13930 4490 13950
rect 4490 13930 4510 13950
rect 4510 13930 4515 13950
rect 4485 13925 4515 13930
rect 4485 13870 4515 13875
rect 4485 13850 4490 13870
rect 4490 13850 4510 13870
rect 4510 13850 4515 13870
rect 4485 13845 4515 13850
rect 4485 13790 4515 13795
rect 4485 13770 4490 13790
rect 4490 13770 4510 13790
rect 4510 13770 4515 13790
rect 4485 13765 4515 13770
rect 4485 13710 4515 13715
rect 4485 13690 4490 13710
rect 4490 13690 4510 13710
rect 4510 13690 4515 13710
rect 4485 13685 4515 13690
rect 4485 13630 4515 13635
rect 4485 13610 4490 13630
rect 4490 13610 4510 13630
rect 4510 13610 4515 13630
rect 4485 13605 4515 13610
rect 4485 13550 4515 13555
rect 4485 13530 4490 13550
rect 4490 13530 4510 13550
rect 4510 13530 4515 13550
rect 4485 13525 4515 13530
rect 4485 13470 4515 13475
rect 4485 13450 4490 13470
rect 4490 13450 4510 13470
rect 4510 13450 4515 13470
rect 4485 13445 4515 13450
rect 4485 13070 4515 13075
rect 4485 13050 4490 13070
rect 4490 13050 4510 13070
rect 4510 13050 4515 13070
rect 4485 13045 4515 13050
rect 4485 12990 4515 12995
rect 4485 12970 4490 12990
rect 4490 12970 4510 12990
rect 4510 12970 4515 12990
rect 4485 12965 4515 12970
rect 4485 12910 4515 12915
rect 4485 12890 4490 12910
rect 4490 12890 4510 12910
rect 4510 12890 4515 12910
rect 4485 12885 4515 12890
rect 4485 12830 4515 12835
rect 4485 12810 4490 12830
rect 4490 12810 4510 12830
rect 4510 12810 4515 12830
rect 4485 12805 4515 12810
rect 4485 12750 4515 12755
rect 4485 12730 4490 12750
rect 4490 12730 4510 12750
rect 4510 12730 4515 12750
rect 4485 12725 4515 12730
rect 4485 12670 4515 12675
rect 4485 12650 4490 12670
rect 4490 12650 4510 12670
rect 4510 12650 4515 12670
rect 4485 12645 4515 12650
rect 4485 12590 4515 12595
rect 4485 12570 4490 12590
rect 4490 12570 4510 12590
rect 4510 12570 4515 12590
rect 4485 12565 4515 12570
rect 4485 12510 4515 12515
rect 4485 12490 4490 12510
rect 4490 12490 4510 12510
rect 4510 12490 4515 12510
rect 4485 12485 4515 12490
rect 4485 12350 4515 12355
rect 4485 12330 4490 12350
rect 4490 12330 4510 12350
rect 4510 12330 4515 12350
rect 4485 12325 4515 12330
rect 4485 12270 4515 12275
rect 4485 12250 4490 12270
rect 4490 12250 4510 12270
rect 4510 12250 4515 12270
rect 4485 12245 4515 12250
rect 4485 12190 4515 12195
rect 4485 12170 4490 12190
rect 4490 12170 4510 12190
rect 4510 12170 4515 12190
rect 4485 12165 4515 12170
rect 4485 12110 4515 12115
rect 4485 12090 4490 12110
rect 4490 12090 4510 12110
rect 4510 12090 4515 12110
rect 4485 12085 4515 12090
rect 4485 12030 4515 12035
rect 4485 12010 4490 12030
rect 4490 12010 4510 12030
rect 4510 12010 4515 12030
rect 4485 12005 4515 12010
rect 4485 11950 4515 11955
rect 4485 11930 4490 11950
rect 4490 11930 4510 11950
rect 4510 11930 4515 11950
rect 4485 11925 4515 11930
rect 4485 11870 4515 11875
rect 4485 11850 4490 11870
rect 4490 11850 4510 11870
rect 4510 11850 4515 11870
rect 4485 11845 4515 11850
rect 4485 11790 4515 11795
rect 4485 11770 4490 11790
rect 4490 11770 4510 11790
rect 4510 11770 4515 11790
rect 4485 11765 4515 11770
rect 4485 11710 4515 11715
rect 4485 11690 4490 11710
rect 4490 11690 4510 11710
rect 4510 11690 4515 11710
rect 4485 11685 4515 11690
rect 4485 11630 4515 11635
rect 4485 11610 4490 11630
rect 4490 11610 4510 11630
rect 4510 11610 4515 11630
rect 4485 11605 4515 11610
rect 4485 11550 4515 11555
rect 4485 11530 4490 11550
rect 4490 11530 4510 11550
rect 4510 11530 4515 11550
rect 4485 11525 4515 11530
rect 4485 11470 4515 11475
rect 4485 11450 4490 11470
rect 4490 11450 4510 11470
rect 4510 11450 4515 11470
rect 4485 11445 4515 11450
rect 4485 11390 4515 11395
rect 4485 11370 4490 11390
rect 4490 11370 4510 11390
rect 4510 11370 4515 11390
rect 4485 11365 4515 11370
rect 4485 11310 4515 11315
rect 4485 11290 4490 11310
rect 4490 11290 4510 11310
rect 4510 11290 4515 11310
rect 4485 11285 4515 11290
rect 4485 11230 4515 11235
rect 4485 11210 4490 11230
rect 4490 11210 4510 11230
rect 4510 11210 4515 11230
rect 4485 11205 4515 11210
rect 4485 11150 4515 11155
rect 4485 11130 4490 11150
rect 4490 11130 4510 11150
rect 4510 11130 4515 11150
rect 4485 11125 4515 11130
rect 4485 11070 4515 11075
rect 4485 11050 4490 11070
rect 4490 11050 4510 11070
rect 4510 11050 4515 11070
rect 4485 11045 4515 11050
rect 4485 10910 4515 10915
rect 4485 10890 4490 10910
rect 4490 10890 4510 10910
rect 4510 10890 4515 10910
rect 4485 10885 4515 10890
rect 4485 10830 4515 10835
rect 4485 10810 4490 10830
rect 4490 10810 4510 10830
rect 4510 10810 4515 10830
rect 4485 10805 4515 10810
rect 4485 10750 4515 10755
rect 4485 10730 4490 10750
rect 4490 10730 4510 10750
rect 4510 10730 4515 10750
rect 4485 10725 4515 10730
rect 4485 10670 4515 10675
rect 4485 10650 4490 10670
rect 4490 10650 4510 10670
rect 4510 10650 4515 10670
rect 4485 10645 4515 10650
rect 4485 10590 4515 10595
rect 4485 10570 4490 10590
rect 4490 10570 4510 10590
rect 4510 10570 4515 10590
rect 4485 10565 4515 10570
rect 4485 10510 4515 10515
rect 4485 10490 4490 10510
rect 4490 10490 4510 10510
rect 4510 10490 4515 10510
rect 4485 10485 4515 10490
rect 4485 10430 4515 10435
rect 4485 10410 4490 10430
rect 4490 10410 4510 10430
rect 4510 10410 4515 10430
rect 4485 10405 4515 10410
rect 4485 10350 4515 10355
rect 4485 10330 4490 10350
rect 4490 10330 4510 10350
rect 4510 10330 4515 10350
rect 4485 10325 4515 10330
rect 4485 9950 4515 9955
rect 4485 9930 4490 9950
rect 4490 9930 4510 9950
rect 4510 9930 4515 9950
rect 4485 9925 4515 9930
rect 4485 9870 4515 9875
rect 4485 9850 4490 9870
rect 4490 9850 4510 9870
rect 4510 9850 4515 9870
rect 4485 9845 4515 9850
rect 4485 9790 4515 9795
rect 4485 9770 4490 9790
rect 4490 9770 4510 9790
rect 4510 9770 4515 9790
rect 4485 9765 4515 9770
rect 4485 9710 4515 9715
rect 4485 9690 4490 9710
rect 4490 9690 4510 9710
rect 4510 9690 4515 9710
rect 4485 9685 4515 9690
rect 4485 9630 4515 9635
rect 4485 9610 4490 9630
rect 4490 9610 4510 9630
rect 4510 9610 4515 9630
rect 4485 9605 4515 9610
rect 4485 9550 4515 9555
rect 4485 9530 4490 9550
rect 4490 9530 4510 9550
rect 4510 9530 4515 9550
rect 4485 9525 4515 9530
rect 4485 9470 4515 9475
rect 4485 9450 4490 9470
rect 4490 9450 4510 9470
rect 4510 9450 4515 9470
rect 4485 9445 4515 9450
rect 4485 9390 4515 9395
rect 4485 9370 4490 9390
rect 4490 9370 4510 9390
rect 4510 9370 4515 9390
rect 4485 9365 4515 9370
rect 4485 8990 4515 8995
rect 4485 8970 4490 8990
rect 4490 8970 4510 8990
rect 4510 8970 4515 8990
rect 4485 8965 4515 8970
rect 4485 8910 4515 8915
rect 4485 8890 4490 8910
rect 4490 8890 4510 8910
rect 4510 8890 4515 8910
rect 4485 8885 4515 8890
rect 4485 8830 4515 8835
rect 4485 8810 4490 8830
rect 4490 8810 4510 8830
rect 4510 8810 4515 8830
rect 4485 8805 4515 8810
rect 4485 8750 4515 8755
rect 4485 8730 4490 8750
rect 4490 8730 4510 8750
rect 4510 8730 4515 8750
rect 4485 8725 4515 8730
rect 4485 8670 4515 8675
rect 4485 8650 4490 8670
rect 4490 8650 4510 8670
rect 4510 8650 4515 8670
rect 4485 8645 4515 8650
rect 4485 8590 4515 8595
rect 4485 8570 4490 8590
rect 4490 8570 4510 8590
rect 4510 8570 4515 8590
rect 4485 8565 4515 8570
rect 4485 8510 4515 8515
rect 4485 8490 4490 8510
rect 4490 8490 4510 8510
rect 4510 8490 4515 8510
rect 4485 8485 4515 8490
rect 4485 8430 4515 8435
rect 4485 8410 4490 8430
rect 4490 8410 4510 8430
rect 4510 8410 4515 8430
rect 4485 8405 4515 8410
rect 4485 8270 4515 8275
rect 4485 8250 4490 8270
rect 4490 8250 4510 8270
rect 4510 8250 4515 8270
rect 4485 8245 4515 8250
rect 4485 8190 4515 8195
rect 4485 8170 4490 8190
rect 4490 8170 4510 8190
rect 4510 8170 4515 8190
rect 4485 8165 4515 8170
rect 4485 8110 4515 8115
rect 4485 8090 4490 8110
rect 4490 8090 4510 8110
rect 4510 8090 4515 8110
rect 4485 8085 4515 8090
rect 4485 8030 4515 8035
rect 4485 8010 4490 8030
rect 4490 8010 4510 8030
rect 4510 8010 4515 8030
rect 4485 8005 4515 8010
rect 4485 7950 4515 7955
rect 4485 7930 4490 7950
rect 4490 7930 4510 7950
rect 4510 7930 4515 7950
rect 4485 7925 4515 7930
rect 4485 7870 4515 7875
rect 4485 7850 4490 7870
rect 4490 7850 4510 7870
rect 4510 7850 4515 7870
rect 4485 7845 4515 7850
rect 4485 7790 4515 7795
rect 4485 7770 4490 7790
rect 4490 7770 4510 7790
rect 4510 7770 4515 7790
rect 4485 7765 4515 7770
rect 4485 7710 4515 7715
rect 4485 7690 4490 7710
rect 4490 7690 4510 7710
rect 4510 7690 4515 7710
rect 4485 7685 4515 7690
rect 4485 7630 4515 7635
rect 4485 7610 4490 7630
rect 4490 7610 4510 7630
rect 4510 7610 4515 7630
rect 4485 7605 4515 7610
rect 4485 7550 4515 7555
rect 4485 7530 4490 7550
rect 4490 7530 4510 7550
rect 4510 7530 4515 7550
rect 4485 7525 4515 7530
rect 4485 7470 4515 7475
rect 4485 7450 4490 7470
rect 4490 7450 4510 7470
rect 4510 7450 4515 7470
rect 4485 7445 4515 7450
rect 4485 7390 4515 7395
rect 4485 7370 4490 7390
rect 4490 7370 4510 7390
rect 4510 7370 4515 7390
rect 4485 7365 4515 7370
rect 4485 7310 4515 7315
rect 4485 7290 4490 7310
rect 4490 7290 4510 7310
rect 4510 7290 4515 7310
rect 4485 7285 4515 7290
rect 4485 7230 4515 7235
rect 4485 7210 4490 7230
rect 4490 7210 4510 7230
rect 4510 7210 4515 7230
rect 4485 7205 4515 7210
rect 4485 7150 4515 7155
rect 4485 7130 4490 7150
rect 4490 7130 4510 7150
rect 4510 7130 4515 7150
rect 4485 7125 4515 7130
rect 4485 7070 4515 7075
rect 4485 7050 4490 7070
rect 4490 7050 4510 7070
rect 4510 7050 4515 7070
rect 4485 7045 4515 7050
rect 4485 6990 4515 6995
rect 4485 6970 4490 6990
rect 4490 6970 4510 6990
rect 4510 6970 4515 6990
rect 4485 6965 4515 6970
rect 4485 6830 4515 6835
rect 4485 6810 4490 6830
rect 4490 6810 4510 6830
rect 4510 6810 4515 6830
rect 4485 6805 4515 6810
rect 4485 6750 4515 6755
rect 4485 6730 4490 6750
rect 4490 6730 4510 6750
rect 4510 6730 4515 6750
rect 4485 6725 4515 6730
rect 4485 6670 4515 6675
rect 4485 6650 4490 6670
rect 4490 6650 4510 6670
rect 4510 6650 4515 6670
rect 4485 6645 4515 6650
rect 4485 6590 4515 6595
rect 4485 6570 4490 6590
rect 4490 6570 4510 6590
rect 4510 6570 4515 6590
rect 4485 6565 4515 6570
rect 4485 6510 4515 6515
rect 4485 6490 4490 6510
rect 4490 6490 4510 6510
rect 4510 6490 4515 6510
rect 4485 6485 4515 6490
rect 4485 6430 4515 6435
rect 4485 6410 4490 6430
rect 4490 6410 4510 6430
rect 4510 6410 4515 6430
rect 4485 6405 4515 6410
rect 4485 6350 4515 6355
rect 4485 6330 4490 6350
rect 4490 6330 4510 6350
rect 4510 6330 4515 6350
rect 4485 6325 4515 6330
rect 4485 6270 4515 6275
rect 4485 6250 4490 6270
rect 4490 6250 4510 6270
rect 4510 6250 4515 6270
rect 4485 6245 4515 6250
rect 4485 5870 4515 5875
rect 4485 5850 4490 5870
rect 4490 5850 4510 5870
rect 4510 5850 4515 5870
rect 4485 5845 4515 5850
rect 4485 5790 4515 5795
rect 4485 5770 4490 5790
rect 4490 5770 4510 5790
rect 4510 5770 4515 5790
rect 4485 5765 4515 5770
rect 4485 5710 4515 5715
rect 4485 5690 4490 5710
rect 4490 5690 4510 5710
rect 4510 5690 4515 5710
rect 4485 5685 4515 5690
rect 4485 5630 4515 5635
rect 4485 5610 4490 5630
rect 4490 5610 4510 5630
rect 4510 5610 4515 5630
rect 4485 5605 4515 5610
rect 4485 5550 4515 5555
rect 4485 5530 4490 5550
rect 4490 5530 4510 5550
rect 4510 5530 4515 5550
rect 4485 5525 4515 5530
rect 4485 5470 4515 5475
rect 4485 5450 4490 5470
rect 4490 5450 4510 5470
rect 4510 5450 4515 5470
rect 4485 5445 4515 5450
rect 4485 5390 4515 5395
rect 4485 5370 4490 5390
rect 4490 5370 4510 5390
rect 4510 5370 4515 5390
rect 4485 5365 4515 5370
rect 4485 5310 4515 5315
rect 4485 5290 4490 5310
rect 4490 5290 4510 5310
rect 4510 5290 4515 5310
rect 4485 5285 4515 5290
rect 4485 5230 4515 5235
rect 4485 5210 4490 5230
rect 4490 5210 4510 5230
rect 4510 5210 4515 5230
rect 4485 5205 4515 5210
rect 4485 5150 4515 5155
rect 4485 5130 4490 5150
rect 4490 5130 4510 5150
rect 4510 5130 4515 5150
rect 4485 5125 4515 5130
rect 4485 5070 4515 5075
rect 4485 5050 4490 5070
rect 4490 5050 4510 5070
rect 4510 5050 4515 5070
rect 4485 5045 4515 5050
rect 4485 4990 4515 4995
rect 4485 4970 4490 4990
rect 4490 4970 4510 4990
rect 4510 4970 4515 4990
rect 4485 4965 4515 4970
rect 4485 4910 4515 4915
rect 4485 4890 4490 4910
rect 4490 4890 4510 4910
rect 4510 4890 4515 4910
rect 4485 4885 4515 4890
rect 4485 4750 4515 4755
rect 4485 4730 4490 4750
rect 4490 4730 4510 4750
rect 4510 4730 4515 4750
rect 4485 4725 4515 4730
rect 4485 4670 4515 4675
rect 4485 4650 4490 4670
rect 4490 4650 4510 4670
rect 4510 4650 4515 4670
rect 4485 4645 4515 4650
rect 4485 4510 4515 4515
rect 4485 4490 4490 4510
rect 4490 4490 4510 4510
rect 4510 4490 4515 4510
rect 4485 4485 4515 4490
rect 4485 4430 4515 4435
rect 4485 4410 4490 4430
rect 4490 4410 4510 4430
rect 4510 4410 4515 4430
rect 4485 4405 4515 4410
rect 4485 4350 4515 4355
rect 4485 4330 4490 4350
rect 4490 4330 4510 4350
rect 4510 4330 4515 4350
rect 4485 4325 4515 4330
rect 4485 4270 4515 4275
rect 4485 4250 4490 4270
rect 4490 4250 4510 4270
rect 4510 4250 4515 4270
rect 4485 4245 4515 4250
rect 4485 4190 4515 4195
rect 4485 4170 4490 4190
rect 4490 4170 4510 4190
rect 4510 4170 4515 4190
rect 4485 4165 4515 4170
rect 4485 4110 4515 4115
rect 4485 4090 4490 4110
rect 4490 4090 4510 4110
rect 4510 4090 4515 4110
rect 4485 4085 4515 4090
rect 4485 4030 4515 4035
rect 4485 4010 4490 4030
rect 4490 4010 4510 4030
rect 4510 4010 4515 4030
rect 4485 4005 4515 4010
rect 4485 3950 4515 3955
rect 4485 3930 4490 3950
rect 4490 3930 4510 3950
rect 4510 3930 4515 3950
rect 4485 3925 4515 3930
rect 4485 3870 4515 3875
rect 4485 3850 4490 3870
rect 4490 3850 4510 3870
rect 4510 3850 4515 3870
rect 4485 3845 4515 3850
rect 4485 3710 4515 3715
rect 4485 3690 4490 3710
rect 4490 3690 4510 3710
rect 4510 3690 4515 3710
rect 4485 3685 4515 3690
rect 4485 3630 4515 3635
rect 4485 3610 4490 3630
rect 4490 3610 4510 3630
rect 4510 3610 4515 3630
rect 4485 3605 4515 3610
rect 4485 3470 4515 3475
rect 4485 3450 4490 3470
rect 4490 3450 4510 3470
rect 4510 3450 4515 3470
rect 4485 3445 4515 3450
rect 4485 3390 4515 3395
rect 4485 3370 4490 3390
rect 4490 3370 4510 3390
rect 4510 3370 4515 3390
rect 4485 3365 4515 3370
rect 4485 3230 4515 3235
rect 4485 3210 4490 3230
rect 4490 3210 4510 3230
rect 4510 3210 4515 3230
rect 4485 3205 4515 3210
rect 4485 3150 4515 3155
rect 4485 3130 4490 3150
rect 4490 3130 4510 3150
rect 4510 3130 4515 3150
rect 4485 3125 4515 3130
rect 4485 3070 4515 3075
rect 4485 3050 4490 3070
rect 4490 3050 4510 3070
rect 4510 3050 4515 3070
rect 4485 3045 4515 3050
rect 4485 2990 4515 2995
rect 4485 2970 4490 2990
rect 4490 2970 4510 2990
rect 4510 2970 4515 2990
rect 4485 2965 4515 2970
rect 4485 2910 4515 2915
rect 4485 2890 4490 2910
rect 4490 2890 4510 2910
rect 4510 2890 4515 2910
rect 4485 2885 4515 2890
rect 4485 2830 4515 2835
rect 4485 2810 4490 2830
rect 4490 2810 4510 2830
rect 4510 2810 4515 2830
rect 4485 2805 4515 2810
rect 4485 2750 4515 2755
rect 4485 2730 4490 2750
rect 4490 2730 4510 2750
rect 4510 2730 4515 2750
rect 4485 2725 4515 2730
rect 4485 2670 4515 2675
rect 4485 2650 4490 2670
rect 4490 2650 4510 2670
rect 4510 2650 4515 2670
rect 4485 2645 4515 2650
rect 4485 2590 4515 2595
rect 4485 2570 4490 2590
rect 4490 2570 4510 2590
rect 4510 2570 4515 2590
rect 4485 2565 4515 2570
rect 4485 2510 4515 2515
rect 4485 2490 4490 2510
rect 4490 2490 4510 2510
rect 4510 2490 4515 2510
rect 4485 2485 4515 2490
rect 4485 2430 4515 2435
rect 4485 2410 4490 2430
rect 4490 2410 4510 2430
rect 4510 2410 4515 2430
rect 4485 2405 4515 2410
rect 4485 2350 4515 2355
rect 4485 2330 4490 2350
rect 4490 2330 4510 2350
rect 4510 2330 4515 2350
rect 4485 2325 4515 2330
rect 4485 2270 4515 2275
rect 4485 2250 4490 2270
rect 4490 2250 4510 2270
rect 4510 2250 4515 2270
rect 4485 2245 4515 2250
rect 4485 2190 4515 2195
rect 4485 2170 4490 2190
rect 4490 2170 4510 2190
rect 4510 2170 4515 2190
rect 4485 2165 4515 2170
rect 4485 2110 4515 2115
rect 4485 2090 4490 2110
rect 4490 2090 4510 2110
rect 4510 2090 4515 2110
rect 4485 2085 4515 2090
rect 4485 2030 4515 2035
rect 4485 2010 4490 2030
rect 4490 2010 4510 2030
rect 4510 2010 4515 2030
rect 4485 2005 4515 2010
rect 4485 1950 4515 1955
rect 4485 1930 4490 1950
rect 4490 1930 4510 1950
rect 4510 1930 4515 1950
rect 4485 1925 4515 1930
rect 4485 1710 4515 1715
rect 4485 1690 4490 1710
rect 4490 1690 4510 1710
rect 4510 1690 4515 1710
rect 4485 1685 4515 1690
rect 4485 1630 4515 1635
rect 4485 1610 4490 1630
rect 4490 1610 4510 1630
rect 4510 1610 4515 1630
rect 4485 1605 4515 1610
rect 4485 1550 4515 1555
rect 4485 1530 4490 1550
rect 4490 1530 4510 1550
rect 4510 1530 4515 1550
rect 4485 1525 4515 1530
rect 4485 1470 4515 1475
rect 4485 1450 4490 1470
rect 4490 1450 4510 1470
rect 4510 1450 4515 1470
rect 4485 1445 4515 1450
rect 4485 1390 4515 1395
rect 4485 1370 4490 1390
rect 4490 1370 4510 1390
rect 4510 1370 4515 1390
rect 4485 1365 4515 1370
rect 4485 1310 4515 1315
rect 4485 1290 4490 1310
rect 4490 1290 4510 1310
rect 4510 1290 4515 1310
rect 4485 1285 4515 1290
rect 4485 1230 4515 1235
rect 4485 1210 4490 1230
rect 4490 1210 4510 1230
rect 4510 1210 4515 1230
rect 4485 1205 4515 1210
rect 4485 1150 4515 1155
rect 4485 1130 4490 1150
rect 4490 1130 4510 1150
rect 4510 1130 4515 1150
rect 4485 1125 4515 1130
rect 4485 1070 4515 1075
rect 4485 1050 4490 1070
rect 4490 1050 4510 1070
rect 4510 1050 4515 1070
rect 4485 1045 4515 1050
rect 4485 990 4515 995
rect 4485 970 4490 990
rect 4490 970 4510 990
rect 4510 970 4515 990
rect 4485 965 4515 970
rect 4485 830 4515 835
rect 4485 810 4490 830
rect 4490 810 4510 830
rect 4510 810 4515 830
rect 4485 805 4515 810
rect 4485 750 4515 755
rect 4485 730 4490 750
rect 4490 730 4510 750
rect 4510 730 4515 750
rect 4485 725 4515 730
rect 4485 670 4515 675
rect 4485 650 4490 670
rect 4490 650 4510 670
rect 4510 650 4515 670
rect 4485 645 4515 650
rect 4485 590 4515 595
rect 4485 570 4490 590
rect 4490 570 4510 590
rect 4510 570 4515 590
rect 4485 565 4515 570
rect 4485 510 4515 515
rect 4485 490 4490 510
rect 4490 490 4510 510
rect 4510 490 4515 510
rect 4485 485 4515 490
rect 4485 270 4515 275
rect 4485 250 4490 270
rect 4490 250 4510 270
rect 4510 250 4515 270
rect 4485 245 4515 250
rect 4485 190 4515 195
rect 4485 170 4490 190
rect 4490 170 4510 190
rect 4510 170 4515 190
rect 4485 165 4515 170
rect 4485 110 4515 115
rect 4485 90 4490 110
rect 4490 90 4510 110
rect 4510 90 4515 110
rect 4485 85 4515 90
rect 4485 30 4515 35
rect 4485 10 4490 30
rect 4490 10 4510 30
rect 4510 10 4515 30
rect 4485 5 4515 10
rect 4645 15710 4675 15715
rect 4645 15690 4650 15710
rect 4650 15690 4670 15710
rect 4670 15690 4675 15710
rect 4645 15685 4675 15690
rect 4645 15630 4675 15635
rect 4645 15610 4650 15630
rect 4650 15610 4670 15630
rect 4670 15610 4675 15630
rect 4645 15605 4675 15610
rect 4645 15550 4675 15555
rect 4645 15530 4650 15550
rect 4650 15530 4670 15550
rect 4670 15530 4675 15550
rect 4645 15525 4675 15530
rect 4645 15470 4675 15475
rect 4645 15450 4650 15470
rect 4650 15450 4670 15470
rect 4670 15450 4675 15470
rect 4645 15445 4675 15450
rect 4645 15390 4675 15395
rect 4645 15370 4650 15390
rect 4650 15370 4670 15390
rect 4670 15370 4675 15390
rect 4645 15365 4675 15370
rect 4645 15310 4675 15315
rect 4645 15290 4650 15310
rect 4650 15290 4670 15310
rect 4670 15290 4675 15310
rect 4645 15285 4675 15290
rect 4645 15230 4675 15235
rect 4645 15210 4650 15230
rect 4650 15210 4670 15230
rect 4670 15210 4675 15230
rect 4645 15205 4675 15210
rect 4645 15150 4675 15155
rect 4645 15130 4650 15150
rect 4650 15130 4670 15150
rect 4670 15130 4675 15150
rect 4645 15125 4675 15130
rect 4645 14990 4675 14995
rect 4645 14970 4650 14990
rect 4650 14970 4670 14990
rect 4670 14970 4675 14990
rect 4645 14965 4675 14970
rect 4645 14910 4675 14915
rect 4645 14890 4650 14910
rect 4650 14890 4670 14910
rect 4670 14890 4675 14910
rect 4645 14885 4675 14890
rect 4645 14830 4675 14835
rect 4645 14810 4650 14830
rect 4650 14810 4670 14830
rect 4670 14810 4675 14830
rect 4645 14805 4675 14810
rect 4645 14750 4675 14755
rect 4645 14730 4650 14750
rect 4650 14730 4670 14750
rect 4670 14730 4675 14750
rect 4645 14725 4675 14730
rect 4645 14670 4675 14675
rect 4645 14650 4650 14670
rect 4650 14650 4670 14670
rect 4670 14650 4675 14670
rect 4645 14645 4675 14650
rect 4645 14590 4675 14595
rect 4645 14570 4650 14590
rect 4650 14570 4670 14590
rect 4670 14570 4675 14590
rect 4645 14565 4675 14570
rect 4645 14510 4675 14515
rect 4645 14490 4650 14510
rect 4650 14490 4670 14510
rect 4670 14490 4675 14510
rect 4645 14485 4675 14490
rect 4645 14430 4675 14435
rect 4645 14410 4650 14430
rect 4650 14410 4670 14430
rect 4670 14410 4675 14430
rect 4645 14405 4675 14410
rect 4645 14030 4675 14035
rect 4645 14010 4650 14030
rect 4650 14010 4670 14030
rect 4670 14010 4675 14030
rect 4645 14005 4675 14010
rect 4645 13950 4675 13955
rect 4645 13930 4650 13950
rect 4650 13930 4670 13950
rect 4670 13930 4675 13950
rect 4645 13925 4675 13930
rect 4645 13870 4675 13875
rect 4645 13850 4650 13870
rect 4650 13850 4670 13870
rect 4670 13850 4675 13870
rect 4645 13845 4675 13850
rect 4645 13790 4675 13795
rect 4645 13770 4650 13790
rect 4650 13770 4670 13790
rect 4670 13770 4675 13790
rect 4645 13765 4675 13770
rect 4645 13710 4675 13715
rect 4645 13690 4650 13710
rect 4650 13690 4670 13710
rect 4670 13690 4675 13710
rect 4645 13685 4675 13690
rect 4645 13630 4675 13635
rect 4645 13610 4650 13630
rect 4650 13610 4670 13630
rect 4670 13610 4675 13630
rect 4645 13605 4675 13610
rect 4645 13550 4675 13555
rect 4645 13530 4650 13550
rect 4650 13530 4670 13550
rect 4670 13530 4675 13550
rect 4645 13525 4675 13530
rect 4645 13470 4675 13475
rect 4645 13450 4650 13470
rect 4650 13450 4670 13470
rect 4670 13450 4675 13470
rect 4645 13445 4675 13450
rect 4645 13070 4675 13075
rect 4645 13050 4650 13070
rect 4650 13050 4670 13070
rect 4670 13050 4675 13070
rect 4645 13045 4675 13050
rect 4645 12990 4675 12995
rect 4645 12970 4650 12990
rect 4650 12970 4670 12990
rect 4670 12970 4675 12990
rect 4645 12965 4675 12970
rect 4645 12910 4675 12915
rect 4645 12890 4650 12910
rect 4650 12890 4670 12910
rect 4670 12890 4675 12910
rect 4645 12885 4675 12890
rect 4645 12830 4675 12835
rect 4645 12810 4650 12830
rect 4650 12810 4670 12830
rect 4670 12810 4675 12830
rect 4645 12805 4675 12810
rect 4645 12750 4675 12755
rect 4645 12730 4650 12750
rect 4650 12730 4670 12750
rect 4670 12730 4675 12750
rect 4645 12725 4675 12730
rect 4645 12670 4675 12675
rect 4645 12650 4650 12670
rect 4650 12650 4670 12670
rect 4670 12650 4675 12670
rect 4645 12645 4675 12650
rect 4645 12590 4675 12595
rect 4645 12570 4650 12590
rect 4650 12570 4670 12590
rect 4670 12570 4675 12590
rect 4645 12565 4675 12570
rect 4645 12510 4675 12515
rect 4645 12490 4650 12510
rect 4650 12490 4670 12510
rect 4670 12490 4675 12510
rect 4645 12485 4675 12490
rect 4645 12350 4675 12355
rect 4645 12330 4650 12350
rect 4650 12330 4670 12350
rect 4670 12330 4675 12350
rect 4645 12325 4675 12330
rect 4645 12270 4675 12275
rect 4645 12250 4650 12270
rect 4650 12250 4670 12270
rect 4670 12250 4675 12270
rect 4645 12245 4675 12250
rect 4645 12190 4675 12195
rect 4645 12170 4650 12190
rect 4650 12170 4670 12190
rect 4670 12170 4675 12190
rect 4645 12165 4675 12170
rect 4645 12110 4675 12115
rect 4645 12090 4650 12110
rect 4650 12090 4670 12110
rect 4670 12090 4675 12110
rect 4645 12085 4675 12090
rect 4645 12030 4675 12035
rect 4645 12010 4650 12030
rect 4650 12010 4670 12030
rect 4670 12010 4675 12030
rect 4645 12005 4675 12010
rect 4645 11950 4675 11955
rect 4645 11930 4650 11950
rect 4650 11930 4670 11950
rect 4670 11930 4675 11950
rect 4645 11925 4675 11930
rect 4645 11870 4675 11875
rect 4645 11850 4650 11870
rect 4650 11850 4670 11870
rect 4670 11850 4675 11870
rect 4645 11845 4675 11850
rect 4645 11790 4675 11795
rect 4645 11770 4650 11790
rect 4650 11770 4670 11790
rect 4670 11770 4675 11790
rect 4645 11765 4675 11770
rect 4645 11710 4675 11715
rect 4645 11690 4650 11710
rect 4650 11690 4670 11710
rect 4670 11690 4675 11710
rect 4645 11685 4675 11690
rect 4645 11630 4675 11635
rect 4645 11610 4650 11630
rect 4650 11610 4670 11630
rect 4670 11610 4675 11630
rect 4645 11605 4675 11610
rect 4645 11550 4675 11555
rect 4645 11530 4650 11550
rect 4650 11530 4670 11550
rect 4670 11530 4675 11550
rect 4645 11525 4675 11530
rect 4645 11470 4675 11475
rect 4645 11450 4650 11470
rect 4650 11450 4670 11470
rect 4670 11450 4675 11470
rect 4645 11445 4675 11450
rect 4645 11390 4675 11395
rect 4645 11370 4650 11390
rect 4650 11370 4670 11390
rect 4670 11370 4675 11390
rect 4645 11365 4675 11370
rect 4645 11310 4675 11315
rect 4645 11290 4650 11310
rect 4650 11290 4670 11310
rect 4670 11290 4675 11310
rect 4645 11285 4675 11290
rect 4645 11230 4675 11235
rect 4645 11210 4650 11230
rect 4650 11210 4670 11230
rect 4670 11210 4675 11230
rect 4645 11205 4675 11210
rect 4645 11150 4675 11155
rect 4645 11130 4650 11150
rect 4650 11130 4670 11150
rect 4670 11130 4675 11150
rect 4645 11125 4675 11130
rect 4645 11070 4675 11075
rect 4645 11050 4650 11070
rect 4650 11050 4670 11070
rect 4670 11050 4675 11070
rect 4645 11045 4675 11050
rect 4645 10910 4675 10915
rect 4645 10890 4650 10910
rect 4650 10890 4670 10910
rect 4670 10890 4675 10910
rect 4645 10885 4675 10890
rect 4645 10830 4675 10835
rect 4645 10810 4650 10830
rect 4650 10810 4670 10830
rect 4670 10810 4675 10830
rect 4645 10805 4675 10810
rect 4645 10750 4675 10755
rect 4645 10730 4650 10750
rect 4650 10730 4670 10750
rect 4670 10730 4675 10750
rect 4645 10725 4675 10730
rect 4645 10670 4675 10675
rect 4645 10650 4650 10670
rect 4650 10650 4670 10670
rect 4670 10650 4675 10670
rect 4645 10645 4675 10650
rect 4645 10590 4675 10595
rect 4645 10570 4650 10590
rect 4650 10570 4670 10590
rect 4670 10570 4675 10590
rect 4645 10565 4675 10570
rect 4645 10510 4675 10515
rect 4645 10490 4650 10510
rect 4650 10490 4670 10510
rect 4670 10490 4675 10510
rect 4645 10485 4675 10490
rect 4645 10430 4675 10435
rect 4645 10410 4650 10430
rect 4650 10410 4670 10430
rect 4670 10410 4675 10430
rect 4645 10405 4675 10410
rect 4645 10350 4675 10355
rect 4645 10330 4650 10350
rect 4650 10330 4670 10350
rect 4670 10330 4675 10350
rect 4645 10325 4675 10330
rect 4645 9950 4675 9955
rect 4645 9930 4650 9950
rect 4650 9930 4670 9950
rect 4670 9930 4675 9950
rect 4645 9925 4675 9930
rect 4645 9870 4675 9875
rect 4645 9850 4650 9870
rect 4650 9850 4670 9870
rect 4670 9850 4675 9870
rect 4645 9845 4675 9850
rect 4645 9790 4675 9795
rect 4645 9770 4650 9790
rect 4650 9770 4670 9790
rect 4670 9770 4675 9790
rect 4645 9765 4675 9770
rect 4645 9710 4675 9715
rect 4645 9690 4650 9710
rect 4650 9690 4670 9710
rect 4670 9690 4675 9710
rect 4645 9685 4675 9690
rect 4645 9630 4675 9635
rect 4645 9610 4650 9630
rect 4650 9610 4670 9630
rect 4670 9610 4675 9630
rect 4645 9605 4675 9610
rect 4645 9550 4675 9555
rect 4645 9530 4650 9550
rect 4650 9530 4670 9550
rect 4670 9530 4675 9550
rect 4645 9525 4675 9530
rect 4645 9470 4675 9475
rect 4645 9450 4650 9470
rect 4650 9450 4670 9470
rect 4670 9450 4675 9470
rect 4645 9445 4675 9450
rect 4645 9390 4675 9395
rect 4645 9370 4650 9390
rect 4650 9370 4670 9390
rect 4670 9370 4675 9390
rect 4645 9365 4675 9370
rect 4645 8990 4675 8995
rect 4645 8970 4650 8990
rect 4650 8970 4670 8990
rect 4670 8970 4675 8990
rect 4645 8965 4675 8970
rect 4645 8910 4675 8915
rect 4645 8890 4650 8910
rect 4650 8890 4670 8910
rect 4670 8890 4675 8910
rect 4645 8885 4675 8890
rect 4645 8830 4675 8835
rect 4645 8810 4650 8830
rect 4650 8810 4670 8830
rect 4670 8810 4675 8830
rect 4645 8805 4675 8810
rect 4645 8750 4675 8755
rect 4645 8730 4650 8750
rect 4650 8730 4670 8750
rect 4670 8730 4675 8750
rect 4645 8725 4675 8730
rect 4645 8670 4675 8675
rect 4645 8650 4650 8670
rect 4650 8650 4670 8670
rect 4670 8650 4675 8670
rect 4645 8645 4675 8650
rect 4645 8590 4675 8595
rect 4645 8570 4650 8590
rect 4650 8570 4670 8590
rect 4670 8570 4675 8590
rect 4645 8565 4675 8570
rect 4645 8510 4675 8515
rect 4645 8490 4650 8510
rect 4650 8490 4670 8510
rect 4670 8490 4675 8510
rect 4645 8485 4675 8490
rect 4645 8430 4675 8435
rect 4645 8410 4650 8430
rect 4650 8410 4670 8430
rect 4670 8410 4675 8430
rect 4645 8405 4675 8410
rect 4645 8270 4675 8275
rect 4645 8250 4650 8270
rect 4650 8250 4670 8270
rect 4670 8250 4675 8270
rect 4645 8245 4675 8250
rect 4645 8190 4675 8195
rect 4645 8170 4650 8190
rect 4650 8170 4670 8190
rect 4670 8170 4675 8190
rect 4645 8165 4675 8170
rect 4645 8110 4675 8115
rect 4645 8090 4650 8110
rect 4650 8090 4670 8110
rect 4670 8090 4675 8110
rect 4645 8085 4675 8090
rect 4645 8030 4675 8035
rect 4645 8010 4650 8030
rect 4650 8010 4670 8030
rect 4670 8010 4675 8030
rect 4645 8005 4675 8010
rect 4645 7950 4675 7955
rect 4645 7930 4650 7950
rect 4650 7930 4670 7950
rect 4670 7930 4675 7950
rect 4645 7925 4675 7930
rect 4645 7870 4675 7875
rect 4645 7850 4650 7870
rect 4650 7850 4670 7870
rect 4670 7850 4675 7870
rect 4645 7845 4675 7850
rect 4645 7790 4675 7795
rect 4645 7770 4650 7790
rect 4650 7770 4670 7790
rect 4670 7770 4675 7790
rect 4645 7765 4675 7770
rect 4645 7710 4675 7715
rect 4645 7690 4650 7710
rect 4650 7690 4670 7710
rect 4670 7690 4675 7710
rect 4645 7685 4675 7690
rect 4645 7630 4675 7635
rect 4645 7610 4650 7630
rect 4650 7610 4670 7630
rect 4670 7610 4675 7630
rect 4645 7605 4675 7610
rect 4645 7550 4675 7555
rect 4645 7530 4650 7550
rect 4650 7530 4670 7550
rect 4670 7530 4675 7550
rect 4645 7525 4675 7530
rect 4645 7470 4675 7475
rect 4645 7450 4650 7470
rect 4650 7450 4670 7470
rect 4670 7450 4675 7470
rect 4645 7445 4675 7450
rect 4645 7390 4675 7395
rect 4645 7370 4650 7390
rect 4650 7370 4670 7390
rect 4670 7370 4675 7390
rect 4645 7365 4675 7370
rect 4645 7310 4675 7315
rect 4645 7290 4650 7310
rect 4650 7290 4670 7310
rect 4670 7290 4675 7310
rect 4645 7285 4675 7290
rect 4645 7230 4675 7235
rect 4645 7210 4650 7230
rect 4650 7210 4670 7230
rect 4670 7210 4675 7230
rect 4645 7205 4675 7210
rect 4645 7150 4675 7155
rect 4645 7130 4650 7150
rect 4650 7130 4670 7150
rect 4670 7130 4675 7150
rect 4645 7125 4675 7130
rect 4645 7070 4675 7075
rect 4645 7050 4650 7070
rect 4650 7050 4670 7070
rect 4670 7050 4675 7070
rect 4645 7045 4675 7050
rect 4645 6990 4675 6995
rect 4645 6970 4650 6990
rect 4650 6970 4670 6990
rect 4670 6970 4675 6990
rect 4645 6965 4675 6970
rect 4645 6830 4675 6835
rect 4645 6810 4650 6830
rect 4650 6810 4670 6830
rect 4670 6810 4675 6830
rect 4645 6805 4675 6810
rect 4645 6750 4675 6755
rect 4645 6730 4650 6750
rect 4650 6730 4670 6750
rect 4670 6730 4675 6750
rect 4645 6725 4675 6730
rect 4645 6670 4675 6675
rect 4645 6650 4650 6670
rect 4650 6650 4670 6670
rect 4670 6650 4675 6670
rect 4645 6645 4675 6650
rect 4645 6590 4675 6595
rect 4645 6570 4650 6590
rect 4650 6570 4670 6590
rect 4670 6570 4675 6590
rect 4645 6565 4675 6570
rect 4645 6510 4675 6515
rect 4645 6490 4650 6510
rect 4650 6490 4670 6510
rect 4670 6490 4675 6510
rect 4645 6485 4675 6490
rect 4645 6430 4675 6435
rect 4645 6410 4650 6430
rect 4650 6410 4670 6430
rect 4670 6410 4675 6430
rect 4645 6405 4675 6410
rect 4645 6350 4675 6355
rect 4645 6330 4650 6350
rect 4650 6330 4670 6350
rect 4670 6330 4675 6350
rect 4645 6325 4675 6330
rect 4645 6270 4675 6275
rect 4645 6250 4650 6270
rect 4650 6250 4670 6270
rect 4670 6250 4675 6270
rect 4645 6245 4675 6250
rect 4645 5870 4675 5875
rect 4645 5850 4650 5870
rect 4650 5850 4670 5870
rect 4670 5850 4675 5870
rect 4645 5845 4675 5850
rect 4645 5790 4675 5795
rect 4645 5770 4650 5790
rect 4650 5770 4670 5790
rect 4670 5770 4675 5790
rect 4645 5765 4675 5770
rect 4645 5710 4675 5715
rect 4645 5690 4650 5710
rect 4650 5690 4670 5710
rect 4670 5690 4675 5710
rect 4645 5685 4675 5690
rect 4645 5630 4675 5635
rect 4645 5610 4650 5630
rect 4650 5610 4670 5630
rect 4670 5610 4675 5630
rect 4645 5605 4675 5610
rect 4645 5550 4675 5555
rect 4645 5530 4650 5550
rect 4650 5530 4670 5550
rect 4670 5530 4675 5550
rect 4645 5525 4675 5530
rect 4645 5470 4675 5475
rect 4645 5450 4650 5470
rect 4650 5450 4670 5470
rect 4670 5450 4675 5470
rect 4645 5445 4675 5450
rect 4645 5390 4675 5395
rect 4645 5370 4650 5390
rect 4650 5370 4670 5390
rect 4670 5370 4675 5390
rect 4645 5365 4675 5370
rect 4645 5310 4675 5315
rect 4645 5290 4650 5310
rect 4650 5290 4670 5310
rect 4670 5290 4675 5310
rect 4645 5285 4675 5290
rect 4645 5230 4675 5235
rect 4645 5210 4650 5230
rect 4650 5210 4670 5230
rect 4670 5210 4675 5230
rect 4645 5205 4675 5210
rect 4645 5150 4675 5155
rect 4645 5130 4650 5150
rect 4650 5130 4670 5150
rect 4670 5130 4675 5150
rect 4645 5125 4675 5130
rect 4645 5070 4675 5075
rect 4645 5050 4650 5070
rect 4650 5050 4670 5070
rect 4670 5050 4675 5070
rect 4645 5045 4675 5050
rect 4645 4990 4675 4995
rect 4645 4970 4650 4990
rect 4650 4970 4670 4990
rect 4670 4970 4675 4990
rect 4645 4965 4675 4970
rect 4645 4910 4675 4915
rect 4645 4890 4650 4910
rect 4650 4890 4670 4910
rect 4670 4890 4675 4910
rect 4645 4885 4675 4890
rect 4645 4750 4675 4755
rect 4645 4730 4650 4750
rect 4650 4730 4670 4750
rect 4670 4730 4675 4750
rect 4645 4725 4675 4730
rect 4645 4670 4675 4675
rect 4645 4650 4650 4670
rect 4650 4650 4670 4670
rect 4670 4650 4675 4670
rect 4645 4645 4675 4650
rect 4645 4510 4675 4515
rect 4645 4490 4650 4510
rect 4650 4490 4670 4510
rect 4670 4490 4675 4510
rect 4645 4485 4675 4490
rect 4645 4430 4675 4435
rect 4645 4410 4650 4430
rect 4650 4410 4670 4430
rect 4670 4410 4675 4430
rect 4645 4405 4675 4410
rect 4645 4350 4675 4355
rect 4645 4330 4650 4350
rect 4650 4330 4670 4350
rect 4670 4330 4675 4350
rect 4645 4325 4675 4330
rect 4645 4270 4675 4275
rect 4645 4250 4650 4270
rect 4650 4250 4670 4270
rect 4670 4250 4675 4270
rect 4645 4245 4675 4250
rect 4645 4190 4675 4195
rect 4645 4170 4650 4190
rect 4650 4170 4670 4190
rect 4670 4170 4675 4190
rect 4645 4165 4675 4170
rect 4645 4110 4675 4115
rect 4645 4090 4650 4110
rect 4650 4090 4670 4110
rect 4670 4090 4675 4110
rect 4645 4085 4675 4090
rect 4645 4030 4675 4035
rect 4645 4010 4650 4030
rect 4650 4010 4670 4030
rect 4670 4010 4675 4030
rect 4645 4005 4675 4010
rect 4645 3950 4675 3955
rect 4645 3930 4650 3950
rect 4650 3930 4670 3950
rect 4670 3930 4675 3950
rect 4645 3925 4675 3930
rect 4645 3870 4675 3875
rect 4645 3850 4650 3870
rect 4650 3850 4670 3870
rect 4670 3850 4675 3870
rect 4645 3845 4675 3850
rect 4645 3710 4675 3715
rect 4645 3690 4650 3710
rect 4650 3690 4670 3710
rect 4670 3690 4675 3710
rect 4645 3685 4675 3690
rect 4645 3630 4675 3635
rect 4645 3610 4650 3630
rect 4650 3610 4670 3630
rect 4670 3610 4675 3630
rect 4645 3605 4675 3610
rect 4645 3470 4675 3475
rect 4645 3450 4650 3470
rect 4650 3450 4670 3470
rect 4670 3450 4675 3470
rect 4645 3445 4675 3450
rect 4645 3390 4675 3395
rect 4645 3370 4650 3390
rect 4650 3370 4670 3390
rect 4670 3370 4675 3390
rect 4645 3365 4675 3370
rect 4645 3230 4675 3235
rect 4645 3210 4650 3230
rect 4650 3210 4670 3230
rect 4670 3210 4675 3230
rect 4645 3205 4675 3210
rect 4645 3150 4675 3155
rect 4645 3130 4650 3150
rect 4650 3130 4670 3150
rect 4670 3130 4675 3150
rect 4645 3125 4675 3130
rect 4645 3070 4675 3075
rect 4645 3050 4650 3070
rect 4650 3050 4670 3070
rect 4670 3050 4675 3070
rect 4645 3045 4675 3050
rect 4645 2990 4675 2995
rect 4645 2970 4650 2990
rect 4650 2970 4670 2990
rect 4670 2970 4675 2990
rect 4645 2965 4675 2970
rect 4645 2910 4675 2915
rect 4645 2890 4650 2910
rect 4650 2890 4670 2910
rect 4670 2890 4675 2910
rect 4645 2885 4675 2890
rect 4645 2830 4675 2835
rect 4645 2810 4650 2830
rect 4650 2810 4670 2830
rect 4670 2810 4675 2830
rect 4645 2805 4675 2810
rect 4645 2750 4675 2755
rect 4645 2730 4650 2750
rect 4650 2730 4670 2750
rect 4670 2730 4675 2750
rect 4645 2725 4675 2730
rect 4645 2670 4675 2675
rect 4645 2650 4650 2670
rect 4650 2650 4670 2670
rect 4670 2650 4675 2670
rect 4645 2645 4675 2650
rect 4645 2590 4675 2595
rect 4645 2570 4650 2590
rect 4650 2570 4670 2590
rect 4670 2570 4675 2590
rect 4645 2565 4675 2570
rect 4645 2510 4675 2515
rect 4645 2490 4650 2510
rect 4650 2490 4670 2510
rect 4670 2490 4675 2510
rect 4645 2485 4675 2490
rect 4645 2430 4675 2435
rect 4645 2410 4650 2430
rect 4650 2410 4670 2430
rect 4670 2410 4675 2430
rect 4645 2405 4675 2410
rect 4645 2350 4675 2355
rect 4645 2330 4650 2350
rect 4650 2330 4670 2350
rect 4670 2330 4675 2350
rect 4645 2325 4675 2330
rect 4645 2270 4675 2275
rect 4645 2250 4650 2270
rect 4650 2250 4670 2270
rect 4670 2250 4675 2270
rect 4645 2245 4675 2250
rect 4645 2190 4675 2195
rect 4645 2170 4650 2190
rect 4650 2170 4670 2190
rect 4670 2170 4675 2190
rect 4645 2165 4675 2170
rect 4645 2110 4675 2115
rect 4645 2090 4650 2110
rect 4650 2090 4670 2110
rect 4670 2090 4675 2110
rect 4645 2085 4675 2090
rect 4645 2030 4675 2035
rect 4645 2010 4650 2030
rect 4650 2010 4670 2030
rect 4670 2010 4675 2030
rect 4645 2005 4675 2010
rect 4645 1950 4675 1955
rect 4645 1930 4650 1950
rect 4650 1930 4670 1950
rect 4670 1930 4675 1950
rect 4645 1925 4675 1930
rect 4645 1710 4675 1715
rect 4645 1690 4650 1710
rect 4650 1690 4670 1710
rect 4670 1690 4675 1710
rect 4645 1685 4675 1690
rect 4645 1630 4675 1635
rect 4645 1610 4650 1630
rect 4650 1610 4670 1630
rect 4670 1610 4675 1630
rect 4645 1605 4675 1610
rect 4645 1550 4675 1555
rect 4645 1530 4650 1550
rect 4650 1530 4670 1550
rect 4670 1530 4675 1550
rect 4645 1525 4675 1530
rect 4645 1470 4675 1475
rect 4645 1450 4650 1470
rect 4650 1450 4670 1470
rect 4670 1450 4675 1470
rect 4645 1445 4675 1450
rect 4645 1390 4675 1395
rect 4645 1370 4650 1390
rect 4650 1370 4670 1390
rect 4670 1370 4675 1390
rect 4645 1365 4675 1370
rect 4645 1310 4675 1315
rect 4645 1290 4650 1310
rect 4650 1290 4670 1310
rect 4670 1290 4675 1310
rect 4645 1285 4675 1290
rect 4645 1230 4675 1235
rect 4645 1210 4650 1230
rect 4650 1210 4670 1230
rect 4670 1210 4675 1230
rect 4645 1205 4675 1210
rect 4645 1150 4675 1155
rect 4645 1130 4650 1150
rect 4650 1130 4670 1150
rect 4670 1130 4675 1150
rect 4645 1125 4675 1130
rect 4645 1070 4675 1075
rect 4645 1050 4650 1070
rect 4650 1050 4670 1070
rect 4670 1050 4675 1070
rect 4645 1045 4675 1050
rect 4645 990 4675 995
rect 4645 970 4650 990
rect 4650 970 4670 990
rect 4670 970 4675 990
rect 4645 965 4675 970
rect 4645 830 4675 835
rect 4645 810 4650 830
rect 4650 810 4670 830
rect 4670 810 4675 830
rect 4645 805 4675 810
rect 4645 750 4675 755
rect 4645 730 4650 750
rect 4650 730 4670 750
rect 4670 730 4675 750
rect 4645 725 4675 730
rect 4645 670 4675 675
rect 4645 650 4650 670
rect 4650 650 4670 670
rect 4670 650 4675 670
rect 4645 645 4675 650
rect 4645 590 4675 595
rect 4645 570 4650 590
rect 4650 570 4670 590
rect 4670 570 4675 590
rect 4645 565 4675 570
rect 4645 510 4675 515
rect 4645 490 4650 510
rect 4650 490 4670 510
rect 4670 490 4675 510
rect 4645 485 4675 490
rect 4645 270 4675 275
rect 4645 250 4650 270
rect 4650 250 4670 270
rect 4670 250 4675 270
rect 4645 245 4675 250
rect 4645 190 4675 195
rect 4645 170 4650 190
rect 4650 170 4670 190
rect 4670 170 4675 190
rect 4645 165 4675 170
rect 4645 110 4675 115
rect 4645 90 4650 110
rect 4650 90 4670 110
rect 4670 90 4675 110
rect 4645 85 4675 90
rect 4645 30 4675 35
rect 4645 10 4650 30
rect 4650 10 4670 30
rect 4670 10 4675 30
rect 4645 5 4675 10
rect 4725 15710 4755 15715
rect 4725 15690 4730 15710
rect 4730 15690 4750 15710
rect 4750 15690 4755 15710
rect 4725 15685 4755 15690
rect 4725 15630 4755 15635
rect 4725 15610 4730 15630
rect 4730 15610 4750 15630
rect 4750 15610 4755 15630
rect 4725 15605 4755 15610
rect 4725 15550 4755 15555
rect 4725 15530 4730 15550
rect 4730 15530 4750 15550
rect 4750 15530 4755 15550
rect 4725 15525 4755 15530
rect 4725 15470 4755 15475
rect 4725 15450 4730 15470
rect 4730 15450 4750 15470
rect 4750 15450 4755 15470
rect 4725 15445 4755 15450
rect 4725 15390 4755 15395
rect 4725 15370 4730 15390
rect 4730 15370 4750 15390
rect 4750 15370 4755 15390
rect 4725 15365 4755 15370
rect 4725 15310 4755 15315
rect 4725 15290 4730 15310
rect 4730 15290 4750 15310
rect 4750 15290 4755 15310
rect 4725 15285 4755 15290
rect 4725 15230 4755 15235
rect 4725 15210 4730 15230
rect 4730 15210 4750 15230
rect 4750 15210 4755 15230
rect 4725 15205 4755 15210
rect 4725 15150 4755 15155
rect 4725 15130 4730 15150
rect 4730 15130 4750 15150
rect 4750 15130 4755 15150
rect 4725 15125 4755 15130
rect 4725 14990 4755 14995
rect 4725 14970 4730 14990
rect 4730 14970 4750 14990
rect 4750 14970 4755 14990
rect 4725 14965 4755 14970
rect 4725 14910 4755 14915
rect 4725 14890 4730 14910
rect 4730 14890 4750 14910
rect 4750 14890 4755 14910
rect 4725 14885 4755 14890
rect 4725 14830 4755 14835
rect 4725 14810 4730 14830
rect 4730 14810 4750 14830
rect 4750 14810 4755 14830
rect 4725 14805 4755 14810
rect 4725 14750 4755 14755
rect 4725 14730 4730 14750
rect 4730 14730 4750 14750
rect 4750 14730 4755 14750
rect 4725 14725 4755 14730
rect 4725 14670 4755 14675
rect 4725 14650 4730 14670
rect 4730 14650 4750 14670
rect 4750 14650 4755 14670
rect 4725 14645 4755 14650
rect 4725 14590 4755 14595
rect 4725 14570 4730 14590
rect 4730 14570 4750 14590
rect 4750 14570 4755 14590
rect 4725 14565 4755 14570
rect 4725 14510 4755 14515
rect 4725 14490 4730 14510
rect 4730 14490 4750 14510
rect 4750 14490 4755 14510
rect 4725 14485 4755 14490
rect 4725 14430 4755 14435
rect 4725 14410 4730 14430
rect 4730 14410 4750 14430
rect 4750 14410 4755 14430
rect 4725 14405 4755 14410
rect 4725 14030 4755 14035
rect 4725 14010 4730 14030
rect 4730 14010 4750 14030
rect 4750 14010 4755 14030
rect 4725 14005 4755 14010
rect 4725 13950 4755 13955
rect 4725 13930 4730 13950
rect 4730 13930 4750 13950
rect 4750 13930 4755 13950
rect 4725 13925 4755 13930
rect 4725 13870 4755 13875
rect 4725 13850 4730 13870
rect 4730 13850 4750 13870
rect 4750 13850 4755 13870
rect 4725 13845 4755 13850
rect 4725 13790 4755 13795
rect 4725 13770 4730 13790
rect 4730 13770 4750 13790
rect 4750 13770 4755 13790
rect 4725 13765 4755 13770
rect 4725 13710 4755 13715
rect 4725 13690 4730 13710
rect 4730 13690 4750 13710
rect 4750 13690 4755 13710
rect 4725 13685 4755 13690
rect 4725 13630 4755 13635
rect 4725 13610 4730 13630
rect 4730 13610 4750 13630
rect 4750 13610 4755 13630
rect 4725 13605 4755 13610
rect 4725 13550 4755 13555
rect 4725 13530 4730 13550
rect 4730 13530 4750 13550
rect 4750 13530 4755 13550
rect 4725 13525 4755 13530
rect 4725 13470 4755 13475
rect 4725 13450 4730 13470
rect 4730 13450 4750 13470
rect 4750 13450 4755 13470
rect 4725 13445 4755 13450
rect 4725 13070 4755 13075
rect 4725 13050 4730 13070
rect 4730 13050 4750 13070
rect 4750 13050 4755 13070
rect 4725 13045 4755 13050
rect 4725 12990 4755 12995
rect 4725 12970 4730 12990
rect 4730 12970 4750 12990
rect 4750 12970 4755 12990
rect 4725 12965 4755 12970
rect 4725 12910 4755 12915
rect 4725 12890 4730 12910
rect 4730 12890 4750 12910
rect 4750 12890 4755 12910
rect 4725 12885 4755 12890
rect 4725 12830 4755 12835
rect 4725 12810 4730 12830
rect 4730 12810 4750 12830
rect 4750 12810 4755 12830
rect 4725 12805 4755 12810
rect 4725 12750 4755 12755
rect 4725 12730 4730 12750
rect 4730 12730 4750 12750
rect 4750 12730 4755 12750
rect 4725 12725 4755 12730
rect 4725 12670 4755 12675
rect 4725 12650 4730 12670
rect 4730 12650 4750 12670
rect 4750 12650 4755 12670
rect 4725 12645 4755 12650
rect 4725 12590 4755 12595
rect 4725 12570 4730 12590
rect 4730 12570 4750 12590
rect 4750 12570 4755 12590
rect 4725 12565 4755 12570
rect 4725 12510 4755 12515
rect 4725 12490 4730 12510
rect 4730 12490 4750 12510
rect 4750 12490 4755 12510
rect 4725 12485 4755 12490
rect 4725 12350 4755 12355
rect 4725 12330 4730 12350
rect 4730 12330 4750 12350
rect 4750 12330 4755 12350
rect 4725 12325 4755 12330
rect 4725 12270 4755 12275
rect 4725 12250 4730 12270
rect 4730 12250 4750 12270
rect 4750 12250 4755 12270
rect 4725 12245 4755 12250
rect 4725 12190 4755 12195
rect 4725 12170 4730 12190
rect 4730 12170 4750 12190
rect 4750 12170 4755 12190
rect 4725 12165 4755 12170
rect 4725 12110 4755 12115
rect 4725 12090 4730 12110
rect 4730 12090 4750 12110
rect 4750 12090 4755 12110
rect 4725 12085 4755 12090
rect 4725 12030 4755 12035
rect 4725 12010 4730 12030
rect 4730 12010 4750 12030
rect 4750 12010 4755 12030
rect 4725 12005 4755 12010
rect 4725 11950 4755 11955
rect 4725 11930 4730 11950
rect 4730 11930 4750 11950
rect 4750 11930 4755 11950
rect 4725 11925 4755 11930
rect 4725 11870 4755 11875
rect 4725 11850 4730 11870
rect 4730 11850 4750 11870
rect 4750 11850 4755 11870
rect 4725 11845 4755 11850
rect 4725 11790 4755 11795
rect 4725 11770 4730 11790
rect 4730 11770 4750 11790
rect 4750 11770 4755 11790
rect 4725 11765 4755 11770
rect 4725 11710 4755 11715
rect 4725 11690 4730 11710
rect 4730 11690 4750 11710
rect 4750 11690 4755 11710
rect 4725 11685 4755 11690
rect 4725 11630 4755 11635
rect 4725 11610 4730 11630
rect 4730 11610 4750 11630
rect 4750 11610 4755 11630
rect 4725 11605 4755 11610
rect 4725 11550 4755 11555
rect 4725 11530 4730 11550
rect 4730 11530 4750 11550
rect 4750 11530 4755 11550
rect 4725 11525 4755 11530
rect 4725 11470 4755 11475
rect 4725 11450 4730 11470
rect 4730 11450 4750 11470
rect 4750 11450 4755 11470
rect 4725 11445 4755 11450
rect 4725 11390 4755 11395
rect 4725 11370 4730 11390
rect 4730 11370 4750 11390
rect 4750 11370 4755 11390
rect 4725 11365 4755 11370
rect 4725 11310 4755 11315
rect 4725 11290 4730 11310
rect 4730 11290 4750 11310
rect 4750 11290 4755 11310
rect 4725 11285 4755 11290
rect 4725 11230 4755 11235
rect 4725 11210 4730 11230
rect 4730 11210 4750 11230
rect 4750 11210 4755 11230
rect 4725 11205 4755 11210
rect 4725 11150 4755 11155
rect 4725 11130 4730 11150
rect 4730 11130 4750 11150
rect 4750 11130 4755 11150
rect 4725 11125 4755 11130
rect 4725 11070 4755 11075
rect 4725 11050 4730 11070
rect 4730 11050 4750 11070
rect 4750 11050 4755 11070
rect 4725 11045 4755 11050
rect 4725 10910 4755 10915
rect 4725 10890 4730 10910
rect 4730 10890 4750 10910
rect 4750 10890 4755 10910
rect 4725 10885 4755 10890
rect 4725 10830 4755 10835
rect 4725 10810 4730 10830
rect 4730 10810 4750 10830
rect 4750 10810 4755 10830
rect 4725 10805 4755 10810
rect 4725 10750 4755 10755
rect 4725 10730 4730 10750
rect 4730 10730 4750 10750
rect 4750 10730 4755 10750
rect 4725 10725 4755 10730
rect 4725 10670 4755 10675
rect 4725 10650 4730 10670
rect 4730 10650 4750 10670
rect 4750 10650 4755 10670
rect 4725 10645 4755 10650
rect 4725 10590 4755 10595
rect 4725 10570 4730 10590
rect 4730 10570 4750 10590
rect 4750 10570 4755 10590
rect 4725 10565 4755 10570
rect 4725 10510 4755 10515
rect 4725 10490 4730 10510
rect 4730 10490 4750 10510
rect 4750 10490 4755 10510
rect 4725 10485 4755 10490
rect 4725 10430 4755 10435
rect 4725 10410 4730 10430
rect 4730 10410 4750 10430
rect 4750 10410 4755 10430
rect 4725 10405 4755 10410
rect 4725 10350 4755 10355
rect 4725 10330 4730 10350
rect 4730 10330 4750 10350
rect 4750 10330 4755 10350
rect 4725 10325 4755 10330
rect 4725 9950 4755 9955
rect 4725 9930 4730 9950
rect 4730 9930 4750 9950
rect 4750 9930 4755 9950
rect 4725 9925 4755 9930
rect 4725 9870 4755 9875
rect 4725 9850 4730 9870
rect 4730 9850 4750 9870
rect 4750 9850 4755 9870
rect 4725 9845 4755 9850
rect 4725 9790 4755 9795
rect 4725 9770 4730 9790
rect 4730 9770 4750 9790
rect 4750 9770 4755 9790
rect 4725 9765 4755 9770
rect 4725 9710 4755 9715
rect 4725 9690 4730 9710
rect 4730 9690 4750 9710
rect 4750 9690 4755 9710
rect 4725 9685 4755 9690
rect 4725 9630 4755 9635
rect 4725 9610 4730 9630
rect 4730 9610 4750 9630
rect 4750 9610 4755 9630
rect 4725 9605 4755 9610
rect 4725 9550 4755 9555
rect 4725 9530 4730 9550
rect 4730 9530 4750 9550
rect 4750 9530 4755 9550
rect 4725 9525 4755 9530
rect 4725 9470 4755 9475
rect 4725 9450 4730 9470
rect 4730 9450 4750 9470
rect 4750 9450 4755 9470
rect 4725 9445 4755 9450
rect 4725 9390 4755 9395
rect 4725 9370 4730 9390
rect 4730 9370 4750 9390
rect 4750 9370 4755 9390
rect 4725 9365 4755 9370
rect 4725 8990 4755 8995
rect 4725 8970 4730 8990
rect 4730 8970 4750 8990
rect 4750 8970 4755 8990
rect 4725 8965 4755 8970
rect 4725 8910 4755 8915
rect 4725 8890 4730 8910
rect 4730 8890 4750 8910
rect 4750 8890 4755 8910
rect 4725 8885 4755 8890
rect 4725 8830 4755 8835
rect 4725 8810 4730 8830
rect 4730 8810 4750 8830
rect 4750 8810 4755 8830
rect 4725 8805 4755 8810
rect 4725 8750 4755 8755
rect 4725 8730 4730 8750
rect 4730 8730 4750 8750
rect 4750 8730 4755 8750
rect 4725 8725 4755 8730
rect 4725 8670 4755 8675
rect 4725 8650 4730 8670
rect 4730 8650 4750 8670
rect 4750 8650 4755 8670
rect 4725 8645 4755 8650
rect 4725 8590 4755 8595
rect 4725 8570 4730 8590
rect 4730 8570 4750 8590
rect 4750 8570 4755 8590
rect 4725 8565 4755 8570
rect 4725 8510 4755 8515
rect 4725 8490 4730 8510
rect 4730 8490 4750 8510
rect 4750 8490 4755 8510
rect 4725 8485 4755 8490
rect 4725 8430 4755 8435
rect 4725 8410 4730 8430
rect 4730 8410 4750 8430
rect 4750 8410 4755 8430
rect 4725 8405 4755 8410
rect 4725 8270 4755 8275
rect 4725 8250 4730 8270
rect 4730 8250 4750 8270
rect 4750 8250 4755 8270
rect 4725 8245 4755 8250
rect 4725 8190 4755 8195
rect 4725 8170 4730 8190
rect 4730 8170 4750 8190
rect 4750 8170 4755 8190
rect 4725 8165 4755 8170
rect 4725 8110 4755 8115
rect 4725 8090 4730 8110
rect 4730 8090 4750 8110
rect 4750 8090 4755 8110
rect 4725 8085 4755 8090
rect 4725 8030 4755 8035
rect 4725 8010 4730 8030
rect 4730 8010 4750 8030
rect 4750 8010 4755 8030
rect 4725 8005 4755 8010
rect 4725 7950 4755 7955
rect 4725 7930 4730 7950
rect 4730 7930 4750 7950
rect 4750 7930 4755 7950
rect 4725 7925 4755 7930
rect 4725 7870 4755 7875
rect 4725 7850 4730 7870
rect 4730 7850 4750 7870
rect 4750 7850 4755 7870
rect 4725 7845 4755 7850
rect 4725 7790 4755 7795
rect 4725 7770 4730 7790
rect 4730 7770 4750 7790
rect 4750 7770 4755 7790
rect 4725 7765 4755 7770
rect 4725 7710 4755 7715
rect 4725 7690 4730 7710
rect 4730 7690 4750 7710
rect 4750 7690 4755 7710
rect 4725 7685 4755 7690
rect 4725 7630 4755 7635
rect 4725 7610 4730 7630
rect 4730 7610 4750 7630
rect 4750 7610 4755 7630
rect 4725 7605 4755 7610
rect 4725 7550 4755 7555
rect 4725 7530 4730 7550
rect 4730 7530 4750 7550
rect 4750 7530 4755 7550
rect 4725 7525 4755 7530
rect 4725 7470 4755 7475
rect 4725 7450 4730 7470
rect 4730 7450 4750 7470
rect 4750 7450 4755 7470
rect 4725 7445 4755 7450
rect 4725 7390 4755 7395
rect 4725 7370 4730 7390
rect 4730 7370 4750 7390
rect 4750 7370 4755 7390
rect 4725 7365 4755 7370
rect 4725 7310 4755 7315
rect 4725 7290 4730 7310
rect 4730 7290 4750 7310
rect 4750 7290 4755 7310
rect 4725 7285 4755 7290
rect 4725 7230 4755 7235
rect 4725 7210 4730 7230
rect 4730 7210 4750 7230
rect 4750 7210 4755 7230
rect 4725 7205 4755 7210
rect 4725 7150 4755 7155
rect 4725 7130 4730 7150
rect 4730 7130 4750 7150
rect 4750 7130 4755 7150
rect 4725 7125 4755 7130
rect 4725 7070 4755 7075
rect 4725 7050 4730 7070
rect 4730 7050 4750 7070
rect 4750 7050 4755 7070
rect 4725 7045 4755 7050
rect 4725 6990 4755 6995
rect 4725 6970 4730 6990
rect 4730 6970 4750 6990
rect 4750 6970 4755 6990
rect 4725 6965 4755 6970
rect 4725 6830 4755 6835
rect 4725 6810 4730 6830
rect 4730 6810 4750 6830
rect 4750 6810 4755 6830
rect 4725 6805 4755 6810
rect 4725 6750 4755 6755
rect 4725 6730 4730 6750
rect 4730 6730 4750 6750
rect 4750 6730 4755 6750
rect 4725 6725 4755 6730
rect 4725 6670 4755 6675
rect 4725 6650 4730 6670
rect 4730 6650 4750 6670
rect 4750 6650 4755 6670
rect 4725 6645 4755 6650
rect 4725 6590 4755 6595
rect 4725 6570 4730 6590
rect 4730 6570 4750 6590
rect 4750 6570 4755 6590
rect 4725 6565 4755 6570
rect 4725 6510 4755 6515
rect 4725 6490 4730 6510
rect 4730 6490 4750 6510
rect 4750 6490 4755 6510
rect 4725 6485 4755 6490
rect 4725 6430 4755 6435
rect 4725 6410 4730 6430
rect 4730 6410 4750 6430
rect 4750 6410 4755 6430
rect 4725 6405 4755 6410
rect 4725 6350 4755 6355
rect 4725 6330 4730 6350
rect 4730 6330 4750 6350
rect 4750 6330 4755 6350
rect 4725 6325 4755 6330
rect 4725 6270 4755 6275
rect 4725 6250 4730 6270
rect 4730 6250 4750 6270
rect 4750 6250 4755 6270
rect 4725 6245 4755 6250
rect 4725 5870 4755 5875
rect 4725 5850 4730 5870
rect 4730 5850 4750 5870
rect 4750 5850 4755 5870
rect 4725 5845 4755 5850
rect 4725 5790 4755 5795
rect 4725 5770 4730 5790
rect 4730 5770 4750 5790
rect 4750 5770 4755 5790
rect 4725 5765 4755 5770
rect 4725 5710 4755 5715
rect 4725 5690 4730 5710
rect 4730 5690 4750 5710
rect 4750 5690 4755 5710
rect 4725 5685 4755 5690
rect 4725 5630 4755 5635
rect 4725 5610 4730 5630
rect 4730 5610 4750 5630
rect 4750 5610 4755 5630
rect 4725 5605 4755 5610
rect 4725 5550 4755 5555
rect 4725 5530 4730 5550
rect 4730 5530 4750 5550
rect 4750 5530 4755 5550
rect 4725 5525 4755 5530
rect 4725 5470 4755 5475
rect 4725 5450 4730 5470
rect 4730 5450 4750 5470
rect 4750 5450 4755 5470
rect 4725 5445 4755 5450
rect 4725 5390 4755 5395
rect 4725 5370 4730 5390
rect 4730 5370 4750 5390
rect 4750 5370 4755 5390
rect 4725 5365 4755 5370
rect 4725 5310 4755 5315
rect 4725 5290 4730 5310
rect 4730 5290 4750 5310
rect 4750 5290 4755 5310
rect 4725 5285 4755 5290
rect 4725 5230 4755 5235
rect 4725 5210 4730 5230
rect 4730 5210 4750 5230
rect 4750 5210 4755 5230
rect 4725 5205 4755 5210
rect 4725 5150 4755 5155
rect 4725 5130 4730 5150
rect 4730 5130 4750 5150
rect 4750 5130 4755 5150
rect 4725 5125 4755 5130
rect 4725 5070 4755 5075
rect 4725 5050 4730 5070
rect 4730 5050 4750 5070
rect 4750 5050 4755 5070
rect 4725 5045 4755 5050
rect 4725 4990 4755 4995
rect 4725 4970 4730 4990
rect 4730 4970 4750 4990
rect 4750 4970 4755 4990
rect 4725 4965 4755 4970
rect 4725 4910 4755 4915
rect 4725 4890 4730 4910
rect 4730 4890 4750 4910
rect 4750 4890 4755 4910
rect 4725 4885 4755 4890
rect 4725 4750 4755 4755
rect 4725 4730 4730 4750
rect 4730 4730 4750 4750
rect 4750 4730 4755 4750
rect 4725 4725 4755 4730
rect 4725 4670 4755 4675
rect 4725 4650 4730 4670
rect 4730 4650 4750 4670
rect 4750 4650 4755 4670
rect 4725 4645 4755 4650
rect 4725 4510 4755 4515
rect 4725 4490 4730 4510
rect 4730 4490 4750 4510
rect 4750 4490 4755 4510
rect 4725 4485 4755 4490
rect 4725 4430 4755 4435
rect 4725 4410 4730 4430
rect 4730 4410 4750 4430
rect 4750 4410 4755 4430
rect 4725 4405 4755 4410
rect 4725 4350 4755 4355
rect 4725 4330 4730 4350
rect 4730 4330 4750 4350
rect 4750 4330 4755 4350
rect 4725 4325 4755 4330
rect 4725 4270 4755 4275
rect 4725 4250 4730 4270
rect 4730 4250 4750 4270
rect 4750 4250 4755 4270
rect 4725 4245 4755 4250
rect 4725 4190 4755 4195
rect 4725 4170 4730 4190
rect 4730 4170 4750 4190
rect 4750 4170 4755 4190
rect 4725 4165 4755 4170
rect 4725 4110 4755 4115
rect 4725 4090 4730 4110
rect 4730 4090 4750 4110
rect 4750 4090 4755 4110
rect 4725 4085 4755 4090
rect 4725 4030 4755 4035
rect 4725 4010 4730 4030
rect 4730 4010 4750 4030
rect 4750 4010 4755 4030
rect 4725 4005 4755 4010
rect 4725 3950 4755 3955
rect 4725 3930 4730 3950
rect 4730 3930 4750 3950
rect 4750 3930 4755 3950
rect 4725 3925 4755 3930
rect 4725 3870 4755 3875
rect 4725 3850 4730 3870
rect 4730 3850 4750 3870
rect 4750 3850 4755 3870
rect 4725 3845 4755 3850
rect 4725 3710 4755 3715
rect 4725 3690 4730 3710
rect 4730 3690 4750 3710
rect 4750 3690 4755 3710
rect 4725 3685 4755 3690
rect 4725 3630 4755 3635
rect 4725 3610 4730 3630
rect 4730 3610 4750 3630
rect 4750 3610 4755 3630
rect 4725 3605 4755 3610
rect 4725 3470 4755 3475
rect 4725 3450 4730 3470
rect 4730 3450 4750 3470
rect 4750 3450 4755 3470
rect 4725 3445 4755 3450
rect 4725 3390 4755 3395
rect 4725 3370 4730 3390
rect 4730 3370 4750 3390
rect 4750 3370 4755 3390
rect 4725 3365 4755 3370
rect 4725 3230 4755 3235
rect 4725 3210 4730 3230
rect 4730 3210 4750 3230
rect 4750 3210 4755 3230
rect 4725 3205 4755 3210
rect 4725 3150 4755 3155
rect 4725 3130 4730 3150
rect 4730 3130 4750 3150
rect 4750 3130 4755 3150
rect 4725 3125 4755 3130
rect 4725 3070 4755 3075
rect 4725 3050 4730 3070
rect 4730 3050 4750 3070
rect 4750 3050 4755 3070
rect 4725 3045 4755 3050
rect 4725 2990 4755 2995
rect 4725 2970 4730 2990
rect 4730 2970 4750 2990
rect 4750 2970 4755 2990
rect 4725 2965 4755 2970
rect 4725 2910 4755 2915
rect 4725 2890 4730 2910
rect 4730 2890 4750 2910
rect 4750 2890 4755 2910
rect 4725 2885 4755 2890
rect 4725 2830 4755 2835
rect 4725 2810 4730 2830
rect 4730 2810 4750 2830
rect 4750 2810 4755 2830
rect 4725 2805 4755 2810
rect 4725 2750 4755 2755
rect 4725 2730 4730 2750
rect 4730 2730 4750 2750
rect 4750 2730 4755 2750
rect 4725 2725 4755 2730
rect 4725 2670 4755 2675
rect 4725 2650 4730 2670
rect 4730 2650 4750 2670
rect 4750 2650 4755 2670
rect 4725 2645 4755 2650
rect 4725 2590 4755 2595
rect 4725 2570 4730 2590
rect 4730 2570 4750 2590
rect 4750 2570 4755 2590
rect 4725 2565 4755 2570
rect 4725 2510 4755 2515
rect 4725 2490 4730 2510
rect 4730 2490 4750 2510
rect 4750 2490 4755 2510
rect 4725 2485 4755 2490
rect 4725 2430 4755 2435
rect 4725 2410 4730 2430
rect 4730 2410 4750 2430
rect 4750 2410 4755 2430
rect 4725 2405 4755 2410
rect 4725 2350 4755 2355
rect 4725 2330 4730 2350
rect 4730 2330 4750 2350
rect 4750 2330 4755 2350
rect 4725 2325 4755 2330
rect 4725 2270 4755 2275
rect 4725 2250 4730 2270
rect 4730 2250 4750 2270
rect 4750 2250 4755 2270
rect 4725 2245 4755 2250
rect 4725 2190 4755 2195
rect 4725 2170 4730 2190
rect 4730 2170 4750 2190
rect 4750 2170 4755 2190
rect 4725 2165 4755 2170
rect 4725 2110 4755 2115
rect 4725 2090 4730 2110
rect 4730 2090 4750 2110
rect 4750 2090 4755 2110
rect 4725 2085 4755 2090
rect 4725 2030 4755 2035
rect 4725 2010 4730 2030
rect 4730 2010 4750 2030
rect 4750 2010 4755 2030
rect 4725 2005 4755 2010
rect 4725 1950 4755 1955
rect 4725 1930 4730 1950
rect 4730 1930 4750 1950
rect 4750 1930 4755 1950
rect 4725 1925 4755 1930
rect 4725 1710 4755 1715
rect 4725 1690 4730 1710
rect 4730 1690 4750 1710
rect 4750 1690 4755 1710
rect 4725 1685 4755 1690
rect 4725 1630 4755 1635
rect 4725 1610 4730 1630
rect 4730 1610 4750 1630
rect 4750 1610 4755 1630
rect 4725 1605 4755 1610
rect 4725 1550 4755 1555
rect 4725 1530 4730 1550
rect 4730 1530 4750 1550
rect 4750 1530 4755 1550
rect 4725 1525 4755 1530
rect 4725 1470 4755 1475
rect 4725 1450 4730 1470
rect 4730 1450 4750 1470
rect 4750 1450 4755 1470
rect 4725 1445 4755 1450
rect 4725 1390 4755 1395
rect 4725 1370 4730 1390
rect 4730 1370 4750 1390
rect 4750 1370 4755 1390
rect 4725 1365 4755 1370
rect 4725 1310 4755 1315
rect 4725 1290 4730 1310
rect 4730 1290 4750 1310
rect 4750 1290 4755 1310
rect 4725 1285 4755 1290
rect 4725 1230 4755 1235
rect 4725 1210 4730 1230
rect 4730 1210 4750 1230
rect 4750 1210 4755 1230
rect 4725 1205 4755 1210
rect 4725 1150 4755 1155
rect 4725 1130 4730 1150
rect 4730 1130 4750 1150
rect 4750 1130 4755 1150
rect 4725 1125 4755 1130
rect 4725 1070 4755 1075
rect 4725 1050 4730 1070
rect 4730 1050 4750 1070
rect 4750 1050 4755 1070
rect 4725 1045 4755 1050
rect 4725 990 4755 995
rect 4725 970 4730 990
rect 4730 970 4750 990
rect 4750 970 4755 990
rect 4725 965 4755 970
rect 4725 830 4755 835
rect 4725 810 4730 830
rect 4730 810 4750 830
rect 4750 810 4755 830
rect 4725 805 4755 810
rect 4725 750 4755 755
rect 4725 730 4730 750
rect 4730 730 4750 750
rect 4750 730 4755 750
rect 4725 725 4755 730
rect 4725 670 4755 675
rect 4725 650 4730 670
rect 4730 650 4750 670
rect 4750 650 4755 670
rect 4725 645 4755 650
rect 4725 590 4755 595
rect 4725 570 4730 590
rect 4730 570 4750 590
rect 4750 570 4755 590
rect 4725 565 4755 570
rect 4725 510 4755 515
rect 4725 490 4730 510
rect 4730 490 4750 510
rect 4750 490 4755 510
rect 4725 485 4755 490
rect 4725 270 4755 275
rect 4725 250 4730 270
rect 4730 250 4750 270
rect 4750 250 4755 270
rect 4725 245 4755 250
rect 4725 190 4755 195
rect 4725 170 4730 190
rect 4730 170 4750 190
rect 4750 170 4755 190
rect 4725 165 4755 170
rect 4725 110 4755 115
rect 4725 90 4730 110
rect 4730 90 4750 110
rect 4750 90 4755 110
rect 4725 85 4755 90
rect 4725 30 4755 35
rect 4725 10 4730 30
rect 4730 10 4750 30
rect 4750 10 4755 30
rect 4725 5 4755 10
rect 4885 15710 4915 15715
rect 4885 15690 4890 15710
rect 4890 15690 4910 15710
rect 4910 15690 4915 15710
rect 4885 15685 4915 15690
rect 4885 15630 4915 15635
rect 4885 15610 4890 15630
rect 4890 15610 4910 15630
rect 4910 15610 4915 15630
rect 4885 15605 4915 15610
rect 4885 15550 4915 15555
rect 4885 15530 4890 15550
rect 4890 15530 4910 15550
rect 4910 15530 4915 15550
rect 4885 15525 4915 15530
rect 4885 15470 4915 15475
rect 4885 15450 4890 15470
rect 4890 15450 4910 15470
rect 4910 15450 4915 15470
rect 4885 15445 4915 15450
rect 4885 15390 4915 15395
rect 4885 15370 4890 15390
rect 4890 15370 4910 15390
rect 4910 15370 4915 15390
rect 4885 15365 4915 15370
rect 4885 15310 4915 15315
rect 4885 15290 4890 15310
rect 4890 15290 4910 15310
rect 4910 15290 4915 15310
rect 4885 15285 4915 15290
rect 4885 15230 4915 15235
rect 4885 15210 4890 15230
rect 4890 15210 4910 15230
rect 4910 15210 4915 15230
rect 4885 15205 4915 15210
rect 4885 15150 4915 15155
rect 4885 15130 4890 15150
rect 4890 15130 4910 15150
rect 4910 15130 4915 15150
rect 4885 15125 4915 15130
rect 4885 14990 4915 14995
rect 4885 14970 4890 14990
rect 4890 14970 4910 14990
rect 4910 14970 4915 14990
rect 4885 14965 4915 14970
rect 4885 14910 4915 14915
rect 4885 14890 4890 14910
rect 4890 14890 4910 14910
rect 4910 14890 4915 14910
rect 4885 14885 4915 14890
rect 4885 14830 4915 14835
rect 4885 14810 4890 14830
rect 4890 14810 4910 14830
rect 4910 14810 4915 14830
rect 4885 14805 4915 14810
rect 4885 14750 4915 14755
rect 4885 14730 4890 14750
rect 4890 14730 4910 14750
rect 4910 14730 4915 14750
rect 4885 14725 4915 14730
rect 4885 14670 4915 14675
rect 4885 14650 4890 14670
rect 4890 14650 4910 14670
rect 4910 14650 4915 14670
rect 4885 14645 4915 14650
rect 4885 14590 4915 14595
rect 4885 14570 4890 14590
rect 4890 14570 4910 14590
rect 4910 14570 4915 14590
rect 4885 14565 4915 14570
rect 4885 14510 4915 14515
rect 4885 14490 4890 14510
rect 4890 14490 4910 14510
rect 4910 14490 4915 14510
rect 4885 14485 4915 14490
rect 4885 14430 4915 14435
rect 4885 14410 4890 14430
rect 4890 14410 4910 14430
rect 4910 14410 4915 14430
rect 4885 14405 4915 14410
rect 4885 14030 4915 14035
rect 4885 14010 4890 14030
rect 4890 14010 4910 14030
rect 4910 14010 4915 14030
rect 4885 14005 4915 14010
rect 4885 13950 4915 13955
rect 4885 13930 4890 13950
rect 4890 13930 4910 13950
rect 4910 13930 4915 13950
rect 4885 13925 4915 13930
rect 4885 13870 4915 13875
rect 4885 13850 4890 13870
rect 4890 13850 4910 13870
rect 4910 13850 4915 13870
rect 4885 13845 4915 13850
rect 4885 13790 4915 13795
rect 4885 13770 4890 13790
rect 4890 13770 4910 13790
rect 4910 13770 4915 13790
rect 4885 13765 4915 13770
rect 4885 13710 4915 13715
rect 4885 13690 4890 13710
rect 4890 13690 4910 13710
rect 4910 13690 4915 13710
rect 4885 13685 4915 13690
rect 4885 13630 4915 13635
rect 4885 13610 4890 13630
rect 4890 13610 4910 13630
rect 4910 13610 4915 13630
rect 4885 13605 4915 13610
rect 4885 13550 4915 13555
rect 4885 13530 4890 13550
rect 4890 13530 4910 13550
rect 4910 13530 4915 13550
rect 4885 13525 4915 13530
rect 4885 13470 4915 13475
rect 4885 13450 4890 13470
rect 4890 13450 4910 13470
rect 4910 13450 4915 13470
rect 4885 13445 4915 13450
rect 4885 13070 4915 13075
rect 4885 13050 4890 13070
rect 4890 13050 4910 13070
rect 4910 13050 4915 13070
rect 4885 13045 4915 13050
rect 4885 12990 4915 12995
rect 4885 12970 4890 12990
rect 4890 12970 4910 12990
rect 4910 12970 4915 12990
rect 4885 12965 4915 12970
rect 4885 12910 4915 12915
rect 4885 12890 4890 12910
rect 4890 12890 4910 12910
rect 4910 12890 4915 12910
rect 4885 12885 4915 12890
rect 4885 12830 4915 12835
rect 4885 12810 4890 12830
rect 4890 12810 4910 12830
rect 4910 12810 4915 12830
rect 4885 12805 4915 12810
rect 4885 12750 4915 12755
rect 4885 12730 4890 12750
rect 4890 12730 4910 12750
rect 4910 12730 4915 12750
rect 4885 12725 4915 12730
rect 4885 12670 4915 12675
rect 4885 12650 4890 12670
rect 4890 12650 4910 12670
rect 4910 12650 4915 12670
rect 4885 12645 4915 12650
rect 4885 12590 4915 12595
rect 4885 12570 4890 12590
rect 4890 12570 4910 12590
rect 4910 12570 4915 12590
rect 4885 12565 4915 12570
rect 4885 12510 4915 12515
rect 4885 12490 4890 12510
rect 4890 12490 4910 12510
rect 4910 12490 4915 12510
rect 4885 12485 4915 12490
rect 4885 12350 4915 12355
rect 4885 12330 4890 12350
rect 4890 12330 4910 12350
rect 4910 12330 4915 12350
rect 4885 12325 4915 12330
rect 4885 12270 4915 12275
rect 4885 12250 4890 12270
rect 4890 12250 4910 12270
rect 4910 12250 4915 12270
rect 4885 12245 4915 12250
rect 4885 12190 4915 12195
rect 4885 12170 4890 12190
rect 4890 12170 4910 12190
rect 4910 12170 4915 12190
rect 4885 12165 4915 12170
rect 4885 12110 4915 12115
rect 4885 12090 4890 12110
rect 4890 12090 4910 12110
rect 4910 12090 4915 12110
rect 4885 12085 4915 12090
rect 4885 12030 4915 12035
rect 4885 12010 4890 12030
rect 4890 12010 4910 12030
rect 4910 12010 4915 12030
rect 4885 12005 4915 12010
rect 4885 11950 4915 11955
rect 4885 11930 4890 11950
rect 4890 11930 4910 11950
rect 4910 11930 4915 11950
rect 4885 11925 4915 11930
rect 4885 11870 4915 11875
rect 4885 11850 4890 11870
rect 4890 11850 4910 11870
rect 4910 11850 4915 11870
rect 4885 11845 4915 11850
rect 4885 11790 4915 11795
rect 4885 11770 4890 11790
rect 4890 11770 4910 11790
rect 4910 11770 4915 11790
rect 4885 11765 4915 11770
rect 4885 11710 4915 11715
rect 4885 11690 4890 11710
rect 4890 11690 4910 11710
rect 4910 11690 4915 11710
rect 4885 11685 4915 11690
rect 4885 11630 4915 11635
rect 4885 11610 4890 11630
rect 4890 11610 4910 11630
rect 4910 11610 4915 11630
rect 4885 11605 4915 11610
rect 4885 11550 4915 11555
rect 4885 11530 4890 11550
rect 4890 11530 4910 11550
rect 4910 11530 4915 11550
rect 4885 11525 4915 11530
rect 4885 11470 4915 11475
rect 4885 11450 4890 11470
rect 4890 11450 4910 11470
rect 4910 11450 4915 11470
rect 4885 11445 4915 11450
rect 4885 11390 4915 11395
rect 4885 11370 4890 11390
rect 4890 11370 4910 11390
rect 4910 11370 4915 11390
rect 4885 11365 4915 11370
rect 4885 11310 4915 11315
rect 4885 11290 4890 11310
rect 4890 11290 4910 11310
rect 4910 11290 4915 11310
rect 4885 11285 4915 11290
rect 4885 11230 4915 11235
rect 4885 11210 4890 11230
rect 4890 11210 4910 11230
rect 4910 11210 4915 11230
rect 4885 11205 4915 11210
rect 4885 11150 4915 11155
rect 4885 11130 4890 11150
rect 4890 11130 4910 11150
rect 4910 11130 4915 11150
rect 4885 11125 4915 11130
rect 4885 11070 4915 11075
rect 4885 11050 4890 11070
rect 4890 11050 4910 11070
rect 4910 11050 4915 11070
rect 4885 11045 4915 11050
rect 4885 10910 4915 10915
rect 4885 10890 4890 10910
rect 4890 10890 4910 10910
rect 4910 10890 4915 10910
rect 4885 10885 4915 10890
rect 4885 10830 4915 10835
rect 4885 10810 4890 10830
rect 4890 10810 4910 10830
rect 4910 10810 4915 10830
rect 4885 10805 4915 10810
rect 4885 10750 4915 10755
rect 4885 10730 4890 10750
rect 4890 10730 4910 10750
rect 4910 10730 4915 10750
rect 4885 10725 4915 10730
rect 4885 10670 4915 10675
rect 4885 10650 4890 10670
rect 4890 10650 4910 10670
rect 4910 10650 4915 10670
rect 4885 10645 4915 10650
rect 4885 10590 4915 10595
rect 4885 10570 4890 10590
rect 4890 10570 4910 10590
rect 4910 10570 4915 10590
rect 4885 10565 4915 10570
rect 4885 10510 4915 10515
rect 4885 10490 4890 10510
rect 4890 10490 4910 10510
rect 4910 10490 4915 10510
rect 4885 10485 4915 10490
rect 4885 10430 4915 10435
rect 4885 10410 4890 10430
rect 4890 10410 4910 10430
rect 4910 10410 4915 10430
rect 4885 10405 4915 10410
rect 4885 10350 4915 10355
rect 4885 10330 4890 10350
rect 4890 10330 4910 10350
rect 4910 10330 4915 10350
rect 4885 10325 4915 10330
rect 4885 9950 4915 9955
rect 4885 9930 4890 9950
rect 4890 9930 4910 9950
rect 4910 9930 4915 9950
rect 4885 9925 4915 9930
rect 4885 9870 4915 9875
rect 4885 9850 4890 9870
rect 4890 9850 4910 9870
rect 4910 9850 4915 9870
rect 4885 9845 4915 9850
rect 4885 9790 4915 9795
rect 4885 9770 4890 9790
rect 4890 9770 4910 9790
rect 4910 9770 4915 9790
rect 4885 9765 4915 9770
rect 4885 9710 4915 9715
rect 4885 9690 4890 9710
rect 4890 9690 4910 9710
rect 4910 9690 4915 9710
rect 4885 9685 4915 9690
rect 4885 9630 4915 9635
rect 4885 9610 4890 9630
rect 4890 9610 4910 9630
rect 4910 9610 4915 9630
rect 4885 9605 4915 9610
rect 4885 9550 4915 9555
rect 4885 9530 4890 9550
rect 4890 9530 4910 9550
rect 4910 9530 4915 9550
rect 4885 9525 4915 9530
rect 4885 9470 4915 9475
rect 4885 9450 4890 9470
rect 4890 9450 4910 9470
rect 4910 9450 4915 9470
rect 4885 9445 4915 9450
rect 4885 9390 4915 9395
rect 4885 9370 4890 9390
rect 4890 9370 4910 9390
rect 4910 9370 4915 9390
rect 4885 9365 4915 9370
rect 4885 8990 4915 8995
rect 4885 8970 4890 8990
rect 4890 8970 4910 8990
rect 4910 8970 4915 8990
rect 4885 8965 4915 8970
rect 4885 8910 4915 8915
rect 4885 8890 4890 8910
rect 4890 8890 4910 8910
rect 4910 8890 4915 8910
rect 4885 8885 4915 8890
rect 4885 8830 4915 8835
rect 4885 8810 4890 8830
rect 4890 8810 4910 8830
rect 4910 8810 4915 8830
rect 4885 8805 4915 8810
rect 4885 8750 4915 8755
rect 4885 8730 4890 8750
rect 4890 8730 4910 8750
rect 4910 8730 4915 8750
rect 4885 8725 4915 8730
rect 4885 8670 4915 8675
rect 4885 8650 4890 8670
rect 4890 8650 4910 8670
rect 4910 8650 4915 8670
rect 4885 8645 4915 8650
rect 4885 8590 4915 8595
rect 4885 8570 4890 8590
rect 4890 8570 4910 8590
rect 4910 8570 4915 8590
rect 4885 8565 4915 8570
rect 4885 8510 4915 8515
rect 4885 8490 4890 8510
rect 4890 8490 4910 8510
rect 4910 8490 4915 8510
rect 4885 8485 4915 8490
rect 4885 8430 4915 8435
rect 4885 8410 4890 8430
rect 4890 8410 4910 8430
rect 4910 8410 4915 8430
rect 4885 8405 4915 8410
rect 4885 8270 4915 8275
rect 4885 8250 4890 8270
rect 4890 8250 4910 8270
rect 4910 8250 4915 8270
rect 4885 8245 4915 8250
rect 4885 8190 4915 8195
rect 4885 8170 4890 8190
rect 4890 8170 4910 8190
rect 4910 8170 4915 8190
rect 4885 8165 4915 8170
rect 4885 8110 4915 8115
rect 4885 8090 4890 8110
rect 4890 8090 4910 8110
rect 4910 8090 4915 8110
rect 4885 8085 4915 8090
rect 4885 8030 4915 8035
rect 4885 8010 4890 8030
rect 4890 8010 4910 8030
rect 4910 8010 4915 8030
rect 4885 8005 4915 8010
rect 4885 7950 4915 7955
rect 4885 7930 4890 7950
rect 4890 7930 4910 7950
rect 4910 7930 4915 7950
rect 4885 7925 4915 7930
rect 4885 7870 4915 7875
rect 4885 7850 4890 7870
rect 4890 7850 4910 7870
rect 4910 7850 4915 7870
rect 4885 7845 4915 7850
rect 4885 7790 4915 7795
rect 4885 7770 4890 7790
rect 4890 7770 4910 7790
rect 4910 7770 4915 7790
rect 4885 7765 4915 7770
rect 4885 7710 4915 7715
rect 4885 7690 4890 7710
rect 4890 7690 4910 7710
rect 4910 7690 4915 7710
rect 4885 7685 4915 7690
rect 4885 7630 4915 7635
rect 4885 7610 4890 7630
rect 4890 7610 4910 7630
rect 4910 7610 4915 7630
rect 4885 7605 4915 7610
rect 4885 7550 4915 7555
rect 4885 7530 4890 7550
rect 4890 7530 4910 7550
rect 4910 7530 4915 7550
rect 4885 7525 4915 7530
rect 4885 7470 4915 7475
rect 4885 7450 4890 7470
rect 4890 7450 4910 7470
rect 4910 7450 4915 7470
rect 4885 7445 4915 7450
rect 4885 7390 4915 7395
rect 4885 7370 4890 7390
rect 4890 7370 4910 7390
rect 4910 7370 4915 7390
rect 4885 7365 4915 7370
rect 4885 7310 4915 7315
rect 4885 7290 4890 7310
rect 4890 7290 4910 7310
rect 4910 7290 4915 7310
rect 4885 7285 4915 7290
rect 4885 7230 4915 7235
rect 4885 7210 4890 7230
rect 4890 7210 4910 7230
rect 4910 7210 4915 7230
rect 4885 7205 4915 7210
rect 4885 7150 4915 7155
rect 4885 7130 4890 7150
rect 4890 7130 4910 7150
rect 4910 7130 4915 7150
rect 4885 7125 4915 7130
rect 4885 7070 4915 7075
rect 4885 7050 4890 7070
rect 4890 7050 4910 7070
rect 4910 7050 4915 7070
rect 4885 7045 4915 7050
rect 4885 6990 4915 6995
rect 4885 6970 4890 6990
rect 4890 6970 4910 6990
rect 4910 6970 4915 6990
rect 4885 6965 4915 6970
rect 4885 6830 4915 6835
rect 4885 6810 4890 6830
rect 4890 6810 4910 6830
rect 4910 6810 4915 6830
rect 4885 6805 4915 6810
rect 4885 6750 4915 6755
rect 4885 6730 4890 6750
rect 4890 6730 4910 6750
rect 4910 6730 4915 6750
rect 4885 6725 4915 6730
rect 4885 6670 4915 6675
rect 4885 6650 4890 6670
rect 4890 6650 4910 6670
rect 4910 6650 4915 6670
rect 4885 6645 4915 6650
rect 4885 6590 4915 6595
rect 4885 6570 4890 6590
rect 4890 6570 4910 6590
rect 4910 6570 4915 6590
rect 4885 6565 4915 6570
rect 4885 6510 4915 6515
rect 4885 6490 4890 6510
rect 4890 6490 4910 6510
rect 4910 6490 4915 6510
rect 4885 6485 4915 6490
rect 4885 6430 4915 6435
rect 4885 6410 4890 6430
rect 4890 6410 4910 6430
rect 4910 6410 4915 6430
rect 4885 6405 4915 6410
rect 4885 6350 4915 6355
rect 4885 6330 4890 6350
rect 4890 6330 4910 6350
rect 4910 6330 4915 6350
rect 4885 6325 4915 6330
rect 4885 6270 4915 6275
rect 4885 6250 4890 6270
rect 4890 6250 4910 6270
rect 4910 6250 4915 6270
rect 4885 6245 4915 6250
rect 4885 5870 4915 5875
rect 4885 5850 4890 5870
rect 4890 5850 4910 5870
rect 4910 5850 4915 5870
rect 4885 5845 4915 5850
rect 4885 5790 4915 5795
rect 4885 5770 4890 5790
rect 4890 5770 4910 5790
rect 4910 5770 4915 5790
rect 4885 5765 4915 5770
rect 4885 5710 4915 5715
rect 4885 5690 4890 5710
rect 4890 5690 4910 5710
rect 4910 5690 4915 5710
rect 4885 5685 4915 5690
rect 4885 5630 4915 5635
rect 4885 5610 4890 5630
rect 4890 5610 4910 5630
rect 4910 5610 4915 5630
rect 4885 5605 4915 5610
rect 4885 5550 4915 5555
rect 4885 5530 4890 5550
rect 4890 5530 4910 5550
rect 4910 5530 4915 5550
rect 4885 5525 4915 5530
rect 4885 5470 4915 5475
rect 4885 5450 4890 5470
rect 4890 5450 4910 5470
rect 4910 5450 4915 5470
rect 4885 5445 4915 5450
rect 4885 5390 4915 5395
rect 4885 5370 4890 5390
rect 4890 5370 4910 5390
rect 4910 5370 4915 5390
rect 4885 5365 4915 5370
rect 4885 5310 4915 5315
rect 4885 5290 4890 5310
rect 4890 5290 4910 5310
rect 4910 5290 4915 5310
rect 4885 5285 4915 5290
rect 4885 5230 4915 5235
rect 4885 5210 4890 5230
rect 4890 5210 4910 5230
rect 4910 5210 4915 5230
rect 4885 5205 4915 5210
rect 4885 5150 4915 5155
rect 4885 5130 4890 5150
rect 4890 5130 4910 5150
rect 4910 5130 4915 5150
rect 4885 5125 4915 5130
rect 4885 5070 4915 5075
rect 4885 5050 4890 5070
rect 4890 5050 4910 5070
rect 4910 5050 4915 5070
rect 4885 5045 4915 5050
rect 4885 4990 4915 4995
rect 4885 4970 4890 4990
rect 4890 4970 4910 4990
rect 4910 4970 4915 4990
rect 4885 4965 4915 4970
rect 4885 4910 4915 4915
rect 4885 4890 4890 4910
rect 4890 4890 4910 4910
rect 4910 4890 4915 4910
rect 4885 4885 4915 4890
rect 4885 4750 4915 4755
rect 4885 4730 4890 4750
rect 4890 4730 4910 4750
rect 4910 4730 4915 4750
rect 4885 4725 4915 4730
rect 4885 4670 4915 4675
rect 4885 4650 4890 4670
rect 4890 4650 4910 4670
rect 4910 4650 4915 4670
rect 4885 4645 4915 4650
rect 4885 4510 4915 4515
rect 4885 4490 4890 4510
rect 4890 4490 4910 4510
rect 4910 4490 4915 4510
rect 4885 4485 4915 4490
rect 4885 4430 4915 4435
rect 4885 4410 4890 4430
rect 4890 4410 4910 4430
rect 4910 4410 4915 4430
rect 4885 4405 4915 4410
rect 4885 4350 4915 4355
rect 4885 4330 4890 4350
rect 4890 4330 4910 4350
rect 4910 4330 4915 4350
rect 4885 4325 4915 4330
rect 4885 4270 4915 4275
rect 4885 4250 4890 4270
rect 4890 4250 4910 4270
rect 4910 4250 4915 4270
rect 4885 4245 4915 4250
rect 4885 4190 4915 4195
rect 4885 4170 4890 4190
rect 4890 4170 4910 4190
rect 4910 4170 4915 4190
rect 4885 4165 4915 4170
rect 4885 4110 4915 4115
rect 4885 4090 4890 4110
rect 4890 4090 4910 4110
rect 4910 4090 4915 4110
rect 4885 4085 4915 4090
rect 4885 4030 4915 4035
rect 4885 4010 4890 4030
rect 4890 4010 4910 4030
rect 4910 4010 4915 4030
rect 4885 4005 4915 4010
rect 4885 3950 4915 3955
rect 4885 3930 4890 3950
rect 4890 3930 4910 3950
rect 4910 3930 4915 3950
rect 4885 3925 4915 3930
rect 4885 3870 4915 3875
rect 4885 3850 4890 3870
rect 4890 3850 4910 3870
rect 4910 3850 4915 3870
rect 4885 3845 4915 3850
rect 4885 3710 4915 3715
rect 4885 3690 4890 3710
rect 4890 3690 4910 3710
rect 4910 3690 4915 3710
rect 4885 3685 4915 3690
rect 4885 3630 4915 3635
rect 4885 3610 4890 3630
rect 4890 3610 4910 3630
rect 4910 3610 4915 3630
rect 4885 3605 4915 3610
rect 4885 3470 4915 3475
rect 4885 3450 4890 3470
rect 4890 3450 4910 3470
rect 4910 3450 4915 3470
rect 4885 3445 4915 3450
rect 4885 3390 4915 3395
rect 4885 3370 4890 3390
rect 4890 3370 4910 3390
rect 4910 3370 4915 3390
rect 4885 3365 4915 3370
rect 4885 3230 4915 3235
rect 4885 3210 4890 3230
rect 4890 3210 4910 3230
rect 4910 3210 4915 3230
rect 4885 3205 4915 3210
rect 4885 3150 4915 3155
rect 4885 3130 4890 3150
rect 4890 3130 4910 3150
rect 4910 3130 4915 3150
rect 4885 3125 4915 3130
rect 4885 3070 4915 3075
rect 4885 3050 4890 3070
rect 4890 3050 4910 3070
rect 4910 3050 4915 3070
rect 4885 3045 4915 3050
rect 4885 2990 4915 2995
rect 4885 2970 4890 2990
rect 4890 2970 4910 2990
rect 4910 2970 4915 2990
rect 4885 2965 4915 2970
rect 4885 2910 4915 2915
rect 4885 2890 4890 2910
rect 4890 2890 4910 2910
rect 4910 2890 4915 2910
rect 4885 2885 4915 2890
rect 4885 2830 4915 2835
rect 4885 2810 4890 2830
rect 4890 2810 4910 2830
rect 4910 2810 4915 2830
rect 4885 2805 4915 2810
rect 4885 2750 4915 2755
rect 4885 2730 4890 2750
rect 4890 2730 4910 2750
rect 4910 2730 4915 2750
rect 4885 2725 4915 2730
rect 4885 2670 4915 2675
rect 4885 2650 4890 2670
rect 4890 2650 4910 2670
rect 4910 2650 4915 2670
rect 4885 2645 4915 2650
rect 4885 2590 4915 2595
rect 4885 2570 4890 2590
rect 4890 2570 4910 2590
rect 4910 2570 4915 2590
rect 4885 2565 4915 2570
rect 4885 2510 4915 2515
rect 4885 2490 4890 2510
rect 4890 2490 4910 2510
rect 4910 2490 4915 2510
rect 4885 2485 4915 2490
rect 4885 2430 4915 2435
rect 4885 2410 4890 2430
rect 4890 2410 4910 2430
rect 4910 2410 4915 2430
rect 4885 2405 4915 2410
rect 4885 2350 4915 2355
rect 4885 2330 4890 2350
rect 4890 2330 4910 2350
rect 4910 2330 4915 2350
rect 4885 2325 4915 2330
rect 4885 2270 4915 2275
rect 4885 2250 4890 2270
rect 4890 2250 4910 2270
rect 4910 2250 4915 2270
rect 4885 2245 4915 2250
rect 4885 2190 4915 2195
rect 4885 2170 4890 2190
rect 4890 2170 4910 2190
rect 4910 2170 4915 2190
rect 4885 2165 4915 2170
rect 4885 2110 4915 2115
rect 4885 2090 4890 2110
rect 4890 2090 4910 2110
rect 4910 2090 4915 2110
rect 4885 2085 4915 2090
rect 4885 2030 4915 2035
rect 4885 2010 4890 2030
rect 4890 2010 4910 2030
rect 4910 2010 4915 2030
rect 4885 2005 4915 2010
rect 4885 1950 4915 1955
rect 4885 1930 4890 1950
rect 4890 1930 4910 1950
rect 4910 1930 4915 1950
rect 4885 1925 4915 1930
rect 4885 1710 4915 1715
rect 4885 1690 4890 1710
rect 4890 1690 4910 1710
rect 4910 1690 4915 1710
rect 4885 1685 4915 1690
rect 4885 1630 4915 1635
rect 4885 1610 4890 1630
rect 4890 1610 4910 1630
rect 4910 1610 4915 1630
rect 4885 1605 4915 1610
rect 4885 1550 4915 1555
rect 4885 1530 4890 1550
rect 4890 1530 4910 1550
rect 4910 1530 4915 1550
rect 4885 1525 4915 1530
rect 4885 1470 4915 1475
rect 4885 1450 4890 1470
rect 4890 1450 4910 1470
rect 4910 1450 4915 1470
rect 4885 1445 4915 1450
rect 4885 1390 4915 1395
rect 4885 1370 4890 1390
rect 4890 1370 4910 1390
rect 4910 1370 4915 1390
rect 4885 1365 4915 1370
rect 4885 1310 4915 1315
rect 4885 1290 4890 1310
rect 4890 1290 4910 1310
rect 4910 1290 4915 1310
rect 4885 1285 4915 1290
rect 4885 1230 4915 1235
rect 4885 1210 4890 1230
rect 4890 1210 4910 1230
rect 4910 1210 4915 1230
rect 4885 1205 4915 1210
rect 4885 1150 4915 1155
rect 4885 1130 4890 1150
rect 4890 1130 4910 1150
rect 4910 1130 4915 1150
rect 4885 1125 4915 1130
rect 4885 1070 4915 1075
rect 4885 1050 4890 1070
rect 4890 1050 4910 1070
rect 4910 1050 4915 1070
rect 4885 1045 4915 1050
rect 4885 990 4915 995
rect 4885 970 4890 990
rect 4890 970 4910 990
rect 4910 970 4915 990
rect 4885 965 4915 970
rect 4885 830 4915 835
rect 4885 810 4890 830
rect 4890 810 4910 830
rect 4910 810 4915 830
rect 4885 805 4915 810
rect 4885 750 4915 755
rect 4885 730 4890 750
rect 4890 730 4910 750
rect 4910 730 4915 750
rect 4885 725 4915 730
rect 4885 670 4915 675
rect 4885 650 4890 670
rect 4890 650 4910 670
rect 4910 650 4915 670
rect 4885 645 4915 650
rect 4885 590 4915 595
rect 4885 570 4890 590
rect 4890 570 4910 590
rect 4910 570 4915 590
rect 4885 565 4915 570
rect 4885 510 4915 515
rect 4885 490 4890 510
rect 4890 490 4910 510
rect 4910 490 4915 510
rect 4885 485 4915 490
rect 4885 270 4915 275
rect 4885 250 4890 270
rect 4890 250 4910 270
rect 4910 250 4915 270
rect 4885 245 4915 250
rect 4885 190 4915 195
rect 4885 170 4890 190
rect 4890 170 4910 190
rect 4910 170 4915 190
rect 4885 165 4915 170
rect 4885 110 4915 115
rect 4885 90 4890 110
rect 4890 90 4910 110
rect 4910 90 4915 110
rect 4885 85 4915 90
rect 4885 30 4915 35
rect 4885 10 4890 30
rect 4890 10 4910 30
rect 4910 10 4915 30
rect 4885 5 4915 10
rect 5045 15710 5075 15715
rect 5045 15690 5050 15710
rect 5050 15690 5070 15710
rect 5070 15690 5075 15710
rect 5045 15685 5075 15690
rect 5045 15630 5075 15635
rect 5045 15610 5050 15630
rect 5050 15610 5070 15630
rect 5070 15610 5075 15630
rect 5045 15605 5075 15610
rect 5045 15550 5075 15555
rect 5045 15530 5050 15550
rect 5050 15530 5070 15550
rect 5070 15530 5075 15550
rect 5045 15525 5075 15530
rect 5045 15470 5075 15475
rect 5045 15450 5050 15470
rect 5050 15450 5070 15470
rect 5070 15450 5075 15470
rect 5045 15445 5075 15450
rect 5045 15390 5075 15395
rect 5045 15370 5050 15390
rect 5050 15370 5070 15390
rect 5070 15370 5075 15390
rect 5045 15365 5075 15370
rect 5045 15310 5075 15315
rect 5045 15290 5050 15310
rect 5050 15290 5070 15310
rect 5070 15290 5075 15310
rect 5045 15285 5075 15290
rect 5045 15230 5075 15235
rect 5045 15210 5050 15230
rect 5050 15210 5070 15230
rect 5070 15210 5075 15230
rect 5045 15205 5075 15210
rect 5045 15150 5075 15155
rect 5045 15130 5050 15150
rect 5050 15130 5070 15150
rect 5070 15130 5075 15150
rect 5045 15125 5075 15130
rect 5045 14990 5075 14995
rect 5045 14970 5050 14990
rect 5050 14970 5070 14990
rect 5070 14970 5075 14990
rect 5045 14965 5075 14970
rect 5045 14910 5075 14915
rect 5045 14890 5050 14910
rect 5050 14890 5070 14910
rect 5070 14890 5075 14910
rect 5045 14885 5075 14890
rect 5045 14830 5075 14835
rect 5045 14810 5050 14830
rect 5050 14810 5070 14830
rect 5070 14810 5075 14830
rect 5045 14805 5075 14810
rect 5045 14750 5075 14755
rect 5045 14730 5050 14750
rect 5050 14730 5070 14750
rect 5070 14730 5075 14750
rect 5045 14725 5075 14730
rect 5045 14670 5075 14675
rect 5045 14650 5050 14670
rect 5050 14650 5070 14670
rect 5070 14650 5075 14670
rect 5045 14645 5075 14650
rect 5045 14590 5075 14595
rect 5045 14570 5050 14590
rect 5050 14570 5070 14590
rect 5070 14570 5075 14590
rect 5045 14565 5075 14570
rect 5045 14510 5075 14515
rect 5045 14490 5050 14510
rect 5050 14490 5070 14510
rect 5070 14490 5075 14510
rect 5045 14485 5075 14490
rect 5045 14430 5075 14435
rect 5045 14410 5050 14430
rect 5050 14410 5070 14430
rect 5070 14410 5075 14430
rect 5045 14405 5075 14410
rect 5045 14030 5075 14035
rect 5045 14010 5050 14030
rect 5050 14010 5070 14030
rect 5070 14010 5075 14030
rect 5045 14005 5075 14010
rect 5045 13950 5075 13955
rect 5045 13930 5050 13950
rect 5050 13930 5070 13950
rect 5070 13930 5075 13950
rect 5045 13925 5075 13930
rect 5045 13870 5075 13875
rect 5045 13850 5050 13870
rect 5050 13850 5070 13870
rect 5070 13850 5075 13870
rect 5045 13845 5075 13850
rect 5045 13790 5075 13795
rect 5045 13770 5050 13790
rect 5050 13770 5070 13790
rect 5070 13770 5075 13790
rect 5045 13765 5075 13770
rect 5045 13710 5075 13715
rect 5045 13690 5050 13710
rect 5050 13690 5070 13710
rect 5070 13690 5075 13710
rect 5045 13685 5075 13690
rect 5045 13630 5075 13635
rect 5045 13610 5050 13630
rect 5050 13610 5070 13630
rect 5070 13610 5075 13630
rect 5045 13605 5075 13610
rect 5045 13550 5075 13555
rect 5045 13530 5050 13550
rect 5050 13530 5070 13550
rect 5070 13530 5075 13550
rect 5045 13525 5075 13530
rect 5045 13470 5075 13475
rect 5045 13450 5050 13470
rect 5050 13450 5070 13470
rect 5070 13450 5075 13470
rect 5045 13445 5075 13450
rect 5045 13070 5075 13075
rect 5045 13050 5050 13070
rect 5050 13050 5070 13070
rect 5070 13050 5075 13070
rect 5045 13045 5075 13050
rect 5045 12990 5075 12995
rect 5045 12970 5050 12990
rect 5050 12970 5070 12990
rect 5070 12970 5075 12990
rect 5045 12965 5075 12970
rect 5045 12910 5075 12915
rect 5045 12890 5050 12910
rect 5050 12890 5070 12910
rect 5070 12890 5075 12910
rect 5045 12885 5075 12890
rect 5045 12830 5075 12835
rect 5045 12810 5050 12830
rect 5050 12810 5070 12830
rect 5070 12810 5075 12830
rect 5045 12805 5075 12810
rect 5045 12750 5075 12755
rect 5045 12730 5050 12750
rect 5050 12730 5070 12750
rect 5070 12730 5075 12750
rect 5045 12725 5075 12730
rect 5045 12670 5075 12675
rect 5045 12650 5050 12670
rect 5050 12650 5070 12670
rect 5070 12650 5075 12670
rect 5045 12645 5075 12650
rect 5045 12590 5075 12595
rect 5045 12570 5050 12590
rect 5050 12570 5070 12590
rect 5070 12570 5075 12590
rect 5045 12565 5075 12570
rect 5045 12510 5075 12515
rect 5045 12490 5050 12510
rect 5050 12490 5070 12510
rect 5070 12490 5075 12510
rect 5045 12485 5075 12490
rect 5045 12350 5075 12355
rect 5045 12330 5050 12350
rect 5050 12330 5070 12350
rect 5070 12330 5075 12350
rect 5045 12325 5075 12330
rect 5045 12270 5075 12275
rect 5045 12250 5050 12270
rect 5050 12250 5070 12270
rect 5070 12250 5075 12270
rect 5045 12245 5075 12250
rect 5045 12190 5075 12195
rect 5045 12170 5050 12190
rect 5050 12170 5070 12190
rect 5070 12170 5075 12190
rect 5045 12165 5075 12170
rect 5045 12110 5075 12115
rect 5045 12090 5050 12110
rect 5050 12090 5070 12110
rect 5070 12090 5075 12110
rect 5045 12085 5075 12090
rect 5045 12030 5075 12035
rect 5045 12010 5050 12030
rect 5050 12010 5070 12030
rect 5070 12010 5075 12030
rect 5045 12005 5075 12010
rect 5045 11950 5075 11955
rect 5045 11930 5050 11950
rect 5050 11930 5070 11950
rect 5070 11930 5075 11950
rect 5045 11925 5075 11930
rect 5045 11870 5075 11875
rect 5045 11850 5050 11870
rect 5050 11850 5070 11870
rect 5070 11850 5075 11870
rect 5045 11845 5075 11850
rect 5045 11790 5075 11795
rect 5045 11770 5050 11790
rect 5050 11770 5070 11790
rect 5070 11770 5075 11790
rect 5045 11765 5075 11770
rect 5045 11710 5075 11715
rect 5045 11690 5050 11710
rect 5050 11690 5070 11710
rect 5070 11690 5075 11710
rect 5045 11685 5075 11690
rect 5045 11630 5075 11635
rect 5045 11610 5050 11630
rect 5050 11610 5070 11630
rect 5070 11610 5075 11630
rect 5045 11605 5075 11610
rect 5045 11550 5075 11555
rect 5045 11530 5050 11550
rect 5050 11530 5070 11550
rect 5070 11530 5075 11550
rect 5045 11525 5075 11530
rect 5045 11470 5075 11475
rect 5045 11450 5050 11470
rect 5050 11450 5070 11470
rect 5070 11450 5075 11470
rect 5045 11445 5075 11450
rect 5045 11390 5075 11395
rect 5045 11370 5050 11390
rect 5050 11370 5070 11390
rect 5070 11370 5075 11390
rect 5045 11365 5075 11370
rect 5045 11310 5075 11315
rect 5045 11290 5050 11310
rect 5050 11290 5070 11310
rect 5070 11290 5075 11310
rect 5045 11285 5075 11290
rect 5045 11230 5075 11235
rect 5045 11210 5050 11230
rect 5050 11210 5070 11230
rect 5070 11210 5075 11230
rect 5045 11205 5075 11210
rect 5045 11150 5075 11155
rect 5045 11130 5050 11150
rect 5050 11130 5070 11150
rect 5070 11130 5075 11150
rect 5045 11125 5075 11130
rect 5045 11070 5075 11075
rect 5045 11050 5050 11070
rect 5050 11050 5070 11070
rect 5070 11050 5075 11070
rect 5045 11045 5075 11050
rect 5045 10910 5075 10915
rect 5045 10890 5050 10910
rect 5050 10890 5070 10910
rect 5070 10890 5075 10910
rect 5045 10885 5075 10890
rect 5045 10830 5075 10835
rect 5045 10810 5050 10830
rect 5050 10810 5070 10830
rect 5070 10810 5075 10830
rect 5045 10805 5075 10810
rect 5045 10750 5075 10755
rect 5045 10730 5050 10750
rect 5050 10730 5070 10750
rect 5070 10730 5075 10750
rect 5045 10725 5075 10730
rect 5045 10670 5075 10675
rect 5045 10650 5050 10670
rect 5050 10650 5070 10670
rect 5070 10650 5075 10670
rect 5045 10645 5075 10650
rect 5045 10590 5075 10595
rect 5045 10570 5050 10590
rect 5050 10570 5070 10590
rect 5070 10570 5075 10590
rect 5045 10565 5075 10570
rect 5045 10510 5075 10515
rect 5045 10490 5050 10510
rect 5050 10490 5070 10510
rect 5070 10490 5075 10510
rect 5045 10485 5075 10490
rect 5045 10430 5075 10435
rect 5045 10410 5050 10430
rect 5050 10410 5070 10430
rect 5070 10410 5075 10430
rect 5045 10405 5075 10410
rect 5045 10350 5075 10355
rect 5045 10330 5050 10350
rect 5050 10330 5070 10350
rect 5070 10330 5075 10350
rect 5045 10325 5075 10330
rect 5045 9950 5075 9955
rect 5045 9930 5050 9950
rect 5050 9930 5070 9950
rect 5070 9930 5075 9950
rect 5045 9925 5075 9930
rect 5045 9870 5075 9875
rect 5045 9850 5050 9870
rect 5050 9850 5070 9870
rect 5070 9850 5075 9870
rect 5045 9845 5075 9850
rect 5045 9790 5075 9795
rect 5045 9770 5050 9790
rect 5050 9770 5070 9790
rect 5070 9770 5075 9790
rect 5045 9765 5075 9770
rect 5045 9710 5075 9715
rect 5045 9690 5050 9710
rect 5050 9690 5070 9710
rect 5070 9690 5075 9710
rect 5045 9685 5075 9690
rect 5045 9630 5075 9635
rect 5045 9610 5050 9630
rect 5050 9610 5070 9630
rect 5070 9610 5075 9630
rect 5045 9605 5075 9610
rect 5045 9550 5075 9555
rect 5045 9530 5050 9550
rect 5050 9530 5070 9550
rect 5070 9530 5075 9550
rect 5045 9525 5075 9530
rect 5045 9470 5075 9475
rect 5045 9450 5050 9470
rect 5050 9450 5070 9470
rect 5070 9450 5075 9470
rect 5045 9445 5075 9450
rect 5045 9390 5075 9395
rect 5045 9370 5050 9390
rect 5050 9370 5070 9390
rect 5070 9370 5075 9390
rect 5045 9365 5075 9370
rect 5045 8990 5075 8995
rect 5045 8970 5050 8990
rect 5050 8970 5070 8990
rect 5070 8970 5075 8990
rect 5045 8965 5075 8970
rect 5045 8910 5075 8915
rect 5045 8890 5050 8910
rect 5050 8890 5070 8910
rect 5070 8890 5075 8910
rect 5045 8885 5075 8890
rect 5045 8830 5075 8835
rect 5045 8810 5050 8830
rect 5050 8810 5070 8830
rect 5070 8810 5075 8830
rect 5045 8805 5075 8810
rect 5045 8750 5075 8755
rect 5045 8730 5050 8750
rect 5050 8730 5070 8750
rect 5070 8730 5075 8750
rect 5045 8725 5075 8730
rect 5045 8670 5075 8675
rect 5045 8650 5050 8670
rect 5050 8650 5070 8670
rect 5070 8650 5075 8670
rect 5045 8645 5075 8650
rect 5045 8590 5075 8595
rect 5045 8570 5050 8590
rect 5050 8570 5070 8590
rect 5070 8570 5075 8590
rect 5045 8565 5075 8570
rect 5045 8510 5075 8515
rect 5045 8490 5050 8510
rect 5050 8490 5070 8510
rect 5070 8490 5075 8510
rect 5045 8485 5075 8490
rect 5045 8430 5075 8435
rect 5045 8410 5050 8430
rect 5050 8410 5070 8430
rect 5070 8410 5075 8430
rect 5045 8405 5075 8410
rect 5045 8270 5075 8275
rect 5045 8250 5050 8270
rect 5050 8250 5070 8270
rect 5070 8250 5075 8270
rect 5045 8245 5075 8250
rect 5045 8190 5075 8195
rect 5045 8170 5050 8190
rect 5050 8170 5070 8190
rect 5070 8170 5075 8190
rect 5045 8165 5075 8170
rect 5045 8110 5075 8115
rect 5045 8090 5050 8110
rect 5050 8090 5070 8110
rect 5070 8090 5075 8110
rect 5045 8085 5075 8090
rect 5045 8030 5075 8035
rect 5045 8010 5050 8030
rect 5050 8010 5070 8030
rect 5070 8010 5075 8030
rect 5045 8005 5075 8010
rect 5045 7950 5075 7955
rect 5045 7930 5050 7950
rect 5050 7930 5070 7950
rect 5070 7930 5075 7950
rect 5045 7925 5075 7930
rect 5045 7870 5075 7875
rect 5045 7850 5050 7870
rect 5050 7850 5070 7870
rect 5070 7850 5075 7870
rect 5045 7845 5075 7850
rect 5045 7790 5075 7795
rect 5045 7770 5050 7790
rect 5050 7770 5070 7790
rect 5070 7770 5075 7790
rect 5045 7765 5075 7770
rect 5045 7710 5075 7715
rect 5045 7690 5050 7710
rect 5050 7690 5070 7710
rect 5070 7690 5075 7710
rect 5045 7685 5075 7690
rect 5045 7630 5075 7635
rect 5045 7610 5050 7630
rect 5050 7610 5070 7630
rect 5070 7610 5075 7630
rect 5045 7605 5075 7610
rect 5045 7550 5075 7555
rect 5045 7530 5050 7550
rect 5050 7530 5070 7550
rect 5070 7530 5075 7550
rect 5045 7525 5075 7530
rect 5045 7470 5075 7475
rect 5045 7450 5050 7470
rect 5050 7450 5070 7470
rect 5070 7450 5075 7470
rect 5045 7445 5075 7450
rect 5045 7390 5075 7395
rect 5045 7370 5050 7390
rect 5050 7370 5070 7390
rect 5070 7370 5075 7390
rect 5045 7365 5075 7370
rect 5045 7310 5075 7315
rect 5045 7290 5050 7310
rect 5050 7290 5070 7310
rect 5070 7290 5075 7310
rect 5045 7285 5075 7290
rect 5045 7230 5075 7235
rect 5045 7210 5050 7230
rect 5050 7210 5070 7230
rect 5070 7210 5075 7230
rect 5045 7205 5075 7210
rect 5045 7150 5075 7155
rect 5045 7130 5050 7150
rect 5050 7130 5070 7150
rect 5070 7130 5075 7150
rect 5045 7125 5075 7130
rect 5045 7070 5075 7075
rect 5045 7050 5050 7070
rect 5050 7050 5070 7070
rect 5070 7050 5075 7070
rect 5045 7045 5075 7050
rect 5045 6990 5075 6995
rect 5045 6970 5050 6990
rect 5050 6970 5070 6990
rect 5070 6970 5075 6990
rect 5045 6965 5075 6970
rect 5045 6830 5075 6835
rect 5045 6810 5050 6830
rect 5050 6810 5070 6830
rect 5070 6810 5075 6830
rect 5045 6805 5075 6810
rect 5045 6750 5075 6755
rect 5045 6730 5050 6750
rect 5050 6730 5070 6750
rect 5070 6730 5075 6750
rect 5045 6725 5075 6730
rect 5045 6670 5075 6675
rect 5045 6650 5050 6670
rect 5050 6650 5070 6670
rect 5070 6650 5075 6670
rect 5045 6645 5075 6650
rect 5045 6590 5075 6595
rect 5045 6570 5050 6590
rect 5050 6570 5070 6590
rect 5070 6570 5075 6590
rect 5045 6565 5075 6570
rect 5045 6510 5075 6515
rect 5045 6490 5050 6510
rect 5050 6490 5070 6510
rect 5070 6490 5075 6510
rect 5045 6485 5075 6490
rect 5045 6430 5075 6435
rect 5045 6410 5050 6430
rect 5050 6410 5070 6430
rect 5070 6410 5075 6430
rect 5045 6405 5075 6410
rect 5045 6350 5075 6355
rect 5045 6330 5050 6350
rect 5050 6330 5070 6350
rect 5070 6330 5075 6350
rect 5045 6325 5075 6330
rect 5045 6270 5075 6275
rect 5045 6250 5050 6270
rect 5050 6250 5070 6270
rect 5070 6250 5075 6270
rect 5045 6245 5075 6250
rect 5045 5870 5075 5875
rect 5045 5850 5050 5870
rect 5050 5850 5070 5870
rect 5070 5850 5075 5870
rect 5045 5845 5075 5850
rect 5045 5790 5075 5795
rect 5045 5770 5050 5790
rect 5050 5770 5070 5790
rect 5070 5770 5075 5790
rect 5045 5765 5075 5770
rect 5045 5710 5075 5715
rect 5045 5690 5050 5710
rect 5050 5690 5070 5710
rect 5070 5690 5075 5710
rect 5045 5685 5075 5690
rect 5045 5630 5075 5635
rect 5045 5610 5050 5630
rect 5050 5610 5070 5630
rect 5070 5610 5075 5630
rect 5045 5605 5075 5610
rect 5045 5550 5075 5555
rect 5045 5530 5050 5550
rect 5050 5530 5070 5550
rect 5070 5530 5075 5550
rect 5045 5525 5075 5530
rect 5045 5470 5075 5475
rect 5045 5450 5050 5470
rect 5050 5450 5070 5470
rect 5070 5450 5075 5470
rect 5045 5445 5075 5450
rect 5045 5390 5075 5395
rect 5045 5370 5050 5390
rect 5050 5370 5070 5390
rect 5070 5370 5075 5390
rect 5045 5365 5075 5370
rect 5045 5310 5075 5315
rect 5045 5290 5050 5310
rect 5050 5290 5070 5310
rect 5070 5290 5075 5310
rect 5045 5285 5075 5290
rect 5045 5230 5075 5235
rect 5045 5210 5050 5230
rect 5050 5210 5070 5230
rect 5070 5210 5075 5230
rect 5045 5205 5075 5210
rect 5045 5150 5075 5155
rect 5045 5130 5050 5150
rect 5050 5130 5070 5150
rect 5070 5130 5075 5150
rect 5045 5125 5075 5130
rect 5045 5070 5075 5075
rect 5045 5050 5050 5070
rect 5050 5050 5070 5070
rect 5070 5050 5075 5070
rect 5045 5045 5075 5050
rect 5045 4990 5075 4995
rect 5045 4970 5050 4990
rect 5050 4970 5070 4990
rect 5070 4970 5075 4990
rect 5045 4965 5075 4970
rect 5045 4910 5075 4915
rect 5045 4890 5050 4910
rect 5050 4890 5070 4910
rect 5070 4890 5075 4910
rect 5045 4885 5075 4890
rect 5045 4750 5075 4755
rect 5045 4730 5050 4750
rect 5050 4730 5070 4750
rect 5070 4730 5075 4750
rect 5045 4725 5075 4730
rect 5045 4670 5075 4675
rect 5045 4650 5050 4670
rect 5050 4650 5070 4670
rect 5070 4650 5075 4670
rect 5045 4645 5075 4650
rect 5045 4510 5075 4515
rect 5045 4490 5050 4510
rect 5050 4490 5070 4510
rect 5070 4490 5075 4510
rect 5045 4485 5075 4490
rect 5045 4430 5075 4435
rect 5045 4410 5050 4430
rect 5050 4410 5070 4430
rect 5070 4410 5075 4430
rect 5045 4405 5075 4410
rect 5045 4350 5075 4355
rect 5045 4330 5050 4350
rect 5050 4330 5070 4350
rect 5070 4330 5075 4350
rect 5045 4325 5075 4330
rect 5045 4270 5075 4275
rect 5045 4250 5050 4270
rect 5050 4250 5070 4270
rect 5070 4250 5075 4270
rect 5045 4245 5075 4250
rect 5045 4190 5075 4195
rect 5045 4170 5050 4190
rect 5050 4170 5070 4190
rect 5070 4170 5075 4190
rect 5045 4165 5075 4170
rect 5045 4110 5075 4115
rect 5045 4090 5050 4110
rect 5050 4090 5070 4110
rect 5070 4090 5075 4110
rect 5045 4085 5075 4090
rect 5045 4030 5075 4035
rect 5045 4010 5050 4030
rect 5050 4010 5070 4030
rect 5070 4010 5075 4030
rect 5045 4005 5075 4010
rect 5045 3950 5075 3955
rect 5045 3930 5050 3950
rect 5050 3930 5070 3950
rect 5070 3930 5075 3950
rect 5045 3925 5075 3930
rect 5045 3870 5075 3875
rect 5045 3850 5050 3870
rect 5050 3850 5070 3870
rect 5070 3850 5075 3870
rect 5045 3845 5075 3850
rect 5045 3710 5075 3715
rect 5045 3690 5050 3710
rect 5050 3690 5070 3710
rect 5070 3690 5075 3710
rect 5045 3685 5075 3690
rect 5045 3630 5075 3635
rect 5045 3610 5050 3630
rect 5050 3610 5070 3630
rect 5070 3610 5075 3630
rect 5045 3605 5075 3610
rect 5045 3470 5075 3475
rect 5045 3450 5050 3470
rect 5050 3450 5070 3470
rect 5070 3450 5075 3470
rect 5045 3445 5075 3450
rect 5045 3390 5075 3395
rect 5045 3370 5050 3390
rect 5050 3370 5070 3390
rect 5070 3370 5075 3390
rect 5045 3365 5075 3370
rect 5045 3230 5075 3235
rect 5045 3210 5050 3230
rect 5050 3210 5070 3230
rect 5070 3210 5075 3230
rect 5045 3205 5075 3210
rect 5045 3150 5075 3155
rect 5045 3130 5050 3150
rect 5050 3130 5070 3150
rect 5070 3130 5075 3150
rect 5045 3125 5075 3130
rect 5045 3070 5075 3075
rect 5045 3050 5050 3070
rect 5050 3050 5070 3070
rect 5070 3050 5075 3070
rect 5045 3045 5075 3050
rect 5045 2990 5075 2995
rect 5045 2970 5050 2990
rect 5050 2970 5070 2990
rect 5070 2970 5075 2990
rect 5045 2965 5075 2970
rect 5045 2910 5075 2915
rect 5045 2890 5050 2910
rect 5050 2890 5070 2910
rect 5070 2890 5075 2910
rect 5045 2885 5075 2890
rect 5045 2830 5075 2835
rect 5045 2810 5050 2830
rect 5050 2810 5070 2830
rect 5070 2810 5075 2830
rect 5045 2805 5075 2810
rect 5045 2750 5075 2755
rect 5045 2730 5050 2750
rect 5050 2730 5070 2750
rect 5070 2730 5075 2750
rect 5045 2725 5075 2730
rect 5045 2670 5075 2675
rect 5045 2650 5050 2670
rect 5050 2650 5070 2670
rect 5070 2650 5075 2670
rect 5045 2645 5075 2650
rect 5045 2590 5075 2595
rect 5045 2570 5050 2590
rect 5050 2570 5070 2590
rect 5070 2570 5075 2590
rect 5045 2565 5075 2570
rect 5045 2510 5075 2515
rect 5045 2490 5050 2510
rect 5050 2490 5070 2510
rect 5070 2490 5075 2510
rect 5045 2485 5075 2490
rect 5045 2430 5075 2435
rect 5045 2410 5050 2430
rect 5050 2410 5070 2430
rect 5070 2410 5075 2430
rect 5045 2405 5075 2410
rect 5045 2350 5075 2355
rect 5045 2330 5050 2350
rect 5050 2330 5070 2350
rect 5070 2330 5075 2350
rect 5045 2325 5075 2330
rect 5045 2270 5075 2275
rect 5045 2250 5050 2270
rect 5050 2250 5070 2270
rect 5070 2250 5075 2270
rect 5045 2245 5075 2250
rect 5045 2190 5075 2195
rect 5045 2170 5050 2190
rect 5050 2170 5070 2190
rect 5070 2170 5075 2190
rect 5045 2165 5075 2170
rect 5045 2110 5075 2115
rect 5045 2090 5050 2110
rect 5050 2090 5070 2110
rect 5070 2090 5075 2110
rect 5045 2085 5075 2090
rect 5045 2030 5075 2035
rect 5045 2010 5050 2030
rect 5050 2010 5070 2030
rect 5070 2010 5075 2030
rect 5045 2005 5075 2010
rect 5045 1950 5075 1955
rect 5045 1930 5050 1950
rect 5050 1930 5070 1950
rect 5070 1930 5075 1950
rect 5045 1925 5075 1930
rect 5045 1710 5075 1715
rect 5045 1690 5050 1710
rect 5050 1690 5070 1710
rect 5070 1690 5075 1710
rect 5045 1685 5075 1690
rect 5045 1630 5075 1635
rect 5045 1610 5050 1630
rect 5050 1610 5070 1630
rect 5070 1610 5075 1630
rect 5045 1605 5075 1610
rect 5045 1550 5075 1555
rect 5045 1530 5050 1550
rect 5050 1530 5070 1550
rect 5070 1530 5075 1550
rect 5045 1525 5075 1530
rect 5045 1470 5075 1475
rect 5045 1450 5050 1470
rect 5050 1450 5070 1470
rect 5070 1450 5075 1470
rect 5045 1445 5075 1450
rect 5045 1390 5075 1395
rect 5045 1370 5050 1390
rect 5050 1370 5070 1390
rect 5070 1370 5075 1390
rect 5045 1365 5075 1370
rect 5045 1310 5075 1315
rect 5045 1290 5050 1310
rect 5050 1290 5070 1310
rect 5070 1290 5075 1310
rect 5045 1285 5075 1290
rect 5045 1230 5075 1235
rect 5045 1210 5050 1230
rect 5050 1210 5070 1230
rect 5070 1210 5075 1230
rect 5045 1205 5075 1210
rect 5045 1150 5075 1155
rect 5045 1130 5050 1150
rect 5050 1130 5070 1150
rect 5070 1130 5075 1150
rect 5045 1125 5075 1130
rect 5045 1070 5075 1075
rect 5045 1050 5050 1070
rect 5050 1050 5070 1070
rect 5070 1050 5075 1070
rect 5045 1045 5075 1050
rect 5045 990 5075 995
rect 5045 970 5050 990
rect 5050 970 5070 990
rect 5070 970 5075 990
rect 5045 965 5075 970
rect 5045 830 5075 835
rect 5045 810 5050 830
rect 5050 810 5070 830
rect 5070 810 5075 830
rect 5045 805 5075 810
rect 5045 750 5075 755
rect 5045 730 5050 750
rect 5050 730 5070 750
rect 5070 730 5075 750
rect 5045 725 5075 730
rect 5045 670 5075 675
rect 5045 650 5050 670
rect 5050 650 5070 670
rect 5070 650 5075 670
rect 5045 645 5075 650
rect 5045 590 5075 595
rect 5045 570 5050 590
rect 5050 570 5070 590
rect 5070 570 5075 590
rect 5045 565 5075 570
rect 5045 510 5075 515
rect 5045 490 5050 510
rect 5050 490 5070 510
rect 5070 490 5075 510
rect 5045 485 5075 490
rect 5045 270 5075 275
rect 5045 250 5050 270
rect 5050 250 5070 270
rect 5070 250 5075 270
rect 5045 245 5075 250
rect 5045 190 5075 195
rect 5045 170 5050 190
rect 5050 170 5070 190
rect 5070 170 5075 190
rect 5045 165 5075 170
rect 5045 110 5075 115
rect 5045 90 5050 110
rect 5050 90 5070 110
rect 5070 90 5075 110
rect 5045 85 5075 90
rect 5045 30 5075 35
rect 5045 10 5050 30
rect 5050 10 5070 30
rect 5070 10 5075 30
rect 5045 5 5075 10
rect 5205 15710 5235 15715
rect 5205 15690 5210 15710
rect 5210 15690 5230 15710
rect 5230 15690 5235 15710
rect 5205 15685 5235 15690
rect 5205 15630 5235 15635
rect 5205 15610 5210 15630
rect 5210 15610 5230 15630
rect 5230 15610 5235 15630
rect 5205 15605 5235 15610
rect 5205 15550 5235 15555
rect 5205 15530 5210 15550
rect 5210 15530 5230 15550
rect 5230 15530 5235 15550
rect 5205 15525 5235 15530
rect 5205 15470 5235 15475
rect 5205 15450 5210 15470
rect 5210 15450 5230 15470
rect 5230 15450 5235 15470
rect 5205 15445 5235 15450
rect 5205 15390 5235 15395
rect 5205 15370 5210 15390
rect 5210 15370 5230 15390
rect 5230 15370 5235 15390
rect 5205 15365 5235 15370
rect 5205 15310 5235 15315
rect 5205 15290 5210 15310
rect 5210 15290 5230 15310
rect 5230 15290 5235 15310
rect 5205 15285 5235 15290
rect 5205 15230 5235 15235
rect 5205 15210 5210 15230
rect 5210 15210 5230 15230
rect 5230 15210 5235 15230
rect 5205 15205 5235 15210
rect 5205 15150 5235 15155
rect 5205 15130 5210 15150
rect 5210 15130 5230 15150
rect 5230 15130 5235 15150
rect 5205 15125 5235 15130
rect 5205 14990 5235 14995
rect 5205 14970 5210 14990
rect 5210 14970 5230 14990
rect 5230 14970 5235 14990
rect 5205 14965 5235 14970
rect 5205 14910 5235 14915
rect 5205 14890 5210 14910
rect 5210 14890 5230 14910
rect 5230 14890 5235 14910
rect 5205 14885 5235 14890
rect 5205 14830 5235 14835
rect 5205 14810 5210 14830
rect 5210 14810 5230 14830
rect 5230 14810 5235 14830
rect 5205 14805 5235 14810
rect 5205 14750 5235 14755
rect 5205 14730 5210 14750
rect 5210 14730 5230 14750
rect 5230 14730 5235 14750
rect 5205 14725 5235 14730
rect 5205 14670 5235 14675
rect 5205 14650 5210 14670
rect 5210 14650 5230 14670
rect 5230 14650 5235 14670
rect 5205 14645 5235 14650
rect 5205 14590 5235 14595
rect 5205 14570 5210 14590
rect 5210 14570 5230 14590
rect 5230 14570 5235 14590
rect 5205 14565 5235 14570
rect 5205 14510 5235 14515
rect 5205 14490 5210 14510
rect 5210 14490 5230 14510
rect 5230 14490 5235 14510
rect 5205 14485 5235 14490
rect 5205 14430 5235 14435
rect 5205 14410 5210 14430
rect 5210 14410 5230 14430
rect 5230 14410 5235 14430
rect 5205 14405 5235 14410
rect 5205 14030 5235 14035
rect 5205 14010 5210 14030
rect 5210 14010 5230 14030
rect 5230 14010 5235 14030
rect 5205 14005 5235 14010
rect 5205 13950 5235 13955
rect 5205 13930 5210 13950
rect 5210 13930 5230 13950
rect 5230 13930 5235 13950
rect 5205 13925 5235 13930
rect 5205 13870 5235 13875
rect 5205 13850 5210 13870
rect 5210 13850 5230 13870
rect 5230 13850 5235 13870
rect 5205 13845 5235 13850
rect 5205 13790 5235 13795
rect 5205 13770 5210 13790
rect 5210 13770 5230 13790
rect 5230 13770 5235 13790
rect 5205 13765 5235 13770
rect 5205 13710 5235 13715
rect 5205 13690 5210 13710
rect 5210 13690 5230 13710
rect 5230 13690 5235 13710
rect 5205 13685 5235 13690
rect 5205 13630 5235 13635
rect 5205 13610 5210 13630
rect 5210 13610 5230 13630
rect 5230 13610 5235 13630
rect 5205 13605 5235 13610
rect 5205 13550 5235 13555
rect 5205 13530 5210 13550
rect 5210 13530 5230 13550
rect 5230 13530 5235 13550
rect 5205 13525 5235 13530
rect 5205 13470 5235 13475
rect 5205 13450 5210 13470
rect 5210 13450 5230 13470
rect 5230 13450 5235 13470
rect 5205 13445 5235 13450
rect 5205 13070 5235 13075
rect 5205 13050 5210 13070
rect 5210 13050 5230 13070
rect 5230 13050 5235 13070
rect 5205 13045 5235 13050
rect 5205 12990 5235 12995
rect 5205 12970 5210 12990
rect 5210 12970 5230 12990
rect 5230 12970 5235 12990
rect 5205 12965 5235 12970
rect 5205 12910 5235 12915
rect 5205 12890 5210 12910
rect 5210 12890 5230 12910
rect 5230 12890 5235 12910
rect 5205 12885 5235 12890
rect 5205 12830 5235 12835
rect 5205 12810 5210 12830
rect 5210 12810 5230 12830
rect 5230 12810 5235 12830
rect 5205 12805 5235 12810
rect 5205 12750 5235 12755
rect 5205 12730 5210 12750
rect 5210 12730 5230 12750
rect 5230 12730 5235 12750
rect 5205 12725 5235 12730
rect 5205 12670 5235 12675
rect 5205 12650 5210 12670
rect 5210 12650 5230 12670
rect 5230 12650 5235 12670
rect 5205 12645 5235 12650
rect 5205 12590 5235 12595
rect 5205 12570 5210 12590
rect 5210 12570 5230 12590
rect 5230 12570 5235 12590
rect 5205 12565 5235 12570
rect 5205 12510 5235 12515
rect 5205 12490 5210 12510
rect 5210 12490 5230 12510
rect 5230 12490 5235 12510
rect 5205 12485 5235 12490
rect 5205 12350 5235 12355
rect 5205 12330 5210 12350
rect 5210 12330 5230 12350
rect 5230 12330 5235 12350
rect 5205 12325 5235 12330
rect 5205 12270 5235 12275
rect 5205 12250 5210 12270
rect 5210 12250 5230 12270
rect 5230 12250 5235 12270
rect 5205 12245 5235 12250
rect 5205 12190 5235 12195
rect 5205 12170 5210 12190
rect 5210 12170 5230 12190
rect 5230 12170 5235 12190
rect 5205 12165 5235 12170
rect 5205 12110 5235 12115
rect 5205 12090 5210 12110
rect 5210 12090 5230 12110
rect 5230 12090 5235 12110
rect 5205 12085 5235 12090
rect 5205 12030 5235 12035
rect 5205 12010 5210 12030
rect 5210 12010 5230 12030
rect 5230 12010 5235 12030
rect 5205 12005 5235 12010
rect 5205 11950 5235 11955
rect 5205 11930 5210 11950
rect 5210 11930 5230 11950
rect 5230 11930 5235 11950
rect 5205 11925 5235 11930
rect 5205 11870 5235 11875
rect 5205 11850 5210 11870
rect 5210 11850 5230 11870
rect 5230 11850 5235 11870
rect 5205 11845 5235 11850
rect 5205 11790 5235 11795
rect 5205 11770 5210 11790
rect 5210 11770 5230 11790
rect 5230 11770 5235 11790
rect 5205 11765 5235 11770
rect 5205 11710 5235 11715
rect 5205 11690 5210 11710
rect 5210 11690 5230 11710
rect 5230 11690 5235 11710
rect 5205 11685 5235 11690
rect 5205 11630 5235 11635
rect 5205 11610 5210 11630
rect 5210 11610 5230 11630
rect 5230 11610 5235 11630
rect 5205 11605 5235 11610
rect 5205 11550 5235 11555
rect 5205 11530 5210 11550
rect 5210 11530 5230 11550
rect 5230 11530 5235 11550
rect 5205 11525 5235 11530
rect 5205 11470 5235 11475
rect 5205 11450 5210 11470
rect 5210 11450 5230 11470
rect 5230 11450 5235 11470
rect 5205 11445 5235 11450
rect 5205 11390 5235 11395
rect 5205 11370 5210 11390
rect 5210 11370 5230 11390
rect 5230 11370 5235 11390
rect 5205 11365 5235 11370
rect 5205 11310 5235 11315
rect 5205 11290 5210 11310
rect 5210 11290 5230 11310
rect 5230 11290 5235 11310
rect 5205 11285 5235 11290
rect 5205 11230 5235 11235
rect 5205 11210 5210 11230
rect 5210 11210 5230 11230
rect 5230 11210 5235 11230
rect 5205 11205 5235 11210
rect 5205 11150 5235 11155
rect 5205 11130 5210 11150
rect 5210 11130 5230 11150
rect 5230 11130 5235 11150
rect 5205 11125 5235 11130
rect 5205 11070 5235 11075
rect 5205 11050 5210 11070
rect 5210 11050 5230 11070
rect 5230 11050 5235 11070
rect 5205 11045 5235 11050
rect 5205 10910 5235 10915
rect 5205 10890 5210 10910
rect 5210 10890 5230 10910
rect 5230 10890 5235 10910
rect 5205 10885 5235 10890
rect 5205 10830 5235 10835
rect 5205 10810 5210 10830
rect 5210 10810 5230 10830
rect 5230 10810 5235 10830
rect 5205 10805 5235 10810
rect 5205 10750 5235 10755
rect 5205 10730 5210 10750
rect 5210 10730 5230 10750
rect 5230 10730 5235 10750
rect 5205 10725 5235 10730
rect 5205 10670 5235 10675
rect 5205 10650 5210 10670
rect 5210 10650 5230 10670
rect 5230 10650 5235 10670
rect 5205 10645 5235 10650
rect 5205 10590 5235 10595
rect 5205 10570 5210 10590
rect 5210 10570 5230 10590
rect 5230 10570 5235 10590
rect 5205 10565 5235 10570
rect 5205 10510 5235 10515
rect 5205 10490 5210 10510
rect 5210 10490 5230 10510
rect 5230 10490 5235 10510
rect 5205 10485 5235 10490
rect 5205 10430 5235 10435
rect 5205 10410 5210 10430
rect 5210 10410 5230 10430
rect 5230 10410 5235 10430
rect 5205 10405 5235 10410
rect 5205 10350 5235 10355
rect 5205 10330 5210 10350
rect 5210 10330 5230 10350
rect 5230 10330 5235 10350
rect 5205 10325 5235 10330
rect 5205 9950 5235 9955
rect 5205 9930 5210 9950
rect 5210 9930 5230 9950
rect 5230 9930 5235 9950
rect 5205 9925 5235 9930
rect 5205 9870 5235 9875
rect 5205 9850 5210 9870
rect 5210 9850 5230 9870
rect 5230 9850 5235 9870
rect 5205 9845 5235 9850
rect 5205 9790 5235 9795
rect 5205 9770 5210 9790
rect 5210 9770 5230 9790
rect 5230 9770 5235 9790
rect 5205 9765 5235 9770
rect 5205 9710 5235 9715
rect 5205 9690 5210 9710
rect 5210 9690 5230 9710
rect 5230 9690 5235 9710
rect 5205 9685 5235 9690
rect 5205 9630 5235 9635
rect 5205 9610 5210 9630
rect 5210 9610 5230 9630
rect 5230 9610 5235 9630
rect 5205 9605 5235 9610
rect 5205 9550 5235 9555
rect 5205 9530 5210 9550
rect 5210 9530 5230 9550
rect 5230 9530 5235 9550
rect 5205 9525 5235 9530
rect 5205 9470 5235 9475
rect 5205 9450 5210 9470
rect 5210 9450 5230 9470
rect 5230 9450 5235 9470
rect 5205 9445 5235 9450
rect 5205 9390 5235 9395
rect 5205 9370 5210 9390
rect 5210 9370 5230 9390
rect 5230 9370 5235 9390
rect 5205 9365 5235 9370
rect 5205 8990 5235 8995
rect 5205 8970 5210 8990
rect 5210 8970 5230 8990
rect 5230 8970 5235 8990
rect 5205 8965 5235 8970
rect 5205 8910 5235 8915
rect 5205 8890 5210 8910
rect 5210 8890 5230 8910
rect 5230 8890 5235 8910
rect 5205 8885 5235 8890
rect 5205 8830 5235 8835
rect 5205 8810 5210 8830
rect 5210 8810 5230 8830
rect 5230 8810 5235 8830
rect 5205 8805 5235 8810
rect 5205 8750 5235 8755
rect 5205 8730 5210 8750
rect 5210 8730 5230 8750
rect 5230 8730 5235 8750
rect 5205 8725 5235 8730
rect 5205 8670 5235 8675
rect 5205 8650 5210 8670
rect 5210 8650 5230 8670
rect 5230 8650 5235 8670
rect 5205 8645 5235 8650
rect 5205 8590 5235 8595
rect 5205 8570 5210 8590
rect 5210 8570 5230 8590
rect 5230 8570 5235 8590
rect 5205 8565 5235 8570
rect 5205 8510 5235 8515
rect 5205 8490 5210 8510
rect 5210 8490 5230 8510
rect 5230 8490 5235 8510
rect 5205 8485 5235 8490
rect 5205 8430 5235 8435
rect 5205 8410 5210 8430
rect 5210 8410 5230 8430
rect 5230 8410 5235 8430
rect 5205 8405 5235 8410
rect 5205 8270 5235 8275
rect 5205 8250 5210 8270
rect 5210 8250 5230 8270
rect 5230 8250 5235 8270
rect 5205 8245 5235 8250
rect 5205 8190 5235 8195
rect 5205 8170 5210 8190
rect 5210 8170 5230 8190
rect 5230 8170 5235 8190
rect 5205 8165 5235 8170
rect 5205 8110 5235 8115
rect 5205 8090 5210 8110
rect 5210 8090 5230 8110
rect 5230 8090 5235 8110
rect 5205 8085 5235 8090
rect 5205 8030 5235 8035
rect 5205 8010 5210 8030
rect 5210 8010 5230 8030
rect 5230 8010 5235 8030
rect 5205 8005 5235 8010
rect 5205 7950 5235 7955
rect 5205 7930 5210 7950
rect 5210 7930 5230 7950
rect 5230 7930 5235 7950
rect 5205 7925 5235 7930
rect 5205 7870 5235 7875
rect 5205 7850 5210 7870
rect 5210 7850 5230 7870
rect 5230 7850 5235 7870
rect 5205 7845 5235 7850
rect 5205 7790 5235 7795
rect 5205 7770 5210 7790
rect 5210 7770 5230 7790
rect 5230 7770 5235 7790
rect 5205 7765 5235 7770
rect 5205 7710 5235 7715
rect 5205 7690 5210 7710
rect 5210 7690 5230 7710
rect 5230 7690 5235 7710
rect 5205 7685 5235 7690
rect 5205 7630 5235 7635
rect 5205 7610 5210 7630
rect 5210 7610 5230 7630
rect 5230 7610 5235 7630
rect 5205 7605 5235 7610
rect 5205 7550 5235 7555
rect 5205 7530 5210 7550
rect 5210 7530 5230 7550
rect 5230 7530 5235 7550
rect 5205 7525 5235 7530
rect 5205 7470 5235 7475
rect 5205 7450 5210 7470
rect 5210 7450 5230 7470
rect 5230 7450 5235 7470
rect 5205 7445 5235 7450
rect 5205 7390 5235 7395
rect 5205 7370 5210 7390
rect 5210 7370 5230 7390
rect 5230 7370 5235 7390
rect 5205 7365 5235 7370
rect 5205 7310 5235 7315
rect 5205 7290 5210 7310
rect 5210 7290 5230 7310
rect 5230 7290 5235 7310
rect 5205 7285 5235 7290
rect 5205 7230 5235 7235
rect 5205 7210 5210 7230
rect 5210 7210 5230 7230
rect 5230 7210 5235 7230
rect 5205 7205 5235 7210
rect 5205 7150 5235 7155
rect 5205 7130 5210 7150
rect 5210 7130 5230 7150
rect 5230 7130 5235 7150
rect 5205 7125 5235 7130
rect 5205 7070 5235 7075
rect 5205 7050 5210 7070
rect 5210 7050 5230 7070
rect 5230 7050 5235 7070
rect 5205 7045 5235 7050
rect 5205 6990 5235 6995
rect 5205 6970 5210 6990
rect 5210 6970 5230 6990
rect 5230 6970 5235 6990
rect 5205 6965 5235 6970
rect 5205 6830 5235 6835
rect 5205 6810 5210 6830
rect 5210 6810 5230 6830
rect 5230 6810 5235 6830
rect 5205 6805 5235 6810
rect 5205 6750 5235 6755
rect 5205 6730 5210 6750
rect 5210 6730 5230 6750
rect 5230 6730 5235 6750
rect 5205 6725 5235 6730
rect 5205 6670 5235 6675
rect 5205 6650 5210 6670
rect 5210 6650 5230 6670
rect 5230 6650 5235 6670
rect 5205 6645 5235 6650
rect 5205 6590 5235 6595
rect 5205 6570 5210 6590
rect 5210 6570 5230 6590
rect 5230 6570 5235 6590
rect 5205 6565 5235 6570
rect 5205 6510 5235 6515
rect 5205 6490 5210 6510
rect 5210 6490 5230 6510
rect 5230 6490 5235 6510
rect 5205 6485 5235 6490
rect 5205 6430 5235 6435
rect 5205 6410 5210 6430
rect 5210 6410 5230 6430
rect 5230 6410 5235 6430
rect 5205 6405 5235 6410
rect 5205 6350 5235 6355
rect 5205 6330 5210 6350
rect 5210 6330 5230 6350
rect 5230 6330 5235 6350
rect 5205 6325 5235 6330
rect 5205 6270 5235 6275
rect 5205 6250 5210 6270
rect 5210 6250 5230 6270
rect 5230 6250 5235 6270
rect 5205 6245 5235 6250
rect 5205 5870 5235 5875
rect 5205 5850 5210 5870
rect 5210 5850 5230 5870
rect 5230 5850 5235 5870
rect 5205 5845 5235 5850
rect 5205 5790 5235 5795
rect 5205 5770 5210 5790
rect 5210 5770 5230 5790
rect 5230 5770 5235 5790
rect 5205 5765 5235 5770
rect 5205 5710 5235 5715
rect 5205 5690 5210 5710
rect 5210 5690 5230 5710
rect 5230 5690 5235 5710
rect 5205 5685 5235 5690
rect 5205 5630 5235 5635
rect 5205 5610 5210 5630
rect 5210 5610 5230 5630
rect 5230 5610 5235 5630
rect 5205 5605 5235 5610
rect 5205 5550 5235 5555
rect 5205 5530 5210 5550
rect 5210 5530 5230 5550
rect 5230 5530 5235 5550
rect 5205 5525 5235 5530
rect 5205 5470 5235 5475
rect 5205 5450 5210 5470
rect 5210 5450 5230 5470
rect 5230 5450 5235 5470
rect 5205 5445 5235 5450
rect 5205 5390 5235 5395
rect 5205 5370 5210 5390
rect 5210 5370 5230 5390
rect 5230 5370 5235 5390
rect 5205 5365 5235 5370
rect 5205 5310 5235 5315
rect 5205 5290 5210 5310
rect 5210 5290 5230 5310
rect 5230 5290 5235 5310
rect 5205 5285 5235 5290
rect 5205 5230 5235 5235
rect 5205 5210 5210 5230
rect 5210 5210 5230 5230
rect 5230 5210 5235 5230
rect 5205 5205 5235 5210
rect 5205 5150 5235 5155
rect 5205 5130 5210 5150
rect 5210 5130 5230 5150
rect 5230 5130 5235 5150
rect 5205 5125 5235 5130
rect 5205 5070 5235 5075
rect 5205 5050 5210 5070
rect 5210 5050 5230 5070
rect 5230 5050 5235 5070
rect 5205 5045 5235 5050
rect 5205 4990 5235 4995
rect 5205 4970 5210 4990
rect 5210 4970 5230 4990
rect 5230 4970 5235 4990
rect 5205 4965 5235 4970
rect 5205 4910 5235 4915
rect 5205 4890 5210 4910
rect 5210 4890 5230 4910
rect 5230 4890 5235 4910
rect 5205 4885 5235 4890
rect 5205 4750 5235 4755
rect 5205 4730 5210 4750
rect 5210 4730 5230 4750
rect 5230 4730 5235 4750
rect 5205 4725 5235 4730
rect 5205 4670 5235 4675
rect 5205 4650 5210 4670
rect 5210 4650 5230 4670
rect 5230 4650 5235 4670
rect 5205 4645 5235 4650
rect 5205 4510 5235 4515
rect 5205 4490 5210 4510
rect 5210 4490 5230 4510
rect 5230 4490 5235 4510
rect 5205 4485 5235 4490
rect 5205 4430 5235 4435
rect 5205 4410 5210 4430
rect 5210 4410 5230 4430
rect 5230 4410 5235 4430
rect 5205 4405 5235 4410
rect 5205 4350 5235 4355
rect 5205 4330 5210 4350
rect 5210 4330 5230 4350
rect 5230 4330 5235 4350
rect 5205 4325 5235 4330
rect 5205 4270 5235 4275
rect 5205 4250 5210 4270
rect 5210 4250 5230 4270
rect 5230 4250 5235 4270
rect 5205 4245 5235 4250
rect 5205 4190 5235 4195
rect 5205 4170 5210 4190
rect 5210 4170 5230 4190
rect 5230 4170 5235 4190
rect 5205 4165 5235 4170
rect 5205 4110 5235 4115
rect 5205 4090 5210 4110
rect 5210 4090 5230 4110
rect 5230 4090 5235 4110
rect 5205 4085 5235 4090
rect 5205 4030 5235 4035
rect 5205 4010 5210 4030
rect 5210 4010 5230 4030
rect 5230 4010 5235 4030
rect 5205 4005 5235 4010
rect 5205 3950 5235 3955
rect 5205 3930 5210 3950
rect 5210 3930 5230 3950
rect 5230 3930 5235 3950
rect 5205 3925 5235 3930
rect 5205 3870 5235 3875
rect 5205 3850 5210 3870
rect 5210 3850 5230 3870
rect 5230 3850 5235 3870
rect 5205 3845 5235 3850
rect 5205 3710 5235 3715
rect 5205 3690 5210 3710
rect 5210 3690 5230 3710
rect 5230 3690 5235 3710
rect 5205 3685 5235 3690
rect 5205 3630 5235 3635
rect 5205 3610 5210 3630
rect 5210 3610 5230 3630
rect 5230 3610 5235 3630
rect 5205 3605 5235 3610
rect 5205 3470 5235 3475
rect 5205 3450 5210 3470
rect 5210 3450 5230 3470
rect 5230 3450 5235 3470
rect 5205 3445 5235 3450
rect 5205 3390 5235 3395
rect 5205 3370 5210 3390
rect 5210 3370 5230 3390
rect 5230 3370 5235 3390
rect 5205 3365 5235 3370
rect 5205 3230 5235 3235
rect 5205 3210 5210 3230
rect 5210 3210 5230 3230
rect 5230 3210 5235 3230
rect 5205 3205 5235 3210
rect 5205 3150 5235 3155
rect 5205 3130 5210 3150
rect 5210 3130 5230 3150
rect 5230 3130 5235 3150
rect 5205 3125 5235 3130
rect 5205 3070 5235 3075
rect 5205 3050 5210 3070
rect 5210 3050 5230 3070
rect 5230 3050 5235 3070
rect 5205 3045 5235 3050
rect 5205 2990 5235 2995
rect 5205 2970 5210 2990
rect 5210 2970 5230 2990
rect 5230 2970 5235 2990
rect 5205 2965 5235 2970
rect 5205 2910 5235 2915
rect 5205 2890 5210 2910
rect 5210 2890 5230 2910
rect 5230 2890 5235 2910
rect 5205 2885 5235 2890
rect 5205 2830 5235 2835
rect 5205 2810 5210 2830
rect 5210 2810 5230 2830
rect 5230 2810 5235 2830
rect 5205 2805 5235 2810
rect 5205 2750 5235 2755
rect 5205 2730 5210 2750
rect 5210 2730 5230 2750
rect 5230 2730 5235 2750
rect 5205 2725 5235 2730
rect 5205 2670 5235 2675
rect 5205 2650 5210 2670
rect 5210 2650 5230 2670
rect 5230 2650 5235 2670
rect 5205 2645 5235 2650
rect 5205 2590 5235 2595
rect 5205 2570 5210 2590
rect 5210 2570 5230 2590
rect 5230 2570 5235 2590
rect 5205 2565 5235 2570
rect 5205 2510 5235 2515
rect 5205 2490 5210 2510
rect 5210 2490 5230 2510
rect 5230 2490 5235 2510
rect 5205 2485 5235 2490
rect 5205 2430 5235 2435
rect 5205 2410 5210 2430
rect 5210 2410 5230 2430
rect 5230 2410 5235 2430
rect 5205 2405 5235 2410
rect 5205 2350 5235 2355
rect 5205 2330 5210 2350
rect 5210 2330 5230 2350
rect 5230 2330 5235 2350
rect 5205 2325 5235 2330
rect 5205 2270 5235 2275
rect 5205 2250 5210 2270
rect 5210 2250 5230 2270
rect 5230 2250 5235 2270
rect 5205 2245 5235 2250
rect 5205 2190 5235 2195
rect 5205 2170 5210 2190
rect 5210 2170 5230 2190
rect 5230 2170 5235 2190
rect 5205 2165 5235 2170
rect 5205 2110 5235 2115
rect 5205 2090 5210 2110
rect 5210 2090 5230 2110
rect 5230 2090 5235 2110
rect 5205 2085 5235 2090
rect 5205 2030 5235 2035
rect 5205 2010 5210 2030
rect 5210 2010 5230 2030
rect 5230 2010 5235 2030
rect 5205 2005 5235 2010
rect 5205 1950 5235 1955
rect 5205 1930 5210 1950
rect 5210 1930 5230 1950
rect 5230 1930 5235 1950
rect 5205 1925 5235 1930
rect 5205 1710 5235 1715
rect 5205 1690 5210 1710
rect 5210 1690 5230 1710
rect 5230 1690 5235 1710
rect 5205 1685 5235 1690
rect 5205 1630 5235 1635
rect 5205 1610 5210 1630
rect 5210 1610 5230 1630
rect 5230 1610 5235 1630
rect 5205 1605 5235 1610
rect 5205 1550 5235 1555
rect 5205 1530 5210 1550
rect 5210 1530 5230 1550
rect 5230 1530 5235 1550
rect 5205 1525 5235 1530
rect 5205 1470 5235 1475
rect 5205 1450 5210 1470
rect 5210 1450 5230 1470
rect 5230 1450 5235 1470
rect 5205 1445 5235 1450
rect 5205 1390 5235 1395
rect 5205 1370 5210 1390
rect 5210 1370 5230 1390
rect 5230 1370 5235 1390
rect 5205 1365 5235 1370
rect 5205 1310 5235 1315
rect 5205 1290 5210 1310
rect 5210 1290 5230 1310
rect 5230 1290 5235 1310
rect 5205 1285 5235 1290
rect 5205 1230 5235 1235
rect 5205 1210 5210 1230
rect 5210 1210 5230 1230
rect 5230 1210 5235 1230
rect 5205 1205 5235 1210
rect 5205 1150 5235 1155
rect 5205 1130 5210 1150
rect 5210 1130 5230 1150
rect 5230 1130 5235 1150
rect 5205 1125 5235 1130
rect 5205 1070 5235 1075
rect 5205 1050 5210 1070
rect 5210 1050 5230 1070
rect 5230 1050 5235 1070
rect 5205 1045 5235 1050
rect 5205 990 5235 995
rect 5205 970 5210 990
rect 5210 970 5230 990
rect 5230 970 5235 990
rect 5205 965 5235 970
rect 5205 830 5235 835
rect 5205 810 5210 830
rect 5210 810 5230 830
rect 5230 810 5235 830
rect 5205 805 5235 810
rect 5205 750 5235 755
rect 5205 730 5210 750
rect 5210 730 5230 750
rect 5230 730 5235 750
rect 5205 725 5235 730
rect 5205 670 5235 675
rect 5205 650 5210 670
rect 5210 650 5230 670
rect 5230 650 5235 670
rect 5205 645 5235 650
rect 5205 590 5235 595
rect 5205 570 5210 590
rect 5210 570 5230 590
rect 5230 570 5235 590
rect 5205 565 5235 570
rect 5205 510 5235 515
rect 5205 490 5210 510
rect 5210 490 5230 510
rect 5230 490 5235 510
rect 5205 485 5235 490
rect 5205 270 5235 275
rect 5205 250 5210 270
rect 5210 250 5230 270
rect 5230 250 5235 270
rect 5205 245 5235 250
rect 5205 190 5235 195
rect 5205 170 5210 190
rect 5210 170 5230 190
rect 5230 170 5235 190
rect 5205 165 5235 170
rect 5205 110 5235 115
rect 5205 90 5210 110
rect 5210 90 5230 110
rect 5230 90 5235 110
rect 5205 85 5235 90
rect 5205 30 5235 35
rect 5205 10 5210 30
rect 5210 10 5230 30
rect 5230 10 5235 30
rect 5205 5 5235 10
rect 5365 15710 5395 15715
rect 5365 15690 5370 15710
rect 5370 15690 5390 15710
rect 5390 15690 5395 15710
rect 5365 15685 5395 15690
rect 5365 15630 5395 15635
rect 5365 15610 5370 15630
rect 5370 15610 5390 15630
rect 5390 15610 5395 15630
rect 5365 15605 5395 15610
rect 5365 15550 5395 15555
rect 5365 15530 5370 15550
rect 5370 15530 5390 15550
rect 5390 15530 5395 15550
rect 5365 15525 5395 15530
rect 5365 15470 5395 15475
rect 5365 15450 5370 15470
rect 5370 15450 5390 15470
rect 5390 15450 5395 15470
rect 5365 15445 5395 15450
rect 5365 15390 5395 15395
rect 5365 15370 5370 15390
rect 5370 15370 5390 15390
rect 5390 15370 5395 15390
rect 5365 15365 5395 15370
rect 5365 15310 5395 15315
rect 5365 15290 5370 15310
rect 5370 15290 5390 15310
rect 5390 15290 5395 15310
rect 5365 15285 5395 15290
rect 5365 15230 5395 15235
rect 5365 15210 5370 15230
rect 5370 15210 5390 15230
rect 5390 15210 5395 15230
rect 5365 15205 5395 15210
rect 5365 15150 5395 15155
rect 5365 15130 5370 15150
rect 5370 15130 5390 15150
rect 5390 15130 5395 15150
rect 5365 15125 5395 15130
rect 5365 14990 5395 14995
rect 5365 14970 5370 14990
rect 5370 14970 5390 14990
rect 5390 14970 5395 14990
rect 5365 14965 5395 14970
rect 5365 14910 5395 14915
rect 5365 14890 5370 14910
rect 5370 14890 5390 14910
rect 5390 14890 5395 14910
rect 5365 14885 5395 14890
rect 5365 14830 5395 14835
rect 5365 14810 5370 14830
rect 5370 14810 5390 14830
rect 5390 14810 5395 14830
rect 5365 14805 5395 14810
rect 5365 14750 5395 14755
rect 5365 14730 5370 14750
rect 5370 14730 5390 14750
rect 5390 14730 5395 14750
rect 5365 14725 5395 14730
rect 5365 14670 5395 14675
rect 5365 14650 5370 14670
rect 5370 14650 5390 14670
rect 5390 14650 5395 14670
rect 5365 14645 5395 14650
rect 5365 14590 5395 14595
rect 5365 14570 5370 14590
rect 5370 14570 5390 14590
rect 5390 14570 5395 14590
rect 5365 14565 5395 14570
rect 5365 14510 5395 14515
rect 5365 14490 5370 14510
rect 5370 14490 5390 14510
rect 5390 14490 5395 14510
rect 5365 14485 5395 14490
rect 5365 14430 5395 14435
rect 5365 14410 5370 14430
rect 5370 14410 5390 14430
rect 5390 14410 5395 14430
rect 5365 14405 5395 14410
rect 5365 14030 5395 14035
rect 5365 14010 5370 14030
rect 5370 14010 5390 14030
rect 5390 14010 5395 14030
rect 5365 14005 5395 14010
rect 5365 13950 5395 13955
rect 5365 13930 5370 13950
rect 5370 13930 5390 13950
rect 5390 13930 5395 13950
rect 5365 13925 5395 13930
rect 5365 13870 5395 13875
rect 5365 13850 5370 13870
rect 5370 13850 5390 13870
rect 5390 13850 5395 13870
rect 5365 13845 5395 13850
rect 5365 13790 5395 13795
rect 5365 13770 5370 13790
rect 5370 13770 5390 13790
rect 5390 13770 5395 13790
rect 5365 13765 5395 13770
rect 5365 13710 5395 13715
rect 5365 13690 5370 13710
rect 5370 13690 5390 13710
rect 5390 13690 5395 13710
rect 5365 13685 5395 13690
rect 5365 13630 5395 13635
rect 5365 13610 5370 13630
rect 5370 13610 5390 13630
rect 5390 13610 5395 13630
rect 5365 13605 5395 13610
rect 5365 13550 5395 13555
rect 5365 13530 5370 13550
rect 5370 13530 5390 13550
rect 5390 13530 5395 13550
rect 5365 13525 5395 13530
rect 5365 13470 5395 13475
rect 5365 13450 5370 13470
rect 5370 13450 5390 13470
rect 5390 13450 5395 13470
rect 5365 13445 5395 13450
rect 5365 13070 5395 13075
rect 5365 13050 5370 13070
rect 5370 13050 5390 13070
rect 5390 13050 5395 13070
rect 5365 13045 5395 13050
rect 5365 12990 5395 12995
rect 5365 12970 5370 12990
rect 5370 12970 5390 12990
rect 5390 12970 5395 12990
rect 5365 12965 5395 12970
rect 5365 12910 5395 12915
rect 5365 12890 5370 12910
rect 5370 12890 5390 12910
rect 5390 12890 5395 12910
rect 5365 12885 5395 12890
rect 5365 12830 5395 12835
rect 5365 12810 5370 12830
rect 5370 12810 5390 12830
rect 5390 12810 5395 12830
rect 5365 12805 5395 12810
rect 5365 12750 5395 12755
rect 5365 12730 5370 12750
rect 5370 12730 5390 12750
rect 5390 12730 5395 12750
rect 5365 12725 5395 12730
rect 5365 12670 5395 12675
rect 5365 12650 5370 12670
rect 5370 12650 5390 12670
rect 5390 12650 5395 12670
rect 5365 12645 5395 12650
rect 5365 12590 5395 12595
rect 5365 12570 5370 12590
rect 5370 12570 5390 12590
rect 5390 12570 5395 12590
rect 5365 12565 5395 12570
rect 5365 12510 5395 12515
rect 5365 12490 5370 12510
rect 5370 12490 5390 12510
rect 5390 12490 5395 12510
rect 5365 12485 5395 12490
rect 5365 12350 5395 12355
rect 5365 12330 5370 12350
rect 5370 12330 5390 12350
rect 5390 12330 5395 12350
rect 5365 12325 5395 12330
rect 5365 12270 5395 12275
rect 5365 12250 5370 12270
rect 5370 12250 5390 12270
rect 5390 12250 5395 12270
rect 5365 12245 5395 12250
rect 5365 12190 5395 12195
rect 5365 12170 5370 12190
rect 5370 12170 5390 12190
rect 5390 12170 5395 12190
rect 5365 12165 5395 12170
rect 5365 12110 5395 12115
rect 5365 12090 5370 12110
rect 5370 12090 5390 12110
rect 5390 12090 5395 12110
rect 5365 12085 5395 12090
rect 5365 12030 5395 12035
rect 5365 12010 5370 12030
rect 5370 12010 5390 12030
rect 5390 12010 5395 12030
rect 5365 12005 5395 12010
rect 5365 11950 5395 11955
rect 5365 11930 5370 11950
rect 5370 11930 5390 11950
rect 5390 11930 5395 11950
rect 5365 11925 5395 11930
rect 5365 11870 5395 11875
rect 5365 11850 5370 11870
rect 5370 11850 5390 11870
rect 5390 11850 5395 11870
rect 5365 11845 5395 11850
rect 5365 11790 5395 11795
rect 5365 11770 5370 11790
rect 5370 11770 5390 11790
rect 5390 11770 5395 11790
rect 5365 11765 5395 11770
rect 5365 11710 5395 11715
rect 5365 11690 5370 11710
rect 5370 11690 5390 11710
rect 5390 11690 5395 11710
rect 5365 11685 5395 11690
rect 5365 11630 5395 11635
rect 5365 11610 5370 11630
rect 5370 11610 5390 11630
rect 5390 11610 5395 11630
rect 5365 11605 5395 11610
rect 5365 11550 5395 11555
rect 5365 11530 5370 11550
rect 5370 11530 5390 11550
rect 5390 11530 5395 11550
rect 5365 11525 5395 11530
rect 5365 11470 5395 11475
rect 5365 11450 5370 11470
rect 5370 11450 5390 11470
rect 5390 11450 5395 11470
rect 5365 11445 5395 11450
rect 5365 11390 5395 11395
rect 5365 11370 5370 11390
rect 5370 11370 5390 11390
rect 5390 11370 5395 11390
rect 5365 11365 5395 11370
rect 5365 11310 5395 11315
rect 5365 11290 5370 11310
rect 5370 11290 5390 11310
rect 5390 11290 5395 11310
rect 5365 11285 5395 11290
rect 5365 11230 5395 11235
rect 5365 11210 5370 11230
rect 5370 11210 5390 11230
rect 5390 11210 5395 11230
rect 5365 11205 5395 11210
rect 5365 11150 5395 11155
rect 5365 11130 5370 11150
rect 5370 11130 5390 11150
rect 5390 11130 5395 11150
rect 5365 11125 5395 11130
rect 5365 11070 5395 11075
rect 5365 11050 5370 11070
rect 5370 11050 5390 11070
rect 5390 11050 5395 11070
rect 5365 11045 5395 11050
rect 5365 10910 5395 10915
rect 5365 10890 5370 10910
rect 5370 10890 5390 10910
rect 5390 10890 5395 10910
rect 5365 10885 5395 10890
rect 5365 10830 5395 10835
rect 5365 10810 5370 10830
rect 5370 10810 5390 10830
rect 5390 10810 5395 10830
rect 5365 10805 5395 10810
rect 5365 10750 5395 10755
rect 5365 10730 5370 10750
rect 5370 10730 5390 10750
rect 5390 10730 5395 10750
rect 5365 10725 5395 10730
rect 5365 10670 5395 10675
rect 5365 10650 5370 10670
rect 5370 10650 5390 10670
rect 5390 10650 5395 10670
rect 5365 10645 5395 10650
rect 5365 10590 5395 10595
rect 5365 10570 5370 10590
rect 5370 10570 5390 10590
rect 5390 10570 5395 10590
rect 5365 10565 5395 10570
rect 5365 10510 5395 10515
rect 5365 10490 5370 10510
rect 5370 10490 5390 10510
rect 5390 10490 5395 10510
rect 5365 10485 5395 10490
rect 5365 10430 5395 10435
rect 5365 10410 5370 10430
rect 5370 10410 5390 10430
rect 5390 10410 5395 10430
rect 5365 10405 5395 10410
rect 5365 10350 5395 10355
rect 5365 10330 5370 10350
rect 5370 10330 5390 10350
rect 5390 10330 5395 10350
rect 5365 10325 5395 10330
rect 5365 9950 5395 9955
rect 5365 9930 5370 9950
rect 5370 9930 5390 9950
rect 5390 9930 5395 9950
rect 5365 9925 5395 9930
rect 5365 9870 5395 9875
rect 5365 9850 5370 9870
rect 5370 9850 5390 9870
rect 5390 9850 5395 9870
rect 5365 9845 5395 9850
rect 5365 9790 5395 9795
rect 5365 9770 5370 9790
rect 5370 9770 5390 9790
rect 5390 9770 5395 9790
rect 5365 9765 5395 9770
rect 5365 9710 5395 9715
rect 5365 9690 5370 9710
rect 5370 9690 5390 9710
rect 5390 9690 5395 9710
rect 5365 9685 5395 9690
rect 5365 9630 5395 9635
rect 5365 9610 5370 9630
rect 5370 9610 5390 9630
rect 5390 9610 5395 9630
rect 5365 9605 5395 9610
rect 5365 9550 5395 9555
rect 5365 9530 5370 9550
rect 5370 9530 5390 9550
rect 5390 9530 5395 9550
rect 5365 9525 5395 9530
rect 5365 9470 5395 9475
rect 5365 9450 5370 9470
rect 5370 9450 5390 9470
rect 5390 9450 5395 9470
rect 5365 9445 5395 9450
rect 5365 9390 5395 9395
rect 5365 9370 5370 9390
rect 5370 9370 5390 9390
rect 5390 9370 5395 9390
rect 5365 9365 5395 9370
rect 5365 8990 5395 8995
rect 5365 8970 5370 8990
rect 5370 8970 5390 8990
rect 5390 8970 5395 8990
rect 5365 8965 5395 8970
rect 5365 8910 5395 8915
rect 5365 8890 5370 8910
rect 5370 8890 5390 8910
rect 5390 8890 5395 8910
rect 5365 8885 5395 8890
rect 5365 8830 5395 8835
rect 5365 8810 5370 8830
rect 5370 8810 5390 8830
rect 5390 8810 5395 8830
rect 5365 8805 5395 8810
rect 5365 8750 5395 8755
rect 5365 8730 5370 8750
rect 5370 8730 5390 8750
rect 5390 8730 5395 8750
rect 5365 8725 5395 8730
rect 5365 8670 5395 8675
rect 5365 8650 5370 8670
rect 5370 8650 5390 8670
rect 5390 8650 5395 8670
rect 5365 8645 5395 8650
rect 5365 8590 5395 8595
rect 5365 8570 5370 8590
rect 5370 8570 5390 8590
rect 5390 8570 5395 8590
rect 5365 8565 5395 8570
rect 5365 8510 5395 8515
rect 5365 8490 5370 8510
rect 5370 8490 5390 8510
rect 5390 8490 5395 8510
rect 5365 8485 5395 8490
rect 5365 8430 5395 8435
rect 5365 8410 5370 8430
rect 5370 8410 5390 8430
rect 5390 8410 5395 8430
rect 5365 8405 5395 8410
rect 5365 8270 5395 8275
rect 5365 8250 5370 8270
rect 5370 8250 5390 8270
rect 5390 8250 5395 8270
rect 5365 8245 5395 8250
rect 5365 8190 5395 8195
rect 5365 8170 5370 8190
rect 5370 8170 5390 8190
rect 5390 8170 5395 8190
rect 5365 8165 5395 8170
rect 5365 8110 5395 8115
rect 5365 8090 5370 8110
rect 5370 8090 5390 8110
rect 5390 8090 5395 8110
rect 5365 8085 5395 8090
rect 5365 8030 5395 8035
rect 5365 8010 5370 8030
rect 5370 8010 5390 8030
rect 5390 8010 5395 8030
rect 5365 8005 5395 8010
rect 5365 7950 5395 7955
rect 5365 7930 5370 7950
rect 5370 7930 5390 7950
rect 5390 7930 5395 7950
rect 5365 7925 5395 7930
rect 5365 7870 5395 7875
rect 5365 7850 5370 7870
rect 5370 7850 5390 7870
rect 5390 7850 5395 7870
rect 5365 7845 5395 7850
rect 5365 7790 5395 7795
rect 5365 7770 5370 7790
rect 5370 7770 5390 7790
rect 5390 7770 5395 7790
rect 5365 7765 5395 7770
rect 5365 7710 5395 7715
rect 5365 7690 5370 7710
rect 5370 7690 5390 7710
rect 5390 7690 5395 7710
rect 5365 7685 5395 7690
rect 5365 7630 5395 7635
rect 5365 7610 5370 7630
rect 5370 7610 5390 7630
rect 5390 7610 5395 7630
rect 5365 7605 5395 7610
rect 5365 7550 5395 7555
rect 5365 7530 5370 7550
rect 5370 7530 5390 7550
rect 5390 7530 5395 7550
rect 5365 7525 5395 7530
rect 5365 7470 5395 7475
rect 5365 7450 5370 7470
rect 5370 7450 5390 7470
rect 5390 7450 5395 7470
rect 5365 7445 5395 7450
rect 5365 7390 5395 7395
rect 5365 7370 5370 7390
rect 5370 7370 5390 7390
rect 5390 7370 5395 7390
rect 5365 7365 5395 7370
rect 5365 7310 5395 7315
rect 5365 7290 5370 7310
rect 5370 7290 5390 7310
rect 5390 7290 5395 7310
rect 5365 7285 5395 7290
rect 5365 7230 5395 7235
rect 5365 7210 5370 7230
rect 5370 7210 5390 7230
rect 5390 7210 5395 7230
rect 5365 7205 5395 7210
rect 5365 7150 5395 7155
rect 5365 7130 5370 7150
rect 5370 7130 5390 7150
rect 5390 7130 5395 7150
rect 5365 7125 5395 7130
rect 5365 7070 5395 7075
rect 5365 7050 5370 7070
rect 5370 7050 5390 7070
rect 5390 7050 5395 7070
rect 5365 7045 5395 7050
rect 5365 6990 5395 6995
rect 5365 6970 5370 6990
rect 5370 6970 5390 6990
rect 5390 6970 5395 6990
rect 5365 6965 5395 6970
rect 5365 6830 5395 6835
rect 5365 6810 5370 6830
rect 5370 6810 5390 6830
rect 5390 6810 5395 6830
rect 5365 6805 5395 6810
rect 5365 6750 5395 6755
rect 5365 6730 5370 6750
rect 5370 6730 5390 6750
rect 5390 6730 5395 6750
rect 5365 6725 5395 6730
rect 5365 6670 5395 6675
rect 5365 6650 5370 6670
rect 5370 6650 5390 6670
rect 5390 6650 5395 6670
rect 5365 6645 5395 6650
rect 5365 6590 5395 6595
rect 5365 6570 5370 6590
rect 5370 6570 5390 6590
rect 5390 6570 5395 6590
rect 5365 6565 5395 6570
rect 5365 6510 5395 6515
rect 5365 6490 5370 6510
rect 5370 6490 5390 6510
rect 5390 6490 5395 6510
rect 5365 6485 5395 6490
rect 5365 6430 5395 6435
rect 5365 6410 5370 6430
rect 5370 6410 5390 6430
rect 5390 6410 5395 6430
rect 5365 6405 5395 6410
rect 5365 6350 5395 6355
rect 5365 6330 5370 6350
rect 5370 6330 5390 6350
rect 5390 6330 5395 6350
rect 5365 6325 5395 6330
rect 5365 6270 5395 6275
rect 5365 6250 5370 6270
rect 5370 6250 5390 6270
rect 5390 6250 5395 6270
rect 5365 6245 5395 6250
rect 5365 5870 5395 5875
rect 5365 5850 5370 5870
rect 5370 5850 5390 5870
rect 5390 5850 5395 5870
rect 5365 5845 5395 5850
rect 5365 5790 5395 5795
rect 5365 5770 5370 5790
rect 5370 5770 5390 5790
rect 5390 5770 5395 5790
rect 5365 5765 5395 5770
rect 5365 5710 5395 5715
rect 5365 5690 5370 5710
rect 5370 5690 5390 5710
rect 5390 5690 5395 5710
rect 5365 5685 5395 5690
rect 5365 5630 5395 5635
rect 5365 5610 5370 5630
rect 5370 5610 5390 5630
rect 5390 5610 5395 5630
rect 5365 5605 5395 5610
rect 5365 5550 5395 5555
rect 5365 5530 5370 5550
rect 5370 5530 5390 5550
rect 5390 5530 5395 5550
rect 5365 5525 5395 5530
rect 5365 5470 5395 5475
rect 5365 5450 5370 5470
rect 5370 5450 5390 5470
rect 5390 5450 5395 5470
rect 5365 5445 5395 5450
rect 5365 5390 5395 5395
rect 5365 5370 5370 5390
rect 5370 5370 5390 5390
rect 5390 5370 5395 5390
rect 5365 5365 5395 5370
rect 5365 5310 5395 5315
rect 5365 5290 5370 5310
rect 5370 5290 5390 5310
rect 5390 5290 5395 5310
rect 5365 5285 5395 5290
rect 5365 5230 5395 5235
rect 5365 5210 5370 5230
rect 5370 5210 5390 5230
rect 5390 5210 5395 5230
rect 5365 5205 5395 5210
rect 5365 5150 5395 5155
rect 5365 5130 5370 5150
rect 5370 5130 5390 5150
rect 5390 5130 5395 5150
rect 5365 5125 5395 5130
rect 5365 5070 5395 5075
rect 5365 5050 5370 5070
rect 5370 5050 5390 5070
rect 5390 5050 5395 5070
rect 5365 5045 5395 5050
rect 5365 4990 5395 4995
rect 5365 4970 5370 4990
rect 5370 4970 5390 4990
rect 5390 4970 5395 4990
rect 5365 4965 5395 4970
rect 5365 4910 5395 4915
rect 5365 4890 5370 4910
rect 5370 4890 5390 4910
rect 5390 4890 5395 4910
rect 5365 4885 5395 4890
rect 5365 4750 5395 4755
rect 5365 4730 5370 4750
rect 5370 4730 5390 4750
rect 5390 4730 5395 4750
rect 5365 4725 5395 4730
rect 5365 4670 5395 4675
rect 5365 4650 5370 4670
rect 5370 4650 5390 4670
rect 5390 4650 5395 4670
rect 5365 4645 5395 4650
rect 5365 4510 5395 4515
rect 5365 4490 5370 4510
rect 5370 4490 5390 4510
rect 5390 4490 5395 4510
rect 5365 4485 5395 4490
rect 5365 4430 5395 4435
rect 5365 4410 5370 4430
rect 5370 4410 5390 4430
rect 5390 4410 5395 4430
rect 5365 4405 5395 4410
rect 5365 4350 5395 4355
rect 5365 4330 5370 4350
rect 5370 4330 5390 4350
rect 5390 4330 5395 4350
rect 5365 4325 5395 4330
rect 5365 4270 5395 4275
rect 5365 4250 5370 4270
rect 5370 4250 5390 4270
rect 5390 4250 5395 4270
rect 5365 4245 5395 4250
rect 5365 4190 5395 4195
rect 5365 4170 5370 4190
rect 5370 4170 5390 4190
rect 5390 4170 5395 4190
rect 5365 4165 5395 4170
rect 5365 4110 5395 4115
rect 5365 4090 5370 4110
rect 5370 4090 5390 4110
rect 5390 4090 5395 4110
rect 5365 4085 5395 4090
rect 5365 4030 5395 4035
rect 5365 4010 5370 4030
rect 5370 4010 5390 4030
rect 5390 4010 5395 4030
rect 5365 4005 5395 4010
rect 5365 3950 5395 3955
rect 5365 3930 5370 3950
rect 5370 3930 5390 3950
rect 5390 3930 5395 3950
rect 5365 3925 5395 3930
rect 5365 3870 5395 3875
rect 5365 3850 5370 3870
rect 5370 3850 5390 3870
rect 5390 3850 5395 3870
rect 5365 3845 5395 3850
rect 5365 3710 5395 3715
rect 5365 3690 5370 3710
rect 5370 3690 5390 3710
rect 5390 3690 5395 3710
rect 5365 3685 5395 3690
rect 5365 3630 5395 3635
rect 5365 3610 5370 3630
rect 5370 3610 5390 3630
rect 5390 3610 5395 3630
rect 5365 3605 5395 3610
rect 5365 3470 5395 3475
rect 5365 3450 5370 3470
rect 5370 3450 5390 3470
rect 5390 3450 5395 3470
rect 5365 3445 5395 3450
rect 5365 3390 5395 3395
rect 5365 3370 5370 3390
rect 5370 3370 5390 3390
rect 5390 3370 5395 3390
rect 5365 3365 5395 3370
rect 5365 3230 5395 3235
rect 5365 3210 5370 3230
rect 5370 3210 5390 3230
rect 5390 3210 5395 3230
rect 5365 3205 5395 3210
rect 5365 3150 5395 3155
rect 5365 3130 5370 3150
rect 5370 3130 5390 3150
rect 5390 3130 5395 3150
rect 5365 3125 5395 3130
rect 5365 3070 5395 3075
rect 5365 3050 5370 3070
rect 5370 3050 5390 3070
rect 5390 3050 5395 3070
rect 5365 3045 5395 3050
rect 5365 2990 5395 2995
rect 5365 2970 5370 2990
rect 5370 2970 5390 2990
rect 5390 2970 5395 2990
rect 5365 2965 5395 2970
rect 5365 2910 5395 2915
rect 5365 2890 5370 2910
rect 5370 2890 5390 2910
rect 5390 2890 5395 2910
rect 5365 2885 5395 2890
rect 5365 2830 5395 2835
rect 5365 2810 5370 2830
rect 5370 2810 5390 2830
rect 5390 2810 5395 2830
rect 5365 2805 5395 2810
rect 5365 2750 5395 2755
rect 5365 2730 5370 2750
rect 5370 2730 5390 2750
rect 5390 2730 5395 2750
rect 5365 2725 5395 2730
rect 5365 2670 5395 2675
rect 5365 2650 5370 2670
rect 5370 2650 5390 2670
rect 5390 2650 5395 2670
rect 5365 2645 5395 2650
rect 5365 2590 5395 2595
rect 5365 2570 5370 2590
rect 5370 2570 5390 2590
rect 5390 2570 5395 2590
rect 5365 2565 5395 2570
rect 5365 2510 5395 2515
rect 5365 2490 5370 2510
rect 5370 2490 5390 2510
rect 5390 2490 5395 2510
rect 5365 2485 5395 2490
rect 5365 2430 5395 2435
rect 5365 2410 5370 2430
rect 5370 2410 5390 2430
rect 5390 2410 5395 2430
rect 5365 2405 5395 2410
rect 5365 2350 5395 2355
rect 5365 2330 5370 2350
rect 5370 2330 5390 2350
rect 5390 2330 5395 2350
rect 5365 2325 5395 2330
rect 5365 2270 5395 2275
rect 5365 2250 5370 2270
rect 5370 2250 5390 2270
rect 5390 2250 5395 2270
rect 5365 2245 5395 2250
rect 5365 2190 5395 2195
rect 5365 2170 5370 2190
rect 5370 2170 5390 2190
rect 5390 2170 5395 2190
rect 5365 2165 5395 2170
rect 5365 2110 5395 2115
rect 5365 2090 5370 2110
rect 5370 2090 5390 2110
rect 5390 2090 5395 2110
rect 5365 2085 5395 2090
rect 5365 2030 5395 2035
rect 5365 2010 5370 2030
rect 5370 2010 5390 2030
rect 5390 2010 5395 2030
rect 5365 2005 5395 2010
rect 5365 1950 5395 1955
rect 5365 1930 5370 1950
rect 5370 1930 5390 1950
rect 5390 1930 5395 1950
rect 5365 1925 5395 1930
rect 5365 1710 5395 1715
rect 5365 1690 5370 1710
rect 5370 1690 5390 1710
rect 5390 1690 5395 1710
rect 5365 1685 5395 1690
rect 5365 1630 5395 1635
rect 5365 1610 5370 1630
rect 5370 1610 5390 1630
rect 5390 1610 5395 1630
rect 5365 1605 5395 1610
rect 5365 1550 5395 1555
rect 5365 1530 5370 1550
rect 5370 1530 5390 1550
rect 5390 1530 5395 1550
rect 5365 1525 5395 1530
rect 5365 1470 5395 1475
rect 5365 1450 5370 1470
rect 5370 1450 5390 1470
rect 5390 1450 5395 1470
rect 5365 1445 5395 1450
rect 5365 1390 5395 1395
rect 5365 1370 5370 1390
rect 5370 1370 5390 1390
rect 5390 1370 5395 1390
rect 5365 1365 5395 1370
rect 5365 1310 5395 1315
rect 5365 1290 5370 1310
rect 5370 1290 5390 1310
rect 5390 1290 5395 1310
rect 5365 1285 5395 1290
rect 5365 1230 5395 1235
rect 5365 1210 5370 1230
rect 5370 1210 5390 1230
rect 5390 1210 5395 1230
rect 5365 1205 5395 1210
rect 5365 1150 5395 1155
rect 5365 1130 5370 1150
rect 5370 1130 5390 1150
rect 5390 1130 5395 1150
rect 5365 1125 5395 1130
rect 5365 1070 5395 1075
rect 5365 1050 5370 1070
rect 5370 1050 5390 1070
rect 5390 1050 5395 1070
rect 5365 1045 5395 1050
rect 5365 990 5395 995
rect 5365 970 5370 990
rect 5370 970 5390 990
rect 5390 970 5395 990
rect 5365 965 5395 970
rect 5365 830 5395 835
rect 5365 810 5370 830
rect 5370 810 5390 830
rect 5390 810 5395 830
rect 5365 805 5395 810
rect 5365 750 5395 755
rect 5365 730 5370 750
rect 5370 730 5390 750
rect 5390 730 5395 750
rect 5365 725 5395 730
rect 5365 670 5395 675
rect 5365 650 5370 670
rect 5370 650 5390 670
rect 5390 650 5395 670
rect 5365 645 5395 650
rect 5365 590 5395 595
rect 5365 570 5370 590
rect 5370 570 5390 590
rect 5390 570 5395 590
rect 5365 565 5395 570
rect 5365 510 5395 515
rect 5365 490 5370 510
rect 5370 490 5390 510
rect 5390 490 5395 510
rect 5365 485 5395 490
rect 5365 270 5395 275
rect 5365 250 5370 270
rect 5370 250 5390 270
rect 5390 250 5395 270
rect 5365 245 5395 250
rect 5365 190 5395 195
rect 5365 170 5370 190
rect 5370 170 5390 190
rect 5390 170 5395 190
rect 5365 165 5395 170
rect 5365 110 5395 115
rect 5365 90 5370 110
rect 5370 90 5390 110
rect 5390 90 5395 110
rect 5365 85 5395 90
rect 5365 30 5395 35
rect 5365 10 5370 30
rect 5370 10 5390 30
rect 5390 10 5395 30
rect 5365 5 5395 10
rect 5525 15710 5555 15715
rect 5525 15690 5530 15710
rect 5530 15690 5550 15710
rect 5550 15690 5555 15710
rect 5525 15685 5555 15690
rect 5525 15630 5555 15635
rect 5525 15610 5530 15630
rect 5530 15610 5550 15630
rect 5550 15610 5555 15630
rect 5525 15605 5555 15610
rect 5525 15550 5555 15555
rect 5525 15530 5530 15550
rect 5530 15530 5550 15550
rect 5550 15530 5555 15550
rect 5525 15525 5555 15530
rect 5525 15470 5555 15475
rect 5525 15450 5530 15470
rect 5530 15450 5550 15470
rect 5550 15450 5555 15470
rect 5525 15445 5555 15450
rect 5525 15390 5555 15395
rect 5525 15370 5530 15390
rect 5530 15370 5550 15390
rect 5550 15370 5555 15390
rect 5525 15365 5555 15370
rect 5525 15310 5555 15315
rect 5525 15290 5530 15310
rect 5530 15290 5550 15310
rect 5550 15290 5555 15310
rect 5525 15285 5555 15290
rect 5525 15230 5555 15235
rect 5525 15210 5530 15230
rect 5530 15210 5550 15230
rect 5550 15210 5555 15230
rect 5525 15205 5555 15210
rect 5525 15150 5555 15155
rect 5525 15130 5530 15150
rect 5530 15130 5550 15150
rect 5550 15130 5555 15150
rect 5525 15125 5555 15130
rect 5525 14990 5555 14995
rect 5525 14970 5530 14990
rect 5530 14970 5550 14990
rect 5550 14970 5555 14990
rect 5525 14965 5555 14970
rect 5525 14910 5555 14915
rect 5525 14890 5530 14910
rect 5530 14890 5550 14910
rect 5550 14890 5555 14910
rect 5525 14885 5555 14890
rect 5525 14830 5555 14835
rect 5525 14810 5530 14830
rect 5530 14810 5550 14830
rect 5550 14810 5555 14830
rect 5525 14805 5555 14810
rect 5525 14750 5555 14755
rect 5525 14730 5530 14750
rect 5530 14730 5550 14750
rect 5550 14730 5555 14750
rect 5525 14725 5555 14730
rect 5525 14670 5555 14675
rect 5525 14650 5530 14670
rect 5530 14650 5550 14670
rect 5550 14650 5555 14670
rect 5525 14645 5555 14650
rect 5525 14590 5555 14595
rect 5525 14570 5530 14590
rect 5530 14570 5550 14590
rect 5550 14570 5555 14590
rect 5525 14565 5555 14570
rect 5525 14510 5555 14515
rect 5525 14490 5530 14510
rect 5530 14490 5550 14510
rect 5550 14490 5555 14510
rect 5525 14485 5555 14490
rect 5525 14430 5555 14435
rect 5525 14410 5530 14430
rect 5530 14410 5550 14430
rect 5550 14410 5555 14430
rect 5525 14405 5555 14410
rect 5525 14030 5555 14035
rect 5525 14010 5530 14030
rect 5530 14010 5550 14030
rect 5550 14010 5555 14030
rect 5525 14005 5555 14010
rect 5525 13950 5555 13955
rect 5525 13930 5530 13950
rect 5530 13930 5550 13950
rect 5550 13930 5555 13950
rect 5525 13925 5555 13930
rect 5525 13870 5555 13875
rect 5525 13850 5530 13870
rect 5530 13850 5550 13870
rect 5550 13850 5555 13870
rect 5525 13845 5555 13850
rect 5525 13790 5555 13795
rect 5525 13770 5530 13790
rect 5530 13770 5550 13790
rect 5550 13770 5555 13790
rect 5525 13765 5555 13770
rect 5525 13710 5555 13715
rect 5525 13690 5530 13710
rect 5530 13690 5550 13710
rect 5550 13690 5555 13710
rect 5525 13685 5555 13690
rect 5525 13630 5555 13635
rect 5525 13610 5530 13630
rect 5530 13610 5550 13630
rect 5550 13610 5555 13630
rect 5525 13605 5555 13610
rect 5525 13550 5555 13555
rect 5525 13530 5530 13550
rect 5530 13530 5550 13550
rect 5550 13530 5555 13550
rect 5525 13525 5555 13530
rect 5525 13470 5555 13475
rect 5525 13450 5530 13470
rect 5530 13450 5550 13470
rect 5550 13450 5555 13470
rect 5525 13445 5555 13450
rect 5525 13070 5555 13075
rect 5525 13050 5530 13070
rect 5530 13050 5550 13070
rect 5550 13050 5555 13070
rect 5525 13045 5555 13050
rect 5525 12990 5555 12995
rect 5525 12970 5530 12990
rect 5530 12970 5550 12990
rect 5550 12970 5555 12990
rect 5525 12965 5555 12970
rect 5525 12910 5555 12915
rect 5525 12890 5530 12910
rect 5530 12890 5550 12910
rect 5550 12890 5555 12910
rect 5525 12885 5555 12890
rect 5525 12830 5555 12835
rect 5525 12810 5530 12830
rect 5530 12810 5550 12830
rect 5550 12810 5555 12830
rect 5525 12805 5555 12810
rect 5525 12750 5555 12755
rect 5525 12730 5530 12750
rect 5530 12730 5550 12750
rect 5550 12730 5555 12750
rect 5525 12725 5555 12730
rect 5525 12670 5555 12675
rect 5525 12650 5530 12670
rect 5530 12650 5550 12670
rect 5550 12650 5555 12670
rect 5525 12645 5555 12650
rect 5525 12590 5555 12595
rect 5525 12570 5530 12590
rect 5530 12570 5550 12590
rect 5550 12570 5555 12590
rect 5525 12565 5555 12570
rect 5525 12510 5555 12515
rect 5525 12490 5530 12510
rect 5530 12490 5550 12510
rect 5550 12490 5555 12510
rect 5525 12485 5555 12490
rect 5525 12350 5555 12355
rect 5525 12330 5530 12350
rect 5530 12330 5550 12350
rect 5550 12330 5555 12350
rect 5525 12325 5555 12330
rect 5525 12270 5555 12275
rect 5525 12250 5530 12270
rect 5530 12250 5550 12270
rect 5550 12250 5555 12270
rect 5525 12245 5555 12250
rect 5525 12190 5555 12195
rect 5525 12170 5530 12190
rect 5530 12170 5550 12190
rect 5550 12170 5555 12190
rect 5525 12165 5555 12170
rect 5525 12110 5555 12115
rect 5525 12090 5530 12110
rect 5530 12090 5550 12110
rect 5550 12090 5555 12110
rect 5525 12085 5555 12090
rect 5525 12030 5555 12035
rect 5525 12010 5530 12030
rect 5530 12010 5550 12030
rect 5550 12010 5555 12030
rect 5525 12005 5555 12010
rect 5525 11950 5555 11955
rect 5525 11930 5530 11950
rect 5530 11930 5550 11950
rect 5550 11930 5555 11950
rect 5525 11925 5555 11930
rect 5525 11870 5555 11875
rect 5525 11850 5530 11870
rect 5530 11850 5550 11870
rect 5550 11850 5555 11870
rect 5525 11845 5555 11850
rect 5525 11790 5555 11795
rect 5525 11770 5530 11790
rect 5530 11770 5550 11790
rect 5550 11770 5555 11790
rect 5525 11765 5555 11770
rect 5525 11710 5555 11715
rect 5525 11690 5530 11710
rect 5530 11690 5550 11710
rect 5550 11690 5555 11710
rect 5525 11685 5555 11690
rect 5525 11630 5555 11635
rect 5525 11610 5530 11630
rect 5530 11610 5550 11630
rect 5550 11610 5555 11630
rect 5525 11605 5555 11610
rect 5525 11550 5555 11555
rect 5525 11530 5530 11550
rect 5530 11530 5550 11550
rect 5550 11530 5555 11550
rect 5525 11525 5555 11530
rect 5525 11470 5555 11475
rect 5525 11450 5530 11470
rect 5530 11450 5550 11470
rect 5550 11450 5555 11470
rect 5525 11445 5555 11450
rect 5525 11390 5555 11395
rect 5525 11370 5530 11390
rect 5530 11370 5550 11390
rect 5550 11370 5555 11390
rect 5525 11365 5555 11370
rect 5525 11310 5555 11315
rect 5525 11290 5530 11310
rect 5530 11290 5550 11310
rect 5550 11290 5555 11310
rect 5525 11285 5555 11290
rect 5525 11230 5555 11235
rect 5525 11210 5530 11230
rect 5530 11210 5550 11230
rect 5550 11210 5555 11230
rect 5525 11205 5555 11210
rect 5525 11150 5555 11155
rect 5525 11130 5530 11150
rect 5530 11130 5550 11150
rect 5550 11130 5555 11150
rect 5525 11125 5555 11130
rect 5525 11070 5555 11075
rect 5525 11050 5530 11070
rect 5530 11050 5550 11070
rect 5550 11050 5555 11070
rect 5525 11045 5555 11050
rect 5525 10910 5555 10915
rect 5525 10890 5530 10910
rect 5530 10890 5550 10910
rect 5550 10890 5555 10910
rect 5525 10885 5555 10890
rect 5525 10830 5555 10835
rect 5525 10810 5530 10830
rect 5530 10810 5550 10830
rect 5550 10810 5555 10830
rect 5525 10805 5555 10810
rect 5525 10750 5555 10755
rect 5525 10730 5530 10750
rect 5530 10730 5550 10750
rect 5550 10730 5555 10750
rect 5525 10725 5555 10730
rect 5525 10670 5555 10675
rect 5525 10650 5530 10670
rect 5530 10650 5550 10670
rect 5550 10650 5555 10670
rect 5525 10645 5555 10650
rect 5525 10590 5555 10595
rect 5525 10570 5530 10590
rect 5530 10570 5550 10590
rect 5550 10570 5555 10590
rect 5525 10565 5555 10570
rect 5525 10510 5555 10515
rect 5525 10490 5530 10510
rect 5530 10490 5550 10510
rect 5550 10490 5555 10510
rect 5525 10485 5555 10490
rect 5525 10430 5555 10435
rect 5525 10410 5530 10430
rect 5530 10410 5550 10430
rect 5550 10410 5555 10430
rect 5525 10405 5555 10410
rect 5525 10350 5555 10355
rect 5525 10330 5530 10350
rect 5530 10330 5550 10350
rect 5550 10330 5555 10350
rect 5525 10325 5555 10330
rect 5525 9950 5555 9955
rect 5525 9930 5530 9950
rect 5530 9930 5550 9950
rect 5550 9930 5555 9950
rect 5525 9925 5555 9930
rect 5525 9870 5555 9875
rect 5525 9850 5530 9870
rect 5530 9850 5550 9870
rect 5550 9850 5555 9870
rect 5525 9845 5555 9850
rect 5525 9790 5555 9795
rect 5525 9770 5530 9790
rect 5530 9770 5550 9790
rect 5550 9770 5555 9790
rect 5525 9765 5555 9770
rect 5525 9710 5555 9715
rect 5525 9690 5530 9710
rect 5530 9690 5550 9710
rect 5550 9690 5555 9710
rect 5525 9685 5555 9690
rect 5525 9630 5555 9635
rect 5525 9610 5530 9630
rect 5530 9610 5550 9630
rect 5550 9610 5555 9630
rect 5525 9605 5555 9610
rect 5525 9550 5555 9555
rect 5525 9530 5530 9550
rect 5530 9530 5550 9550
rect 5550 9530 5555 9550
rect 5525 9525 5555 9530
rect 5525 9470 5555 9475
rect 5525 9450 5530 9470
rect 5530 9450 5550 9470
rect 5550 9450 5555 9470
rect 5525 9445 5555 9450
rect 5525 9390 5555 9395
rect 5525 9370 5530 9390
rect 5530 9370 5550 9390
rect 5550 9370 5555 9390
rect 5525 9365 5555 9370
rect 5525 8990 5555 8995
rect 5525 8970 5530 8990
rect 5530 8970 5550 8990
rect 5550 8970 5555 8990
rect 5525 8965 5555 8970
rect 5525 8910 5555 8915
rect 5525 8890 5530 8910
rect 5530 8890 5550 8910
rect 5550 8890 5555 8910
rect 5525 8885 5555 8890
rect 5525 8830 5555 8835
rect 5525 8810 5530 8830
rect 5530 8810 5550 8830
rect 5550 8810 5555 8830
rect 5525 8805 5555 8810
rect 5525 8750 5555 8755
rect 5525 8730 5530 8750
rect 5530 8730 5550 8750
rect 5550 8730 5555 8750
rect 5525 8725 5555 8730
rect 5525 8670 5555 8675
rect 5525 8650 5530 8670
rect 5530 8650 5550 8670
rect 5550 8650 5555 8670
rect 5525 8645 5555 8650
rect 5525 8590 5555 8595
rect 5525 8570 5530 8590
rect 5530 8570 5550 8590
rect 5550 8570 5555 8590
rect 5525 8565 5555 8570
rect 5525 8510 5555 8515
rect 5525 8490 5530 8510
rect 5530 8490 5550 8510
rect 5550 8490 5555 8510
rect 5525 8485 5555 8490
rect 5525 8430 5555 8435
rect 5525 8410 5530 8430
rect 5530 8410 5550 8430
rect 5550 8410 5555 8430
rect 5525 8405 5555 8410
rect 5525 8270 5555 8275
rect 5525 8250 5530 8270
rect 5530 8250 5550 8270
rect 5550 8250 5555 8270
rect 5525 8245 5555 8250
rect 5525 8190 5555 8195
rect 5525 8170 5530 8190
rect 5530 8170 5550 8190
rect 5550 8170 5555 8190
rect 5525 8165 5555 8170
rect 5525 8110 5555 8115
rect 5525 8090 5530 8110
rect 5530 8090 5550 8110
rect 5550 8090 5555 8110
rect 5525 8085 5555 8090
rect 5525 8030 5555 8035
rect 5525 8010 5530 8030
rect 5530 8010 5550 8030
rect 5550 8010 5555 8030
rect 5525 8005 5555 8010
rect 5525 7950 5555 7955
rect 5525 7930 5530 7950
rect 5530 7930 5550 7950
rect 5550 7930 5555 7950
rect 5525 7925 5555 7930
rect 5525 7870 5555 7875
rect 5525 7850 5530 7870
rect 5530 7850 5550 7870
rect 5550 7850 5555 7870
rect 5525 7845 5555 7850
rect 5525 7790 5555 7795
rect 5525 7770 5530 7790
rect 5530 7770 5550 7790
rect 5550 7770 5555 7790
rect 5525 7765 5555 7770
rect 5525 7710 5555 7715
rect 5525 7690 5530 7710
rect 5530 7690 5550 7710
rect 5550 7690 5555 7710
rect 5525 7685 5555 7690
rect 5525 7630 5555 7635
rect 5525 7610 5530 7630
rect 5530 7610 5550 7630
rect 5550 7610 5555 7630
rect 5525 7605 5555 7610
rect 5525 7550 5555 7555
rect 5525 7530 5530 7550
rect 5530 7530 5550 7550
rect 5550 7530 5555 7550
rect 5525 7525 5555 7530
rect 5525 7470 5555 7475
rect 5525 7450 5530 7470
rect 5530 7450 5550 7470
rect 5550 7450 5555 7470
rect 5525 7445 5555 7450
rect 5525 7390 5555 7395
rect 5525 7370 5530 7390
rect 5530 7370 5550 7390
rect 5550 7370 5555 7390
rect 5525 7365 5555 7370
rect 5525 7310 5555 7315
rect 5525 7290 5530 7310
rect 5530 7290 5550 7310
rect 5550 7290 5555 7310
rect 5525 7285 5555 7290
rect 5525 7230 5555 7235
rect 5525 7210 5530 7230
rect 5530 7210 5550 7230
rect 5550 7210 5555 7230
rect 5525 7205 5555 7210
rect 5525 7150 5555 7155
rect 5525 7130 5530 7150
rect 5530 7130 5550 7150
rect 5550 7130 5555 7150
rect 5525 7125 5555 7130
rect 5525 7070 5555 7075
rect 5525 7050 5530 7070
rect 5530 7050 5550 7070
rect 5550 7050 5555 7070
rect 5525 7045 5555 7050
rect 5525 6990 5555 6995
rect 5525 6970 5530 6990
rect 5530 6970 5550 6990
rect 5550 6970 5555 6990
rect 5525 6965 5555 6970
rect 5525 6830 5555 6835
rect 5525 6810 5530 6830
rect 5530 6810 5550 6830
rect 5550 6810 5555 6830
rect 5525 6805 5555 6810
rect 5525 6750 5555 6755
rect 5525 6730 5530 6750
rect 5530 6730 5550 6750
rect 5550 6730 5555 6750
rect 5525 6725 5555 6730
rect 5525 6670 5555 6675
rect 5525 6650 5530 6670
rect 5530 6650 5550 6670
rect 5550 6650 5555 6670
rect 5525 6645 5555 6650
rect 5525 6590 5555 6595
rect 5525 6570 5530 6590
rect 5530 6570 5550 6590
rect 5550 6570 5555 6590
rect 5525 6565 5555 6570
rect 5525 6510 5555 6515
rect 5525 6490 5530 6510
rect 5530 6490 5550 6510
rect 5550 6490 5555 6510
rect 5525 6485 5555 6490
rect 5525 6430 5555 6435
rect 5525 6410 5530 6430
rect 5530 6410 5550 6430
rect 5550 6410 5555 6430
rect 5525 6405 5555 6410
rect 5525 6350 5555 6355
rect 5525 6330 5530 6350
rect 5530 6330 5550 6350
rect 5550 6330 5555 6350
rect 5525 6325 5555 6330
rect 5525 6270 5555 6275
rect 5525 6250 5530 6270
rect 5530 6250 5550 6270
rect 5550 6250 5555 6270
rect 5525 6245 5555 6250
rect 5525 5870 5555 5875
rect 5525 5850 5530 5870
rect 5530 5850 5550 5870
rect 5550 5850 5555 5870
rect 5525 5845 5555 5850
rect 5525 5790 5555 5795
rect 5525 5770 5530 5790
rect 5530 5770 5550 5790
rect 5550 5770 5555 5790
rect 5525 5765 5555 5770
rect 5525 5710 5555 5715
rect 5525 5690 5530 5710
rect 5530 5690 5550 5710
rect 5550 5690 5555 5710
rect 5525 5685 5555 5690
rect 5525 5630 5555 5635
rect 5525 5610 5530 5630
rect 5530 5610 5550 5630
rect 5550 5610 5555 5630
rect 5525 5605 5555 5610
rect 5525 5550 5555 5555
rect 5525 5530 5530 5550
rect 5530 5530 5550 5550
rect 5550 5530 5555 5550
rect 5525 5525 5555 5530
rect 5525 5470 5555 5475
rect 5525 5450 5530 5470
rect 5530 5450 5550 5470
rect 5550 5450 5555 5470
rect 5525 5445 5555 5450
rect 5525 5390 5555 5395
rect 5525 5370 5530 5390
rect 5530 5370 5550 5390
rect 5550 5370 5555 5390
rect 5525 5365 5555 5370
rect 5525 5310 5555 5315
rect 5525 5290 5530 5310
rect 5530 5290 5550 5310
rect 5550 5290 5555 5310
rect 5525 5285 5555 5290
rect 5525 5230 5555 5235
rect 5525 5210 5530 5230
rect 5530 5210 5550 5230
rect 5550 5210 5555 5230
rect 5525 5205 5555 5210
rect 5525 5150 5555 5155
rect 5525 5130 5530 5150
rect 5530 5130 5550 5150
rect 5550 5130 5555 5150
rect 5525 5125 5555 5130
rect 5525 5070 5555 5075
rect 5525 5050 5530 5070
rect 5530 5050 5550 5070
rect 5550 5050 5555 5070
rect 5525 5045 5555 5050
rect 5525 4990 5555 4995
rect 5525 4970 5530 4990
rect 5530 4970 5550 4990
rect 5550 4970 5555 4990
rect 5525 4965 5555 4970
rect 5525 4910 5555 4915
rect 5525 4890 5530 4910
rect 5530 4890 5550 4910
rect 5550 4890 5555 4910
rect 5525 4885 5555 4890
rect 5525 4750 5555 4755
rect 5525 4730 5530 4750
rect 5530 4730 5550 4750
rect 5550 4730 5555 4750
rect 5525 4725 5555 4730
rect 5525 4670 5555 4675
rect 5525 4650 5530 4670
rect 5530 4650 5550 4670
rect 5550 4650 5555 4670
rect 5525 4645 5555 4650
rect 5525 4510 5555 4515
rect 5525 4490 5530 4510
rect 5530 4490 5550 4510
rect 5550 4490 5555 4510
rect 5525 4485 5555 4490
rect 5525 4430 5555 4435
rect 5525 4410 5530 4430
rect 5530 4410 5550 4430
rect 5550 4410 5555 4430
rect 5525 4405 5555 4410
rect 5525 4350 5555 4355
rect 5525 4330 5530 4350
rect 5530 4330 5550 4350
rect 5550 4330 5555 4350
rect 5525 4325 5555 4330
rect 5525 4270 5555 4275
rect 5525 4250 5530 4270
rect 5530 4250 5550 4270
rect 5550 4250 5555 4270
rect 5525 4245 5555 4250
rect 5525 4190 5555 4195
rect 5525 4170 5530 4190
rect 5530 4170 5550 4190
rect 5550 4170 5555 4190
rect 5525 4165 5555 4170
rect 5525 4110 5555 4115
rect 5525 4090 5530 4110
rect 5530 4090 5550 4110
rect 5550 4090 5555 4110
rect 5525 4085 5555 4090
rect 5525 4030 5555 4035
rect 5525 4010 5530 4030
rect 5530 4010 5550 4030
rect 5550 4010 5555 4030
rect 5525 4005 5555 4010
rect 5525 3950 5555 3955
rect 5525 3930 5530 3950
rect 5530 3930 5550 3950
rect 5550 3930 5555 3950
rect 5525 3925 5555 3930
rect 5525 3870 5555 3875
rect 5525 3850 5530 3870
rect 5530 3850 5550 3870
rect 5550 3850 5555 3870
rect 5525 3845 5555 3850
rect 5525 3710 5555 3715
rect 5525 3690 5530 3710
rect 5530 3690 5550 3710
rect 5550 3690 5555 3710
rect 5525 3685 5555 3690
rect 5525 3630 5555 3635
rect 5525 3610 5530 3630
rect 5530 3610 5550 3630
rect 5550 3610 5555 3630
rect 5525 3605 5555 3610
rect 5525 3470 5555 3475
rect 5525 3450 5530 3470
rect 5530 3450 5550 3470
rect 5550 3450 5555 3470
rect 5525 3445 5555 3450
rect 5525 3390 5555 3395
rect 5525 3370 5530 3390
rect 5530 3370 5550 3390
rect 5550 3370 5555 3390
rect 5525 3365 5555 3370
rect 5525 3230 5555 3235
rect 5525 3210 5530 3230
rect 5530 3210 5550 3230
rect 5550 3210 5555 3230
rect 5525 3205 5555 3210
rect 5525 3150 5555 3155
rect 5525 3130 5530 3150
rect 5530 3130 5550 3150
rect 5550 3130 5555 3150
rect 5525 3125 5555 3130
rect 5525 3070 5555 3075
rect 5525 3050 5530 3070
rect 5530 3050 5550 3070
rect 5550 3050 5555 3070
rect 5525 3045 5555 3050
rect 5525 2990 5555 2995
rect 5525 2970 5530 2990
rect 5530 2970 5550 2990
rect 5550 2970 5555 2990
rect 5525 2965 5555 2970
rect 5525 2910 5555 2915
rect 5525 2890 5530 2910
rect 5530 2890 5550 2910
rect 5550 2890 5555 2910
rect 5525 2885 5555 2890
rect 5525 2830 5555 2835
rect 5525 2810 5530 2830
rect 5530 2810 5550 2830
rect 5550 2810 5555 2830
rect 5525 2805 5555 2810
rect 5525 2750 5555 2755
rect 5525 2730 5530 2750
rect 5530 2730 5550 2750
rect 5550 2730 5555 2750
rect 5525 2725 5555 2730
rect 5525 2670 5555 2675
rect 5525 2650 5530 2670
rect 5530 2650 5550 2670
rect 5550 2650 5555 2670
rect 5525 2645 5555 2650
rect 5525 2590 5555 2595
rect 5525 2570 5530 2590
rect 5530 2570 5550 2590
rect 5550 2570 5555 2590
rect 5525 2565 5555 2570
rect 5525 2510 5555 2515
rect 5525 2490 5530 2510
rect 5530 2490 5550 2510
rect 5550 2490 5555 2510
rect 5525 2485 5555 2490
rect 5525 2430 5555 2435
rect 5525 2410 5530 2430
rect 5530 2410 5550 2430
rect 5550 2410 5555 2430
rect 5525 2405 5555 2410
rect 5525 2350 5555 2355
rect 5525 2330 5530 2350
rect 5530 2330 5550 2350
rect 5550 2330 5555 2350
rect 5525 2325 5555 2330
rect 5525 2270 5555 2275
rect 5525 2250 5530 2270
rect 5530 2250 5550 2270
rect 5550 2250 5555 2270
rect 5525 2245 5555 2250
rect 5525 2190 5555 2195
rect 5525 2170 5530 2190
rect 5530 2170 5550 2190
rect 5550 2170 5555 2190
rect 5525 2165 5555 2170
rect 5525 2110 5555 2115
rect 5525 2090 5530 2110
rect 5530 2090 5550 2110
rect 5550 2090 5555 2110
rect 5525 2085 5555 2090
rect 5525 2030 5555 2035
rect 5525 2010 5530 2030
rect 5530 2010 5550 2030
rect 5550 2010 5555 2030
rect 5525 2005 5555 2010
rect 5525 1950 5555 1955
rect 5525 1930 5530 1950
rect 5530 1930 5550 1950
rect 5550 1930 5555 1950
rect 5525 1925 5555 1930
rect 5525 1710 5555 1715
rect 5525 1690 5530 1710
rect 5530 1690 5550 1710
rect 5550 1690 5555 1710
rect 5525 1685 5555 1690
rect 5525 1630 5555 1635
rect 5525 1610 5530 1630
rect 5530 1610 5550 1630
rect 5550 1610 5555 1630
rect 5525 1605 5555 1610
rect 5525 1550 5555 1555
rect 5525 1530 5530 1550
rect 5530 1530 5550 1550
rect 5550 1530 5555 1550
rect 5525 1525 5555 1530
rect 5525 1470 5555 1475
rect 5525 1450 5530 1470
rect 5530 1450 5550 1470
rect 5550 1450 5555 1470
rect 5525 1445 5555 1450
rect 5525 1390 5555 1395
rect 5525 1370 5530 1390
rect 5530 1370 5550 1390
rect 5550 1370 5555 1390
rect 5525 1365 5555 1370
rect 5525 1310 5555 1315
rect 5525 1290 5530 1310
rect 5530 1290 5550 1310
rect 5550 1290 5555 1310
rect 5525 1285 5555 1290
rect 5525 1230 5555 1235
rect 5525 1210 5530 1230
rect 5530 1210 5550 1230
rect 5550 1210 5555 1230
rect 5525 1205 5555 1210
rect 5525 1150 5555 1155
rect 5525 1130 5530 1150
rect 5530 1130 5550 1150
rect 5550 1130 5555 1150
rect 5525 1125 5555 1130
rect 5525 1070 5555 1075
rect 5525 1050 5530 1070
rect 5530 1050 5550 1070
rect 5550 1050 5555 1070
rect 5525 1045 5555 1050
rect 5525 990 5555 995
rect 5525 970 5530 990
rect 5530 970 5550 990
rect 5550 970 5555 990
rect 5525 965 5555 970
rect 5525 830 5555 835
rect 5525 810 5530 830
rect 5530 810 5550 830
rect 5550 810 5555 830
rect 5525 805 5555 810
rect 5525 750 5555 755
rect 5525 730 5530 750
rect 5530 730 5550 750
rect 5550 730 5555 750
rect 5525 725 5555 730
rect 5525 670 5555 675
rect 5525 650 5530 670
rect 5530 650 5550 670
rect 5550 650 5555 670
rect 5525 645 5555 650
rect 5525 590 5555 595
rect 5525 570 5530 590
rect 5530 570 5550 590
rect 5550 570 5555 590
rect 5525 565 5555 570
rect 5525 510 5555 515
rect 5525 490 5530 510
rect 5530 490 5550 510
rect 5550 490 5555 510
rect 5525 485 5555 490
rect 5525 270 5555 275
rect 5525 250 5530 270
rect 5530 250 5550 270
rect 5550 250 5555 270
rect 5525 245 5555 250
rect 5525 190 5555 195
rect 5525 170 5530 190
rect 5530 170 5550 190
rect 5550 170 5555 190
rect 5525 165 5555 170
rect 5525 110 5555 115
rect 5525 90 5530 110
rect 5530 90 5550 110
rect 5550 90 5555 110
rect 5525 85 5555 90
rect 5525 30 5555 35
rect 5525 10 5530 30
rect 5530 10 5550 30
rect 5550 10 5555 30
rect 5525 5 5555 10
rect 5685 15710 5715 15715
rect 5685 15690 5690 15710
rect 5690 15690 5710 15710
rect 5710 15690 5715 15710
rect 5685 15685 5715 15690
rect 5685 15630 5715 15635
rect 5685 15610 5690 15630
rect 5690 15610 5710 15630
rect 5710 15610 5715 15630
rect 5685 15605 5715 15610
rect 5685 15550 5715 15555
rect 5685 15530 5690 15550
rect 5690 15530 5710 15550
rect 5710 15530 5715 15550
rect 5685 15525 5715 15530
rect 5685 15470 5715 15475
rect 5685 15450 5690 15470
rect 5690 15450 5710 15470
rect 5710 15450 5715 15470
rect 5685 15445 5715 15450
rect 5685 15390 5715 15395
rect 5685 15370 5690 15390
rect 5690 15370 5710 15390
rect 5710 15370 5715 15390
rect 5685 15365 5715 15370
rect 5685 15310 5715 15315
rect 5685 15290 5690 15310
rect 5690 15290 5710 15310
rect 5710 15290 5715 15310
rect 5685 15285 5715 15290
rect 5685 15230 5715 15235
rect 5685 15210 5690 15230
rect 5690 15210 5710 15230
rect 5710 15210 5715 15230
rect 5685 15205 5715 15210
rect 5685 15150 5715 15155
rect 5685 15130 5690 15150
rect 5690 15130 5710 15150
rect 5710 15130 5715 15150
rect 5685 15125 5715 15130
rect 5685 14990 5715 14995
rect 5685 14970 5690 14990
rect 5690 14970 5710 14990
rect 5710 14970 5715 14990
rect 5685 14965 5715 14970
rect 5685 14910 5715 14915
rect 5685 14890 5690 14910
rect 5690 14890 5710 14910
rect 5710 14890 5715 14910
rect 5685 14885 5715 14890
rect 5685 14830 5715 14835
rect 5685 14810 5690 14830
rect 5690 14810 5710 14830
rect 5710 14810 5715 14830
rect 5685 14805 5715 14810
rect 5685 14750 5715 14755
rect 5685 14730 5690 14750
rect 5690 14730 5710 14750
rect 5710 14730 5715 14750
rect 5685 14725 5715 14730
rect 5685 14670 5715 14675
rect 5685 14650 5690 14670
rect 5690 14650 5710 14670
rect 5710 14650 5715 14670
rect 5685 14645 5715 14650
rect 5685 14590 5715 14595
rect 5685 14570 5690 14590
rect 5690 14570 5710 14590
rect 5710 14570 5715 14590
rect 5685 14565 5715 14570
rect 5685 14510 5715 14515
rect 5685 14490 5690 14510
rect 5690 14490 5710 14510
rect 5710 14490 5715 14510
rect 5685 14485 5715 14490
rect 5685 14430 5715 14435
rect 5685 14410 5690 14430
rect 5690 14410 5710 14430
rect 5710 14410 5715 14430
rect 5685 14405 5715 14410
rect 5685 14030 5715 14035
rect 5685 14010 5690 14030
rect 5690 14010 5710 14030
rect 5710 14010 5715 14030
rect 5685 14005 5715 14010
rect 5685 13950 5715 13955
rect 5685 13930 5690 13950
rect 5690 13930 5710 13950
rect 5710 13930 5715 13950
rect 5685 13925 5715 13930
rect 5685 13870 5715 13875
rect 5685 13850 5690 13870
rect 5690 13850 5710 13870
rect 5710 13850 5715 13870
rect 5685 13845 5715 13850
rect 5685 13790 5715 13795
rect 5685 13770 5690 13790
rect 5690 13770 5710 13790
rect 5710 13770 5715 13790
rect 5685 13765 5715 13770
rect 5685 13710 5715 13715
rect 5685 13690 5690 13710
rect 5690 13690 5710 13710
rect 5710 13690 5715 13710
rect 5685 13685 5715 13690
rect 5685 13630 5715 13635
rect 5685 13610 5690 13630
rect 5690 13610 5710 13630
rect 5710 13610 5715 13630
rect 5685 13605 5715 13610
rect 5685 13550 5715 13555
rect 5685 13530 5690 13550
rect 5690 13530 5710 13550
rect 5710 13530 5715 13550
rect 5685 13525 5715 13530
rect 5685 13470 5715 13475
rect 5685 13450 5690 13470
rect 5690 13450 5710 13470
rect 5710 13450 5715 13470
rect 5685 13445 5715 13450
rect 5685 13070 5715 13075
rect 5685 13050 5690 13070
rect 5690 13050 5710 13070
rect 5710 13050 5715 13070
rect 5685 13045 5715 13050
rect 5685 12990 5715 12995
rect 5685 12970 5690 12990
rect 5690 12970 5710 12990
rect 5710 12970 5715 12990
rect 5685 12965 5715 12970
rect 5685 12910 5715 12915
rect 5685 12890 5690 12910
rect 5690 12890 5710 12910
rect 5710 12890 5715 12910
rect 5685 12885 5715 12890
rect 5685 12830 5715 12835
rect 5685 12810 5690 12830
rect 5690 12810 5710 12830
rect 5710 12810 5715 12830
rect 5685 12805 5715 12810
rect 5685 12750 5715 12755
rect 5685 12730 5690 12750
rect 5690 12730 5710 12750
rect 5710 12730 5715 12750
rect 5685 12725 5715 12730
rect 5685 12670 5715 12675
rect 5685 12650 5690 12670
rect 5690 12650 5710 12670
rect 5710 12650 5715 12670
rect 5685 12645 5715 12650
rect 5685 12590 5715 12595
rect 5685 12570 5690 12590
rect 5690 12570 5710 12590
rect 5710 12570 5715 12590
rect 5685 12565 5715 12570
rect 5685 12510 5715 12515
rect 5685 12490 5690 12510
rect 5690 12490 5710 12510
rect 5710 12490 5715 12510
rect 5685 12485 5715 12490
rect 5685 12350 5715 12355
rect 5685 12330 5690 12350
rect 5690 12330 5710 12350
rect 5710 12330 5715 12350
rect 5685 12325 5715 12330
rect 5685 12270 5715 12275
rect 5685 12250 5690 12270
rect 5690 12250 5710 12270
rect 5710 12250 5715 12270
rect 5685 12245 5715 12250
rect 5685 12190 5715 12195
rect 5685 12170 5690 12190
rect 5690 12170 5710 12190
rect 5710 12170 5715 12190
rect 5685 12165 5715 12170
rect 5685 12110 5715 12115
rect 5685 12090 5690 12110
rect 5690 12090 5710 12110
rect 5710 12090 5715 12110
rect 5685 12085 5715 12090
rect 5685 12030 5715 12035
rect 5685 12010 5690 12030
rect 5690 12010 5710 12030
rect 5710 12010 5715 12030
rect 5685 12005 5715 12010
rect 5685 11950 5715 11955
rect 5685 11930 5690 11950
rect 5690 11930 5710 11950
rect 5710 11930 5715 11950
rect 5685 11925 5715 11930
rect 5685 11870 5715 11875
rect 5685 11850 5690 11870
rect 5690 11850 5710 11870
rect 5710 11850 5715 11870
rect 5685 11845 5715 11850
rect 5685 11790 5715 11795
rect 5685 11770 5690 11790
rect 5690 11770 5710 11790
rect 5710 11770 5715 11790
rect 5685 11765 5715 11770
rect 5685 11710 5715 11715
rect 5685 11690 5690 11710
rect 5690 11690 5710 11710
rect 5710 11690 5715 11710
rect 5685 11685 5715 11690
rect 5685 11630 5715 11635
rect 5685 11610 5690 11630
rect 5690 11610 5710 11630
rect 5710 11610 5715 11630
rect 5685 11605 5715 11610
rect 5685 11550 5715 11555
rect 5685 11530 5690 11550
rect 5690 11530 5710 11550
rect 5710 11530 5715 11550
rect 5685 11525 5715 11530
rect 5685 11470 5715 11475
rect 5685 11450 5690 11470
rect 5690 11450 5710 11470
rect 5710 11450 5715 11470
rect 5685 11445 5715 11450
rect 5685 11390 5715 11395
rect 5685 11370 5690 11390
rect 5690 11370 5710 11390
rect 5710 11370 5715 11390
rect 5685 11365 5715 11370
rect 5685 11310 5715 11315
rect 5685 11290 5690 11310
rect 5690 11290 5710 11310
rect 5710 11290 5715 11310
rect 5685 11285 5715 11290
rect 5685 11230 5715 11235
rect 5685 11210 5690 11230
rect 5690 11210 5710 11230
rect 5710 11210 5715 11230
rect 5685 11205 5715 11210
rect 5685 11150 5715 11155
rect 5685 11130 5690 11150
rect 5690 11130 5710 11150
rect 5710 11130 5715 11150
rect 5685 11125 5715 11130
rect 5685 11070 5715 11075
rect 5685 11050 5690 11070
rect 5690 11050 5710 11070
rect 5710 11050 5715 11070
rect 5685 11045 5715 11050
rect 5685 10910 5715 10915
rect 5685 10890 5690 10910
rect 5690 10890 5710 10910
rect 5710 10890 5715 10910
rect 5685 10885 5715 10890
rect 5685 10830 5715 10835
rect 5685 10810 5690 10830
rect 5690 10810 5710 10830
rect 5710 10810 5715 10830
rect 5685 10805 5715 10810
rect 5685 10750 5715 10755
rect 5685 10730 5690 10750
rect 5690 10730 5710 10750
rect 5710 10730 5715 10750
rect 5685 10725 5715 10730
rect 5685 10670 5715 10675
rect 5685 10650 5690 10670
rect 5690 10650 5710 10670
rect 5710 10650 5715 10670
rect 5685 10645 5715 10650
rect 5685 10590 5715 10595
rect 5685 10570 5690 10590
rect 5690 10570 5710 10590
rect 5710 10570 5715 10590
rect 5685 10565 5715 10570
rect 5685 10510 5715 10515
rect 5685 10490 5690 10510
rect 5690 10490 5710 10510
rect 5710 10490 5715 10510
rect 5685 10485 5715 10490
rect 5685 10430 5715 10435
rect 5685 10410 5690 10430
rect 5690 10410 5710 10430
rect 5710 10410 5715 10430
rect 5685 10405 5715 10410
rect 5685 10350 5715 10355
rect 5685 10330 5690 10350
rect 5690 10330 5710 10350
rect 5710 10330 5715 10350
rect 5685 10325 5715 10330
rect 5685 9950 5715 9955
rect 5685 9930 5690 9950
rect 5690 9930 5710 9950
rect 5710 9930 5715 9950
rect 5685 9925 5715 9930
rect 5685 9870 5715 9875
rect 5685 9850 5690 9870
rect 5690 9850 5710 9870
rect 5710 9850 5715 9870
rect 5685 9845 5715 9850
rect 5685 9790 5715 9795
rect 5685 9770 5690 9790
rect 5690 9770 5710 9790
rect 5710 9770 5715 9790
rect 5685 9765 5715 9770
rect 5685 9710 5715 9715
rect 5685 9690 5690 9710
rect 5690 9690 5710 9710
rect 5710 9690 5715 9710
rect 5685 9685 5715 9690
rect 5685 9630 5715 9635
rect 5685 9610 5690 9630
rect 5690 9610 5710 9630
rect 5710 9610 5715 9630
rect 5685 9605 5715 9610
rect 5685 9550 5715 9555
rect 5685 9530 5690 9550
rect 5690 9530 5710 9550
rect 5710 9530 5715 9550
rect 5685 9525 5715 9530
rect 5685 9470 5715 9475
rect 5685 9450 5690 9470
rect 5690 9450 5710 9470
rect 5710 9450 5715 9470
rect 5685 9445 5715 9450
rect 5685 9390 5715 9395
rect 5685 9370 5690 9390
rect 5690 9370 5710 9390
rect 5710 9370 5715 9390
rect 5685 9365 5715 9370
rect 5685 8990 5715 8995
rect 5685 8970 5690 8990
rect 5690 8970 5710 8990
rect 5710 8970 5715 8990
rect 5685 8965 5715 8970
rect 5685 8910 5715 8915
rect 5685 8890 5690 8910
rect 5690 8890 5710 8910
rect 5710 8890 5715 8910
rect 5685 8885 5715 8890
rect 5685 8830 5715 8835
rect 5685 8810 5690 8830
rect 5690 8810 5710 8830
rect 5710 8810 5715 8830
rect 5685 8805 5715 8810
rect 5685 8750 5715 8755
rect 5685 8730 5690 8750
rect 5690 8730 5710 8750
rect 5710 8730 5715 8750
rect 5685 8725 5715 8730
rect 5685 8670 5715 8675
rect 5685 8650 5690 8670
rect 5690 8650 5710 8670
rect 5710 8650 5715 8670
rect 5685 8645 5715 8650
rect 5685 8590 5715 8595
rect 5685 8570 5690 8590
rect 5690 8570 5710 8590
rect 5710 8570 5715 8590
rect 5685 8565 5715 8570
rect 5685 8510 5715 8515
rect 5685 8490 5690 8510
rect 5690 8490 5710 8510
rect 5710 8490 5715 8510
rect 5685 8485 5715 8490
rect 5685 8430 5715 8435
rect 5685 8410 5690 8430
rect 5690 8410 5710 8430
rect 5710 8410 5715 8430
rect 5685 8405 5715 8410
rect 5685 8270 5715 8275
rect 5685 8250 5690 8270
rect 5690 8250 5710 8270
rect 5710 8250 5715 8270
rect 5685 8245 5715 8250
rect 5685 8190 5715 8195
rect 5685 8170 5690 8190
rect 5690 8170 5710 8190
rect 5710 8170 5715 8190
rect 5685 8165 5715 8170
rect 5685 8110 5715 8115
rect 5685 8090 5690 8110
rect 5690 8090 5710 8110
rect 5710 8090 5715 8110
rect 5685 8085 5715 8090
rect 5685 8030 5715 8035
rect 5685 8010 5690 8030
rect 5690 8010 5710 8030
rect 5710 8010 5715 8030
rect 5685 8005 5715 8010
rect 5685 7950 5715 7955
rect 5685 7930 5690 7950
rect 5690 7930 5710 7950
rect 5710 7930 5715 7950
rect 5685 7925 5715 7930
rect 5685 7870 5715 7875
rect 5685 7850 5690 7870
rect 5690 7850 5710 7870
rect 5710 7850 5715 7870
rect 5685 7845 5715 7850
rect 5685 7790 5715 7795
rect 5685 7770 5690 7790
rect 5690 7770 5710 7790
rect 5710 7770 5715 7790
rect 5685 7765 5715 7770
rect 5685 7710 5715 7715
rect 5685 7690 5690 7710
rect 5690 7690 5710 7710
rect 5710 7690 5715 7710
rect 5685 7685 5715 7690
rect 5685 7630 5715 7635
rect 5685 7610 5690 7630
rect 5690 7610 5710 7630
rect 5710 7610 5715 7630
rect 5685 7605 5715 7610
rect 5685 7550 5715 7555
rect 5685 7530 5690 7550
rect 5690 7530 5710 7550
rect 5710 7530 5715 7550
rect 5685 7525 5715 7530
rect 5685 7470 5715 7475
rect 5685 7450 5690 7470
rect 5690 7450 5710 7470
rect 5710 7450 5715 7470
rect 5685 7445 5715 7450
rect 5685 7390 5715 7395
rect 5685 7370 5690 7390
rect 5690 7370 5710 7390
rect 5710 7370 5715 7390
rect 5685 7365 5715 7370
rect 5685 7310 5715 7315
rect 5685 7290 5690 7310
rect 5690 7290 5710 7310
rect 5710 7290 5715 7310
rect 5685 7285 5715 7290
rect 5685 7230 5715 7235
rect 5685 7210 5690 7230
rect 5690 7210 5710 7230
rect 5710 7210 5715 7230
rect 5685 7205 5715 7210
rect 5685 7150 5715 7155
rect 5685 7130 5690 7150
rect 5690 7130 5710 7150
rect 5710 7130 5715 7150
rect 5685 7125 5715 7130
rect 5685 7070 5715 7075
rect 5685 7050 5690 7070
rect 5690 7050 5710 7070
rect 5710 7050 5715 7070
rect 5685 7045 5715 7050
rect 5685 6990 5715 6995
rect 5685 6970 5690 6990
rect 5690 6970 5710 6990
rect 5710 6970 5715 6990
rect 5685 6965 5715 6970
rect 5685 6830 5715 6835
rect 5685 6810 5690 6830
rect 5690 6810 5710 6830
rect 5710 6810 5715 6830
rect 5685 6805 5715 6810
rect 5685 6750 5715 6755
rect 5685 6730 5690 6750
rect 5690 6730 5710 6750
rect 5710 6730 5715 6750
rect 5685 6725 5715 6730
rect 5685 6670 5715 6675
rect 5685 6650 5690 6670
rect 5690 6650 5710 6670
rect 5710 6650 5715 6670
rect 5685 6645 5715 6650
rect 5685 6590 5715 6595
rect 5685 6570 5690 6590
rect 5690 6570 5710 6590
rect 5710 6570 5715 6590
rect 5685 6565 5715 6570
rect 5685 6510 5715 6515
rect 5685 6490 5690 6510
rect 5690 6490 5710 6510
rect 5710 6490 5715 6510
rect 5685 6485 5715 6490
rect 5685 6430 5715 6435
rect 5685 6410 5690 6430
rect 5690 6410 5710 6430
rect 5710 6410 5715 6430
rect 5685 6405 5715 6410
rect 5685 6350 5715 6355
rect 5685 6330 5690 6350
rect 5690 6330 5710 6350
rect 5710 6330 5715 6350
rect 5685 6325 5715 6330
rect 5685 6270 5715 6275
rect 5685 6250 5690 6270
rect 5690 6250 5710 6270
rect 5710 6250 5715 6270
rect 5685 6245 5715 6250
rect 5685 5870 5715 5875
rect 5685 5850 5690 5870
rect 5690 5850 5710 5870
rect 5710 5850 5715 5870
rect 5685 5845 5715 5850
rect 5685 5790 5715 5795
rect 5685 5770 5690 5790
rect 5690 5770 5710 5790
rect 5710 5770 5715 5790
rect 5685 5765 5715 5770
rect 5685 5710 5715 5715
rect 5685 5690 5690 5710
rect 5690 5690 5710 5710
rect 5710 5690 5715 5710
rect 5685 5685 5715 5690
rect 5685 5630 5715 5635
rect 5685 5610 5690 5630
rect 5690 5610 5710 5630
rect 5710 5610 5715 5630
rect 5685 5605 5715 5610
rect 5685 5550 5715 5555
rect 5685 5530 5690 5550
rect 5690 5530 5710 5550
rect 5710 5530 5715 5550
rect 5685 5525 5715 5530
rect 5685 5470 5715 5475
rect 5685 5450 5690 5470
rect 5690 5450 5710 5470
rect 5710 5450 5715 5470
rect 5685 5445 5715 5450
rect 5685 5390 5715 5395
rect 5685 5370 5690 5390
rect 5690 5370 5710 5390
rect 5710 5370 5715 5390
rect 5685 5365 5715 5370
rect 5685 5310 5715 5315
rect 5685 5290 5690 5310
rect 5690 5290 5710 5310
rect 5710 5290 5715 5310
rect 5685 5285 5715 5290
rect 5685 5230 5715 5235
rect 5685 5210 5690 5230
rect 5690 5210 5710 5230
rect 5710 5210 5715 5230
rect 5685 5205 5715 5210
rect 5685 5150 5715 5155
rect 5685 5130 5690 5150
rect 5690 5130 5710 5150
rect 5710 5130 5715 5150
rect 5685 5125 5715 5130
rect 5685 5070 5715 5075
rect 5685 5050 5690 5070
rect 5690 5050 5710 5070
rect 5710 5050 5715 5070
rect 5685 5045 5715 5050
rect 5685 4990 5715 4995
rect 5685 4970 5690 4990
rect 5690 4970 5710 4990
rect 5710 4970 5715 4990
rect 5685 4965 5715 4970
rect 5685 4910 5715 4915
rect 5685 4890 5690 4910
rect 5690 4890 5710 4910
rect 5710 4890 5715 4910
rect 5685 4885 5715 4890
rect 5685 4750 5715 4755
rect 5685 4730 5690 4750
rect 5690 4730 5710 4750
rect 5710 4730 5715 4750
rect 5685 4725 5715 4730
rect 5685 4670 5715 4675
rect 5685 4650 5690 4670
rect 5690 4650 5710 4670
rect 5710 4650 5715 4670
rect 5685 4645 5715 4650
rect 5685 4510 5715 4515
rect 5685 4490 5690 4510
rect 5690 4490 5710 4510
rect 5710 4490 5715 4510
rect 5685 4485 5715 4490
rect 5685 4430 5715 4435
rect 5685 4410 5690 4430
rect 5690 4410 5710 4430
rect 5710 4410 5715 4430
rect 5685 4405 5715 4410
rect 5685 4350 5715 4355
rect 5685 4330 5690 4350
rect 5690 4330 5710 4350
rect 5710 4330 5715 4350
rect 5685 4325 5715 4330
rect 5685 4270 5715 4275
rect 5685 4250 5690 4270
rect 5690 4250 5710 4270
rect 5710 4250 5715 4270
rect 5685 4245 5715 4250
rect 5685 4190 5715 4195
rect 5685 4170 5690 4190
rect 5690 4170 5710 4190
rect 5710 4170 5715 4190
rect 5685 4165 5715 4170
rect 5685 4110 5715 4115
rect 5685 4090 5690 4110
rect 5690 4090 5710 4110
rect 5710 4090 5715 4110
rect 5685 4085 5715 4090
rect 5685 4030 5715 4035
rect 5685 4010 5690 4030
rect 5690 4010 5710 4030
rect 5710 4010 5715 4030
rect 5685 4005 5715 4010
rect 5685 3950 5715 3955
rect 5685 3930 5690 3950
rect 5690 3930 5710 3950
rect 5710 3930 5715 3950
rect 5685 3925 5715 3930
rect 5685 3870 5715 3875
rect 5685 3850 5690 3870
rect 5690 3850 5710 3870
rect 5710 3850 5715 3870
rect 5685 3845 5715 3850
rect 5685 3710 5715 3715
rect 5685 3690 5690 3710
rect 5690 3690 5710 3710
rect 5710 3690 5715 3710
rect 5685 3685 5715 3690
rect 5685 3630 5715 3635
rect 5685 3610 5690 3630
rect 5690 3610 5710 3630
rect 5710 3610 5715 3630
rect 5685 3605 5715 3610
rect 5685 3470 5715 3475
rect 5685 3450 5690 3470
rect 5690 3450 5710 3470
rect 5710 3450 5715 3470
rect 5685 3445 5715 3450
rect 5685 3390 5715 3395
rect 5685 3370 5690 3390
rect 5690 3370 5710 3390
rect 5710 3370 5715 3390
rect 5685 3365 5715 3370
rect 5685 3230 5715 3235
rect 5685 3210 5690 3230
rect 5690 3210 5710 3230
rect 5710 3210 5715 3230
rect 5685 3205 5715 3210
rect 5685 3150 5715 3155
rect 5685 3130 5690 3150
rect 5690 3130 5710 3150
rect 5710 3130 5715 3150
rect 5685 3125 5715 3130
rect 5685 3070 5715 3075
rect 5685 3050 5690 3070
rect 5690 3050 5710 3070
rect 5710 3050 5715 3070
rect 5685 3045 5715 3050
rect 5685 2990 5715 2995
rect 5685 2970 5690 2990
rect 5690 2970 5710 2990
rect 5710 2970 5715 2990
rect 5685 2965 5715 2970
rect 5685 2910 5715 2915
rect 5685 2890 5690 2910
rect 5690 2890 5710 2910
rect 5710 2890 5715 2910
rect 5685 2885 5715 2890
rect 5685 2830 5715 2835
rect 5685 2810 5690 2830
rect 5690 2810 5710 2830
rect 5710 2810 5715 2830
rect 5685 2805 5715 2810
rect 5685 2750 5715 2755
rect 5685 2730 5690 2750
rect 5690 2730 5710 2750
rect 5710 2730 5715 2750
rect 5685 2725 5715 2730
rect 5685 2670 5715 2675
rect 5685 2650 5690 2670
rect 5690 2650 5710 2670
rect 5710 2650 5715 2670
rect 5685 2645 5715 2650
rect 5685 2590 5715 2595
rect 5685 2570 5690 2590
rect 5690 2570 5710 2590
rect 5710 2570 5715 2590
rect 5685 2565 5715 2570
rect 5685 2510 5715 2515
rect 5685 2490 5690 2510
rect 5690 2490 5710 2510
rect 5710 2490 5715 2510
rect 5685 2485 5715 2490
rect 5685 2430 5715 2435
rect 5685 2410 5690 2430
rect 5690 2410 5710 2430
rect 5710 2410 5715 2430
rect 5685 2405 5715 2410
rect 5685 2350 5715 2355
rect 5685 2330 5690 2350
rect 5690 2330 5710 2350
rect 5710 2330 5715 2350
rect 5685 2325 5715 2330
rect 5685 2270 5715 2275
rect 5685 2250 5690 2270
rect 5690 2250 5710 2270
rect 5710 2250 5715 2270
rect 5685 2245 5715 2250
rect 5685 2190 5715 2195
rect 5685 2170 5690 2190
rect 5690 2170 5710 2190
rect 5710 2170 5715 2190
rect 5685 2165 5715 2170
rect 5685 2110 5715 2115
rect 5685 2090 5690 2110
rect 5690 2090 5710 2110
rect 5710 2090 5715 2110
rect 5685 2085 5715 2090
rect 5685 2030 5715 2035
rect 5685 2010 5690 2030
rect 5690 2010 5710 2030
rect 5710 2010 5715 2030
rect 5685 2005 5715 2010
rect 5685 1950 5715 1955
rect 5685 1930 5690 1950
rect 5690 1930 5710 1950
rect 5710 1930 5715 1950
rect 5685 1925 5715 1930
rect 5685 1710 5715 1715
rect 5685 1690 5690 1710
rect 5690 1690 5710 1710
rect 5710 1690 5715 1710
rect 5685 1685 5715 1690
rect 5685 1630 5715 1635
rect 5685 1610 5690 1630
rect 5690 1610 5710 1630
rect 5710 1610 5715 1630
rect 5685 1605 5715 1610
rect 5685 1550 5715 1555
rect 5685 1530 5690 1550
rect 5690 1530 5710 1550
rect 5710 1530 5715 1550
rect 5685 1525 5715 1530
rect 5685 1470 5715 1475
rect 5685 1450 5690 1470
rect 5690 1450 5710 1470
rect 5710 1450 5715 1470
rect 5685 1445 5715 1450
rect 5685 1390 5715 1395
rect 5685 1370 5690 1390
rect 5690 1370 5710 1390
rect 5710 1370 5715 1390
rect 5685 1365 5715 1370
rect 5685 1310 5715 1315
rect 5685 1290 5690 1310
rect 5690 1290 5710 1310
rect 5710 1290 5715 1310
rect 5685 1285 5715 1290
rect 5685 1230 5715 1235
rect 5685 1210 5690 1230
rect 5690 1210 5710 1230
rect 5710 1210 5715 1230
rect 5685 1205 5715 1210
rect 5685 1150 5715 1155
rect 5685 1130 5690 1150
rect 5690 1130 5710 1150
rect 5710 1130 5715 1150
rect 5685 1125 5715 1130
rect 5685 1070 5715 1075
rect 5685 1050 5690 1070
rect 5690 1050 5710 1070
rect 5710 1050 5715 1070
rect 5685 1045 5715 1050
rect 5685 990 5715 995
rect 5685 970 5690 990
rect 5690 970 5710 990
rect 5710 970 5715 990
rect 5685 965 5715 970
rect 5685 830 5715 835
rect 5685 810 5690 830
rect 5690 810 5710 830
rect 5710 810 5715 830
rect 5685 805 5715 810
rect 5685 750 5715 755
rect 5685 730 5690 750
rect 5690 730 5710 750
rect 5710 730 5715 750
rect 5685 725 5715 730
rect 5685 670 5715 675
rect 5685 650 5690 670
rect 5690 650 5710 670
rect 5710 650 5715 670
rect 5685 645 5715 650
rect 5685 590 5715 595
rect 5685 570 5690 590
rect 5690 570 5710 590
rect 5710 570 5715 590
rect 5685 565 5715 570
rect 5685 510 5715 515
rect 5685 490 5690 510
rect 5690 490 5710 510
rect 5710 490 5715 510
rect 5685 485 5715 490
rect 5685 270 5715 275
rect 5685 250 5690 270
rect 5690 250 5710 270
rect 5710 250 5715 270
rect 5685 245 5715 250
rect 5685 190 5715 195
rect 5685 170 5690 190
rect 5690 170 5710 190
rect 5710 170 5715 190
rect 5685 165 5715 170
rect 5685 110 5715 115
rect 5685 90 5690 110
rect 5690 90 5710 110
rect 5710 90 5715 110
rect 5685 85 5715 90
rect 5685 30 5715 35
rect 5685 10 5690 30
rect 5690 10 5710 30
rect 5710 10 5715 30
rect 5685 5 5715 10
rect 5765 15710 5795 15715
rect 5765 15690 5770 15710
rect 5770 15690 5790 15710
rect 5790 15690 5795 15710
rect 5765 15685 5795 15690
rect 5765 15630 5795 15635
rect 5765 15610 5770 15630
rect 5770 15610 5790 15630
rect 5790 15610 5795 15630
rect 5765 15605 5795 15610
rect 5765 15550 5795 15555
rect 5765 15530 5770 15550
rect 5770 15530 5790 15550
rect 5790 15530 5795 15550
rect 5765 15525 5795 15530
rect 5765 15470 5795 15475
rect 5765 15450 5770 15470
rect 5770 15450 5790 15470
rect 5790 15450 5795 15470
rect 5765 15445 5795 15450
rect 5765 15390 5795 15395
rect 5765 15370 5770 15390
rect 5770 15370 5790 15390
rect 5790 15370 5795 15390
rect 5765 15365 5795 15370
rect 5765 15310 5795 15315
rect 5765 15290 5770 15310
rect 5770 15290 5790 15310
rect 5790 15290 5795 15310
rect 5765 15285 5795 15290
rect 5765 15230 5795 15235
rect 5765 15210 5770 15230
rect 5770 15210 5790 15230
rect 5790 15210 5795 15230
rect 5765 15205 5795 15210
rect 5765 15150 5795 15155
rect 5765 15130 5770 15150
rect 5770 15130 5790 15150
rect 5790 15130 5795 15150
rect 5765 15125 5795 15130
rect 5765 14990 5795 14995
rect 5765 14970 5770 14990
rect 5770 14970 5790 14990
rect 5790 14970 5795 14990
rect 5765 14965 5795 14970
rect 5765 14910 5795 14915
rect 5765 14890 5770 14910
rect 5770 14890 5790 14910
rect 5790 14890 5795 14910
rect 5765 14885 5795 14890
rect 5765 14830 5795 14835
rect 5765 14810 5770 14830
rect 5770 14810 5790 14830
rect 5790 14810 5795 14830
rect 5765 14805 5795 14810
rect 5765 14750 5795 14755
rect 5765 14730 5770 14750
rect 5770 14730 5790 14750
rect 5790 14730 5795 14750
rect 5765 14725 5795 14730
rect 5765 14670 5795 14675
rect 5765 14650 5770 14670
rect 5770 14650 5790 14670
rect 5790 14650 5795 14670
rect 5765 14645 5795 14650
rect 5765 14590 5795 14595
rect 5765 14570 5770 14590
rect 5770 14570 5790 14590
rect 5790 14570 5795 14590
rect 5765 14565 5795 14570
rect 5765 14510 5795 14515
rect 5765 14490 5770 14510
rect 5770 14490 5790 14510
rect 5790 14490 5795 14510
rect 5765 14485 5795 14490
rect 5765 14430 5795 14435
rect 5765 14410 5770 14430
rect 5770 14410 5790 14430
rect 5790 14410 5795 14430
rect 5765 14405 5795 14410
rect 5765 14030 5795 14035
rect 5765 14010 5770 14030
rect 5770 14010 5790 14030
rect 5790 14010 5795 14030
rect 5765 14005 5795 14010
rect 5765 13950 5795 13955
rect 5765 13930 5770 13950
rect 5770 13930 5790 13950
rect 5790 13930 5795 13950
rect 5765 13925 5795 13930
rect 5765 13870 5795 13875
rect 5765 13850 5770 13870
rect 5770 13850 5790 13870
rect 5790 13850 5795 13870
rect 5765 13845 5795 13850
rect 5765 13790 5795 13795
rect 5765 13770 5770 13790
rect 5770 13770 5790 13790
rect 5790 13770 5795 13790
rect 5765 13765 5795 13770
rect 5765 13710 5795 13715
rect 5765 13690 5770 13710
rect 5770 13690 5790 13710
rect 5790 13690 5795 13710
rect 5765 13685 5795 13690
rect 5765 13630 5795 13635
rect 5765 13610 5770 13630
rect 5770 13610 5790 13630
rect 5790 13610 5795 13630
rect 5765 13605 5795 13610
rect 5765 13550 5795 13555
rect 5765 13530 5770 13550
rect 5770 13530 5790 13550
rect 5790 13530 5795 13550
rect 5765 13525 5795 13530
rect 5765 13470 5795 13475
rect 5765 13450 5770 13470
rect 5770 13450 5790 13470
rect 5790 13450 5795 13470
rect 5765 13445 5795 13450
rect 5765 13070 5795 13075
rect 5765 13050 5770 13070
rect 5770 13050 5790 13070
rect 5790 13050 5795 13070
rect 5765 13045 5795 13050
rect 5765 12990 5795 12995
rect 5765 12970 5770 12990
rect 5770 12970 5790 12990
rect 5790 12970 5795 12990
rect 5765 12965 5795 12970
rect 5765 12910 5795 12915
rect 5765 12890 5770 12910
rect 5770 12890 5790 12910
rect 5790 12890 5795 12910
rect 5765 12885 5795 12890
rect 5765 12830 5795 12835
rect 5765 12810 5770 12830
rect 5770 12810 5790 12830
rect 5790 12810 5795 12830
rect 5765 12805 5795 12810
rect 5765 12750 5795 12755
rect 5765 12730 5770 12750
rect 5770 12730 5790 12750
rect 5790 12730 5795 12750
rect 5765 12725 5795 12730
rect 5765 12670 5795 12675
rect 5765 12650 5770 12670
rect 5770 12650 5790 12670
rect 5790 12650 5795 12670
rect 5765 12645 5795 12650
rect 5765 12590 5795 12595
rect 5765 12570 5770 12590
rect 5770 12570 5790 12590
rect 5790 12570 5795 12590
rect 5765 12565 5795 12570
rect 5765 12510 5795 12515
rect 5765 12490 5770 12510
rect 5770 12490 5790 12510
rect 5790 12490 5795 12510
rect 5765 12485 5795 12490
rect 5765 12350 5795 12355
rect 5765 12330 5770 12350
rect 5770 12330 5790 12350
rect 5790 12330 5795 12350
rect 5765 12325 5795 12330
rect 5765 12270 5795 12275
rect 5765 12250 5770 12270
rect 5770 12250 5790 12270
rect 5790 12250 5795 12270
rect 5765 12245 5795 12250
rect 5765 12190 5795 12195
rect 5765 12170 5770 12190
rect 5770 12170 5790 12190
rect 5790 12170 5795 12190
rect 5765 12165 5795 12170
rect 5765 12110 5795 12115
rect 5765 12090 5770 12110
rect 5770 12090 5790 12110
rect 5790 12090 5795 12110
rect 5765 12085 5795 12090
rect 5765 12030 5795 12035
rect 5765 12010 5770 12030
rect 5770 12010 5790 12030
rect 5790 12010 5795 12030
rect 5765 12005 5795 12010
rect 5765 11950 5795 11955
rect 5765 11930 5770 11950
rect 5770 11930 5790 11950
rect 5790 11930 5795 11950
rect 5765 11925 5795 11930
rect 5765 11870 5795 11875
rect 5765 11850 5770 11870
rect 5770 11850 5790 11870
rect 5790 11850 5795 11870
rect 5765 11845 5795 11850
rect 5765 11790 5795 11795
rect 5765 11770 5770 11790
rect 5770 11770 5790 11790
rect 5790 11770 5795 11790
rect 5765 11765 5795 11770
rect 5765 11710 5795 11715
rect 5765 11690 5770 11710
rect 5770 11690 5790 11710
rect 5790 11690 5795 11710
rect 5765 11685 5795 11690
rect 5765 11630 5795 11635
rect 5765 11610 5770 11630
rect 5770 11610 5790 11630
rect 5790 11610 5795 11630
rect 5765 11605 5795 11610
rect 5765 11550 5795 11555
rect 5765 11530 5770 11550
rect 5770 11530 5790 11550
rect 5790 11530 5795 11550
rect 5765 11525 5795 11530
rect 5765 11470 5795 11475
rect 5765 11450 5770 11470
rect 5770 11450 5790 11470
rect 5790 11450 5795 11470
rect 5765 11445 5795 11450
rect 5765 11390 5795 11395
rect 5765 11370 5770 11390
rect 5770 11370 5790 11390
rect 5790 11370 5795 11390
rect 5765 11365 5795 11370
rect 5765 11310 5795 11315
rect 5765 11290 5770 11310
rect 5770 11290 5790 11310
rect 5790 11290 5795 11310
rect 5765 11285 5795 11290
rect 5765 11230 5795 11235
rect 5765 11210 5770 11230
rect 5770 11210 5790 11230
rect 5790 11210 5795 11230
rect 5765 11205 5795 11210
rect 5765 11150 5795 11155
rect 5765 11130 5770 11150
rect 5770 11130 5790 11150
rect 5790 11130 5795 11150
rect 5765 11125 5795 11130
rect 5765 11070 5795 11075
rect 5765 11050 5770 11070
rect 5770 11050 5790 11070
rect 5790 11050 5795 11070
rect 5765 11045 5795 11050
rect 5765 10910 5795 10915
rect 5765 10890 5770 10910
rect 5770 10890 5790 10910
rect 5790 10890 5795 10910
rect 5765 10885 5795 10890
rect 5765 10830 5795 10835
rect 5765 10810 5770 10830
rect 5770 10810 5790 10830
rect 5790 10810 5795 10830
rect 5765 10805 5795 10810
rect 5765 10750 5795 10755
rect 5765 10730 5770 10750
rect 5770 10730 5790 10750
rect 5790 10730 5795 10750
rect 5765 10725 5795 10730
rect 5765 10670 5795 10675
rect 5765 10650 5770 10670
rect 5770 10650 5790 10670
rect 5790 10650 5795 10670
rect 5765 10645 5795 10650
rect 5765 10590 5795 10595
rect 5765 10570 5770 10590
rect 5770 10570 5790 10590
rect 5790 10570 5795 10590
rect 5765 10565 5795 10570
rect 5765 10510 5795 10515
rect 5765 10490 5770 10510
rect 5770 10490 5790 10510
rect 5790 10490 5795 10510
rect 5765 10485 5795 10490
rect 5765 10430 5795 10435
rect 5765 10410 5770 10430
rect 5770 10410 5790 10430
rect 5790 10410 5795 10430
rect 5765 10405 5795 10410
rect 5765 10350 5795 10355
rect 5765 10330 5770 10350
rect 5770 10330 5790 10350
rect 5790 10330 5795 10350
rect 5765 10325 5795 10330
rect 5765 9950 5795 9955
rect 5765 9930 5770 9950
rect 5770 9930 5790 9950
rect 5790 9930 5795 9950
rect 5765 9925 5795 9930
rect 5765 9870 5795 9875
rect 5765 9850 5770 9870
rect 5770 9850 5790 9870
rect 5790 9850 5795 9870
rect 5765 9845 5795 9850
rect 5765 9790 5795 9795
rect 5765 9770 5770 9790
rect 5770 9770 5790 9790
rect 5790 9770 5795 9790
rect 5765 9765 5795 9770
rect 5765 9710 5795 9715
rect 5765 9690 5770 9710
rect 5770 9690 5790 9710
rect 5790 9690 5795 9710
rect 5765 9685 5795 9690
rect 5765 9630 5795 9635
rect 5765 9610 5770 9630
rect 5770 9610 5790 9630
rect 5790 9610 5795 9630
rect 5765 9605 5795 9610
rect 5765 9550 5795 9555
rect 5765 9530 5770 9550
rect 5770 9530 5790 9550
rect 5790 9530 5795 9550
rect 5765 9525 5795 9530
rect 5765 9470 5795 9475
rect 5765 9450 5770 9470
rect 5770 9450 5790 9470
rect 5790 9450 5795 9470
rect 5765 9445 5795 9450
rect 5765 9390 5795 9395
rect 5765 9370 5770 9390
rect 5770 9370 5790 9390
rect 5790 9370 5795 9390
rect 5765 9365 5795 9370
rect 5765 8990 5795 8995
rect 5765 8970 5770 8990
rect 5770 8970 5790 8990
rect 5790 8970 5795 8990
rect 5765 8965 5795 8970
rect 5765 8910 5795 8915
rect 5765 8890 5770 8910
rect 5770 8890 5790 8910
rect 5790 8890 5795 8910
rect 5765 8885 5795 8890
rect 5765 8830 5795 8835
rect 5765 8810 5770 8830
rect 5770 8810 5790 8830
rect 5790 8810 5795 8830
rect 5765 8805 5795 8810
rect 5765 8750 5795 8755
rect 5765 8730 5770 8750
rect 5770 8730 5790 8750
rect 5790 8730 5795 8750
rect 5765 8725 5795 8730
rect 5765 8670 5795 8675
rect 5765 8650 5770 8670
rect 5770 8650 5790 8670
rect 5790 8650 5795 8670
rect 5765 8645 5795 8650
rect 5765 8590 5795 8595
rect 5765 8570 5770 8590
rect 5770 8570 5790 8590
rect 5790 8570 5795 8590
rect 5765 8565 5795 8570
rect 5765 8510 5795 8515
rect 5765 8490 5770 8510
rect 5770 8490 5790 8510
rect 5790 8490 5795 8510
rect 5765 8485 5795 8490
rect 5765 8430 5795 8435
rect 5765 8410 5770 8430
rect 5770 8410 5790 8430
rect 5790 8410 5795 8430
rect 5765 8405 5795 8410
rect 5765 8270 5795 8275
rect 5765 8250 5770 8270
rect 5770 8250 5790 8270
rect 5790 8250 5795 8270
rect 5765 8245 5795 8250
rect 5765 8190 5795 8195
rect 5765 8170 5770 8190
rect 5770 8170 5790 8190
rect 5790 8170 5795 8190
rect 5765 8165 5795 8170
rect 5765 8110 5795 8115
rect 5765 8090 5770 8110
rect 5770 8090 5790 8110
rect 5790 8090 5795 8110
rect 5765 8085 5795 8090
rect 5765 8030 5795 8035
rect 5765 8010 5770 8030
rect 5770 8010 5790 8030
rect 5790 8010 5795 8030
rect 5765 8005 5795 8010
rect 5765 7950 5795 7955
rect 5765 7930 5770 7950
rect 5770 7930 5790 7950
rect 5790 7930 5795 7950
rect 5765 7925 5795 7930
rect 5765 7870 5795 7875
rect 5765 7850 5770 7870
rect 5770 7850 5790 7870
rect 5790 7850 5795 7870
rect 5765 7845 5795 7850
rect 5765 7790 5795 7795
rect 5765 7770 5770 7790
rect 5770 7770 5790 7790
rect 5790 7770 5795 7790
rect 5765 7765 5795 7770
rect 5765 7710 5795 7715
rect 5765 7690 5770 7710
rect 5770 7690 5790 7710
rect 5790 7690 5795 7710
rect 5765 7685 5795 7690
rect 5765 7630 5795 7635
rect 5765 7610 5770 7630
rect 5770 7610 5790 7630
rect 5790 7610 5795 7630
rect 5765 7605 5795 7610
rect 5765 7550 5795 7555
rect 5765 7530 5770 7550
rect 5770 7530 5790 7550
rect 5790 7530 5795 7550
rect 5765 7525 5795 7530
rect 5765 7470 5795 7475
rect 5765 7450 5770 7470
rect 5770 7450 5790 7470
rect 5790 7450 5795 7470
rect 5765 7445 5795 7450
rect 5765 7390 5795 7395
rect 5765 7370 5770 7390
rect 5770 7370 5790 7390
rect 5790 7370 5795 7390
rect 5765 7365 5795 7370
rect 5765 7310 5795 7315
rect 5765 7290 5770 7310
rect 5770 7290 5790 7310
rect 5790 7290 5795 7310
rect 5765 7285 5795 7290
rect 5765 7230 5795 7235
rect 5765 7210 5770 7230
rect 5770 7210 5790 7230
rect 5790 7210 5795 7230
rect 5765 7205 5795 7210
rect 5765 7150 5795 7155
rect 5765 7130 5770 7150
rect 5770 7130 5790 7150
rect 5790 7130 5795 7150
rect 5765 7125 5795 7130
rect 5765 7070 5795 7075
rect 5765 7050 5770 7070
rect 5770 7050 5790 7070
rect 5790 7050 5795 7070
rect 5765 7045 5795 7050
rect 5765 6990 5795 6995
rect 5765 6970 5770 6990
rect 5770 6970 5790 6990
rect 5790 6970 5795 6990
rect 5765 6965 5795 6970
rect 5765 6830 5795 6835
rect 5765 6810 5770 6830
rect 5770 6810 5790 6830
rect 5790 6810 5795 6830
rect 5765 6805 5795 6810
rect 5765 6750 5795 6755
rect 5765 6730 5770 6750
rect 5770 6730 5790 6750
rect 5790 6730 5795 6750
rect 5765 6725 5795 6730
rect 5765 6670 5795 6675
rect 5765 6650 5770 6670
rect 5770 6650 5790 6670
rect 5790 6650 5795 6670
rect 5765 6645 5795 6650
rect 5765 6590 5795 6595
rect 5765 6570 5770 6590
rect 5770 6570 5790 6590
rect 5790 6570 5795 6590
rect 5765 6565 5795 6570
rect 5765 6510 5795 6515
rect 5765 6490 5770 6510
rect 5770 6490 5790 6510
rect 5790 6490 5795 6510
rect 5765 6485 5795 6490
rect 5765 6430 5795 6435
rect 5765 6410 5770 6430
rect 5770 6410 5790 6430
rect 5790 6410 5795 6430
rect 5765 6405 5795 6410
rect 5765 6350 5795 6355
rect 5765 6330 5770 6350
rect 5770 6330 5790 6350
rect 5790 6330 5795 6350
rect 5765 6325 5795 6330
rect 5765 6270 5795 6275
rect 5765 6250 5770 6270
rect 5770 6250 5790 6270
rect 5790 6250 5795 6270
rect 5765 6245 5795 6250
rect 5765 5870 5795 5875
rect 5765 5850 5770 5870
rect 5770 5850 5790 5870
rect 5790 5850 5795 5870
rect 5765 5845 5795 5850
rect 5765 5790 5795 5795
rect 5765 5770 5770 5790
rect 5770 5770 5790 5790
rect 5790 5770 5795 5790
rect 5765 5765 5795 5770
rect 5765 5710 5795 5715
rect 5765 5690 5770 5710
rect 5770 5690 5790 5710
rect 5790 5690 5795 5710
rect 5765 5685 5795 5690
rect 5765 5630 5795 5635
rect 5765 5610 5770 5630
rect 5770 5610 5790 5630
rect 5790 5610 5795 5630
rect 5765 5605 5795 5610
rect 5765 5550 5795 5555
rect 5765 5530 5770 5550
rect 5770 5530 5790 5550
rect 5790 5530 5795 5550
rect 5765 5525 5795 5530
rect 5765 5470 5795 5475
rect 5765 5450 5770 5470
rect 5770 5450 5790 5470
rect 5790 5450 5795 5470
rect 5765 5445 5795 5450
rect 5765 5390 5795 5395
rect 5765 5370 5770 5390
rect 5770 5370 5790 5390
rect 5790 5370 5795 5390
rect 5765 5365 5795 5370
rect 5765 5310 5795 5315
rect 5765 5290 5770 5310
rect 5770 5290 5790 5310
rect 5790 5290 5795 5310
rect 5765 5285 5795 5290
rect 5765 5230 5795 5235
rect 5765 5210 5770 5230
rect 5770 5210 5790 5230
rect 5790 5210 5795 5230
rect 5765 5205 5795 5210
rect 5765 5150 5795 5155
rect 5765 5130 5770 5150
rect 5770 5130 5790 5150
rect 5790 5130 5795 5150
rect 5765 5125 5795 5130
rect 5765 5070 5795 5075
rect 5765 5050 5770 5070
rect 5770 5050 5790 5070
rect 5790 5050 5795 5070
rect 5765 5045 5795 5050
rect 5765 4990 5795 4995
rect 5765 4970 5770 4990
rect 5770 4970 5790 4990
rect 5790 4970 5795 4990
rect 5765 4965 5795 4970
rect 5765 4910 5795 4915
rect 5765 4890 5770 4910
rect 5770 4890 5790 4910
rect 5790 4890 5795 4910
rect 5765 4885 5795 4890
rect 5765 4750 5795 4755
rect 5765 4730 5770 4750
rect 5770 4730 5790 4750
rect 5790 4730 5795 4750
rect 5765 4725 5795 4730
rect 5765 4670 5795 4675
rect 5765 4650 5770 4670
rect 5770 4650 5790 4670
rect 5790 4650 5795 4670
rect 5765 4645 5795 4650
rect 5765 4510 5795 4515
rect 5765 4490 5770 4510
rect 5770 4490 5790 4510
rect 5790 4490 5795 4510
rect 5765 4485 5795 4490
rect 5765 4430 5795 4435
rect 5765 4410 5770 4430
rect 5770 4410 5790 4430
rect 5790 4410 5795 4430
rect 5765 4405 5795 4410
rect 5765 4350 5795 4355
rect 5765 4330 5770 4350
rect 5770 4330 5790 4350
rect 5790 4330 5795 4350
rect 5765 4325 5795 4330
rect 5765 4270 5795 4275
rect 5765 4250 5770 4270
rect 5770 4250 5790 4270
rect 5790 4250 5795 4270
rect 5765 4245 5795 4250
rect 5765 4190 5795 4195
rect 5765 4170 5770 4190
rect 5770 4170 5790 4190
rect 5790 4170 5795 4190
rect 5765 4165 5795 4170
rect 5765 4110 5795 4115
rect 5765 4090 5770 4110
rect 5770 4090 5790 4110
rect 5790 4090 5795 4110
rect 5765 4085 5795 4090
rect 5765 4030 5795 4035
rect 5765 4010 5770 4030
rect 5770 4010 5790 4030
rect 5790 4010 5795 4030
rect 5765 4005 5795 4010
rect 5765 3950 5795 3955
rect 5765 3930 5770 3950
rect 5770 3930 5790 3950
rect 5790 3930 5795 3950
rect 5765 3925 5795 3930
rect 5765 3870 5795 3875
rect 5765 3850 5770 3870
rect 5770 3850 5790 3870
rect 5790 3850 5795 3870
rect 5765 3845 5795 3850
rect 5765 3710 5795 3715
rect 5765 3690 5770 3710
rect 5770 3690 5790 3710
rect 5790 3690 5795 3710
rect 5765 3685 5795 3690
rect 5765 3630 5795 3635
rect 5765 3610 5770 3630
rect 5770 3610 5790 3630
rect 5790 3610 5795 3630
rect 5765 3605 5795 3610
rect 5765 3470 5795 3475
rect 5765 3450 5770 3470
rect 5770 3450 5790 3470
rect 5790 3450 5795 3470
rect 5765 3445 5795 3450
rect 5765 3390 5795 3395
rect 5765 3370 5770 3390
rect 5770 3370 5790 3390
rect 5790 3370 5795 3390
rect 5765 3365 5795 3370
rect 5765 3230 5795 3235
rect 5765 3210 5770 3230
rect 5770 3210 5790 3230
rect 5790 3210 5795 3230
rect 5765 3205 5795 3210
rect 5765 3150 5795 3155
rect 5765 3130 5770 3150
rect 5770 3130 5790 3150
rect 5790 3130 5795 3150
rect 5765 3125 5795 3130
rect 5765 3070 5795 3075
rect 5765 3050 5770 3070
rect 5770 3050 5790 3070
rect 5790 3050 5795 3070
rect 5765 3045 5795 3050
rect 5765 2990 5795 2995
rect 5765 2970 5770 2990
rect 5770 2970 5790 2990
rect 5790 2970 5795 2990
rect 5765 2965 5795 2970
rect 5765 2910 5795 2915
rect 5765 2890 5770 2910
rect 5770 2890 5790 2910
rect 5790 2890 5795 2910
rect 5765 2885 5795 2890
rect 5765 2830 5795 2835
rect 5765 2810 5770 2830
rect 5770 2810 5790 2830
rect 5790 2810 5795 2830
rect 5765 2805 5795 2810
rect 5765 2750 5795 2755
rect 5765 2730 5770 2750
rect 5770 2730 5790 2750
rect 5790 2730 5795 2750
rect 5765 2725 5795 2730
rect 5765 2670 5795 2675
rect 5765 2650 5770 2670
rect 5770 2650 5790 2670
rect 5790 2650 5795 2670
rect 5765 2645 5795 2650
rect 5765 2590 5795 2595
rect 5765 2570 5770 2590
rect 5770 2570 5790 2590
rect 5790 2570 5795 2590
rect 5765 2565 5795 2570
rect 5765 2510 5795 2515
rect 5765 2490 5770 2510
rect 5770 2490 5790 2510
rect 5790 2490 5795 2510
rect 5765 2485 5795 2490
rect 5765 2430 5795 2435
rect 5765 2410 5770 2430
rect 5770 2410 5790 2430
rect 5790 2410 5795 2430
rect 5765 2405 5795 2410
rect 5765 2350 5795 2355
rect 5765 2330 5770 2350
rect 5770 2330 5790 2350
rect 5790 2330 5795 2350
rect 5765 2325 5795 2330
rect 5765 2270 5795 2275
rect 5765 2250 5770 2270
rect 5770 2250 5790 2270
rect 5790 2250 5795 2270
rect 5765 2245 5795 2250
rect 5765 2190 5795 2195
rect 5765 2170 5770 2190
rect 5770 2170 5790 2190
rect 5790 2170 5795 2190
rect 5765 2165 5795 2170
rect 5765 2110 5795 2115
rect 5765 2090 5770 2110
rect 5770 2090 5790 2110
rect 5790 2090 5795 2110
rect 5765 2085 5795 2090
rect 5765 2030 5795 2035
rect 5765 2010 5770 2030
rect 5770 2010 5790 2030
rect 5790 2010 5795 2030
rect 5765 2005 5795 2010
rect 5765 1950 5795 1955
rect 5765 1930 5770 1950
rect 5770 1930 5790 1950
rect 5790 1930 5795 1950
rect 5765 1925 5795 1930
rect 5765 1710 5795 1715
rect 5765 1690 5770 1710
rect 5770 1690 5790 1710
rect 5790 1690 5795 1710
rect 5765 1685 5795 1690
rect 5765 1630 5795 1635
rect 5765 1610 5770 1630
rect 5770 1610 5790 1630
rect 5790 1610 5795 1630
rect 5765 1605 5795 1610
rect 5765 1550 5795 1555
rect 5765 1530 5770 1550
rect 5770 1530 5790 1550
rect 5790 1530 5795 1550
rect 5765 1525 5795 1530
rect 5765 1470 5795 1475
rect 5765 1450 5770 1470
rect 5770 1450 5790 1470
rect 5790 1450 5795 1470
rect 5765 1445 5795 1450
rect 5765 1390 5795 1395
rect 5765 1370 5770 1390
rect 5770 1370 5790 1390
rect 5790 1370 5795 1390
rect 5765 1365 5795 1370
rect 5765 1310 5795 1315
rect 5765 1290 5770 1310
rect 5770 1290 5790 1310
rect 5790 1290 5795 1310
rect 5765 1285 5795 1290
rect 5765 1230 5795 1235
rect 5765 1210 5770 1230
rect 5770 1210 5790 1230
rect 5790 1210 5795 1230
rect 5765 1205 5795 1210
rect 5765 1150 5795 1155
rect 5765 1130 5770 1150
rect 5770 1130 5790 1150
rect 5790 1130 5795 1150
rect 5765 1125 5795 1130
rect 5765 1070 5795 1075
rect 5765 1050 5770 1070
rect 5770 1050 5790 1070
rect 5790 1050 5795 1070
rect 5765 1045 5795 1050
rect 5765 990 5795 995
rect 5765 970 5770 990
rect 5770 970 5790 990
rect 5790 970 5795 990
rect 5765 965 5795 970
rect 5765 830 5795 835
rect 5765 810 5770 830
rect 5770 810 5790 830
rect 5790 810 5795 830
rect 5765 805 5795 810
rect 5765 750 5795 755
rect 5765 730 5770 750
rect 5770 730 5790 750
rect 5790 730 5795 750
rect 5765 725 5795 730
rect 5765 670 5795 675
rect 5765 650 5770 670
rect 5770 650 5790 670
rect 5790 650 5795 670
rect 5765 645 5795 650
rect 5765 590 5795 595
rect 5765 570 5770 590
rect 5770 570 5790 590
rect 5790 570 5795 590
rect 5765 565 5795 570
rect 5765 510 5795 515
rect 5765 490 5770 510
rect 5770 490 5790 510
rect 5790 490 5795 510
rect 5765 485 5795 490
rect 5765 270 5795 275
rect 5765 250 5770 270
rect 5770 250 5790 270
rect 5790 250 5795 270
rect 5765 245 5795 250
rect 5765 190 5795 195
rect 5765 170 5770 190
rect 5770 170 5790 190
rect 5790 170 5795 190
rect 5765 165 5795 170
rect 5765 110 5795 115
rect 5765 90 5770 110
rect 5770 90 5790 110
rect 5790 90 5795 110
rect 5765 85 5795 90
rect 5765 30 5795 35
rect 5765 10 5770 30
rect 5770 10 5790 30
rect 5790 10 5795 30
rect 5765 5 5795 10
rect 5925 15710 5955 15715
rect 5925 15690 5930 15710
rect 5930 15690 5950 15710
rect 5950 15690 5955 15710
rect 5925 15685 5955 15690
rect 5925 15630 5955 15635
rect 5925 15610 5930 15630
rect 5930 15610 5950 15630
rect 5950 15610 5955 15630
rect 5925 15605 5955 15610
rect 5925 15550 5955 15555
rect 5925 15530 5930 15550
rect 5930 15530 5950 15550
rect 5950 15530 5955 15550
rect 5925 15525 5955 15530
rect 5925 15470 5955 15475
rect 5925 15450 5930 15470
rect 5930 15450 5950 15470
rect 5950 15450 5955 15470
rect 5925 15445 5955 15450
rect 5925 15390 5955 15395
rect 5925 15370 5930 15390
rect 5930 15370 5950 15390
rect 5950 15370 5955 15390
rect 5925 15365 5955 15370
rect 5925 15310 5955 15315
rect 5925 15290 5930 15310
rect 5930 15290 5950 15310
rect 5950 15290 5955 15310
rect 5925 15285 5955 15290
rect 5925 15230 5955 15235
rect 5925 15210 5930 15230
rect 5930 15210 5950 15230
rect 5950 15210 5955 15230
rect 5925 15205 5955 15210
rect 5925 15150 5955 15155
rect 5925 15130 5930 15150
rect 5930 15130 5950 15150
rect 5950 15130 5955 15150
rect 5925 15125 5955 15130
rect 5925 14990 5955 14995
rect 5925 14970 5930 14990
rect 5930 14970 5950 14990
rect 5950 14970 5955 14990
rect 5925 14965 5955 14970
rect 5925 14910 5955 14915
rect 5925 14890 5930 14910
rect 5930 14890 5950 14910
rect 5950 14890 5955 14910
rect 5925 14885 5955 14890
rect 5925 14830 5955 14835
rect 5925 14810 5930 14830
rect 5930 14810 5950 14830
rect 5950 14810 5955 14830
rect 5925 14805 5955 14810
rect 5925 14750 5955 14755
rect 5925 14730 5930 14750
rect 5930 14730 5950 14750
rect 5950 14730 5955 14750
rect 5925 14725 5955 14730
rect 5925 14670 5955 14675
rect 5925 14650 5930 14670
rect 5930 14650 5950 14670
rect 5950 14650 5955 14670
rect 5925 14645 5955 14650
rect 5925 14590 5955 14595
rect 5925 14570 5930 14590
rect 5930 14570 5950 14590
rect 5950 14570 5955 14590
rect 5925 14565 5955 14570
rect 5925 14510 5955 14515
rect 5925 14490 5930 14510
rect 5930 14490 5950 14510
rect 5950 14490 5955 14510
rect 5925 14485 5955 14490
rect 5925 14430 5955 14435
rect 5925 14410 5930 14430
rect 5930 14410 5950 14430
rect 5950 14410 5955 14430
rect 5925 14405 5955 14410
rect 5925 14030 5955 14035
rect 5925 14010 5930 14030
rect 5930 14010 5950 14030
rect 5950 14010 5955 14030
rect 5925 14005 5955 14010
rect 5925 13950 5955 13955
rect 5925 13930 5930 13950
rect 5930 13930 5950 13950
rect 5950 13930 5955 13950
rect 5925 13925 5955 13930
rect 5925 13870 5955 13875
rect 5925 13850 5930 13870
rect 5930 13850 5950 13870
rect 5950 13850 5955 13870
rect 5925 13845 5955 13850
rect 5925 13790 5955 13795
rect 5925 13770 5930 13790
rect 5930 13770 5950 13790
rect 5950 13770 5955 13790
rect 5925 13765 5955 13770
rect 5925 13710 5955 13715
rect 5925 13690 5930 13710
rect 5930 13690 5950 13710
rect 5950 13690 5955 13710
rect 5925 13685 5955 13690
rect 5925 13630 5955 13635
rect 5925 13610 5930 13630
rect 5930 13610 5950 13630
rect 5950 13610 5955 13630
rect 5925 13605 5955 13610
rect 5925 13550 5955 13555
rect 5925 13530 5930 13550
rect 5930 13530 5950 13550
rect 5950 13530 5955 13550
rect 5925 13525 5955 13530
rect 5925 13470 5955 13475
rect 5925 13450 5930 13470
rect 5930 13450 5950 13470
rect 5950 13450 5955 13470
rect 5925 13445 5955 13450
rect 5925 13070 5955 13075
rect 5925 13050 5930 13070
rect 5930 13050 5950 13070
rect 5950 13050 5955 13070
rect 5925 13045 5955 13050
rect 5925 12990 5955 12995
rect 5925 12970 5930 12990
rect 5930 12970 5950 12990
rect 5950 12970 5955 12990
rect 5925 12965 5955 12970
rect 5925 12910 5955 12915
rect 5925 12890 5930 12910
rect 5930 12890 5950 12910
rect 5950 12890 5955 12910
rect 5925 12885 5955 12890
rect 5925 12830 5955 12835
rect 5925 12810 5930 12830
rect 5930 12810 5950 12830
rect 5950 12810 5955 12830
rect 5925 12805 5955 12810
rect 5925 12750 5955 12755
rect 5925 12730 5930 12750
rect 5930 12730 5950 12750
rect 5950 12730 5955 12750
rect 5925 12725 5955 12730
rect 5925 12670 5955 12675
rect 5925 12650 5930 12670
rect 5930 12650 5950 12670
rect 5950 12650 5955 12670
rect 5925 12645 5955 12650
rect 5925 12590 5955 12595
rect 5925 12570 5930 12590
rect 5930 12570 5950 12590
rect 5950 12570 5955 12590
rect 5925 12565 5955 12570
rect 5925 12510 5955 12515
rect 5925 12490 5930 12510
rect 5930 12490 5950 12510
rect 5950 12490 5955 12510
rect 5925 12485 5955 12490
rect 5925 12350 5955 12355
rect 5925 12330 5930 12350
rect 5930 12330 5950 12350
rect 5950 12330 5955 12350
rect 5925 12325 5955 12330
rect 5925 12270 5955 12275
rect 5925 12250 5930 12270
rect 5930 12250 5950 12270
rect 5950 12250 5955 12270
rect 5925 12245 5955 12250
rect 5925 12190 5955 12195
rect 5925 12170 5930 12190
rect 5930 12170 5950 12190
rect 5950 12170 5955 12190
rect 5925 12165 5955 12170
rect 5925 12110 5955 12115
rect 5925 12090 5930 12110
rect 5930 12090 5950 12110
rect 5950 12090 5955 12110
rect 5925 12085 5955 12090
rect 5925 12030 5955 12035
rect 5925 12010 5930 12030
rect 5930 12010 5950 12030
rect 5950 12010 5955 12030
rect 5925 12005 5955 12010
rect 5925 11950 5955 11955
rect 5925 11930 5930 11950
rect 5930 11930 5950 11950
rect 5950 11930 5955 11950
rect 5925 11925 5955 11930
rect 5925 11870 5955 11875
rect 5925 11850 5930 11870
rect 5930 11850 5950 11870
rect 5950 11850 5955 11870
rect 5925 11845 5955 11850
rect 5925 11790 5955 11795
rect 5925 11770 5930 11790
rect 5930 11770 5950 11790
rect 5950 11770 5955 11790
rect 5925 11765 5955 11770
rect 5925 11710 5955 11715
rect 5925 11690 5930 11710
rect 5930 11690 5950 11710
rect 5950 11690 5955 11710
rect 5925 11685 5955 11690
rect 5925 11630 5955 11635
rect 5925 11610 5930 11630
rect 5930 11610 5950 11630
rect 5950 11610 5955 11630
rect 5925 11605 5955 11610
rect 5925 11550 5955 11555
rect 5925 11530 5930 11550
rect 5930 11530 5950 11550
rect 5950 11530 5955 11550
rect 5925 11525 5955 11530
rect 5925 11470 5955 11475
rect 5925 11450 5930 11470
rect 5930 11450 5950 11470
rect 5950 11450 5955 11470
rect 5925 11445 5955 11450
rect 5925 11390 5955 11395
rect 5925 11370 5930 11390
rect 5930 11370 5950 11390
rect 5950 11370 5955 11390
rect 5925 11365 5955 11370
rect 5925 11310 5955 11315
rect 5925 11290 5930 11310
rect 5930 11290 5950 11310
rect 5950 11290 5955 11310
rect 5925 11285 5955 11290
rect 5925 11230 5955 11235
rect 5925 11210 5930 11230
rect 5930 11210 5950 11230
rect 5950 11210 5955 11230
rect 5925 11205 5955 11210
rect 5925 11150 5955 11155
rect 5925 11130 5930 11150
rect 5930 11130 5950 11150
rect 5950 11130 5955 11150
rect 5925 11125 5955 11130
rect 5925 11070 5955 11075
rect 5925 11050 5930 11070
rect 5930 11050 5950 11070
rect 5950 11050 5955 11070
rect 5925 11045 5955 11050
rect 5925 10910 5955 10915
rect 5925 10890 5930 10910
rect 5930 10890 5950 10910
rect 5950 10890 5955 10910
rect 5925 10885 5955 10890
rect 5925 10830 5955 10835
rect 5925 10810 5930 10830
rect 5930 10810 5950 10830
rect 5950 10810 5955 10830
rect 5925 10805 5955 10810
rect 5925 10750 5955 10755
rect 5925 10730 5930 10750
rect 5930 10730 5950 10750
rect 5950 10730 5955 10750
rect 5925 10725 5955 10730
rect 5925 10670 5955 10675
rect 5925 10650 5930 10670
rect 5930 10650 5950 10670
rect 5950 10650 5955 10670
rect 5925 10645 5955 10650
rect 5925 10590 5955 10595
rect 5925 10570 5930 10590
rect 5930 10570 5950 10590
rect 5950 10570 5955 10590
rect 5925 10565 5955 10570
rect 5925 10510 5955 10515
rect 5925 10490 5930 10510
rect 5930 10490 5950 10510
rect 5950 10490 5955 10510
rect 5925 10485 5955 10490
rect 5925 10430 5955 10435
rect 5925 10410 5930 10430
rect 5930 10410 5950 10430
rect 5950 10410 5955 10430
rect 5925 10405 5955 10410
rect 5925 10350 5955 10355
rect 5925 10330 5930 10350
rect 5930 10330 5950 10350
rect 5950 10330 5955 10350
rect 5925 10325 5955 10330
rect 5925 9950 5955 9955
rect 5925 9930 5930 9950
rect 5930 9930 5950 9950
rect 5950 9930 5955 9950
rect 5925 9925 5955 9930
rect 5925 9870 5955 9875
rect 5925 9850 5930 9870
rect 5930 9850 5950 9870
rect 5950 9850 5955 9870
rect 5925 9845 5955 9850
rect 5925 9790 5955 9795
rect 5925 9770 5930 9790
rect 5930 9770 5950 9790
rect 5950 9770 5955 9790
rect 5925 9765 5955 9770
rect 5925 9710 5955 9715
rect 5925 9690 5930 9710
rect 5930 9690 5950 9710
rect 5950 9690 5955 9710
rect 5925 9685 5955 9690
rect 5925 9630 5955 9635
rect 5925 9610 5930 9630
rect 5930 9610 5950 9630
rect 5950 9610 5955 9630
rect 5925 9605 5955 9610
rect 5925 9550 5955 9555
rect 5925 9530 5930 9550
rect 5930 9530 5950 9550
rect 5950 9530 5955 9550
rect 5925 9525 5955 9530
rect 5925 9470 5955 9475
rect 5925 9450 5930 9470
rect 5930 9450 5950 9470
rect 5950 9450 5955 9470
rect 5925 9445 5955 9450
rect 5925 9390 5955 9395
rect 5925 9370 5930 9390
rect 5930 9370 5950 9390
rect 5950 9370 5955 9390
rect 5925 9365 5955 9370
rect 5925 8990 5955 8995
rect 5925 8970 5930 8990
rect 5930 8970 5950 8990
rect 5950 8970 5955 8990
rect 5925 8965 5955 8970
rect 5925 8910 5955 8915
rect 5925 8890 5930 8910
rect 5930 8890 5950 8910
rect 5950 8890 5955 8910
rect 5925 8885 5955 8890
rect 5925 8830 5955 8835
rect 5925 8810 5930 8830
rect 5930 8810 5950 8830
rect 5950 8810 5955 8830
rect 5925 8805 5955 8810
rect 5925 8750 5955 8755
rect 5925 8730 5930 8750
rect 5930 8730 5950 8750
rect 5950 8730 5955 8750
rect 5925 8725 5955 8730
rect 5925 8670 5955 8675
rect 5925 8650 5930 8670
rect 5930 8650 5950 8670
rect 5950 8650 5955 8670
rect 5925 8645 5955 8650
rect 5925 8590 5955 8595
rect 5925 8570 5930 8590
rect 5930 8570 5950 8590
rect 5950 8570 5955 8590
rect 5925 8565 5955 8570
rect 5925 8510 5955 8515
rect 5925 8490 5930 8510
rect 5930 8490 5950 8510
rect 5950 8490 5955 8510
rect 5925 8485 5955 8490
rect 5925 8430 5955 8435
rect 5925 8410 5930 8430
rect 5930 8410 5950 8430
rect 5950 8410 5955 8430
rect 5925 8405 5955 8410
rect 5925 8270 5955 8275
rect 5925 8250 5930 8270
rect 5930 8250 5950 8270
rect 5950 8250 5955 8270
rect 5925 8245 5955 8250
rect 5925 8190 5955 8195
rect 5925 8170 5930 8190
rect 5930 8170 5950 8190
rect 5950 8170 5955 8190
rect 5925 8165 5955 8170
rect 5925 8110 5955 8115
rect 5925 8090 5930 8110
rect 5930 8090 5950 8110
rect 5950 8090 5955 8110
rect 5925 8085 5955 8090
rect 5925 8030 5955 8035
rect 5925 8010 5930 8030
rect 5930 8010 5950 8030
rect 5950 8010 5955 8030
rect 5925 8005 5955 8010
rect 5925 7950 5955 7955
rect 5925 7930 5930 7950
rect 5930 7930 5950 7950
rect 5950 7930 5955 7950
rect 5925 7925 5955 7930
rect 5925 7870 5955 7875
rect 5925 7850 5930 7870
rect 5930 7850 5950 7870
rect 5950 7850 5955 7870
rect 5925 7845 5955 7850
rect 5925 7790 5955 7795
rect 5925 7770 5930 7790
rect 5930 7770 5950 7790
rect 5950 7770 5955 7790
rect 5925 7765 5955 7770
rect 5925 7710 5955 7715
rect 5925 7690 5930 7710
rect 5930 7690 5950 7710
rect 5950 7690 5955 7710
rect 5925 7685 5955 7690
rect 5925 7630 5955 7635
rect 5925 7610 5930 7630
rect 5930 7610 5950 7630
rect 5950 7610 5955 7630
rect 5925 7605 5955 7610
rect 5925 7550 5955 7555
rect 5925 7530 5930 7550
rect 5930 7530 5950 7550
rect 5950 7530 5955 7550
rect 5925 7525 5955 7530
rect 5925 7470 5955 7475
rect 5925 7450 5930 7470
rect 5930 7450 5950 7470
rect 5950 7450 5955 7470
rect 5925 7445 5955 7450
rect 5925 7390 5955 7395
rect 5925 7370 5930 7390
rect 5930 7370 5950 7390
rect 5950 7370 5955 7390
rect 5925 7365 5955 7370
rect 5925 7310 5955 7315
rect 5925 7290 5930 7310
rect 5930 7290 5950 7310
rect 5950 7290 5955 7310
rect 5925 7285 5955 7290
rect 5925 7230 5955 7235
rect 5925 7210 5930 7230
rect 5930 7210 5950 7230
rect 5950 7210 5955 7230
rect 5925 7205 5955 7210
rect 5925 7150 5955 7155
rect 5925 7130 5930 7150
rect 5930 7130 5950 7150
rect 5950 7130 5955 7150
rect 5925 7125 5955 7130
rect 5925 7070 5955 7075
rect 5925 7050 5930 7070
rect 5930 7050 5950 7070
rect 5950 7050 5955 7070
rect 5925 7045 5955 7050
rect 5925 6990 5955 6995
rect 5925 6970 5930 6990
rect 5930 6970 5950 6990
rect 5950 6970 5955 6990
rect 5925 6965 5955 6970
rect 5925 6830 5955 6835
rect 5925 6810 5930 6830
rect 5930 6810 5950 6830
rect 5950 6810 5955 6830
rect 5925 6805 5955 6810
rect 5925 6750 5955 6755
rect 5925 6730 5930 6750
rect 5930 6730 5950 6750
rect 5950 6730 5955 6750
rect 5925 6725 5955 6730
rect 5925 6670 5955 6675
rect 5925 6650 5930 6670
rect 5930 6650 5950 6670
rect 5950 6650 5955 6670
rect 5925 6645 5955 6650
rect 5925 6590 5955 6595
rect 5925 6570 5930 6590
rect 5930 6570 5950 6590
rect 5950 6570 5955 6590
rect 5925 6565 5955 6570
rect 5925 6510 5955 6515
rect 5925 6490 5930 6510
rect 5930 6490 5950 6510
rect 5950 6490 5955 6510
rect 5925 6485 5955 6490
rect 5925 6430 5955 6435
rect 5925 6410 5930 6430
rect 5930 6410 5950 6430
rect 5950 6410 5955 6430
rect 5925 6405 5955 6410
rect 5925 6350 5955 6355
rect 5925 6330 5930 6350
rect 5930 6330 5950 6350
rect 5950 6330 5955 6350
rect 5925 6325 5955 6330
rect 5925 6270 5955 6275
rect 5925 6250 5930 6270
rect 5930 6250 5950 6270
rect 5950 6250 5955 6270
rect 5925 6245 5955 6250
rect 5925 5870 5955 5875
rect 5925 5850 5930 5870
rect 5930 5850 5950 5870
rect 5950 5850 5955 5870
rect 5925 5845 5955 5850
rect 5925 5790 5955 5795
rect 5925 5770 5930 5790
rect 5930 5770 5950 5790
rect 5950 5770 5955 5790
rect 5925 5765 5955 5770
rect 5925 5710 5955 5715
rect 5925 5690 5930 5710
rect 5930 5690 5950 5710
rect 5950 5690 5955 5710
rect 5925 5685 5955 5690
rect 5925 5630 5955 5635
rect 5925 5610 5930 5630
rect 5930 5610 5950 5630
rect 5950 5610 5955 5630
rect 5925 5605 5955 5610
rect 5925 5550 5955 5555
rect 5925 5530 5930 5550
rect 5930 5530 5950 5550
rect 5950 5530 5955 5550
rect 5925 5525 5955 5530
rect 5925 5470 5955 5475
rect 5925 5450 5930 5470
rect 5930 5450 5950 5470
rect 5950 5450 5955 5470
rect 5925 5445 5955 5450
rect 5925 5390 5955 5395
rect 5925 5370 5930 5390
rect 5930 5370 5950 5390
rect 5950 5370 5955 5390
rect 5925 5365 5955 5370
rect 5925 5310 5955 5315
rect 5925 5290 5930 5310
rect 5930 5290 5950 5310
rect 5950 5290 5955 5310
rect 5925 5285 5955 5290
rect 5925 5230 5955 5235
rect 5925 5210 5930 5230
rect 5930 5210 5950 5230
rect 5950 5210 5955 5230
rect 5925 5205 5955 5210
rect 5925 5150 5955 5155
rect 5925 5130 5930 5150
rect 5930 5130 5950 5150
rect 5950 5130 5955 5150
rect 5925 5125 5955 5130
rect 5925 5070 5955 5075
rect 5925 5050 5930 5070
rect 5930 5050 5950 5070
rect 5950 5050 5955 5070
rect 5925 5045 5955 5050
rect 5925 4990 5955 4995
rect 5925 4970 5930 4990
rect 5930 4970 5950 4990
rect 5950 4970 5955 4990
rect 5925 4965 5955 4970
rect 5925 4910 5955 4915
rect 5925 4890 5930 4910
rect 5930 4890 5950 4910
rect 5950 4890 5955 4910
rect 5925 4885 5955 4890
rect 5925 4750 5955 4755
rect 5925 4730 5930 4750
rect 5930 4730 5950 4750
rect 5950 4730 5955 4750
rect 5925 4725 5955 4730
rect 5925 4670 5955 4675
rect 5925 4650 5930 4670
rect 5930 4650 5950 4670
rect 5950 4650 5955 4670
rect 5925 4645 5955 4650
rect 5925 4510 5955 4515
rect 5925 4490 5930 4510
rect 5930 4490 5950 4510
rect 5950 4490 5955 4510
rect 5925 4485 5955 4490
rect 5925 4430 5955 4435
rect 5925 4410 5930 4430
rect 5930 4410 5950 4430
rect 5950 4410 5955 4430
rect 5925 4405 5955 4410
rect 5925 4350 5955 4355
rect 5925 4330 5930 4350
rect 5930 4330 5950 4350
rect 5950 4330 5955 4350
rect 5925 4325 5955 4330
rect 5925 4270 5955 4275
rect 5925 4250 5930 4270
rect 5930 4250 5950 4270
rect 5950 4250 5955 4270
rect 5925 4245 5955 4250
rect 5925 4190 5955 4195
rect 5925 4170 5930 4190
rect 5930 4170 5950 4190
rect 5950 4170 5955 4190
rect 5925 4165 5955 4170
rect 5925 4110 5955 4115
rect 5925 4090 5930 4110
rect 5930 4090 5950 4110
rect 5950 4090 5955 4110
rect 5925 4085 5955 4090
rect 5925 4030 5955 4035
rect 5925 4010 5930 4030
rect 5930 4010 5950 4030
rect 5950 4010 5955 4030
rect 5925 4005 5955 4010
rect 5925 3950 5955 3955
rect 5925 3930 5930 3950
rect 5930 3930 5950 3950
rect 5950 3930 5955 3950
rect 5925 3925 5955 3930
rect 5925 3870 5955 3875
rect 5925 3850 5930 3870
rect 5930 3850 5950 3870
rect 5950 3850 5955 3870
rect 5925 3845 5955 3850
rect 5925 3710 5955 3715
rect 5925 3690 5930 3710
rect 5930 3690 5950 3710
rect 5950 3690 5955 3710
rect 5925 3685 5955 3690
rect 5925 3630 5955 3635
rect 5925 3610 5930 3630
rect 5930 3610 5950 3630
rect 5950 3610 5955 3630
rect 5925 3605 5955 3610
rect 5925 3470 5955 3475
rect 5925 3450 5930 3470
rect 5930 3450 5950 3470
rect 5950 3450 5955 3470
rect 5925 3445 5955 3450
rect 5925 3390 5955 3395
rect 5925 3370 5930 3390
rect 5930 3370 5950 3390
rect 5950 3370 5955 3390
rect 5925 3365 5955 3370
rect 5925 3230 5955 3235
rect 5925 3210 5930 3230
rect 5930 3210 5950 3230
rect 5950 3210 5955 3230
rect 5925 3205 5955 3210
rect 5925 3150 5955 3155
rect 5925 3130 5930 3150
rect 5930 3130 5950 3150
rect 5950 3130 5955 3150
rect 5925 3125 5955 3130
rect 5925 3070 5955 3075
rect 5925 3050 5930 3070
rect 5930 3050 5950 3070
rect 5950 3050 5955 3070
rect 5925 3045 5955 3050
rect 5925 2990 5955 2995
rect 5925 2970 5930 2990
rect 5930 2970 5950 2990
rect 5950 2970 5955 2990
rect 5925 2965 5955 2970
rect 5925 2910 5955 2915
rect 5925 2890 5930 2910
rect 5930 2890 5950 2910
rect 5950 2890 5955 2910
rect 5925 2885 5955 2890
rect 5925 2830 5955 2835
rect 5925 2810 5930 2830
rect 5930 2810 5950 2830
rect 5950 2810 5955 2830
rect 5925 2805 5955 2810
rect 5925 2750 5955 2755
rect 5925 2730 5930 2750
rect 5930 2730 5950 2750
rect 5950 2730 5955 2750
rect 5925 2725 5955 2730
rect 5925 2670 5955 2675
rect 5925 2650 5930 2670
rect 5930 2650 5950 2670
rect 5950 2650 5955 2670
rect 5925 2645 5955 2650
rect 5925 2590 5955 2595
rect 5925 2570 5930 2590
rect 5930 2570 5950 2590
rect 5950 2570 5955 2590
rect 5925 2565 5955 2570
rect 5925 2510 5955 2515
rect 5925 2490 5930 2510
rect 5930 2490 5950 2510
rect 5950 2490 5955 2510
rect 5925 2485 5955 2490
rect 5925 2430 5955 2435
rect 5925 2410 5930 2430
rect 5930 2410 5950 2430
rect 5950 2410 5955 2430
rect 5925 2405 5955 2410
rect 5925 2350 5955 2355
rect 5925 2330 5930 2350
rect 5930 2330 5950 2350
rect 5950 2330 5955 2350
rect 5925 2325 5955 2330
rect 5925 2270 5955 2275
rect 5925 2250 5930 2270
rect 5930 2250 5950 2270
rect 5950 2250 5955 2270
rect 5925 2245 5955 2250
rect 5925 2190 5955 2195
rect 5925 2170 5930 2190
rect 5930 2170 5950 2190
rect 5950 2170 5955 2190
rect 5925 2165 5955 2170
rect 5925 2110 5955 2115
rect 5925 2090 5930 2110
rect 5930 2090 5950 2110
rect 5950 2090 5955 2110
rect 5925 2085 5955 2090
rect 5925 2030 5955 2035
rect 5925 2010 5930 2030
rect 5930 2010 5950 2030
rect 5950 2010 5955 2030
rect 5925 2005 5955 2010
rect 5925 1950 5955 1955
rect 5925 1930 5930 1950
rect 5930 1930 5950 1950
rect 5950 1930 5955 1950
rect 5925 1925 5955 1930
rect 5925 1710 5955 1715
rect 5925 1690 5930 1710
rect 5930 1690 5950 1710
rect 5950 1690 5955 1710
rect 5925 1685 5955 1690
rect 5925 1630 5955 1635
rect 5925 1610 5930 1630
rect 5930 1610 5950 1630
rect 5950 1610 5955 1630
rect 5925 1605 5955 1610
rect 5925 1550 5955 1555
rect 5925 1530 5930 1550
rect 5930 1530 5950 1550
rect 5950 1530 5955 1550
rect 5925 1525 5955 1530
rect 5925 1470 5955 1475
rect 5925 1450 5930 1470
rect 5930 1450 5950 1470
rect 5950 1450 5955 1470
rect 5925 1445 5955 1450
rect 5925 1390 5955 1395
rect 5925 1370 5930 1390
rect 5930 1370 5950 1390
rect 5950 1370 5955 1390
rect 5925 1365 5955 1370
rect 5925 1310 5955 1315
rect 5925 1290 5930 1310
rect 5930 1290 5950 1310
rect 5950 1290 5955 1310
rect 5925 1285 5955 1290
rect 5925 1230 5955 1235
rect 5925 1210 5930 1230
rect 5930 1210 5950 1230
rect 5950 1210 5955 1230
rect 5925 1205 5955 1210
rect 5925 1150 5955 1155
rect 5925 1130 5930 1150
rect 5930 1130 5950 1150
rect 5950 1130 5955 1150
rect 5925 1125 5955 1130
rect 5925 1070 5955 1075
rect 5925 1050 5930 1070
rect 5930 1050 5950 1070
rect 5950 1050 5955 1070
rect 5925 1045 5955 1050
rect 5925 990 5955 995
rect 5925 970 5930 990
rect 5930 970 5950 990
rect 5950 970 5955 990
rect 5925 965 5955 970
rect 5925 830 5955 835
rect 5925 810 5930 830
rect 5930 810 5950 830
rect 5950 810 5955 830
rect 5925 805 5955 810
rect 5925 750 5955 755
rect 5925 730 5930 750
rect 5930 730 5950 750
rect 5950 730 5955 750
rect 5925 725 5955 730
rect 5925 670 5955 675
rect 5925 650 5930 670
rect 5930 650 5950 670
rect 5950 650 5955 670
rect 5925 645 5955 650
rect 5925 590 5955 595
rect 5925 570 5930 590
rect 5930 570 5950 590
rect 5950 570 5955 590
rect 5925 565 5955 570
rect 5925 510 5955 515
rect 5925 490 5930 510
rect 5930 490 5950 510
rect 5950 490 5955 510
rect 5925 485 5955 490
rect 5925 270 5955 275
rect 5925 250 5930 270
rect 5930 250 5950 270
rect 5950 250 5955 270
rect 5925 245 5955 250
rect 5925 190 5955 195
rect 5925 170 5930 190
rect 5930 170 5950 190
rect 5950 170 5955 190
rect 5925 165 5955 170
rect 5925 110 5955 115
rect 5925 90 5930 110
rect 5930 90 5950 110
rect 5950 90 5955 110
rect 5925 85 5955 90
rect 5925 30 5955 35
rect 5925 10 5930 30
rect 5930 10 5950 30
rect 5950 10 5955 30
rect 5925 5 5955 10
rect 6005 15710 6035 15715
rect 6005 15690 6010 15710
rect 6010 15690 6030 15710
rect 6030 15690 6035 15710
rect 6005 15685 6035 15690
rect 6005 15630 6035 15635
rect 6005 15610 6010 15630
rect 6010 15610 6030 15630
rect 6030 15610 6035 15630
rect 6005 15605 6035 15610
rect 6005 15550 6035 15555
rect 6005 15530 6010 15550
rect 6010 15530 6030 15550
rect 6030 15530 6035 15550
rect 6005 15525 6035 15530
rect 6005 15470 6035 15475
rect 6005 15450 6010 15470
rect 6010 15450 6030 15470
rect 6030 15450 6035 15470
rect 6005 15445 6035 15450
rect 6005 15390 6035 15395
rect 6005 15370 6010 15390
rect 6010 15370 6030 15390
rect 6030 15370 6035 15390
rect 6005 15365 6035 15370
rect 6005 15310 6035 15315
rect 6005 15290 6010 15310
rect 6010 15290 6030 15310
rect 6030 15290 6035 15310
rect 6005 15285 6035 15290
rect 6005 15230 6035 15235
rect 6005 15210 6010 15230
rect 6010 15210 6030 15230
rect 6030 15210 6035 15230
rect 6005 15205 6035 15210
rect 6005 15150 6035 15155
rect 6005 15130 6010 15150
rect 6010 15130 6030 15150
rect 6030 15130 6035 15150
rect 6005 15125 6035 15130
rect 6005 14990 6035 14995
rect 6005 14970 6010 14990
rect 6010 14970 6030 14990
rect 6030 14970 6035 14990
rect 6005 14965 6035 14970
rect 6005 14910 6035 14915
rect 6005 14890 6010 14910
rect 6010 14890 6030 14910
rect 6030 14890 6035 14910
rect 6005 14885 6035 14890
rect 6005 14830 6035 14835
rect 6005 14810 6010 14830
rect 6010 14810 6030 14830
rect 6030 14810 6035 14830
rect 6005 14805 6035 14810
rect 6005 14750 6035 14755
rect 6005 14730 6010 14750
rect 6010 14730 6030 14750
rect 6030 14730 6035 14750
rect 6005 14725 6035 14730
rect 6005 14670 6035 14675
rect 6005 14650 6010 14670
rect 6010 14650 6030 14670
rect 6030 14650 6035 14670
rect 6005 14645 6035 14650
rect 6005 14590 6035 14595
rect 6005 14570 6010 14590
rect 6010 14570 6030 14590
rect 6030 14570 6035 14590
rect 6005 14565 6035 14570
rect 6005 14510 6035 14515
rect 6005 14490 6010 14510
rect 6010 14490 6030 14510
rect 6030 14490 6035 14510
rect 6005 14485 6035 14490
rect 6005 14430 6035 14435
rect 6005 14410 6010 14430
rect 6010 14410 6030 14430
rect 6030 14410 6035 14430
rect 6005 14405 6035 14410
rect 6005 14030 6035 14035
rect 6005 14010 6010 14030
rect 6010 14010 6030 14030
rect 6030 14010 6035 14030
rect 6005 14005 6035 14010
rect 6005 13950 6035 13955
rect 6005 13930 6010 13950
rect 6010 13930 6030 13950
rect 6030 13930 6035 13950
rect 6005 13925 6035 13930
rect 6005 13870 6035 13875
rect 6005 13850 6010 13870
rect 6010 13850 6030 13870
rect 6030 13850 6035 13870
rect 6005 13845 6035 13850
rect 6005 13790 6035 13795
rect 6005 13770 6010 13790
rect 6010 13770 6030 13790
rect 6030 13770 6035 13790
rect 6005 13765 6035 13770
rect 6005 13710 6035 13715
rect 6005 13690 6010 13710
rect 6010 13690 6030 13710
rect 6030 13690 6035 13710
rect 6005 13685 6035 13690
rect 6005 13630 6035 13635
rect 6005 13610 6010 13630
rect 6010 13610 6030 13630
rect 6030 13610 6035 13630
rect 6005 13605 6035 13610
rect 6005 13550 6035 13555
rect 6005 13530 6010 13550
rect 6010 13530 6030 13550
rect 6030 13530 6035 13550
rect 6005 13525 6035 13530
rect 6005 13470 6035 13475
rect 6005 13450 6010 13470
rect 6010 13450 6030 13470
rect 6030 13450 6035 13470
rect 6005 13445 6035 13450
rect 6005 13070 6035 13075
rect 6005 13050 6010 13070
rect 6010 13050 6030 13070
rect 6030 13050 6035 13070
rect 6005 13045 6035 13050
rect 6005 12990 6035 12995
rect 6005 12970 6010 12990
rect 6010 12970 6030 12990
rect 6030 12970 6035 12990
rect 6005 12965 6035 12970
rect 6005 12910 6035 12915
rect 6005 12890 6010 12910
rect 6010 12890 6030 12910
rect 6030 12890 6035 12910
rect 6005 12885 6035 12890
rect 6005 12830 6035 12835
rect 6005 12810 6010 12830
rect 6010 12810 6030 12830
rect 6030 12810 6035 12830
rect 6005 12805 6035 12810
rect 6005 12750 6035 12755
rect 6005 12730 6010 12750
rect 6010 12730 6030 12750
rect 6030 12730 6035 12750
rect 6005 12725 6035 12730
rect 6005 12670 6035 12675
rect 6005 12650 6010 12670
rect 6010 12650 6030 12670
rect 6030 12650 6035 12670
rect 6005 12645 6035 12650
rect 6005 12590 6035 12595
rect 6005 12570 6010 12590
rect 6010 12570 6030 12590
rect 6030 12570 6035 12590
rect 6005 12565 6035 12570
rect 6005 12510 6035 12515
rect 6005 12490 6010 12510
rect 6010 12490 6030 12510
rect 6030 12490 6035 12510
rect 6005 12485 6035 12490
rect 6005 12350 6035 12355
rect 6005 12330 6010 12350
rect 6010 12330 6030 12350
rect 6030 12330 6035 12350
rect 6005 12325 6035 12330
rect 6005 12270 6035 12275
rect 6005 12250 6010 12270
rect 6010 12250 6030 12270
rect 6030 12250 6035 12270
rect 6005 12245 6035 12250
rect 6005 12190 6035 12195
rect 6005 12170 6010 12190
rect 6010 12170 6030 12190
rect 6030 12170 6035 12190
rect 6005 12165 6035 12170
rect 6005 12110 6035 12115
rect 6005 12090 6010 12110
rect 6010 12090 6030 12110
rect 6030 12090 6035 12110
rect 6005 12085 6035 12090
rect 6005 12030 6035 12035
rect 6005 12010 6010 12030
rect 6010 12010 6030 12030
rect 6030 12010 6035 12030
rect 6005 12005 6035 12010
rect 6005 11950 6035 11955
rect 6005 11930 6010 11950
rect 6010 11930 6030 11950
rect 6030 11930 6035 11950
rect 6005 11925 6035 11930
rect 6005 11870 6035 11875
rect 6005 11850 6010 11870
rect 6010 11850 6030 11870
rect 6030 11850 6035 11870
rect 6005 11845 6035 11850
rect 6005 11790 6035 11795
rect 6005 11770 6010 11790
rect 6010 11770 6030 11790
rect 6030 11770 6035 11790
rect 6005 11765 6035 11770
rect 6005 11710 6035 11715
rect 6005 11690 6010 11710
rect 6010 11690 6030 11710
rect 6030 11690 6035 11710
rect 6005 11685 6035 11690
rect 6005 11630 6035 11635
rect 6005 11610 6010 11630
rect 6010 11610 6030 11630
rect 6030 11610 6035 11630
rect 6005 11605 6035 11610
rect 6005 11550 6035 11555
rect 6005 11530 6010 11550
rect 6010 11530 6030 11550
rect 6030 11530 6035 11550
rect 6005 11525 6035 11530
rect 6005 11470 6035 11475
rect 6005 11450 6010 11470
rect 6010 11450 6030 11470
rect 6030 11450 6035 11470
rect 6005 11445 6035 11450
rect 6005 11390 6035 11395
rect 6005 11370 6010 11390
rect 6010 11370 6030 11390
rect 6030 11370 6035 11390
rect 6005 11365 6035 11370
rect 6005 11310 6035 11315
rect 6005 11290 6010 11310
rect 6010 11290 6030 11310
rect 6030 11290 6035 11310
rect 6005 11285 6035 11290
rect 6005 11230 6035 11235
rect 6005 11210 6010 11230
rect 6010 11210 6030 11230
rect 6030 11210 6035 11230
rect 6005 11205 6035 11210
rect 6005 11150 6035 11155
rect 6005 11130 6010 11150
rect 6010 11130 6030 11150
rect 6030 11130 6035 11150
rect 6005 11125 6035 11130
rect 6005 11070 6035 11075
rect 6005 11050 6010 11070
rect 6010 11050 6030 11070
rect 6030 11050 6035 11070
rect 6005 11045 6035 11050
rect 6005 10910 6035 10915
rect 6005 10890 6010 10910
rect 6010 10890 6030 10910
rect 6030 10890 6035 10910
rect 6005 10885 6035 10890
rect 6005 10830 6035 10835
rect 6005 10810 6010 10830
rect 6010 10810 6030 10830
rect 6030 10810 6035 10830
rect 6005 10805 6035 10810
rect 6005 10750 6035 10755
rect 6005 10730 6010 10750
rect 6010 10730 6030 10750
rect 6030 10730 6035 10750
rect 6005 10725 6035 10730
rect 6005 10670 6035 10675
rect 6005 10650 6010 10670
rect 6010 10650 6030 10670
rect 6030 10650 6035 10670
rect 6005 10645 6035 10650
rect 6005 10590 6035 10595
rect 6005 10570 6010 10590
rect 6010 10570 6030 10590
rect 6030 10570 6035 10590
rect 6005 10565 6035 10570
rect 6005 10510 6035 10515
rect 6005 10490 6010 10510
rect 6010 10490 6030 10510
rect 6030 10490 6035 10510
rect 6005 10485 6035 10490
rect 6005 10430 6035 10435
rect 6005 10410 6010 10430
rect 6010 10410 6030 10430
rect 6030 10410 6035 10430
rect 6005 10405 6035 10410
rect 6005 10350 6035 10355
rect 6005 10330 6010 10350
rect 6010 10330 6030 10350
rect 6030 10330 6035 10350
rect 6005 10325 6035 10330
rect 6005 9950 6035 9955
rect 6005 9930 6010 9950
rect 6010 9930 6030 9950
rect 6030 9930 6035 9950
rect 6005 9925 6035 9930
rect 6005 9870 6035 9875
rect 6005 9850 6010 9870
rect 6010 9850 6030 9870
rect 6030 9850 6035 9870
rect 6005 9845 6035 9850
rect 6005 9790 6035 9795
rect 6005 9770 6010 9790
rect 6010 9770 6030 9790
rect 6030 9770 6035 9790
rect 6005 9765 6035 9770
rect 6005 9710 6035 9715
rect 6005 9690 6010 9710
rect 6010 9690 6030 9710
rect 6030 9690 6035 9710
rect 6005 9685 6035 9690
rect 6005 9630 6035 9635
rect 6005 9610 6010 9630
rect 6010 9610 6030 9630
rect 6030 9610 6035 9630
rect 6005 9605 6035 9610
rect 6005 9550 6035 9555
rect 6005 9530 6010 9550
rect 6010 9530 6030 9550
rect 6030 9530 6035 9550
rect 6005 9525 6035 9530
rect 6005 9470 6035 9475
rect 6005 9450 6010 9470
rect 6010 9450 6030 9470
rect 6030 9450 6035 9470
rect 6005 9445 6035 9450
rect 6005 9390 6035 9395
rect 6005 9370 6010 9390
rect 6010 9370 6030 9390
rect 6030 9370 6035 9390
rect 6005 9365 6035 9370
rect 6005 8990 6035 8995
rect 6005 8970 6010 8990
rect 6010 8970 6030 8990
rect 6030 8970 6035 8990
rect 6005 8965 6035 8970
rect 6005 8910 6035 8915
rect 6005 8890 6010 8910
rect 6010 8890 6030 8910
rect 6030 8890 6035 8910
rect 6005 8885 6035 8890
rect 6005 8830 6035 8835
rect 6005 8810 6010 8830
rect 6010 8810 6030 8830
rect 6030 8810 6035 8830
rect 6005 8805 6035 8810
rect 6005 8750 6035 8755
rect 6005 8730 6010 8750
rect 6010 8730 6030 8750
rect 6030 8730 6035 8750
rect 6005 8725 6035 8730
rect 6005 8670 6035 8675
rect 6005 8650 6010 8670
rect 6010 8650 6030 8670
rect 6030 8650 6035 8670
rect 6005 8645 6035 8650
rect 6005 8590 6035 8595
rect 6005 8570 6010 8590
rect 6010 8570 6030 8590
rect 6030 8570 6035 8590
rect 6005 8565 6035 8570
rect 6005 8510 6035 8515
rect 6005 8490 6010 8510
rect 6010 8490 6030 8510
rect 6030 8490 6035 8510
rect 6005 8485 6035 8490
rect 6005 8430 6035 8435
rect 6005 8410 6010 8430
rect 6010 8410 6030 8430
rect 6030 8410 6035 8430
rect 6005 8405 6035 8410
rect 6005 8270 6035 8275
rect 6005 8250 6010 8270
rect 6010 8250 6030 8270
rect 6030 8250 6035 8270
rect 6005 8245 6035 8250
rect 6005 8190 6035 8195
rect 6005 8170 6010 8190
rect 6010 8170 6030 8190
rect 6030 8170 6035 8190
rect 6005 8165 6035 8170
rect 6005 8110 6035 8115
rect 6005 8090 6010 8110
rect 6010 8090 6030 8110
rect 6030 8090 6035 8110
rect 6005 8085 6035 8090
rect 6005 8030 6035 8035
rect 6005 8010 6010 8030
rect 6010 8010 6030 8030
rect 6030 8010 6035 8030
rect 6005 8005 6035 8010
rect 6005 7950 6035 7955
rect 6005 7930 6010 7950
rect 6010 7930 6030 7950
rect 6030 7930 6035 7950
rect 6005 7925 6035 7930
rect 6005 7870 6035 7875
rect 6005 7850 6010 7870
rect 6010 7850 6030 7870
rect 6030 7850 6035 7870
rect 6005 7845 6035 7850
rect 6005 7790 6035 7795
rect 6005 7770 6010 7790
rect 6010 7770 6030 7790
rect 6030 7770 6035 7790
rect 6005 7765 6035 7770
rect 6005 7710 6035 7715
rect 6005 7690 6010 7710
rect 6010 7690 6030 7710
rect 6030 7690 6035 7710
rect 6005 7685 6035 7690
rect 6005 7630 6035 7635
rect 6005 7610 6010 7630
rect 6010 7610 6030 7630
rect 6030 7610 6035 7630
rect 6005 7605 6035 7610
rect 6005 7550 6035 7555
rect 6005 7530 6010 7550
rect 6010 7530 6030 7550
rect 6030 7530 6035 7550
rect 6005 7525 6035 7530
rect 6005 7470 6035 7475
rect 6005 7450 6010 7470
rect 6010 7450 6030 7470
rect 6030 7450 6035 7470
rect 6005 7445 6035 7450
rect 6005 7390 6035 7395
rect 6005 7370 6010 7390
rect 6010 7370 6030 7390
rect 6030 7370 6035 7390
rect 6005 7365 6035 7370
rect 6005 7310 6035 7315
rect 6005 7290 6010 7310
rect 6010 7290 6030 7310
rect 6030 7290 6035 7310
rect 6005 7285 6035 7290
rect 6005 7230 6035 7235
rect 6005 7210 6010 7230
rect 6010 7210 6030 7230
rect 6030 7210 6035 7230
rect 6005 7205 6035 7210
rect 6005 7150 6035 7155
rect 6005 7130 6010 7150
rect 6010 7130 6030 7150
rect 6030 7130 6035 7150
rect 6005 7125 6035 7130
rect 6005 7070 6035 7075
rect 6005 7050 6010 7070
rect 6010 7050 6030 7070
rect 6030 7050 6035 7070
rect 6005 7045 6035 7050
rect 6005 6990 6035 6995
rect 6005 6970 6010 6990
rect 6010 6970 6030 6990
rect 6030 6970 6035 6990
rect 6005 6965 6035 6970
rect 6005 6830 6035 6835
rect 6005 6810 6010 6830
rect 6010 6810 6030 6830
rect 6030 6810 6035 6830
rect 6005 6805 6035 6810
rect 6005 6750 6035 6755
rect 6005 6730 6010 6750
rect 6010 6730 6030 6750
rect 6030 6730 6035 6750
rect 6005 6725 6035 6730
rect 6005 6670 6035 6675
rect 6005 6650 6010 6670
rect 6010 6650 6030 6670
rect 6030 6650 6035 6670
rect 6005 6645 6035 6650
rect 6005 6590 6035 6595
rect 6005 6570 6010 6590
rect 6010 6570 6030 6590
rect 6030 6570 6035 6590
rect 6005 6565 6035 6570
rect 6005 6510 6035 6515
rect 6005 6490 6010 6510
rect 6010 6490 6030 6510
rect 6030 6490 6035 6510
rect 6005 6485 6035 6490
rect 6005 6430 6035 6435
rect 6005 6410 6010 6430
rect 6010 6410 6030 6430
rect 6030 6410 6035 6430
rect 6005 6405 6035 6410
rect 6005 6350 6035 6355
rect 6005 6330 6010 6350
rect 6010 6330 6030 6350
rect 6030 6330 6035 6350
rect 6005 6325 6035 6330
rect 6005 6270 6035 6275
rect 6005 6250 6010 6270
rect 6010 6250 6030 6270
rect 6030 6250 6035 6270
rect 6005 6245 6035 6250
rect 6005 5870 6035 5875
rect 6005 5850 6010 5870
rect 6010 5850 6030 5870
rect 6030 5850 6035 5870
rect 6005 5845 6035 5850
rect 6005 5790 6035 5795
rect 6005 5770 6010 5790
rect 6010 5770 6030 5790
rect 6030 5770 6035 5790
rect 6005 5765 6035 5770
rect 6005 5710 6035 5715
rect 6005 5690 6010 5710
rect 6010 5690 6030 5710
rect 6030 5690 6035 5710
rect 6005 5685 6035 5690
rect 6005 5630 6035 5635
rect 6005 5610 6010 5630
rect 6010 5610 6030 5630
rect 6030 5610 6035 5630
rect 6005 5605 6035 5610
rect 6005 5550 6035 5555
rect 6005 5530 6010 5550
rect 6010 5530 6030 5550
rect 6030 5530 6035 5550
rect 6005 5525 6035 5530
rect 6005 5470 6035 5475
rect 6005 5450 6010 5470
rect 6010 5450 6030 5470
rect 6030 5450 6035 5470
rect 6005 5445 6035 5450
rect 6005 5390 6035 5395
rect 6005 5370 6010 5390
rect 6010 5370 6030 5390
rect 6030 5370 6035 5390
rect 6005 5365 6035 5370
rect 6005 5310 6035 5315
rect 6005 5290 6010 5310
rect 6010 5290 6030 5310
rect 6030 5290 6035 5310
rect 6005 5285 6035 5290
rect 6005 5230 6035 5235
rect 6005 5210 6010 5230
rect 6010 5210 6030 5230
rect 6030 5210 6035 5230
rect 6005 5205 6035 5210
rect 6005 5150 6035 5155
rect 6005 5130 6010 5150
rect 6010 5130 6030 5150
rect 6030 5130 6035 5150
rect 6005 5125 6035 5130
rect 6005 5070 6035 5075
rect 6005 5050 6010 5070
rect 6010 5050 6030 5070
rect 6030 5050 6035 5070
rect 6005 5045 6035 5050
rect 6005 4990 6035 4995
rect 6005 4970 6010 4990
rect 6010 4970 6030 4990
rect 6030 4970 6035 4990
rect 6005 4965 6035 4970
rect 6005 4910 6035 4915
rect 6005 4890 6010 4910
rect 6010 4890 6030 4910
rect 6030 4890 6035 4910
rect 6005 4885 6035 4890
rect 6005 4750 6035 4755
rect 6005 4730 6010 4750
rect 6010 4730 6030 4750
rect 6030 4730 6035 4750
rect 6005 4725 6035 4730
rect 6005 4670 6035 4675
rect 6005 4650 6010 4670
rect 6010 4650 6030 4670
rect 6030 4650 6035 4670
rect 6005 4645 6035 4650
rect 6005 4510 6035 4515
rect 6005 4490 6010 4510
rect 6010 4490 6030 4510
rect 6030 4490 6035 4510
rect 6005 4485 6035 4490
rect 6005 4430 6035 4435
rect 6005 4410 6010 4430
rect 6010 4410 6030 4430
rect 6030 4410 6035 4430
rect 6005 4405 6035 4410
rect 6005 4350 6035 4355
rect 6005 4330 6010 4350
rect 6010 4330 6030 4350
rect 6030 4330 6035 4350
rect 6005 4325 6035 4330
rect 6005 4270 6035 4275
rect 6005 4250 6010 4270
rect 6010 4250 6030 4270
rect 6030 4250 6035 4270
rect 6005 4245 6035 4250
rect 6005 4190 6035 4195
rect 6005 4170 6010 4190
rect 6010 4170 6030 4190
rect 6030 4170 6035 4190
rect 6005 4165 6035 4170
rect 6005 4110 6035 4115
rect 6005 4090 6010 4110
rect 6010 4090 6030 4110
rect 6030 4090 6035 4110
rect 6005 4085 6035 4090
rect 6005 4030 6035 4035
rect 6005 4010 6010 4030
rect 6010 4010 6030 4030
rect 6030 4010 6035 4030
rect 6005 4005 6035 4010
rect 6005 3950 6035 3955
rect 6005 3930 6010 3950
rect 6010 3930 6030 3950
rect 6030 3930 6035 3950
rect 6005 3925 6035 3930
rect 6005 3870 6035 3875
rect 6005 3850 6010 3870
rect 6010 3850 6030 3870
rect 6030 3850 6035 3870
rect 6005 3845 6035 3850
rect 6005 3710 6035 3715
rect 6005 3690 6010 3710
rect 6010 3690 6030 3710
rect 6030 3690 6035 3710
rect 6005 3685 6035 3690
rect 6005 3630 6035 3635
rect 6005 3610 6010 3630
rect 6010 3610 6030 3630
rect 6030 3610 6035 3630
rect 6005 3605 6035 3610
rect 6005 3470 6035 3475
rect 6005 3450 6010 3470
rect 6010 3450 6030 3470
rect 6030 3450 6035 3470
rect 6005 3445 6035 3450
rect 6005 3390 6035 3395
rect 6005 3370 6010 3390
rect 6010 3370 6030 3390
rect 6030 3370 6035 3390
rect 6005 3365 6035 3370
rect 6005 3230 6035 3235
rect 6005 3210 6010 3230
rect 6010 3210 6030 3230
rect 6030 3210 6035 3230
rect 6005 3205 6035 3210
rect 6005 3150 6035 3155
rect 6005 3130 6010 3150
rect 6010 3130 6030 3150
rect 6030 3130 6035 3150
rect 6005 3125 6035 3130
rect 6005 3070 6035 3075
rect 6005 3050 6010 3070
rect 6010 3050 6030 3070
rect 6030 3050 6035 3070
rect 6005 3045 6035 3050
rect 6005 2990 6035 2995
rect 6005 2970 6010 2990
rect 6010 2970 6030 2990
rect 6030 2970 6035 2990
rect 6005 2965 6035 2970
rect 6005 2910 6035 2915
rect 6005 2890 6010 2910
rect 6010 2890 6030 2910
rect 6030 2890 6035 2910
rect 6005 2885 6035 2890
rect 6005 2830 6035 2835
rect 6005 2810 6010 2830
rect 6010 2810 6030 2830
rect 6030 2810 6035 2830
rect 6005 2805 6035 2810
rect 6005 2750 6035 2755
rect 6005 2730 6010 2750
rect 6010 2730 6030 2750
rect 6030 2730 6035 2750
rect 6005 2725 6035 2730
rect 6005 2670 6035 2675
rect 6005 2650 6010 2670
rect 6010 2650 6030 2670
rect 6030 2650 6035 2670
rect 6005 2645 6035 2650
rect 6005 2590 6035 2595
rect 6005 2570 6010 2590
rect 6010 2570 6030 2590
rect 6030 2570 6035 2590
rect 6005 2565 6035 2570
rect 6005 2510 6035 2515
rect 6005 2490 6010 2510
rect 6010 2490 6030 2510
rect 6030 2490 6035 2510
rect 6005 2485 6035 2490
rect 6005 2430 6035 2435
rect 6005 2410 6010 2430
rect 6010 2410 6030 2430
rect 6030 2410 6035 2430
rect 6005 2405 6035 2410
rect 6005 2350 6035 2355
rect 6005 2330 6010 2350
rect 6010 2330 6030 2350
rect 6030 2330 6035 2350
rect 6005 2325 6035 2330
rect 6005 2270 6035 2275
rect 6005 2250 6010 2270
rect 6010 2250 6030 2270
rect 6030 2250 6035 2270
rect 6005 2245 6035 2250
rect 6005 2190 6035 2195
rect 6005 2170 6010 2190
rect 6010 2170 6030 2190
rect 6030 2170 6035 2190
rect 6005 2165 6035 2170
rect 6005 2110 6035 2115
rect 6005 2090 6010 2110
rect 6010 2090 6030 2110
rect 6030 2090 6035 2110
rect 6005 2085 6035 2090
rect 6005 2030 6035 2035
rect 6005 2010 6010 2030
rect 6010 2010 6030 2030
rect 6030 2010 6035 2030
rect 6005 2005 6035 2010
rect 6005 1950 6035 1955
rect 6005 1930 6010 1950
rect 6010 1930 6030 1950
rect 6030 1930 6035 1950
rect 6005 1925 6035 1930
rect 6005 1710 6035 1715
rect 6005 1690 6010 1710
rect 6010 1690 6030 1710
rect 6030 1690 6035 1710
rect 6005 1685 6035 1690
rect 6005 1630 6035 1635
rect 6005 1610 6010 1630
rect 6010 1610 6030 1630
rect 6030 1610 6035 1630
rect 6005 1605 6035 1610
rect 6005 1550 6035 1555
rect 6005 1530 6010 1550
rect 6010 1530 6030 1550
rect 6030 1530 6035 1550
rect 6005 1525 6035 1530
rect 6005 1470 6035 1475
rect 6005 1450 6010 1470
rect 6010 1450 6030 1470
rect 6030 1450 6035 1470
rect 6005 1445 6035 1450
rect 6005 1390 6035 1395
rect 6005 1370 6010 1390
rect 6010 1370 6030 1390
rect 6030 1370 6035 1390
rect 6005 1365 6035 1370
rect 6005 1310 6035 1315
rect 6005 1290 6010 1310
rect 6010 1290 6030 1310
rect 6030 1290 6035 1310
rect 6005 1285 6035 1290
rect 6005 1230 6035 1235
rect 6005 1210 6010 1230
rect 6010 1210 6030 1230
rect 6030 1210 6035 1230
rect 6005 1205 6035 1210
rect 6005 1150 6035 1155
rect 6005 1130 6010 1150
rect 6010 1130 6030 1150
rect 6030 1130 6035 1150
rect 6005 1125 6035 1130
rect 6005 1070 6035 1075
rect 6005 1050 6010 1070
rect 6010 1050 6030 1070
rect 6030 1050 6035 1070
rect 6005 1045 6035 1050
rect 6005 990 6035 995
rect 6005 970 6010 990
rect 6010 970 6030 990
rect 6030 970 6035 990
rect 6005 965 6035 970
rect 6005 830 6035 835
rect 6005 810 6010 830
rect 6010 810 6030 830
rect 6030 810 6035 830
rect 6005 805 6035 810
rect 6005 750 6035 755
rect 6005 730 6010 750
rect 6010 730 6030 750
rect 6030 730 6035 750
rect 6005 725 6035 730
rect 6005 670 6035 675
rect 6005 650 6010 670
rect 6010 650 6030 670
rect 6030 650 6035 670
rect 6005 645 6035 650
rect 6005 590 6035 595
rect 6005 570 6010 590
rect 6010 570 6030 590
rect 6030 570 6035 590
rect 6005 565 6035 570
rect 6005 510 6035 515
rect 6005 490 6010 510
rect 6010 490 6030 510
rect 6030 490 6035 510
rect 6005 485 6035 490
rect 6005 270 6035 275
rect 6005 250 6010 270
rect 6010 250 6030 270
rect 6030 250 6035 270
rect 6005 245 6035 250
rect 6005 190 6035 195
rect 6005 170 6010 190
rect 6010 170 6030 190
rect 6030 170 6035 190
rect 6005 165 6035 170
rect 6005 110 6035 115
rect 6005 90 6010 110
rect 6010 90 6030 110
rect 6030 90 6035 110
rect 6005 85 6035 90
rect 6005 30 6035 35
rect 6005 10 6010 30
rect 6010 10 6030 30
rect 6030 10 6035 30
rect 6005 5 6035 10
rect 6165 15710 6195 15715
rect 6165 15690 6170 15710
rect 6170 15690 6190 15710
rect 6190 15690 6195 15710
rect 6165 15685 6195 15690
rect 6165 15630 6195 15635
rect 6165 15610 6170 15630
rect 6170 15610 6190 15630
rect 6190 15610 6195 15630
rect 6165 15605 6195 15610
rect 6165 15550 6195 15555
rect 6165 15530 6170 15550
rect 6170 15530 6190 15550
rect 6190 15530 6195 15550
rect 6165 15525 6195 15530
rect 6165 15470 6195 15475
rect 6165 15450 6170 15470
rect 6170 15450 6190 15470
rect 6190 15450 6195 15470
rect 6165 15445 6195 15450
rect 6165 15390 6195 15395
rect 6165 15370 6170 15390
rect 6170 15370 6190 15390
rect 6190 15370 6195 15390
rect 6165 15365 6195 15370
rect 6165 15310 6195 15315
rect 6165 15290 6170 15310
rect 6170 15290 6190 15310
rect 6190 15290 6195 15310
rect 6165 15285 6195 15290
rect 6165 15230 6195 15235
rect 6165 15210 6170 15230
rect 6170 15210 6190 15230
rect 6190 15210 6195 15230
rect 6165 15205 6195 15210
rect 6165 15150 6195 15155
rect 6165 15130 6170 15150
rect 6170 15130 6190 15150
rect 6190 15130 6195 15150
rect 6165 15125 6195 15130
rect 6165 14990 6195 14995
rect 6165 14970 6170 14990
rect 6170 14970 6190 14990
rect 6190 14970 6195 14990
rect 6165 14965 6195 14970
rect 6165 14910 6195 14915
rect 6165 14890 6170 14910
rect 6170 14890 6190 14910
rect 6190 14890 6195 14910
rect 6165 14885 6195 14890
rect 6165 14830 6195 14835
rect 6165 14810 6170 14830
rect 6170 14810 6190 14830
rect 6190 14810 6195 14830
rect 6165 14805 6195 14810
rect 6165 14750 6195 14755
rect 6165 14730 6170 14750
rect 6170 14730 6190 14750
rect 6190 14730 6195 14750
rect 6165 14725 6195 14730
rect 6165 14670 6195 14675
rect 6165 14650 6170 14670
rect 6170 14650 6190 14670
rect 6190 14650 6195 14670
rect 6165 14645 6195 14650
rect 6165 14590 6195 14595
rect 6165 14570 6170 14590
rect 6170 14570 6190 14590
rect 6190 14570 6195 14590
rect 6165 14565 6195 14570
rect 6165 14510 6195 14515
rect 6165 14490 6170 14510
rect 6170 14490 6190 14510
rect 6190 14490 6195 14510
rect 6165 14485 6195 14490
rect 6165 14430 6195 14435
rect 6165 14410 6170 14430
rect 6170 14410 6190 14430
rect 6190 14410 6195 14430
rect 6165 14405 6195 14410
rect 6165 14030 6195 14035
rect 6165 14010 6170 14030
rect 6170 14010 6190 14030
rect 6190 14010 6195 14030
rect 6165 14005 6195 14010
rect 6165 13950 6195 13955
rect 6165 13930 6170 13950
rect 6170 13930 6190 13950
rect 6190 13930 6195 13950
rect 6165 13925 6195 13930
rect 6165 13870 6195 13875
rect 6165 13850 6170 13870
rect 6170 13850 6190 13870
rect 6190 13850 6195 13870
rect 6165 13845 6195 13850
rect 6165 13790 6195 13795
rect 6165 13770 6170 13790
rect 6170 13770 6190 13790
rect 6190 13770 6195 13790
rect 6165 13765 6195 13770
rect 6165 13710 6195 13715
rect 6165 13690 6170 13710
rect 6170 13690 6190 13710
rect 6190 13690 6195 13710
rect 6165 13685 6195 13690
rect 6165 13630 6195 13635
rect 6165 13610 6170 13630
rect 6170 13610 6190 13630
rect 6190 13610 6195 13630
rect 6165 13605 6195 13610
rect 6165 13550 6195 13555
rect 6165 13530 6170 13550
rect 6170 13530 6190 13550
rect 6190 13530 6195 13550
rect 6165 13525 6195 13530
rect 6165 13470 6195 13475
rect 6165 13450 6170 13470
rect 6170 13450 6190 13470
rect 6190 13450 6195 13470
rect 6165 13445 6195 13450
rect 6165 13070 6195 13075
rect 6165 13050 6170 13070
rect 6170 13050 6190 13070
rect 6190 13050 6195 13070
rect 6165 13045 6195 13050
rect 6165 12990 6195 12995
rect 6165 12970 6170 12990
rect 6170 12970 6190 12990
rect 6190 12970 6195 12990
rect 6165 12965 6195 12970
rect 6165 12910 6195 12915
rect 6165 12890 6170 12910
rect 6170 12890 6190 12910
rect 6190 12890 6195 12910
rect 6165 12885 6195 12890
rect 6165 12830 6195 12835
rect 6165 12810 6170 12830
rect 6170 12810 6190 12830
rect 6190 12810 6195 12830
rect 6165 12805 6195 12810
rect 6165 12750 6195 12755
rect 6165 12730 6170 12750
rect 6170 12730 6190 12750
rect 6190 12730 6195 12750
rect 6165 12725 6195 12730
rect 6165 12670 6195 12675
rect 6165 12650 6170 12670
rect 6170 12650 6190 12670
rect 6190 12650 6195 12670
rect 6165 12645 6195 12650
rect 6165 12590 6195 12595
rect 6165 12570 6170 12590
rect 6170 12570 6190 12590
rect 6190 12570 6195 12590
rect 6165 12565 6195 12570
rect 6165 12510 6195 12515
rect 6165 12490 6170 12510
rect 6170 12490 6190 12510
rect 6190 12490 6195 12510
rect 6165 12485 6195 12490
rect 6165 12350 6195 12355
rect 6165 12330 6170 12350
rect 6170 12330 6190 12350
rect 6190 12330 6195 12350
rect 6165 12325 6195 12330
rect 6165 12270 6195 12275
rect 6165 12250 6170 12270
rect 6170 12250 6190 12270
rect 6190 12250 6195 12270
rect 6165 12245 6195 12250
rect 6165 12190 6195 12195
rect 6165 12170 6170 12190
rect 6170 12170 6190 12190
rect 6190 12170 6195 12190
rect 6165 12165 6195 12170
rect 6165 12110 6195 12115
rect 6165 12090 6170 12110
rect 6170 12090 6190 12110
rect 6190 12090 6195 12110
rect 6165 12085 6195 12090
rect 6165 12030 6195 12035
rect 6165 12010 6170 12030
rect 6170 12010 6190 12030
rect 6190 12010 6195 12030
rect 6165 12005 6195 12010
rect 6165 11950 6195 11955
rect 6165 11930 6170 11950
rect 6170 11930 6190 11950
rect 6190 11930 6195 11950
rect 6165 11925 6195 11930
rect 6165 11870 6195 11875
rect 6165 11850 6170 11870
rect 6170 11850 6190 11870
rect 6190 11850 6195 11870
rect 6165 11845 6195 11850
rect 6165 11790 6195 11795
rect 6165 11770 6170 11790
rect 6170 11770 6190 11790
rect 6190 11770 6195 11790
rect 6165 11765 6195 11770
rect 6165 11710 6195 11715
rect 6165 11690 6170 11710
rect 6170 11690 6190 11710
rect 6190 11690 6195 11710
rect 6165 11685 6195 11690
rect 6165 11630 6195 11635
rect 6165 11610 6170 11630
rect 6170 11610 6190 11630
rect 6190 11610 6195 11630
rect 6165 11605 6195 11610
rect 6165 11550 6195 11555
rect 6165 11530 6170 11550
rect 6170 11530 6190 11550
rect 6190 11530 6195 11550
rect 6165 11525 6195 11530
rect 6165 11470 6195 11475
rect 6165 11450 6170 11470
rect 6170 11450 6190 11470
rect 6190 11450 6195 11470
rect 6165 11445 6195 11450
rect 6165 11390 6195 11395
rect 6165 11370 6170 11390
rect 6170 11370 6190 11390
rect 6190 11370 6195 11390
rect 6165 11365 6195 11370
rect 6165 11310 6195 11315
rect 6165 11290 6170 11310
rect 6170 11290 6190 11310
rect 6190 11290 6195 11310
rect 6165 11285 6195 11290
rect 6165 11230 6195 11235
rect 6165 11210 6170 11230
rect 6170 11210 6190 11230
rect 6190 11210 6195 11230
rect 6165 11205 6195 11210
rect 6165 11150 6195 11155
rect 6165 11130 6170 11150
rect 6170 11130 6190 11150
rect 6190 11130 6195 11150
rect 6165 11125 6195 11130
rect 6165 11070 6195 11075
rect 6165 11050 6170 11070
rect 6170 11050 6190 11070
rect 6190 11050 6195 11070
rect 6165 11045 6195 11050
rect 6165 10910 6195 10915
rect 6165 10890 6170 10910
rect 6170 10890 6190 10910
rect 6190 10890 6195 10910
rect 6165 10885 6195 10890
rect 6165 10830 6195 10835
rect 6165 10810 6170 10830
rect 6170 10810 6190 10830
rect 6190 10810 6195 10830
rect 6165 10805 6195 10810
rect 6165 10750 6195 10755
rect 6165 10730 6170 10750
rect 6170 10730 6190 10750
rect 6190 10730 6195 10750
rect 6165 10725 6195 10730
rect 6165 10670 6195 10675
rect 6165 10650 6170 10670
rect 6170 10650 6190 10670
rect 6190 10650 6195 10670
rect 6165 10645 6195 10650
rect 6165 10590 6195 10595
rect 6165 10570 6170 10590
rect 6170 10570 6190 10590
rect 6190 10570 6195 10590
rect 6165 10565 6195 10570
rect 6165 10510 6195 10515
rect 6165 10490 6170 10510
rect 6170 10490 6190 10510
rect 6190 10490 6195 10510
rect 6165 10485 6195 10490
rect 6165 10430 6195 10435
rect 6165 10410 6170 10430
rect 6170 10410 6190 10430
rect 6190 10410 6195 10430
rect 6165 10405 6195 10410
rect 6165 10350 6195 10355
rect 6165 10330 6170 10350
rect 6170 10330 6190 10350
rect 6190 10330 6195 10350
rect 6165 10325 6195 10330
rect 6165 9950 6195 9955
rect 6165 9930 6170 9950
rect 6170 9930 6190 9950
rect 6190 9930 6195 9950
rect 6165 9925 6195 9930
rect 6165 9870 6195 9875
rect 6165 9850 6170 9870
rect 6170 9850 6190 9870
rect 6190 9850 6195 9870
rect 6165 9845 6195 9850
rect 6165 9790 6195 9795
rect 6165 9770 6170 9790
rect 6170 9770 6190 9790
rect 6190 9770 6195 9790
rect 6165 9765 6195 9770
rect 6165 9710 6195 9715
rect 6165 9690 6170 9710
rect 6170 9690 6190 9710
rect 6190 9690 6195 9710
rect 6165 9685 6195 9690
rect 6165 9630 6195 9635
rect 6165 9610 6170 9630
rect 6170 9610 6190 9630
rect 6190 9610 6195 9630
rect 6165 9605 6195 9610
rect 6165 9550 6195 9555
rect 6165 9530 6170 9550
rect 6170 9530 6190 9550
rect 6190 9530 6195 9550
rect 6165 9525 6195 9530
rect 6165 9470 6195 9475
rect 6165 9450 6170 9470
rect 6170 9450 6190 9470
rect 6190 9450 6195 9470
rect 6165 9445 6195 9450
rect 6165 9390 6195 9395
rect 6165 9370 6170 9390
rect 6170 9370 6190 9390
rect 6190 9370 6195 9390
rect 6165 9365 6195 9370
rect 6165 8990 6195 8995
rect 6165 8970 6170 8990
rect 6170 8970 6190 8990
rect 6190 8970 6195 8990
rect 6165 8965 6195 8970
rect 6165 8910 6195 8915
rect 6165 8890 6170 8910
rect 6170 8890 6190 8910
rect 6190 8890 6195 8910
rect 6165 8885 6195 8890
rect 6165 8830 6195 8835
rect 6165 8810 6170 8830
rect 6170 8810 6190 8830
rect 6190 8810 6195 8830
rect 6165 8805 6195 8810
rect 6165 8750 6195 8755
rect 6165 8730 6170 8750
rect 6170 8730 6190 8750
rect 6190 8730 6195 8750
rect 6165 8725 6195 8730
rect 6165 8670 6195 8675
rect 6165 8650 6170 8670
rect 6170 8650 6190 8670
rect 6190 8650 6195 8670
rect 6165 8645 6195 8650
rect 6165 8590 6195 8595
rect 6165 8570 6170 8590
rect 6170 8570 6190 8590
rect 6190 8570 6195 8590
rect 6165 8565 6195 8570
rect 6165 8510 6195 8515
rect 6165 8490 6170 8510
rect 6170 8490 6190 8510
rect 6190 8490 6195 8510
rect 6165 8485 6195 8490
rect 6165 8430 6195 8435
rect 6165 8410 6170 8430
rect 6170 8410 6190 8430
rect 6190 8410 6195 8430
rect 6165 8405 6195 8410
rect 6165 8270 6195 8275
rect 6165 8250 6170 8270
rect 6170 8250 6190 8270
rect 6190 8250 6195 8270
rect 6165 8245 6195 8250
rect 6165 8190 6195 8195
rect 6165 8170 6170 8190
rect 6170 8170 6190 8190
rect 6190 8170 6195 8190
rect 6165 8165 6195 8170
rect 6165 8110 6195 8115
rect 6165 8090 6170 8110
rect 6170 8090 6190 8110
rect 6190 8090 6195 8110
rect 6165 8085 6195 8090
rect 6165 8030 6195 8035
rect 6165 8010 6170 8030
rect 6170 8010 6190 8030
rect 6190 8010 6195 8030
rect 6165 8005 6195 8010
rect 6165 7950 6195 7955
rect 6165 7930 6170 7950
rect 6170 7930 6190 7950
rect 6190 7930 6195 7950
rect 6165 7925 6195 7930
rect 6165 7870 6195 7875
rect 6165 7850 6170 7870
rect 6170 7850 6190 7870
rect 6190 7850 6195 7870
rect 6165 7845 6195 7850
rect 6165 7790 6195 7795
rect 6165 7770 6170 7790
rect 6170 7770 6190 7790
rect 6190 7770 6195 7790
rect 6165 7765 6195 7770
rect 6165 7710 6195 7715
rect 6165 7690 6170 7710
rect 6170 7690 6190 7710
rect 6190 7690 6195 7710
rect 6165 7685 6195 7690
rect 6165 7630 6195 7635
rect 6165 7610 6170 7630
rect 6170 7610 6190 7630
rect 6190 7610 6195 7630
rect 6165 7605 6195 7610
rect 6165 7550 6195 7555
rect 6165 7530 6170 7550
rect 6170 7530 6190 7550
rect 6190 7530 6195 7550
rect 6165 7525 6195 7530
rect 6165 7470 6195 7475
rect 6165 7450 6170 7470
rect 6170 7450 6190 7470
rect 6190 7450 6195 7470
rect 6165 7445 6195 7450
rect 6165 7390 6195 7395
rect 6165 7370 6170 7390
rect 6170 7370 6190 7390
rect 6190 7370 6195 7390
rect 6165 7365 6195 7370
rect 6165 7310 6195 7315
rect 6165 7290 6170 7310
rect 6170 7290 6190 7310
rect 6190 7290 6195 7310
rect 6165 7285 6195 7290
rect 6165 7230 6195 7235
rect 6165 7210 6170 7230
rect 6170 7210 6190 7230
rect 6190 7210 6195 7230
rect 6165 7205 6195 7210
rect 6165 7150 6195 7155
rect 6165 7130 6170 7150
rect 6170 7130 6190 7150
rect 6190 7130 6195 7150
rect 6165 7125 6195 7130
rect 6165 7070 6195 7075
rect 6165 7050 6170 7070
rect 6170 7050 6190 7070
rect 6190 7050 6195 7070
rect 6165 7045 6195 7050
rect 6165 6990 6195 6995
rect 6165 6970 6170 6990
rect 6170 6970 6190 6990
rect 6190 6970 6195 6990
rect 6165 6965 6195 6970
rect 6165 6830 6195 6835
rect 6165 6810 6170 6830
rect 6170 6810 6190 6830
rect 6190 6810 6195 6830
rect 6165 6805 6195 6810
rect 6165 6750 6195 6755
rect 6165 6730 6170 6750
rect 6170 6730 6190 6750
rect 6190 6730 6195 6750
rect 6165 6725 6195 6730
rect 6165 6670 6195 6675
rect 6165 6650 6170 6670
rect 6170 6650 6190 6670
rect 6190 6650 6195 6670
rect 6165 6645 6195 6650
rect 6165 6590 6195 6595
rect 6165 6570 6170 6590
rect 6170 6570 6190 6590
rect 6190 6570 6195 6590
rect 6165 6565 6195 6570
rect 6165 6510 6195 6515
rect 6165 6490 6170 6510
rect 6170 6490 6190 6510
rect 6190 6490 6195 6510
rect 6165 6485 6195 6490
rect 6165 6430 6195 6435
rect 6165 6410 6170 6430
rect 6170 6410 6190 6430
rect 6190 6410 6195 6430
rect 6165 6405 6195 6410
rect 6165 6350 6195 6355
rect 6165 6330 6170 6350
rect 6170 6330 6190 6350
rect 6190 6330 6195 6350
rect 6165 6325 6195 6330
rect 6165 6270 6195 6275
rect 6165 6250 6170 6270
rect 6170 6250 6190 6270
rect 6190 6250 6195 6270
rect 6165 6245 6195 6250
rect 6165 5870 6195 5875
rect 6165 5850 6170 5870
rect 6170 5850 6190 5870
rect 6190 5850 6195 5870
rect 6165 5845 6195 5850
rect 6165 5790 6195 5795
rect 6165 5770 6170 5790
rect 6170 5770 6190 5790
rect 6190 5770 6195 5790
rect 6165 5765 6195 5770
rect 6165 5710 6195 5715
rect 6165 5690 6170 5710
rect 6170 5690 6190 5710
rect 6190 5690 6195 5710
rect 6165 5685 6195 5690
rect 6165 5630 6195 5635
rect 6165 5610 6170 5630
rect 6170 5610 6190 5630
rect 6190 5610 6195 5630
rect 6165 5605 6195 5610
rect 6165 5550 6195 5555
rect 6165 5530 6170 5550
rect 6170 5530 6190 5550
rect 6190 5530 6195 5550
rect 6165 5525 6195 5530
rect 6165 5470 6195 5475
rect 6165 5450 6170 5470
rect 6170 5450 6190 5470
rect 6190 5450 6195 5470
rect 6165 5445 6195 5450
rect 6165 5390 6195 5395
rect 6165 5370 6170 5390
rect 6170 5370 6190 5390
rect 6190 5370 6195 5390
rect 6165 5365 6195 5370
rect 6165 5310 6195 5315
rect 6165 5290 6170 5310
rect 6170 5290 6190 5310
rect 6190 5290 6195 5310
rect 6165 5285 6195 5290
rect 6165 5230 6195 5235
rect 6165 5210 6170 5230
rect 6170 5210 6190 5230
rect 6190 5210 6195 5230
rect 6165 5205 6195 5210
rect 6165 5150 6195 5155
rect 6165 5130 6170 5150
rect 6170 5130 6190 5150
rect 6190 5130 6195 5150
rect 6165 5125 6195 5130
rect 6165 5070 6195 5075
rect 6165 5050 6170 5070
rect 6170 5050 6190 5070
rect 6190 5050 6195 5070
rect 6165 5045 6195 5050
rect 6165 4990 6195 4995
rect 6165 4970 6170 4990
rect 6170 4970 6190 4990
rect 6190 4970 6195 4990
rect 6165 4965 6195 4970
rect 6165 4910 6195 4915
rect 6165 4890 6170 4910
rect 6170 4890 6190 4910
rect 6190 4890 6195 4910
rect 6165 4885 6195 4890
rect 6165 4750 6195 4755
rect 6165 4730 6170 4750
rect 6170 4730 6190 4750
rect 6190 4730 6195 4750
rect 6165 4725 6195 4730
rect 6165 4670 6195 4675
rect 6165 4650 6170 4670
rect 6170 4650 6190 4670
rect 6190 4650 6195 4670
rect 6165 4645 6195 4650
rect 6165 4510 6195 4515
rect 6165 4490 6170 4510
rect 6170 4490 6190 4510
rect 6190 4490 6195 4510
rect 6165 4485 6195 4490
rect 6165 4430 6195 4435
rect 6165 4410 6170 4430
rect 6170 4410 6190 4430
rect 6190 4410 6195 4430
rect 6165 4405 6195 4410
rect 6165 4350 6195 4355
rect 6165 4330 6170 4350
rect 6170 4330 6190 4350
rect 6190 4330 6195 4350
rect 6165 4325 6195 4330
rect 6165 4270 6195 4275
rect 6165 4250 6170 4270
rect 6170 4250 6190 4270
rect 6190 4250 6195 4270
rect 6165 4245 6195 4250
rect 6165 4190 6195 4195
rect 6165 4170 6170 4190
rect 6170 4170 6190 4190
rect 6190 4170 6195 4190
rect 6165 4165 6195 4170
rect 6165 4110 6195 4115
rect 6165 4090 6170 4110
rect 6170 4090 6190 4110
rect 6190 4090 6195 4110
rect 6165 4085 6195 4090
rect 6165 4030 6195 4035
rect 6165 4010 6170 4030
rect 6170 4010 6190 4030
rect 6190 4010 6195 4030
rect 6165 4005 6195 4010
rect 6165 3950 6195 3955
rect 6165 3930 6170 3950
rect 6170 3930 6190 3950
rect 6190 3930 6195 3950
rect 6165 3925 6195 3930
rect 6165 3870 6195 3875
rect 6165 3850 6170 3870
rect 6170 3850 6190 3870
rect 6190 3850 6195 3870
rect 6165 3845 6195 3850
rect 6165 3710 6195 3715
rect 6165 3690 6170 3710
rect 6170 3690 6190 3710
rect 6190 3690 6195 3710
rect 6165 3685 6195 3690
rect 6165 3630 6195 3635
rect 6165 3610 6170 3630
rect 6170 3610 6190 3630
rect 6190 3610 6195 3630
rect 6165 3605 6195 3610
rect 6165 3470 6195 3475
rect 6165 3450 6170 3470
rect 6170 3450 6190 3470
rect 6190 3450 6195 3470
rect 6165 3445 6195 3450
rect 6165 3390 6195 3395
rect 6165 3370 6170 3390
rect 6170 3370 6190 3390
rect 6190 3370 6195 3390
rect 6165 3365 6195 3370
rect 6165 3230 6195 3235
rect 6165 3210 6170 3230
rect 6170 3210 6190 3230
rect 6190 3210 6195 3230
rect 6165 3205 6195 3210
rect 6165 3150 6195 3155
rect 6165 3130 6170 3150
rect 6170 3130 6190 3150
rect 6190 3130 6195 3150
rect 6165 3125 6195 3130
rect 6165 3070 6195 3075
rect 6165 3050 6170 3070
rect 6170 3050 6190 3070
rect 6190 3050 6195 3070
rect 6165 3045 6195 3050
rect 6165 2990 6195 2995
rect 6165 2970 6170 2990
rect 6170 2970 6190 2990
rect 6190 2970 6195 2990
rect 6165 2965 6195 2970
rect 6165 2910 6195 2915
rect 6165 2890 6170 2910
rect 6170 2890 6190 2910
rect 6190 2890 6195 2910
rect 6165 2885 6195 2890
rect 6165 2830 6195 2835
rect 6165 2810 6170 2830
rect 6170 2810 6190 2830
rect 6190 2810 6195 2830
rect 6165 2805 6195 2810
rect 6165 2750 6195 2755
rect 6165 2730 6170 2750
rect 6170 2730 6190 2750
rect 6190 2730 6195 2750
rect 6165 2725 6195 2730
rect 6165 2670 6195 2675
rect 6165 2650 6170 2670
rect 6170 2650 6190 2670
rect 6190 2650 6195 2670
rect 6165 2645 6195 2650
rect 6165 2590 6195 2595
rect 6165 2570 6170 2590
rect 6170 2570 6190 2590
rect 6190 2570 6195 2590
rect 6165 2565 6195 2570
rect 6165 2510 6195 2515
rect 6165 2490 6170 2510
rect 6170 2490 6190 2510
rect 6190 2490 6195 2510
rect 6165 2485 6195 2490
rect 6165 2430 6195 2435
rect 6165 2410 6170 2430
rect 6170 2410 6190 2430
rect 6190 2410 6195 2430
rect 6165 2405 6195 2410
rect 6165 2350 6195 2355
rect 6165 2330 6170 2350
rect 6170 2330 6190 2350
rect 6190 2330 6195 2350
rect 6165 2325 6195 2330
rect 6165 2270 6195 2275
rect 6165 2250 6170 2270
rect 6170 2250 6190 2270
rect 6190 2250 6195 2270
rect 6165 2245 6195 2250
rect 6165 2190 6195 2195
rect 6165 2170 6170 2190
rect 6170 2170 6190 2190
rect 6190 2170 6195 2190
rect 6165 2165 6195 2170
rect 6165 2110 6195 2115
rect 6165 2090 6170 2110
rect 6170 2090 6190 2110
rect 6190 2090 6195 2110
rect 6165 2085 6195 2090
rect 6165 2030 6195 2035
rect 6165 2010 6170 2030
rect 6170 2010 6190 2030
rect 6190 2010 6195 2030
rect 6165 2005 6195 2010
rect 6165 1950 6195 1955
rect 6165 1930 6170 1950
rect 6170 1930 6190 1950
rect 6190 1930 6195 1950
rect 6165 1925 6195 1930
rect 6165 1710 6195 1715
rect 6165 1690 6170 1710
rect 6170 1690 6190 1710
rect 6190 1690 6195 1710
rect 6165 1685 6195 1690
rect 6165 1630 6195 1635
rect 6165 1610 6170 1630
rect 6170 1610 6190 1630
rect 6190 1610 6195 1630
rect 6165 1605 6195 1610
rect 6165 1550 6195 1555
rect 6165 1530 6170 1550
rect 6170 1530 6190 1550
rect 6190 1530 6195 1550
rect 6165 1525 6195 1530
rect 6165 1470 6195 1475
rect 6165 1450 6170 1470
rect 6170 1450 6190 1470
rect 6190 1450 6195 1470
rect 6165 1445 6195 1450
rect 6165 1390 6195 1395
rect 6165 1370 6170 1390
rect 6170 1370 6190 1390
rect 6190 1370 6195 1390
rect 6165 1365 6195 1370
rect 6165 1310 6195 1315
rect 6165 1290 6170 1310
rect 6170 1290 6190 1310
rect 6190 1290 6195 1310
rect 6165 1285 6195 1290
rect 6165 1230 6195 1235
rect 6165 1210 6170 1230
rect 6170 1210 6190 1230
rect 6190 1210 6195 1230
rect 6165 1205 6195 1210
rect 6165 1150 6195 1155
rect 6165 1130 6170 1150
rect 6170 1130 6190 1150
rect 6190 1130 6195 1150
rect 6165 1125 6195 1130
rect 6165 1070 6195 1075
rect 6165 1050 6170 1070
rect 6170 1050 6190 1070
rect 6190 1050 6195 1070
rect 6165 1045 6195 1050
rect 6165 990 6195 995
rect 6165 970 6170 990
rect 6170 970 6190 990
rect 6190 970 6195 990
rect 6165 965 6195 970
rect 6165 830 6195 835
rect 6165 810 6170 830
rect 6170 810 6190 830
rect 6190 810 6195 830
rect 6165 805 6195 810
rect 6165 750 6195 755
rect 6165 730 6170 750
rect 6170 730 6190 750
rect 6190 730 6195 750
rect 6165 725 6195 730
rect 6165 670 6195 675
rect 6165 650 6170 670
rect 6170 650 6190 670
rect 6190 650 6195 670
rect 6165 645 6195 650
rect 6165 590 6195 595
rect 6165 570 6170 590
rect 6170 570 6190 590
rect 6190 570 6195 590
rect 6165 565 6195 570
rect 6165 510 6195 515
rect 6165 490 6170 510
rect 6170 490 6190 510
rect 6190 490 6195 510
rect 6165 485 6195 490
rect 6165 270 6195 275
rect 6165 250 6170 270
rect 6170 250 6190 270
rect 6190 250 6195 270
rect 6165 245 6195 250
rect 6165 190 6195 195
rect 6165 170 6170 190
rect 6170 170 6190 190
rect 6190 170 6195 190
rect 6165 165 6195 170
rect 6165 110 6195 115
rect 6165 90 6170 110
rect 6170 90 6190 110
rect 6190 90 6195 110
rect 6165 85 6195 90
rect 6165 30 6195 35
rect 6165 10 6170 30
rect 6170 10 6190 30
rect 6190 10 6195 30
rect 6165 5 6195 10
<< metal2 >>
rect 4240 15715 4440 15720
rect 4240 15685 4245 15715
rect 4275 15685 4405 15715
rect 4435 15685 4440 15715
rect 4240 15680 4440 15685
rect 4480 15715 4680 15720
rect 4480 15685 4485 15715
rect 4515 15685 4645 15715
rect 4675 15685 4680 15715
rect 4480 15680 4680 15685
rect 4720 15715 5720 15720
rect 4720 15685 4725 15715
rect 4755 15685 4885 15715
rect 4915 15685 5045 15715
rect 5075 15685 5205 15715
rect 5235 15685 5365 15715
rect 5395 15685 5525 15715
rect 5555 15685 5685 15715
rect 5715 15685 5720 15715
rect 4720 15680 5720 15685
rect 5760 15715 5960 15720
rect 5760 15685 5765 15715
rect 5795 15685 5925 15715
rect 5955 15685 5960 15715
rect 5760 15680 5960 15685
rect 6000 15715 6200 15720
rect 6000 15685 6005 15715
rect 6035 15685 6165 15715
rect 6195 15685 6200 15715
rect 6000 15680 6200 15685
rect 4240 15635 4440 15640
rect 4240 15605 4245 15635
rect 4275 15605 4405 15635
rect 4435 15605 4440 15635
rect 4240 15600 4440 15605
rect 4480 15635 4680 15640
rect 4480 15605 4485 15635
rect 4515 15605 4645 15635
rect 4675 15605 4680 15635
rect 4480 15600 4680 15605
rect 4720 15635 5720 15640
rect 4720 15605 4725 15635
rect 4755 15605 4885 15635
rect 4915 15605 5045 15635
rect 5075 15605 5205 15635
rect 5235 15605 5365 15635
rect 5395 15605 5525 15635
rect 5555 15605 5685 15635
rect 5715 15605 5720 15635
rect 4720 15600 5720 15605
rect 5760 15635 5960 15640
rect 5760 15605 5765 15635
rect 5795 15605 5925 15635
rect 5955 15605 5960 15635
rect 5760 15600 5960 15605
rect 6000 15635 6200 15640
rect 6000 15605 6005 15635
rect 6035 15605 6165 15635
rect 6195 15605 6200 15635
rect 6000 15600 6200 15605
rect 4240 15555 4440 15560
rect 4240 15525 4245 15555
rect 4275 15525 4405 15555
rect 4435 15525 4440 15555
rect 4240 15520 4440 15525
rect 4480 15555 4680 15560
rect 4480 15525 4485 15555
rect 4515 15525 4645 15555
rect 4675 15525 4680 15555
rect 4480 15520 4680 15525
rect 4720 15555 5720 15560
rect 4720 15525 4725 15555
rect 4755 15525 4885 15555
rect 4915 15525 5045 15555
rect 5075 15525 5205 15555
rect 5235 15525 5365 15555
rect 5395 15525 5525 15555
rect 5555 15525 5685 15555
rect 5715 15525 5720 15555
rect 4720 15520 5720 15525
rect 5760 15555 5960 15560
rect 5760 15525 5765 15555
rect 5795 15525 5925 15555
rect 5955 15525 5960 15555
rect 5760 15520 5960 15525
rect 6000 15555 6200 15560
rect 6000 15525 6005 15555
rect 6035 15525 6165 15555
rect 6195 15525 6200 15555
rect 6000 15520 6200 15525
rect 4240 15475 4440 15480
rect 4240 15445 4245 15475
rect 4275 15445 4405 15475
rect 4435 15445 4440 15475
rect 4240 15440 4440 15445
rect 4480 15475 4680 15480
rect 4480 15445 4485 15475
rect 4515 15445 4645 15475
rect 4675 15445 4680 15475
rect 4480 15440 4680 15445
rect 4720 15475 5720 15480
rect 4720 15445 4725 15475
rect 4755 15445 4885 15475
rect 4915 15445 5045 15475
rect 5075 15445 5205 15475
rect 5235 15445 5365 15475
rect 5395 15445 5525 15475
rect 5555 15445 5685 15475
rect 5715 15445 5720 15475
rect 4720 15440 5720 15445
rect 5760 15475 5960 15480
rect 5760 15445 5765 15475
rect 5795 15445 5925 15475
rect 5955 15445 5960 15475
rect 5760 15440 5960 15445
rect 6000 15475 6200 15480
rect 6000 15445 6005 15475
rect 6035 15445 6165 15475
rect 6195 15445 6200 15475
rect 6000 15440 6200 15445
rect 4240 15395 4440 15400
rect 4240 15365 4245 15395
rect 4275 15365 4405 15395
rect 4435 15365 4440 15395
rect 4240 15360 4440 15365
rect 4480 15395 4680 15400
rect 4480 15365 4485 15395
rect 4515 15365 4645 15395
rect 4675 15365 4680 15395
rect 4480 15360 4680 15365
rect 4720 15395 5720 15400
rect 4720 15365 4725 15395
rect 4755 15365 4885 15395
rect 4915 15365 5045 15395
rect 5075 15365 5205 15395
rect 5235 15365 5365 15395
rect 5395 15365 5525 15395
rect 5555 15365 5685 15395
rect 5715 15365 5720 15395
rect 4720 15360 5720 15365
rect 5760 15395 5960 15400
rect 5760 15365 5765 15395
rect 5795 15365 5925 15395
rect 5955 15365 5960 15395
rect 5760 15360 5960 15365
rect 6000 15395 6200 15400
rect 6000 15365 6005 15395
rect 6035 15365 6165 15395
rect 6195 15365 6200 15395
rect 6000 15360 6200 15365
rect 4240 15315 4440 15320
rect 4240 15285 4245 15315
rect 4275 15285 4405 15315
rect 4435 15285 4440 15315
rect 4240 15280 4440 15285
rect 4480 15315 4680 15320
rect 4480 15285 4485 15315
rect 4515 15285 4645 15315
rect 4675 15285 4680 15315
rect 4480 15280 4680 15285
rect 4720 15315 5720 15320
rect 4720 15285 4725 15315
rect 4755 15285 4885 15315
rect 4915 15285 5045 15315
rect 5075 15285 5205 15315
rect 5235 15285 5365 15315
rect 5395 15285 5525 15315
rect 5555 15285 5685 15315
rect 5715 15285 5720 15315
rect 4720 15280 5720 15285
rect 5760 15315 5960 15320
rect 5760 15285 5765 15315
rect 5795 15285 5925 15315
rect 5955 15285 5960 15315
rect 5760 15280 5960 15285
rect 6000 15315 6200 15320
rect 6000 15285 6005 15315
rect 6035 15285 6165 15315
rect 6195 15285 6200 15315
rect 6000 15280 6200 15285
rect 4240 15235 4440 15240
rect 4240 15205 4245 15235
rect 4275 15205 4405 15235
rect 4435 15205 4440 15235
rect 4240 15200 4440 15205
rect 4480 15235 4680 15240
rect 4480 15205 4485 15235
rect 4515 15205 4645 15235
rect 4675 15205 4680 15235
rect 4480 15200 4680 15205
rect 4720 15235 5720 15240
rect 4720 15205 4725 15235
rect 4755 15205 4885 15235
rect 4915 15205 5045 15235
rect 5075 15205 5205 15235
rect 5235 15205 5365 15235
rect 5395 15205 5525 15235
rect 5555 15205 5685 15235
rect 5715 15205 5720 15235
rect 4720 15200 5720 15205
rect 5760 15235 5960 15240
rect 5760 15205 5765 15235
rect 5795 15205 5925 15235
rect 5955 15205 5960 15235
rect 5760 15200 5960 15205
rect 6000 15235 6200 15240
rect 6000 15205 6005 15235
rect 6035 15205 6165 15235
rect 6195 15205 6200 15235
rect 6000 15200 6200 15205
rect 4240 15155 4440 15160
rect 4240 15125 4245 15155
rect 4275 15125 4405 15155
rect 4435 15125 4440 15155
rect 4240 15120 4440 15125
rect 4480 15155 4680 15160
rect 4480 15125 4485 15155
rect 4515 15125 4645 15155
rect 4675 15125 4680 15155
rect 4480 15120 4680 15125
rect 4720 15155 5720 15160
rect 4720 15125 4725 15155
rect 4755 15125 4885 15155
rect 4915 15125 5045 15155
rect 5075 15125 5205 15155
rect 5235 15125 5365 15155
rect 5395 15125 5525 15155
rect 5555 15125 5685 15155
rect 5715 15125 5720 15155
rect 4720 15120 5720 15125
rect 5760 15155 5960 15160
rect 5760 15125 5765 15155
rect 5795 15125 5925 15155
rect 5955 15125 5960 15155
rect 5760 15120 5960 15125
rect 6000 15155 6200 15160
rect 6000 15125 6005 15155
rect 6035 15125 6165 15155
rect 6195 15125 6200 15155
rect 6000 15120 6200 15125
rect 0 15075 10440 15080
rect 0 15045 4565 15075
rect 4595 15045 10440 15075
rect 0 15040 10440 15045
rect 4240 14995 4440 15000
rect 4240 14965 4245 14995
rect 4275 14965 4405 14995
rect 4435 14965 4440 14995
rect 4240 14960 4440 14965
rect 4480 14995 4680 15000
rect 4480 14965 4485 14995
rect 4515 14965 4645 14995
rect 4675 14965 4680 14995
rect 4480 14960 4680 14965
rect 4720 14995 5720 15000
rect 4720 14965 4725 14995
rect 4755 14965 4885 14995
rect 4915 14965 5045 14995
rect 5075 14965 5205 14995
rect 5235 14965 5365 14995
rect 5395 14965 5525 14995
rect 5555 14965 5685 14995
rect 5715 14965 5720 14995
rect 4720 14960 5720 14965
rect 5760 14995 5960 15000
rect 5760 14965 5765 14995
rect 5795 14965 5925 14995
rect 5955 14965 5960 14995
rect 5760 14960 5960 14965
rect 6000 14995 6200 15000
rect 6000 14965 6005 14995
rect 6035 14965 6165 14995
rect 6195 14965 6200 14995
rect 6000 14960 6200 14965
rect 4240 14915 4440 14920
rect 4240 14885 4245 14915
rect 4275 14885 4405 14915
rect 4435 14885 4440 14915
rect 4240 14880 4440 14885
rect 4480 14915 4680 14920
rect 4480 14885 4485 14915
rect 4515 14885 4645 14915
rect 4675 14885 4680 14915
rect 4480 14880 4680 14885
rect 4720 14915 5720 14920
rect 4720 14885 4725 14915
rect 4755 14885 4885 14915
rect 4915 14885 5045 14915
rect 5075 14885 5205 14915
rect 5235 14885 5365 14915
rect 5395 14885 5525 14915
rect 5555 14885 5685 14915
rect 5715 14885 5720 14915
rect 4720 14880 5720 14885
rect 5760 14915 5960 14920
rect 5760 14885 5765 14915
rect 5795 14885 5925 14915
rect 5955 14885 5960 14915
rect 5760 14880 5960 14885
rect 6000 14915 6200 14920
rect 6000 14885 6005 14915
rect 6035 14885 6165 14915
rect 6195 14885 6200 14915
rect 6000 14880 6200 14885
rect 4240 14835 4440 14840
rect 4240 14805 4245 14835
rect 4275 14805 4405 14835
rect 4435 14805 4440 14835
rect 4240 14800 4440 14805
rect 4480 14835 4680 14840
rect 4480 14805 4485 14835
rect 4515 14805 4645 14835
rect 4675 14805 4680 14835
rect 4480 14800 4680 14805
rect 4720 14835 5720 14840
rect 4720 14805 4725 14835
rect 4755 14805 4885 14835
rect 4915 14805 5045 14835
rect 5075 14805 5205 14835
rect 5235 14805 5365 14835
rect 5395 14805 5525 14835
rect 5555 14805 5685 14835
rect 5715 14805 5720 14835
rect 4720 14800 5720 14805
rect 5760 14835 5960 14840
rect 5760 14805 5765 14835
rect 5795 14805 5925 14835
rect 5955 14805 5960 14835
rect 5760 14800 5960 14805
rect 6000 14835 6200 14840
rect 6000 14805 6005 14835
rect 6035 14805 6165 14835
rect 6195 14805 6200 14835
rect 6000 14800 6200 14805
rect 4240 14755 4440 14760
rect 4240 14725 4245 14755
rect 4275 14725 4405 14755
rect 4435 14725 4440 14755
rect 4240 14720 4440 14725
rect 4480 14755 4680 14760
rect 4480 14725 4485 14755
rect 4515 14725 4645 14755
rect 4675 14725 4680 14755
rect 4480 14720 4680 14725
rect 4720 14755 5720 14760
rect 4720 14725 4725 14755
rect 4755 14725 4885 14755
rect 4915 14725 5045 14755
rect 5075 14725 5205 14755
rect 5235 14725 5365 14755
rect 5395 14725 5525 14755
rect 5555 14725 5685 14755
rect 5715 14725 5720 14755
rect 4720 14720 5720 14725
rect 5760 14755 5960 14760
rect 5760 14725 5765 14755
rect 5795 14725 5925 14755
rect 5955 14725 5960 14755
rect 5760 14720 5960 14725
rect 6000 14755 6200 14760
rect 6000 14725 6005 14755
rect 6035 14725 6165 14755
rect 6195 14725 6200 14755
rect 6000 14720 6200 14725
rect 4240 14675 4440 14680
rect 4240 14645 4245 14675
rect 4275 14645 4405 14675
rect 4435 14645 4440 14675
rect 4240 14640 4440 14645
rect 4480 14675 4680 14680
rect 4480 14645 4485 14675
rect 4515 14645 4645 14675
rect 4675 14645 4680 14675
rect 4480 14640 4680 14645
rect 4720 14675 5720 14680
rect 4720 14645 4725 14675
rect 4755 14645 4885 14675
rect 4915 14645 5045 14675
rect 5075 14645 5205 14675
rect 5235 14645 5365 14675
rect 5395 14645 5525 14675
rect 5555 14645 5685 14675
rect 5715 14645 5720 14675
rect 4720 14640 5720 14645
rect 5760 14675 5960 14680
rect 5760 14645 5765 14675
rect 5795 14645 5925 14675
rect 5955 14645 5960 14675
rect 5760 14640 5960 14645
rect 6000 14675 6200 14680
rect 6000 14645 6005 14675
rect 6035 14645 6165 14675
rect 6195 14645 6200 14675
rect 6000 14640 6200 14645
rect 4240 14595 4440 14600
rect 4240 14565 4245 14595
rect 4275 14565 4405 14595
rect 4435 14565 4440 14595
rect 4240 14560 4440 14565
rect 4480 14595 4680 14600
rect 4480 14565 4485 14595
rect 4515 14565 4645 14595
rect 4675 14565 4680 14595
rect 4480 14560 4680 14565
rect 4720 14595 5720 14600
rect 4720 14565 4725 14595
rect 4755 14565 4885 14595
rect 4915 14565 5045 14595
rect 5075 14565 5205 14595
rect 5235 14565 5365 14595
rect 5395 14565 5525 14595
rect 5555 14565 5685 14595
rect 5715 14565 5720 14595
rect 4720 14560 5720 14565
rect 5760 14595 5960 14600
rect 5760 14565 5765 14595
rect 5795 14565 5925 14595
rect 5955 14565 5960 14595
rect 5760 14560 5960 14565
rect 6000 14595 6200 14600
rect 6000 14565 6005 14595
rect 6035 14565 6165 14595
rect 6195 14565 6200 14595
rect 6000 14560 6200 14565
rect 4240 14515 4440 14520
rect 4240 14485 4245 14515
rect 4275 14485 4405 14515
rect 4435 14485 4440 14515
rect 4240 14480 4440 14485
rect 4480 14515 4680 14520
rect 4480 14485 4485 14515
rect 4515 14485 4645 14515
rect 4675 14485 4680 14515
rect 4480 14480 4680 14485
rect 4720 14515 5720 14520
rect 4720 14485 4725 14515
rect 4755 14485 4885 14515
rect 4915 14485 5045 14515
rect 5075 14485 5205 14515
rect 5235 14485 5365 14515
rect 5395 14485 5525 14515
rect 5555 14485 5685 14515
rect 5715 14485 5720 14515
rect 4720 14480 5720 14485
rect 5760 14515 5960 14520
rect 5760 14485 5765 14515
rect 5795 14485 5925 14515
rect 5955 14485 5960 14515
rect 5760 14480 5960 14485
rect 6000 14515 6200 14520
rect 6000 14485 6005 14515
rect 6035 14485 6165 14515
rect 6195 14485 6200 14515
rect 6000 14480 6200 14485
rect 4240 14435 4440 14440
rect 4240 14405 4245 14435
rect 4275 14405 4405 14435
rect 4435 14405 4440 14435
rect 4240 14400 4440 14405
rect 4480 14435 4680 14440
rect 4480 14405 4485 14435
rect 4515 14405 4645 14435
rect 4675 14405 4680 14435
rect 4480 14400 4680 14405
rect 4720 14435 5720 14440
rect 4720 14405 4725 14435
rect 4755 14405 4885 14435
rect 4915 14405 5045 14435
rect 5075 14405 5205 14435
rect 5235 14405 5365 14435
rect 5395 14405 5525 14435
rect 5555 14405 5685 14435
rect 5715 14405 5720 14435
rect 4720 14400 5720 14405
rect 5760 14435 5960 14440
rect 5760 14405 5765 14435
rect 5795 14405 5925 14435
rect 5955 14405 5960 14435
rect 5760 14400 5960 14405
rect 6000 14435 6200 14440
rect 6000 14405 6005 14435
rect 6035 14405 6165 14435
rect 6195 14405 6200 14435
rect 6000 14400 6200 14405
rect 0 14315 10440 14320
rect 0 14285 5285 14315
rect 5315 14285 10440 14315
rect 0 14280 10440 14285
rect 0 14155 5000 14160
rect 0 14125 4965 14155
rect 4995 14125 5000 14155
rect 0 14120 5000 14125
rect 5440 14155 10440 14160
rect 5440 14125 5445 14155
rect 5475 14125 10440 14155
rect 5440 14120 10440 14125
rect 4240 14035 4440 14040
rect 4240 14005 4245 14035
rect 4275 14005 4405 14035
rect 4435 14005 4440 14035
rect 4240 14000 4440 14005
rect 4480 14035 4680 14040
rect 4480 14005 4485 14035
rect 4515 14005 4645 14035
rect 4675 14005 4680 14035
rect 4480 14000 4680 14005
rect 4720 14035 5720 14040
rect 4720 14005 4725 14035
rect 4755 14005 4885 14035
rect 4915 14005 5045 14035
rect 5075 14005 5205 14035
rect 5235 14005 5365 14035
rect 5395 14005 5525 14035
rect 5555 14005 5685 14035
rect 5715 14005 5720 14035
rect 4720 14000 5720 14005
rect 5760 14035 5960 14040
rect 5760 14005 5765 14035
rect 5795 14005 5925 14035
rect 5955 14005 5960 14035
rect 5760 14000 5960 14005
rect 6000 14035 6200 14040
rect 6000 14005 6005 14035
rect 6035 14005 6165 14035
rect 6195 14005 6200 14035
rect 6000 14000 6200 14005
rect 4240 13955 4440 13960
rect 4240 13925 4245 13955
rect 4275 13925 4405 13955
rect 4435 13925 4440 13955
rect 4240 13920 4440 13925
rect 4480 13955 4680 13960
rect 4480 13925 4485 13955
rect 4515 13925 4645 13955
rect 4675 13925 4680 13955
rect 4480 13920 4680 13925
rect 4720 13955 5720 13960
rect 4720 13925 4725 13955
rect 4755 13925 4885 13955
rect 4915 13925 5045 13955
rect 5075 13925 5205 13955
rect 5235 13925 5365 13955
rect 5395 13925 5525 13955
rect 5555 13925 5685 13955
rect 5715 13925 5720 13955
rect 4720 13920 5720 13925
rect 5760 13955 5960 13960
rect 5760 13925 5765 13955
rect 5795 13925 5925 13955
rect 5955 13925 5960 13955
rect 5760 13920 5960 13925
rect 6000 13955 6200 13960
rect 6000 13925 6005 13955
rect 6035 13925 6165 13955
rect 6195 13925 6200 13955
rect 6000 13920 6200 13925
rect 4240 13875 4440 13880
rect 4240 13845 4245 13875
rect 4275 13845 4405 13875
rect 4435 13845 4440 13875
rect 4240 13840 4440 13845
rect 4480 13875 4680 13880
rect 4480 13845 4485 13875
rect 4515 13845 4645 13875
rect 4675 13845 4680 13875
rect 4480 13840 4680 13845
rect 4720 13875 5720 13880
rect 4720 13845 4725 13875
rect 4755 13845 4885 13875
rect 4915 13845 5045 13875
rect 5075 13845 5205 13875
rect 5235 13845 5365 13875
rect 5395 13845 5525 13875
rect 5555 13845 5685 13875
rect 5715 13845 5720 13875
rect 4720 13840 5720 13845
rect 5760 13875 5960 13880
rect 5760 13845 5765 13875
rect 5795 13845 5925 13875
rect 5955 13845 5960 13875
rect 5760 13840 5960 13845
rect 6000 13875 6200 13880
rect 6000 13845 6005 13875
rect 6035 13845 6165 13875
rect 6195 13845 6200 13875
rect 6000 13840 6200 13845
rect 4240 13795 4440 13800
rect 4240 13765 4245 13795
rect 4275 13765 4405 13795
rect 4435 13765 4440 13795
rect 4240 13760 4440 13765
rect 4480 13795 4680 13800
rect 4480 13765 4485 13795
rect 4515 13765 4645 13795
rect 4675 13765 4680 13795
rect 4480 13760 4680 13765
rect 4720 13795 5720 13800
rect 4720 13765 4725 13795
rect 4755 13765 4885 13795
rect 4915 13765 5045 13795
rect 5075 13765 5205 13795
rect 5235 13765 5365 13795
rect 5395 13765 5525 13795
rect 5555 13765 5685 13795
rect 5715 13765 5720 13795
rect 4720 13760 5720 13765
rect 5760 13795 5960 13800
rect 5760 13765 5765 13795
rect 5795 13765 5925 13795
rect 5955 13765 5960 13795
rect 5760 13760 5960 13765
rect 6000 13795 6200 13800
rect 6000 13765 6005 13795
rect 6035 13765 6165 13795
rect 6195 13765 6200 13795
rect 6000 13760 6200 13765
rect 4240 13715 4440 13720
rect 4240 13685 4245 13715
rect 4275 13685 4405 13715
rect 4435 13685 4440 13715
rect 4240 13680 4440 13685
rect 4480 13715 4680 13720
rect 4480 13685 4485 13715
rect 4515 13685 4645 13715
rect 4675 13685 4680 13715
rect 4480 13680 4680 13685
rect 4720 13715 5720 13720
rect 4720 13685 4725 13715
rect 4755 13685 4885 13715
rect 4915 13685 5045 13715
rect 5075 13685 5205 13715
rect 5235 13685 5365 13715
rect 5395 13685 5525 13715
rect 5555 13685 5685 13715
rect 5715 13685 5720 13715
rect 4720 13680 5720 13685
rect 5760 13715 5960 13720
rect 5760 13685 5765 13715
rect 5795 13685 5925 13715
rect 5955 13685 5960 13715
rect 5760 13680 5960 13685
rect 6000 13715 6200 13720
rect 6000 13685 6005 13715
rect 6035 13685 6165 13715
rect 6195 13685 6200 13715
rect 6000 13680 6200 13685
rect 4240 13635 4440 13640
rect 4240 13605 4245 13635
rect 4275 13605 4405 13635
rect 4435 13605 4440 13635
rect 4240 13600 4440 13605
rect 4480 13635 4680 13640
rect 4480 13605 4485 13635
rect 4515 13605 4645 13635
rect 4675 13605 4680 13635
rect 4480 13600 4680 13605
rect 4720 13635 5720 13640
rect 4720 13605 4725 13635
rect 4755 13605 4885 13635
rect 4915 13605 5045 13635
rect 5075 13605 5205 13635
rect 5235 13605 5365 13635
rect 5395 13605 5525 13635
rect 5555 13605 5685 13635
rect 5715 13605 5720 13635
rect 4720 13600 5720 13605
rect 5760 13635 5960 13640
rect 5760 13605 5765 13635
rect 5795 13605 5925 13635
rect 5955 13605 5960 13635
rect 5760 13600 5960 13605
rect 6000 13635 6200 13640
rect 6000 13605 6005 13635
rect 6035 13605 6165 13635
rect 6195 13605 6200 13635
rect 6000 13600 6200 13605
rect 4240 13555 4440 13560
rect 4240 13525 4245 13555
rect 4275 13525 4405 13555
rect 4435 13525 4440 13555
rect 4240 13520 4440 13525
rect 4480 13555 4680 13560
rect 4480 13525 4485 13555
rect 4515 13525 4645 13555
rect 4675 13525 4680 13555
rect 4480 13520 4680 13525
rect 4720 13555 5720 13560
rect 4720 13525 4725 13555
rect 4755 13525 4885 13555
rect 4915 13525 5045 13555
rect 5075 13525 5205 13555
rect 5235 13525 5365 13555
rect 5395 13525 5525 13555
rect 5555 13525 5685 13555
rect 5715 13525 5720 13555
rect 4720 13520 5720 13525
rect 5760 13555 5960 13560
rect 5760 13525 5765 13555
rect 5795 13525 5925 13555
rect 5955 13525 5960 13555
rect 5760 13520 5960 13525
rect 6000 13555 6200 13560
rect 6000 13525 6005 13555
rect 6035 13525 6165 13555
rect 6195 13525 6200 13555
rect 6000 13520 6200 13525
rect 4240 13475 4440 13480
rect 4240 13445 4245 13475
rect 4275 13445 4405 13475
rect 4435 13445 4440 13475
rect 4240 13440 4440 13445
rect 4480 13475 4680 13480
rect 4480 13445 4485 13475
rect 4515 13445 4645 13475
rect 4675 13445 4680 13475
rect 4480 13440 4680 13445
rect 4720 13475 5720 13480
rect 4720 13445 4725 13475
rect 4755 13445 4885 13475
rect 4915 13445 5045 13475
rect 5075 13445 5205 13475
rect 5235 13445 5365 13475
rect 5395 13445 5525 13475
rect 5555 13445 5685 13475
rect 5715 13445 5720 13475
rect 4720 13440 5720 13445
rect 5760 13475 5960 13480
rect 5760 13445 5765 13475
rect 5795 13445 5925 13475
rect 5955 13445 5960 13475
rect 5760 13440 5960 13445
rect 6000 13475 6200 13480
rect 6000 13445 6005 13475
rect 6035 13445 6165 13475
rect 6195 13445 6200 13475
rect 6000 13440 6200 13445
rect 0 13355 10440 13360
rect 0 13325 5285 13355
rect 5315 13325 10440 13355
rect 0 13320 10440 13325
rect 0 13195 5160 13200
rect 0 13165 5125 13195
rect 5155 13165 5160 13195
rect 0 13160 5160 13165
rect 5280 13195 10440 13200
rect 5280 13165 5285 13195
rect 5315 13165 10440 13195
rect 5280 13160 10440 13165
rect 4240 13075 4440 13080
rect 4240 13045 4245 13075
rect 4275 13045 4405 13075
rect 4435 13045 4440 13075
rect 4240 13040 4440 13045
rect 4480 13075 4680 13080
rect 4480 13045 4485 13075
rect 4515 13045 4645 13075
rect 4675 13045 4680 13075
rect 4480 13040 4680 13045
rect 4720 13075 5720 13080
rect 4720 13045 4725 13075
rect 4755 13045 4885 13075
rect 4915 13045 5045 13075
rect 5075 13045 5205 13075
rect 5235 13045 5365 13075
rect 5395 13045 5525 13075
rect 5555 13045 5685 13075
rect 5715 13045 5720 13075
rect 4720 13040 5720 13045
rect 5760 13075 5960 13080
rect 5760 13045 5765 13075
rect 5795 13045 5925 13075
rect 5955 13045 5960 13075
rect 5760 13040 5960 13045
rect 6000 13075 6200 13080
rect 6000 13045 6005 13075
rect 6035 13045 6165 13075
rect 6195 13045 6200 13075
rect 6000 13040 6200 13045
rect 4240 12995 4440 13000
rect 4240 12965 4245 12995
rect 4275 12965 4405 12995
rect 4435 12965 4440 12995
rect 4240 12960 4440 12965
rect 4480 12995 4680 13000
rect 4480 12965 4485 12995
rect 4515 12965 4645 12995
rect 4675 12965 4680 12995
rect 4480 12960 4680 12965
rect 4720 12995 5720 13000
rect 4720 12965 4725 12995
rect 4755 12965 4885 12995
rect 4915 12965 5045 12995
rect 5075 12965 5205 12995
rect 5235 12965 5365 12995
rect 5395 12965 5525 12995
rect 5555 12965 5685 12995
rect 5715 12965 5720 12995
rect 4720 12960 5720 12965
rect 5760 12995 5960 13000
rect 5760 12965 5765 12995
rect 5795 12965 5925 12995
rect 5955 12965 5960 12995
rect 5760 12960 5960 12965
rect 6000 12995 6200 13000
rect 6000 12965 6005 12995
rect 6035 12965 6165 12995
rect 6195 12965 6200 12995
rect 6000 12960 6200 12965
rect 4240 12915 4440 12920
rect 4240 12885 4245 12915
rect 4275 12885 4405 12915
rect 4435 12885 4440 12915
rect 4240 12880 4440 12885
rect 4480 12915 4680 12920
rect 4480 12885 4485 12915
rect 4515 12885 4645 12915
rect 4675 12885 4680 12915
rect 4480 12880 4680 12885
rect 4720 12915 5720 12920
rect 4720 12885 4725 12915
rect 4755 12885 4885 12915
rect 4915 12885 5045 12915
rect 5075 12885 5205 12915
rect 5235 12885 5365 12915
rect 5395 12885 5525 12915
rect 5555 12885 5685 12915
rect 5715 12885 5720 12915
rect 4720 12880 5720 12885
rect 5760 12915 5960 12920
rect 5760 12885 5765 12915
rect 5795 12885 5925 12915
rect 5955 12885 5960 12915
rect 5760 12880 5960 12885
rect 6000 12915 6200 12920
rect 6000 12885 6005 12915
rect 6035 12885 6165 12915
rect 6195 12885 6200 12915
rect 6000 12880 6200 12885
rect 4240 12835 4440 12840
rect 4240 12805 4245 12835
rect 4275 12805 4405 12835
rect 4435 12805 4440 12835
rect 4240 12800 4440 12805
rect 4480 12835 4680 12840
rect 4480 12805 4485 12835
rect 4515 12805 4645 12835
rect 4675 12805 4680 12835
rect 4480 12800 4680 12805
rect 4720 12835 5720 12840
rect 4720 12805 4725 12835
rect 4755 12805 4885 12835
rect 4915 12805 5045 12835
rect 5075 12805 5205 12835
rect 5235 12805 5365 12835
rect 5395 12805 5525 12835
rect 5555 12805 5685 12835
rect 5715 12805 5720 12835
rect 4720 12800 5720 12805
rect 5760 12835 5960 12840
rect 5760 12805 5765 12835
rect 5795 12805 5925 12835
rect 5955 12805 5960 12835
rect 5760 12800 5960 12805
rect 6000 12835 6200 12840
rect 6000 12805 6005 12835
rect 6035 12805 6165 12835
rect 6195 12805 6200 12835
rect 6000 12800 6200 12805
rect 4240 12755 4440 12760
rect 4240 12725 4245 12755
rect 4275 12725 4405 12755
rect 4435 12725 4440 12755
rect 4240 12720 4440 12725
rect 4480 12755 4680 12760
rect 4480 12725 4485 12755
rect 4515 12725 4645 12755
rect 4675 12725 4680 12755
rect 4480 12720 4680 12725
rect 4720 12755 5720 12760
rect 4720 12725 4725 12755
rect 4755 12725 4885 12755
rect 4915 12725 5045 12755
rect 5075 12725 5205 12755
rect 5235 12725 5365 12755
rect 5395 12725 5525 12755
rect 5555 12725 5685 12755
rect 5715 12725 5720 12755
rect 4720 12720 5720 12725
rect 5760 12755 5960 12760
rect 5760 12725 5765 12755
rect 5795 12725 5925 12755
rect 5955 12725 5960 12755
rect 5760 12720 5960 12725
rect 6000 12755 6200 12760
rect 6000 12725 6005 12755
rect 6035 12725 6165 12755
rect 6195 12725 6200 12755
rect 6000 12720 6200 12725
rect 4240 12675 4440 12680
rect 4240 12645 4245 12675
rect 4275 12645 4405 12675
rect 4435 12645 4440 12675
rect 4240 12640 4440 12645
rect 4480 12675 4680 12680
rect 4480 12645 4485 12675
rect 4515 12645 4645 12675
rect 4675 12645 4680 12675
rect 4480 12640 4680 12645
rect 4720 12675 5720 12680
rect 4720 12645 4725 12675
rect 4755 12645 4885 12675
rect 4915 12645 5045 12675
rect 5075 12645 5205 12675
rect 5235 12645 5365 12675
rect 5395 12645 5525 12675
rect 5555 12645 5685 12675
rect 5715 12645 5720 12675
rect 4720 12640 5720 12645
rect 5760 12675 5960 12680
rect 5760 12645 5765 12675
rect 5795 12645 5925 12675
rect 5955 12645 5960 12675
rect 5760 12640 5960 12645
rect 6000 12675 6200 12680
rect 6000 12645 6005 12675
rect 6035 12645 6165 12675
rect 6195 12645 6200 12675
rect 6000 12640 6200 12645
rect 4240 12595 4440 12600
rect 4240 12565 4245 12595
rect 4275 12565 4405 12595
rect 4435 12565 4440 12595
rect 4240 12560 4440 12565
rect 4480 12595 4680 12600
rect 4480 12565 4485 12595
rect 4515 12565 4645 12595
rect 4675 12565 4680 12595
rect 4480 12560 4680 12565
rect 4720 12595 5720 12600
rect 4720 12565 4725 12595
rect 4755 12565 4885 12595
rect 4915 12565 5045 12595
rect 5075 12565 5205 12595
rect 5235 12565 5365 12595
rect 5395 12565 5525 12595
rect 5555 12565 5685 12595
rect 5715 12565 5720 12595
rect 4720 12560 5720 12565
rect 5760 12595 5960 12600
rect 5760 12565 5765 12595
rect 5795 12565 5925 12595
rect 5955 12565 5960 12595
rect 5760 12560 5960 12565
rect 6000 12595 6200 12600
rect 6000 12565 6005 12595
rect 6035 12565 6165 12595
rect 6195 12565 6200 12595
rect 6000 12560 6200 12565
rect 4240 12515 4440 12520
rect 4240 12485 4245 12515
rect 4275 12485 4405 12515
rect 4435 12485 4440 12515
rect 4240 12480 4440 12485
rect 4480 12515 4680 12520
rect 4480 12485 4485 12515
rect 4515 12485 4645 12515
rect 4675 12485 4680 12515
rect 4480 12480 4680 12485
rect 4720 12515 5720 12520
rect 4720 12485 4725 12515
rect 4755 12485 4885 12515
rect 4915 12485 5045 12515
rect 5075 12485 5205 12515
rect 5235 12485 5365 12515
rect 5395 12485 5525 12515
rect 5555 12485 5685 12515
rect 5715 12485 5720 12515
rect 4720 12480 5720 12485
rect 5760 12515 5960 12520
rect 5760 12485 5765 12515
rect 5795 12485 5925 12515
rect 5955 12485 5960 12515
rect 5760 12480 5960 12485
rect 6000 12515 6200 12520
rect 6000 12485 6005 12515
rect 6035 12485 6165 12515
rect 6195 12485 6200 12515
rect 6000 12480 6200 12485
rect 0 12435 10440 12440
rect 0 12405 4565 12435
rect 4595 12405 10440 12435
rect 0 12400 10440 12405
rect 4240 12355 4440 12360
rect 4240 12325 4245 12355
rect 4275 12325 4405 12355
rect 4435 12325 4440 12355
rect 4240 12320 4440 12325
rect 4480 12355 4680 12360
rect 4480 12325 4485 12355
rect 4515 12325 4645 12355
rect 4675 12325 4680 12355
rect 4480 12320 4680 12325
rect 4720 12355 5720 12360
rect 4720 12325 4725 12355
rect 4755 12325 4885 12355
rect 4915 12325 5045 12355
rect 5075 12325 5205 12355
rect 5235 12325 5365 12355
rect 5395 12325 5525 12355
rect 5555 12325 5685 12355
rect 5715 12325 5720 12355
rect 4720 12320 5720 12325
rect 5760 12355 5960 12360
rect 5760 12325 5765 12355
rect 5795 12325 5925 12355
rect 5955 12325 5960 12355
rect 5760 12320 5960 12325
rect 6000 12355 6200 12360
rect 6000 12325 6005 12355
rect 6035 12325 6165 12355
rect 6195 12325 6200 12355
rect 6000 12320 6200 12325
rect 4240 12275 4440 12280
rect 4240 12245 4245 12275
rect 4275 12245 4405 12275
rect 4435 12245 4440 12275
rect 4240 12240 4440 12245
rect 4480 12275 4680 12280
rect 4480 12245 4485 12275
rect 4515 12245 4645 12275
rect 4675 12245 4680 12275
rect 4480 12240 4680 12245
rect 4720 12275 5720 12280
rect 4720 12245 4725 12275
rect 4755 12245 4885 12275
rect 4915 12245 5045 12275
rect 5075 12245 5205 12275
rect 5235 12245 5365 12275
rect 5395 12245 5525 12275
rect 5555 12245 5685 12275
rect 5715 12245 5720 12275
rect 4720 12240 5720 12245
rect 5760 12275 5960 12280
rect 5760 12245 5765 12275
rect 5795 12245 5925 12275
rect 5955 12245 5960 12275
rect 5760 12240 5960 12245
rect 6000 12275 6200 12280
rect 6000 12245 6005 12275
rect 6035 12245 6165 12275
rect 6195 12245 6200 12275
rect 6000 12240 6200 12245
rect 4240 12195 4440 12200
rect 4240 12165 4245 12195
rect 4275 12165 4405 12195
rect 4435 12165 4440 12195
rect 4240 12160 4440 12165
rect 4480 12195 4680 12200
rect 4480 12165 4485 12195
rect 4515 12165 4645 12195
rect 4675 12165 4680 12195
rect 4480 12160 4680 12165
rect 4720 12195 5720 12200
rect 4720 12165 4725 12195
rect 4755 12165 4885 12195
rect 4915 12165 5045 12195
rect 5075 12165 5205 12195
rect 5235 12165 5365 12195
rect 5395 12165 5525 12195
rect 5555 12165 5685 12195
rect 5715 12165 5720 12195
rect 4720 12160 5720 12165
rect 5760 12195 5960 12200
rect 5760 12165 5765 12195
rect 5795 12165 5925 12195
rect 5955 12165 5960 12195
rect 5760 12160 5960 12165
rect 6000 12195 6200 12200
rect 6000 12165 6005 12195
rect 6035 12165 6165 12195
rect 6195 12165 6200 12195
rect 6000 12160 6200 12165
rect 4240 12115 4440 12120
rect 4240 12085 4245 12115
rect 4275 12085 4405 12115
rect 4435 12085 4440 12115
rect 4240 12080 4440 12085
rect 4480 12115 4680 12120
rect 4480 12085 4485 12115
rect 4515 12085 4645 12115
rect 4675 12085 4680 12115
rect 4480 12080 4680 12085
rect 4720 12115 5720 12120
rect 4720 12085 4725 12115
rect 4755 12085 4885 12115
rect 4915 12085 5045 12115
rect 5075 12085 5205 12115
rect 5235 12085 5365 12115
rect 5395 12085 5525 12115
rect 5555 12085 5685 12115
rect 5715 12085 5720 12115
rect 4720 12080 5720 12085
rect 5760 12115 5960 12120
rect 5760 12085 5765 12115
rect 5795 12085 5925 12115
rect 5955 12085 5960 12115
rect 5760 12080 5960 12085
rect 6000 12115 6200 12120
rect 6000 12085 6005 12115
rect 6035 12085 6165 12115
rect 6195 12085 6200 12115
rect 6000 12080 6200 12085
rect 4240 12035 4440 12040
rect 4240 12005 4245 12035
rect 4275 12005 4405 12035
rect 4435 12005 4440 12035
rect 4240 12000 4440 12005
rect 4480 12035 4680 12040
rect 4480 12005 4485 12035
rect 4515 12005 4645 12035
rect 4675 12005 4680 12035
rect 4480 12000 4680 12005
rect 4720 12035 5720 12040
rect 4720 12005 4725 12035
rect 4755 12005 4885 12035
rect 4915 12005 5045 12035
rect 5075 12005 5205 12035
rect 5235 12005 5365 12035
rect 5395 12005 5525 12035
rect 5555 12005 5685 12035
rect 5715 12005 5720 12035
rect 4720 12000 5720 12005
rect 5760 12035 5960 12040
rect 5760 12005 5765 12035
rect 5795 12005 5925 12035
rect 5955 12005 5960 12035
rect 5760 12000 5960 12005
rect 6000 12035 6200 12040
rect 6000 12005 6005 12035
rect 6035 12005 6165 12035
rect 6195 12005 6200 12035
rect 6000 12000 6200 12005
rect 4240 11955 4440 11960
rect 4240 11925 4245 11955
rect 4275 11925 4405 11955
rect 4435 11925 4440 11955
rect 4240 11920 4440 11925
rect 4480 11955 4680 11960
rect 4480 11925 4485 11955
rect 4515 11925 4645 11955
rect 4675 11925 4680 11955
rect 4480 11920 4680 11925
rect 4720 11955 5720 11960
rect 4720 11925 4725 11955
rect 4755 11925 4885 11955
rect 4915 11925 5045 11955
rect 5075 11925 5205 11955
rect 5235 11925 5365 11955
rect 5395 11925 5525 11955
rect 5555 11925 5685 11955
rect 5715 11925 5720 11955
rect 4720 11920 5720 11925
rect 5760 11955 5960 11960
rect 5760 11925 5765 11955
rect 5795 11925 5925 11955
rect 5955 11925 5960 11955
rect 5760 11920 5960 11925
rect 6000 11955 6200 11960
rect 6000 11925 6005 11955
rect 6035 11925 6165 11955
rect 6195 11925 6200 11955
rect 6000 11920 6200 11925
rect 4240 11875 4440 11880
rect 4240 11845 4245 11875
rect 4275 11845 4405 11875
rect 4435 11845 4440 11875
rect 4240 11840 4440 11845
rect 4480 11875 4680 11880
rect 4480 11845 4485 11875
rect 4515 11845 4645 11875
rect 4675 11845 4680 11875
rect 4480 11840 4680 11845
rect 4720 11875 5720 11880
rect 4720 11845 4725 11875
rect 4755 11845 4885 11875
rect 4915 11845 5045 11875
rect 5075 11845 5205 11875
rect 5235 11845 5365 11875
rect 5395 11845 5525 11875
rect 5555 11845 5685 11875
rect 5715 11845 5720 11875
rect 4720 11840 5720 11845
rect 5760 11875 5960 11880
rect 5760 11845 5765 11875
rect 5795 11845 5925 11875
rect 5955 11845 5960 11875
rect 5760 11840 5960 11845
rect 6000 11875 6200 11880
rect 6000 11845 6005 11875
rect 6035 11845 6165 11875
rect 6195 11845 6200 11875
rect 6000 11840 6200 11845
rect 4240 11795 4440 11800
rect 4240 11765 4245 11795
rect 4275 11765 4405 11795
rect 4435 11765 4440 11795
rect 4240 11760 4440 11765
rect 4480 11795 4680 11800
rect 4480 11765 4485 11795
rect 4515 11765 4645 11795
rect 4675 11765 4680 11795
rect 4480 11760 4680 11765
rect 4720 11795 5720 11800
rect 4720 11765 4725 11795
rect 4755 11765 4885 11795
rect 4915 11765 5045 11795
rect 5075 11765 5205 11795
rect 5235 11765 5365 11795
rect 5395 11765 5525 11795
rect 5555 11765 5685 11795
rect 5715 11765 5720 11795
rect 4720 11760 5720 11765
rect 5760 11795 5960 11800
rect 5760 11765 5765 11795
rect 5795 11765 5925 11795
rect 5955 11765 5960 11795
rect 5760 11760 5960 11765
rect 6000 11795 6200 11800
rect 6000 11765 6005 11795
rect 6035 11765 6165 11795
rect 6195 11765 6200 11795
rect 6000 11760 6200 11765
rect 4240 11715 4440 11720
rect 4240 11685 4245 11715
rect 4275 11685 4405 11715
rect 4435 11685 4440 11715
rect 4240 11680 4440 11685
rect 4480 11715 4680 11720
rect 4480 11685 4485 11715
rect 4515 11685 4645 11715
rect 4675 11685 4680 11715
rect 4480 11680 4680 11685
rect 4720 11715 5720 11720
rect 4720 11685 4725 11715
rect 4755 11685 4885 11715
rect 4915 11685 5045 11715
rect 5075 11685 5205 11715
rect 5235 11685 5365 11715
rect 5395 11685 5525 11715
rect 5555 11685 5685 11715
rect 5715 11685 5720 11715
rect 4720 11680 5720 11685
rect 5760 11715 5960 11720
rect 5760 11685 5765 11715
rect 5795 11685 5925 11715
rect 5955 11685 5960 11715
rect 5760 11680 5960 11685
rect 6000 11715 6200 11720
rect 6000 11685 6005 11715
rect 6035 11685 6165 11715
rect 6195 11685 6200 11715
rect 6000 11680 6200 11685
rect 4240 11635 4440 11640
rect 4240 11605 4245 11635
rect 4275 11605 4405 11635
rect 4435 11605 4440 11635
rect 4240 11600 4440 11605
rect 4480 11635 4680 11640
rect 4480 11605 4485 11635
rect 4515 11605 4645 11635
rect 4675 11605 4680 11635
rect 4480 11600 4680 11605
rect 4720 11635 5720 11640
rect 4720 11605 4725 11635
rect 4755 11605 4885 11635
rect 4915 11605 5045 11635
rect 5075 11605 5205 11635
rect 5235 11605 5365 11635
rect 5395 11605 5525 11635
rect 5555 11605 5685 11635
rect 5715 11605 5720 11635
rect 4720 11600 5720 11605
rect 5760 11635 5960 11640
rect 5760 11605 5765 11635
rect 5795 11605 5925 11635
rect 5955 11605 5960 11635
rect 5760 11600 5960 11605
rect 6000 11635 6200 11640
rect 6000 11605 6005 11635
rect 6035 11605 6165 11635
rect 6195 11605 6200 11635
rect 6000 11600 6200 11605
rect 4240 11555 4440 11560
rect 4240 11525 4245 11555
rect 4275 11525 4405 11555
rect 4435 11525 4440 11555
rect 4240 11520 4440 11525
rect 4480 11555 4680 11560
rect 4480 11525 4485 11555
rect 4515 11525 4645 11555
rect 4675 11525 4680 11555
rect 4480 11520 4680 11525
rect 4720 11555 5720 11560
rect 4720 11525 4725 11555
rect 4755 11525 4885 11555
rect 4915 11525 5045 11555
rect 5075 11525 5205 11555
rect 5235 11525 5365 11555
rect 5395 11525 5525 11555
rect 5555 11525 5685 11555
rect 5715 11525 5720 11555
rect 4720 11520 5720 11525
rect 5760 11555 5960 11560
rect 5760 11525 5765 11555
rect 5795 11525 5925 11555
rect 5955 11525 5960 11555
rect 5760 11520 5960 11525
rect 6000 11555 6200 11560
rect 6000 11525 6005 11555
rect 6035 11525 6165 11555
rect 6195 11525 6200 11555
rect 6000 11520 6200 11525
rect 4240 11475 4440 11480
rect 4240 11445 4245 11475
rect 4275 11445 4405 11475
rect 4435 11445 4440 11475
rect 4240 11440 4440 11445
rect 4480 11475 4680 11480
rect 4480 11445 4485 11475
rect 4515 11445 4645 11475
rect 4675 11445 4680 11475
rect 4480 11440 4680 11445
rect 4720 11475 5720 11480
rect 4720 11445 4725 11475
rect 4755 11445 4885 11475
rect 4915 11445 5045 11475
rect 5075 11445 5205 11475
rect 5235 11445 5365 11475
rect 5395 11445 5525 11475
rect 5555 11445 5685 11475
rect 5715 11445 5720 11475
rect 4720 11440 5720 11445
rect 5760 11475 5960 11480
rect 5760 11445 5765 11475
rect 5795 11445 5925 11475
rect 5955 11445 5960 11475
rect 5760 11440 5960 11445
rect 6000 11475 6200 11480
rect 6000 11445 6005 11475
rect 6035 11445 6165 11475
rect 6195 11445 6200 11475
rect 6000 11440 6200 11445
rect 4240 11395 4440 11400
rect 4240 11365 4245 11395
rect 4275 11365 4405 11395
rect 4435 11365 4440 11395
rect 4240 11360 4440 11365
rect 4480 11395 4680 11400
rect 4480 11365 4485 11395
rect 4515 11365 4645 11395
rect 4675 11365 4680 11395
rect 4480 11360 4680 11365
rect 4720 11395 5720 11400
rect 4720 11365 4725 11395
rect 4755 11365 4885 11395
rect 4915 11365 5045 11395
rect 5075 11365 5205 11395
rect 5235 11365 5365 11395
rect 5395 11365 5525 11395
rect 5555 11365 5685 11395
rect 5715 11365 5720 11395
rect 4720 11360 5720 11365
rect 5760 11395 5960 11400
rect 5760 11365 5765 11395
rect 5795 11365 5925 11395
rect 5955 11365 5960 11395
rect 5760 11360 5960 11365
rect 6000 11395 6200 11400
rect 6000 11365 6005 11395
rect 6035 11365 6165 11395
rect 6195 11365 6200 11395
rect 6000 11360 6200 11365
rect 4240 11315 4440 11320
rect 4240 11285 4245 11315
rect 4275 11285 4405 11315
rect 4435 11285 4440 11315
rect 4240 11280 4440 11285
rect 4480 11315 4680 11320
rect 4480 11285 4485 11315
rect 4515 11285 4645 11315
rect 4675 11285 4680 11315
rect 4480 11280 4680 11285
rect 4720 11315 5720 11320
rect 4720 11285 4725 11315
rect 4755 11285 4885 11315
rect 4915 11285 5045 11315
rect 5075 11285 5205 11315
rect 5235 11285 5365 11315
rect 5395 11285 5525 11315
rect 5555 11285 5685 11315
rect 5715 11285 5720 11315
rect 4720 11280 5720 11285
rect 5760 11315 5960 11320
rect 5760 11285 5765 11315
rect 5795 11285 5925 11315
rect 5955 11285 5960 11315
rect 5760 11280 5960 11285
rect 6000 11315 6200 11320
rect 6000 11285 6005 11315
rect 6035 11285 6165 11315
rect 6195 11285 6200 11315
rect 6000 11280 6200 11285
rect 4240 11235 4440 11240
rect 4240 11205 4245 11235
rect 4275 11205 4405 11235
rect 4435 11205 4440 11235
rect 4240 11200 4440 11205
rect 4480 11235 4680 11240
rect 4480 11205 4485 11235
rect 4515 11205 4645 11235
rect 4675 11205 4680 11235
rect 4480 11200 4680 11205
rect 4720 11235 5720 11240
rect 4720 11205 4725 11235
rect 4755 11205 4885 11235
rect 4915 11205 5045 11235
rect 5075 11205 5205 11235
rect 5235 11205 5365 11235
rect 5395 11205 5525 11235
rect 5555 11205 5685 11235
rect 5715 11205 5720 11235
rect 4720 11200 5720 11205
rect 5760 11235 5960 11240
rect 5760 11205 5765 11235
rect 5795 11205 5925 11235
rect 5955 11205 5960 11235
rect 5760 11200 5960 11205
rect 6000 11235 6200 11240
rect 6000 11205 6005 11235
rect 6035 11205 6165 11235
rect 6195 11205 6200 11235
rect 6000 11200 6200 11205
rect 4240 11155 4440 11160
rect 4240 11125 4245 11155
rect 4275 11125 4405 11155
rect 4435 11125 4440 11155
rect 4240 11120 4440 11125
rect 4480 11155 4680 11160
rect 4480 11125 4485 11155
rect 4515 11125 4645 11155
rect 4675 11125 4680 11155
rect 4480 11120 4680 11125
rect 4720 11155 5720 11160
rect 4720 11125 4725 11155
rect 4755 11125 4885 11155
rect 4915 11125 5045 11155
rect 5075 11125 5205 11155
rect 5235 11125 5365 11155
rect 5395 11125 5525 11155
rect 5555 11125 5685 11155
rect 5715 11125 5720 11155
rect 4720 11120 5720 11125
rect 5760 11155 5960 11160
rect 5760 11125 5765 11155
rect 5795 11125 5925 11155
rect 5955 11125 5960 11155
rect 5760 11120 5960 11125
rect 6000 11155 6200 11160
rect 6000 11125 6005 11155
rect 6035 11125 6165 11155
rect 6195 11125 6200 11155
rect 6000 11120 6200 11125
rect 4240 11075 4440 11080
rect 4240 11045 4245 11075
rect 4275 11045 4405 11075
rect 4435 11045 4440 11075
rect 4240 11040 4440 11045
rect 4480 11075 4680 11080
rect 4480 11045 4485 11075
rect 4515 11045 4645 11075
rect 4675 11045 4680 11075
rect 4480 11040 4680 11045
rect 4720 11075 5720 11080
rect 4720 11045 4725 11075
rect 4755 11045 4885 11075
rect 4915 11045 5045 11075
rect 5075 11045 5205 11075
rect 5235 11045 5365 11075
rect 5395 11045 5525 11075
rect 5555 11045 5685 11075
rect 5715 11045 5720 11075
rect 4720 11040 5720 11045
rect 5760 11075 5960 11080
rect 5760 11045 5765 11075
rect 5795 11045 5925 11075
rect 5955 11045 5960 11075
rect 5760 11040 5960 11045
rect 6000 11075 6200 11080
rect 6000 11045 6005 11075
rect 6035 11045 6165 11075
rect 6195 11045 6200 11075
rect 6000 11040 6200 11045
rect 0 10995 10440 11000
rect 0 10965 4565 10995
rect 4595 10965 10440 10995
rect 0 10960 10440 10965
rect 4240 10915 4440 10920
rect 4240 10885 4245 10915
rect 4275 10885 4405 10915
rect 4435 10885 4440 10915
rect 4240 10880 4440 10885
rect 4480 10915 4680 10920
rect 4480 10885 4485 10915
rect 4515 10885 4645 10915
rect 4675 10885 4680 10915
rect 4480 10880 4680 10885
rect 4720 10915 5720 10920
rect 4720 10885 4725 10915
rect 4755 10885 4885 10915
rect 4915 10885 5045 10915
rect 5075 10885 5205 10915
rect 5235 10885 5365 10915
rect 5395 10885 5525 10915
rect 5555 10885 5685 10915
rect 5715 10885 5720 10915
rect 4720 10880 5720 10885
rect 5760 10915 5960 10920
rect 5760 10885 5765 10915
rect 5795 10885 5925 10915
rect 5955 10885 5960 10915
rect 5760 10880 5960 10885
rect 6000 10915 6200 10920
rect 6000 10885 6005 10915
rect 6035 10885 6165 10915
rect 6195 10885 6200 10915
rect 6000 10880 6200 10885
rect 4240 10835 4440 10840
rect 4240 10805 4245 10835
rect 4275 10805 4405 10835
rect 4435 10805 4440 10835
rect 4240 10800 4440 10805
rect 4480 10835 4680 10840
rect 4480 10805 4485 10835
rect 4515 10805 4645 10835
rect 4675 10805 4680 10835
rect 4480 10800 4680 10805
rect 4720 10835 5720 10840
rect 4720 10805 4725 10835
rect 4755 10805 4885 10835
rect 4915 10805 5045 10835
rect 5075 10805 5205 10835
rect 5235 10805 5365 10835
rect 5395 10805 5525 10835
rect 5555 10805 5685 10835
rect 5715 10805 5720 10835
rect 4720 10800 5720 10805
rect 5760 10835 5960 10840
rect 5760 10805 5765 10835
rect 5795 10805 5925 10835
rect 5955 10805 5960 10835
rect 5760 10800 5960 10805
rect 6000 10835 6200 10840
rect 6000 10805 6005 10835
rect 6035 10805 6165 10835
rect 6195 10805 6200 10835
rect 6000 10800 6200 10805
rect 4240 10755 4440 10760
rect 4240 10725 4245 10755
rect 4275 10725 4405 10755
rect 4435 10725 4440 10755
rect 4240 10720 4440 10725
rect 4480 10755 4680 10760
rect 4480 10725 4485 10755
rect 4515 10725 4645 10755
rect 4675 10725 4680 10755
rect 4480 10720 4680 10725
rect 4720 10755 5720 10760
rect 4720 10725 4725 10755
rect 4755 10725 4885 10755
rect 4915 10725 5045 10755
rect 5075 10725 5205 10755
rect 5235 10725 5365 10755
rect 5395 10725 5525 10755
rect 5555 10725 5685 10755
rect 5715 10725 5720 10755
rect 4720 10720 5720 10725
rect 5760 10755 5960 10760
rect 5760 10725 5765 10755
rect 5795 10725 5925 10755
rect 5955 10725 5960 10755
rect 5760 10720 5960 10725
rect 6000 10755 6200 10760
rect 6000 10725 6005 10755
rect 6035 10725 6165 10755
rect 6195 10725 6200 10755
rect 6000 10720 6200 10725
rect 4240 10675 4440 10680
rect 4240 10645 4245 10675
rect 4275 10645 4405 10675
rect 4435 10645 4440 10675
rect 4240 10640 4440 10645
rect 4480 10675 4680 10680
rect 4480 10645 4485 10675
rect 4515 10645 4645 10675
rect 4675 10645 4680 10675
rect 4480 10640 4680 10645
rect 4720 10675 5720 10680
rect 4720 10645 4725 10675
rect 4755 10645 4885 10675
rect 4915 10645 5045 10675
rect 5075 10645 5205 10675
rect 5235 10645 5365 10675
rect 5395 10645 5525 10675
rect 5555 10645 5685 10675
rect 5715 10645 5720 10675
rect 4720 10640 5720 10645
rect 5760 10675 5960 10680
rect 5760 10645 5765 10675
rect 5795 10645 5925 10675
rect 5955 10645 5960 10675
rect 5760 10640 5960 10645
rect 6000 10675 6200 10680
rect 6000 10645 6005 10675
rect 6035 10645 6165 10675
rect 6195 10645 6200 10675
rect 6000 10640 6200 10645
rect 4240 10595 4440 10600
rect 4240 10565 4245 10595
rect 4275 10565 4405 10595
rect 4435 10565 4440 10595
rect 4240 10560 4440 10565
rect 4480 10595 4680 10600
rect 4480 10565 4485 10595
rect 4515 10565 4645 10595
rect 4675 10565 4680 10595
rect 4480 10560 4680 10565
rect 4720 10595 5720 10600
rect 4720 10565 4725 10595
rect 4755 10565 4885 10595
rect 4915 10565 5045 10595
rect 5075 10565 5205 10595
rect 5235 10565 5365 10595
rect 5395 10565 5525 10595
rect 5555 10565 5685 10595
rect 5715 10565 5720 10595
rect 4720 10560 5720 10565
rect 5760 10595 5960 10600
rect 5760 10565 5765 10595
rect 5795 10565 5925 10595
rect 5955 10565 5960 10595
rect 5760 10560 5960 10565
rect 6000 10595 6200 10600
rect 6000 10565 6005 10595
rect 6035 10565 6165 10595
rect 6195 10565 6200 10595
rect 6000 10560 6200 10565
rect 4240 10515 4440 10520
rect 4240 10485 4245 10515
rect 4275 10485 4405 10515
rect 4435 10485 4440 10515
rect 4240 10480 4440 10485
rect 4480 10515 4680 10520
rect 4480 10485 4485 10515
rect 4515 10485 4645 10515
rect 4675 10485 4680 10515
rect 4480 10480 4680 10485
rect 4720 10515 5720 10520
rect 4720 10485 4725 10515
rect 4755 10485 4885 10515
rect 4915 10485 5045 10515
rect 5075 10485 5205 10515
rect 5235 10485 5365 10515
rect 5395 10485 5525 10515
rect 5555 10485 5685 10515
rect 5715 10485 5720 10515
rect 4720 10480 5720 10485
rect 5760 10515 5960 10520
rect 5760 10485 5765 10515
rect 5795 10485 5925 10515
rect 5955 10485 5960 10515
rect 5760 10480 5960 10485
rect 6000 10515 6200 10520
rect 6000 10485 6005 10515
rect 6035 10485 6165 10515
rect 6195 10485 6200 10515
rect 6000 10480 6200 10485
rect 4240 10435 4440 10440
rect 4240 10405 4245 10435
rect 4275 10405 4405 10435
rect 4435 10405 4440 10435
rect 4240 10400 4440 10405
rect 4480 10435 4680 10440
rect 4480 10405 4485 10435
rect 4515 10405 4645 10435
rect 4675 10405 4680 10435
rect 4480 10400 4680 10405
rect 4720 10435 5720 10440
rect 4720 10405 4725 10435
rect 4755 10405 4885 10435
rect 4915 10405 5045 10435
rect 5075 10405 5205 10435
rect 5235 10405 5365 10435
rect 5395 10405 5525 10435
rect 5555 10405 5685 10435
rect 5715 10405 5720 10435
rect 4720 10400 5720 10405
rect 5760 10435 5960 10440
rect 5760 10405 5765 10435
rect 5795 10405 5925 10435
rect 5955 10405 5960 10435
rect 5760 10400 5960 10405
rect 6000 10435 6200 10440
rect 6000 10405 6005 10435
rect 6035 10405 6165 10435
rect 6195 10405 6200 10435
rect 6000 10400 6200 10405
rect 4240 10355 4440 10360
rect 4240 10325 4245 10355
rect 4275 10325 4405 10355
rect 4435 10325 4440 10355
rect 4240 10320 4440 10325
rect 4480 10355 4680 10360
rect 4480 10325 4485 10355
rect 4515 10325 4645 10355
rect 4675 10325 4680 10355
rect 4480 10320 4680 10325
rect 4720 10355 5720 10360
rect 4720 10325 4725 10355
rect 4755 10325 4885 10355
rect 4915 10325 5045 10355
rect 5075 10325 5205 10355
rect 5235 10325 5365 10355
rect 5395 10325 5525 10355
rect 5555 10325 5685 10355
rect 5715 10325 5720 10355
rect 4720 10320 5720 10325
rect 5760 10355 5960 10360
rect 5760 10325 5765 10355
rect 5795 10325 5925 10355
rect 5955 10325 5960 10355
rect 5760 10320 5960 10325
rect 6000 10355 6200 10360
rect 6000 10325 6005 10355
rect 6035 10325 6165 10355
rect 6195 10325 6200 10355
rect 6000 10320 6200 10325
rect 0 10235 10440 10240
rect 0 10205 5125 10235
rect 5155 10205 10440 10235
rect 0 10200 10440 10205
rect 0 10075 10440 10080
rect 0 10045 5125 10075
rect 5155 10045 10440 10075
rect 0 10040 10440 10045
rect 4240 9955 4440 9960
rect 4240 9925 4245 9955
rect 4275 9925 4405 9955
rect 4435 9925 4440 9955
rect 4240 9920 4440 9925
rect 4480 9955 4680 9960
rect 4480 9925 4485 9955
rect 4515 9925 4645 9955
rect 4675 9925 4680 9955
rect 4480 9920 4680 9925
rect 4720 9955 5720 9960
rect 4720 9925 4725 9955
rect 4755 9925 4885 9955
rect 4915 9925 5045 9955
rect 5075 9925 5205 9955
rect 5235 9925 5365 9955
rect 5395 9925 5525 9955
rect 5555 9925 5685 9955
rect 5715 9925 5720 9955
rect 4720 9920 5720 9925
rect 5760 9955 5960 9960
rect 5760 9925 5765 9955
rect 5795 9925 5925 9955
rect 5955 9925 5960 9955
rect 5760 9920 5960 9925
rect 6000 9955 6200 9960
rect 6000 9925 6005 9955
rect 6035 9925 6165 9955
rect 6195 9925 6200 9955
rect 6000 9920 6200 9925
rect 4240 9875 4440 9880
rect 4240 9845 4245 9875
rect 4275 9845 4405 9875
rect 4435 9845 4440 9875
rect 4240 9840 4440 9845
rect 4480 9875 4680 9880
rect 4480 9845 4485 9875
rect 4515 9845 4645 9875
rect 4675 9845 4680 9875
rect 4480 9840 4680 9845
rect 4720 9875 5720 9880
rect 4720 9845 4725 9875
rect 4755 9845 4885 9875
rect 4915 9845 5045 9875
rect 5075 9845 5205 9875
rect 5235 9845 5365 9875
rect 5395 9845 5525 9875
rect 5555 9845 5685 9875
rect 5715 9845 5720 9875
rect 4720 9840 5720 9845
rect 5760 9875 5960 9880
rect 5760 9845 5765 9875
rect 5795 9845 5925 9875
rect 5955 9845 5960 9875
rect 5760 9840 5960 9845
rect 6000 9875 6200 9880
rect 6000 9845 6005 9875
rect 6035 9845 6165 9875
rect 6195 9845 6200 9875
rect 6000 9840 6200 9845
rect 4240 9795 4440 9800
rect 4240 9765 4245 9795
rect 4275 9765 4405 9795
rect 4435 9765 4440 9795
rect 4240 9760 4440 9765
rect 4480 9795 4680 9800
rect 4480 9765 4485 9795
rect 4515 9765 4645 9795
rect 4675 9765 4680 9795
rect 4480 9760 4680 9765
rect 4720 9795 5720 9800
rect 4720 9765 4725 9795
rect 4755 9765 4885 9795
rect 4915 9765 5045 9795
rect 5075 9765 5205 9795
rect 5235 9765 5365 9795
rect 5395 9765 5525 9795
rect 5555 9765 5685 9795
rect 5715 9765 5720 9795
rect 4720 9760 5720 9765
rect 5760 9795 5960 9800
rect 5760 9765 5765 9795
rect 5795 9765 5925 9795
rect 5955 9765 5960 9795
rect 5760 9760 5960 9765
rect 6000 9795 6200 9800
rect 6000 9765 6005 9795
rect 6035 9765 6165 9795
rect 6195 9765 6200 9795
rect 6000 9760 6200 9765
rect 4240 9715 4440 9720
rect 4240 9685 4245 9715
rect 4275 9685 4405 9715
rect 4435 9685 4440 9715
rect 4240 9680 4440 9685
rect 4480 9715 4680 9720
rect 4480 9685 4485 9715
rect 4515 9685 4645 9715
rect 4675 9685 4680 9715
rect 4480 9680 4680 9685
rect 4720 9715 5720 9720
rect 4720 9685 4725 9715
rect 4755 9685 4885 9715
rect 4915 9685 5045 9715
rect 5075 9685 5205 9715
rect 5235 9685 5365 9715
rect 5395 9685 5525 9715
rect 5555 9685 5685 9715
rect 5715 9685 5720 9715
rect 4720 9680 5720 9685
rect 5760 9715 5960 9720
rect 5760 9685 5765 9715
rect 5795 9685 5925 9715
rect 5955 9685 5960 9715
rect 5760 9680 5960 9685
rect 6000 9715 6200 9720
rect 6000 9685 6005 9715
rect 6035 9685 6165 9715
rect 6195 9685 6200 9715
rect 6000 9680 6200 9685
rect 4240 9635 4440 9640
rect 4240 9605 4245 9635
rect 4275 9605 4405 9635
rect 4435 9605 4440 9635
rect 4240 9600 4440 9605
rect 4480 9635 4680 9640
rect 4480 9605 4485 9635
rect 4515 9605 4645 9635
rect 4675 9605 4680 9635
rect 4480 9600 4680 9605
rect 4720 9635 5720 9640
rect 4720 9605 4725 9635
rect 4755 9605 4885 9635
rect 4915 9605 5045 9635
rect 5075 9605 5205 9635
rect 5235 9605 5365 9635
rect 5395 9605 5525 9635
rect 5555 9605 5685 9635
rect 5715 9605 5720 9635
rect 4720 9600 5720 9605
rect 5760 9635 5960 9640
rect 5760 9605 5765 9635
rect 5795 9605 5925 9635
rect 5955 9605 5960 9635
rect 5760 9600 5960 9605
rect 6000 9635 6200 9640
rect 6000 9605 6005 9635
rect 6035 9605 6165 9635
rect 6195 9605 6200 9635
rect 6000 9600 6200 9605
rect 4240 9555 4440 9560
rect 4240 9525 4245 9555
rect 4275 9525 4405 9555
rect 4435 9525 4440 9555
rect 4240 9520 4440 9525
rect 4480 9555 4680 9560
rect 4480 9525 4485 9555
rect 4515 9525 4645 9555
rect 4675 9525 4680 9555
rect 4480 9520 4680 9525
rect 4720 9555 5720 9560
rect 4720 9525 4725 9555
rect 4755 9525 4885 9555
rect 4915 9525 5045 9555
rect 5075 9525 5205 9555
rect 5235 9525 5365 9555
rect 5395 9525 5525 9555
rect 5555 9525 5685 9555
rect 5715 9525 5720 9555
rect 4720 9520 5720 9525
rect 5760 9555 5960 9560
rect 5760 9525 5765 9555
rect 5795 9525 5925 9555
rect 5955 9525 5960 9555
rect 5760 9520 5960 9525
rect 6000 9555 6200 9560
rect 6000 9525 6005 9555
rect 6035 9525 6165 9555
rect 6195 9525 6200 9555
rect 6000 9520 6200 9525
rect 4240 9475 4440 9480
rect 4240 9445 4245 9475
rect 4275 9445 4405 9475
rect 4435 9445 4440 9475
rect 4240 9440 4440 9445
rect 4480 9475 4680 9480
rect 4480 9445 4485 9475
rect 4515 9445 4645 9475
rect 4675 9445 4680 9475
rect 4480 9440 4680 9445
rect 4720 9475 5720 9480
rect 4720 9445 4725 9475
rect 4755 9445 4885 9475
rect 4915 9445 5045 9475
rect 5075 9445 5205 9475
rect 5235 9445 5365 9475
rect 5395 9445 5525 9475
rect 5555 9445 5685 9475
rect 5715 9445 5720 9475
rect 4720 9440 5720 9445
rect 5760 9475 5960 9480
rect 5760 9445 5765 9475
rect 5795 9445 5925 9475
rect 5955 9445 5960 9475
rect 5760 9440 5960 9445
rect 6000 9475 6200 9480
rect 6000 9445 6005 9475
rect 6035 9445 6165 9475
rect 6195 9445 6200 9475
rect 6000 9440 6200 9445
rect 4240 9395 4440 9400
rect 4240 9365 4245 9395
rect 4275 9365 4405 9395
rect 4435 9365 4440 9395
rect 4240 9360 4440 9365
rect 4480 9395 4680 9400
rect 4480 9365 4485 9395
rect 4515 9365 4645 9395
rect 4675 9365 4680 9395
rect 4480 9360 4680 9365
rect 4720 9395 5720 9400
rect 4720 9365 4725 9395
rect 4755 9365 4885 9395
rect 4915 9365 5045 9395
rect 5075 9365 5205 9395
rect 5235 9365 5365 9395
rect 5395 9365 5525 9395
rect 5555 9365 5685 9395
rect 5715 9365 5720 9395
rect 4720 9360 5720 9365
rect 5760 9395 5960 9400
rect 5760 9365 5765 9395
rect 5795 9365 5925 9395
rect 5955 9365 5960 9395
rect 5760 9360 5960 9365
rect 6000 9395 6200 9400
rect 6000 9365 6005 9395
rect 6035 9365 6165 9395
rect 6195 9365 6200 9395
rect 6000 9360 6200 9365
rect 0 9275 10440 9280
rect 0 9245 5125 9275
rect 5155 9245 10440 9275
rect 0 9240 10440 9245
rect 0 9115 5000 9120
rect 0 9085 4965 9115
rect 4995 9085 5000 9115
rect 0 9080 5000 9085
rect 5440 9115 10440 9120
rect 5440 9085 5445 9115
rect 5475 9085 10440 9115
rect 5440 9080 10440 9085
rect 4240 8995 4440 9000
rect 4240 8965 4245 8995
rect 4275 8965 4405 8995
rect 4435 8965 4440 8995
rect 4240 8960 4440 8965
rect 4480 8995 4680 9000
rect 4480 8965 4485 8995
rect 4515 8965 4645 8995
rect 4675 8965 4680 8995
rect 4480 8960 4680 8965
rect 4720 8995 5720 9000
rect 4720 8965 4725 8995
rect 4755 8965 4885 8995
rect 4915 8965 5045 8995
rect 5075 8965 5205 8995
rect 5235 8965 5365 8995
rect 5395 8965 5525 8995
rect 5555 8965 5685 8995
rect 5715 8965 5720 8995
rect 4720 8960 5720 8965
rect 5760 8995 5960 9000
rect 5760 8965 5765 8995
rect 5795 8965 5925 8995
rect 5955 8965 5960 8995
rect 5760 8960 5960 8965
rect 6000 8995 6200 9000
rect 6000 8965 6005 8995
rect 6035 8965 6165 8995
rect 6195 8965 6200 8995
rect 6000 8960 6200 8965
rect 4240 8915 4440 8920
rect 4240 8885 4245 8915
rect 4275 8885 4405 8915
rect 4435 8885 4440 8915
rect 4240 8880 4440 8885
rect 4480 8915 4680 8920
rect 4480 8885 4485 8915
rect 4515 8885 4645 8915
rect 4675 8885 4680 8915
rect 4480 8880 4680 8885
rect 4720 8915 5720 8920
rect 4720 8885 4725 8915
rect 4755 8885 4885 8915
rect 4915 8885 5045 8915
rect 5075 8885 5205 8915
rect 5235 8885 5365 8915
rect 5395 8885 5525 8915
rect 5555 8885 5685 8915
rect 5715 8885 5720 8915
rect 4720 8880 5720 8885
rect 5760 8915 5960 8920
rect 5760 8885 5765 8915
rect 5795 8885 5925 8915
rect 5955 8885 5960 8915
rect 5760 8880 5960 8885
rect 6000 8915 6200 8920
rect 6000 8885 6005 8915
rect 6035 8885 6165 8915
rect 6195 8885 6200 8915
rect 6000 8880 6200 8885
rect 4240 8835 4440 8840
rect 4240 8805 4245 8835
rect 4275 8805 4405 8835
rect 4435 8805 4440 8835
rect 4240 8800 4440 8805
rect 4480 8835 4680 8840
rect 4480 8805 4485 8835
rect 4515 8805 4645 8835
rect 4675 8805 4680 8835
rect 4480 8800 4680 8805
rect 4720 8835 5720 8840
rect 4720 8805 4725 8835
rect 4755 8805 4885 8835
rect 4915 8805 5045 8835
rect 5075 8805 5205 8835
rect 5235 8805 5365 8835
rect 5395 8805 5525 8835
rect 5555 8805 5685 8835
rect 5715 8805 5720 8835
rect 4720 8800 5720 8805
rect 5760 8835 5960 8840
rect 5760 8805 5765 8835
rect 5795 8805 5925 8835
rect 5955 8805 5960 8835
rect 5760 8800 5960 8805
rect 6000 8835 6200 8840
rect 6000 8805 6005 8835
rect 6035 8805 6165 8835
rect 6195 8805 6200 8835
rect 6000 8800 6200 8805
rect 4240 8755 4440 8760
rect 4240 8725 4245 8755
rect 4275 8725 4405 8755
rect 4435 8725 4440 8755
rect 4240 8720 4440 8725
rect 4480 8755 4680 8760
rect 4480 8725 4485 8755
rect 4515 8725 4645 8755
rect 4675 8725 4680 8755
rect 4480 8720 4680 8725
rect 4720 8755 5720 8760
rect 4720 8725 4725 8755
rect 4755 8725 4885 8755
rect 4915 8725 5045 8755
rect 5075 8725 5205 8755
rect 5235 8725 5365 8755
rect 5395 8725 5525 8755
rect 5555 8725 5685 8755
rect 5715 8725 5720 8755
rect 4720 8720 5720 8725
rect 5760 8755 5960 8760
rect 5760 8725 5765 8755
rect 5795 8725 5925 8755
rect 5955 8725 5960 8755
rect 5760 8720 5960 8725
rect 6000 8755 6200 8760
rect 6000 8725 6005 8755
rect 6035 8725 6165 8755
rect 6195 8725 6200 8755
rect 6000 8720 6200 8725
rect 4240 8675 4440 8680
rect 4240 8645 4245 8675
rect 4275 8645 4405 8675
rect 4435 8645 4440 8675
rect 4240 8640 4440 8645
rect 4480 8675 4680 8680
rect 4480 8645 4485 8675
rect 4515 8645 4645 8675
rect 4675 8645 4680 8675
rect 4480 8640 4680 8645
rect 4720 8675 5720 8680
rect 4720 8645 4725 8675
rect 4755 8645 4885 8675
rect 4915 8645 5045 8675
rect 5075 8645 5205 8675
rect 5235 8645 5365 8675
rect 5395 8645 5525 8675
rect 5555 8645 5685 8675
rect 5715 8645 5720 8675
rect 4720 8640 5720 8645
rect 5760 8675 5960 8680
rect 5760 8645 5765 8675
rect 5795 8645 5925 8675
rect 5955 8645 5960 8675
rect 5760 8640 5960 8645
rect 6000 8675 6200 8680
rect 6000 8645 6005 8675
rect 6035 8645 6165 8675
rect 6195 8645 6200 8675
rect 6000 8640 6200 8645
rect 4240 8595 4440 8600
rect 4240 8565 4245 8595
rect 4275 8565 4405 8595
rect 4435 8565 4440 8595
rect 4240 8560 4440 8565
rect 4480 8595 4680 8600
rect 4480 8565 4485 8595
rect 4515 8565 4645 8595
rect 4675 8565 4680 8595
rect 4480 8560 4680 8565
rect 4720 8595 5720 8600
rect 4720 8565 4725 8595
rect 4755 8565 4885 8595
rect 4915 8565 5045 8595
rect 5075 8565 5205 8595
rect 5235 8565 5365 8595
rect 5395 8565 5525 8595
rect 5555 8565 5685 8595
rect 5715 8565 5720 8595
rect 4720 8560 5720 8565
rect 5760 8595 5960 8600
rect 5760 8565 5765 8595
rect 5795 8565 5925 8595
rect 5955 8565 5960 8595
rect 5760 8560 5960 8565
rect 6000 8595 6200 8600
rect 6000 8565 6005 8595
rect 6035 8565 6165 8595
rect 6195 8565 6200 8595
rect 6000 8560 6200 8565
rect 4240 8515 4440 8520
rect 4240 8485 4245 8515
rect 4275 8485 4405 8515
rect 4435 8485 4440 8515
rect 4240 8480 4440 8485
rect 4480 8515 4680 8520
rect 4480 8485 4485 8515
rect 4515 8485 4645 8515
rect 4675 8485 4680 8515
rect 4480 8480 4680 8485
rect 4720 8515 5720 8520
rect 4720 8485 4725 8515
rect 4755 8485 4885 8515
rect 4915 8485 5045 8515
rect 5075 8485 5205 8515
rect 5235 8485 5365 8515
rect 5395 8485 5525 8515
rect 5555 8485 5685 8515
rect 5715 8485 5720 8515
rect 4720 8480 5720 8485
rect 5760 8515 5960 8520
rect 5760 8485 5765 8515
rect 5795 8485 5925 8515
rect 5955 8485 5960 8515
rect 5760 8480 5960 8485
rect 6000 8515 6200 8520
rect 6000 8485 6005 8515
rect 6035 8485 6165 8515
rect 6195 8485 6200 8515
rect 6000 8480 6200 8485
rect 4240 8435 4440 8440
rect 4240 8405 4245 8435
rect 4275 8405 4405 8435
rect 4435 8405 4440 8435
rect 4240 8400 4440 8405
rect 4480 8435 4680 8440
rect 4480 8405 4485 8435
rect 4515 8405 4645 8435
rect 4675 8405 4680 8435
rect 4480 8400 4680 8405
rect 4720 8435 5720 8440
rect 4720 8405 4725 8435
rect 4755 8405 4885 8435
rect 4915 8405 5045 8435
rect 5075 8405 5205 8435
rect 5235 8405 5365 8435
rect 5395 8405 5525 8435
rect 5555 8405 5685 8435
rect 5715 8405 5720 8435
rect 4720 8400 5720 8405
rect 5760 8435 5960 8440
rect 5760 8405 5765 8435
rect 5795 8405 5925 8435
rect 5955 8405 5960 8435
rect 5760 8400 5960 8405
rect 6000 8435 6200 8440
rect 6000 8405 6005 8435
rect 6035 8405 6165 8435
rect 6195 8405 6200 8435
rect 6000 8400 6200 8405
rect 0 8355 10440 8360
rect 0 8325 4565 8355
rect 4595 8325 10440 8355
rect 0 8320 10440 8325
rect 4240 8275 4440 8280
rect 4240 8245 4245 8275
rect 4275 8245 4405 8275
rect 4435 8245 4440 8275
rect 4240 8240 4440 8245
rect 4480 8275 4680 8280
rect 4480 8245 4485 8275
rect 4515 8245 4645 8275
rect 4675 8245 4680 8275
rect 4480 8240 4680 8245
rect 4720 8275 5720 8280
rect 4720 8245 4725 8275
rect 4755 8245 4885 8275
rect 4915 8245 5045 8275
rect 5075 8245 5205 8275
rect 5235 8245 5365 8275
rect 5395 8245 5525 8275
rect 5555 8245 5685 8275
rect 5715 8245 5720 8275
rect 4720 8240 5720 8245
rect 5760 8275 5960 8280
rect 5760 8245 5765 8275
rect 5795 8245 5925 8275
rect 5955 8245 5960 8275
rect 5760 8240 5960 8245
rect 6000 8275 6200 8280
rect 6000 8245 6005 8275
rect 6035 8245 6165 8275
rect 6195 8245 6200 8275
rect 6000 8240 6200 8245
rect 4240 8195 4440 8200
rect 4240 8165 4245 8195
rect 4275 8165 4405 8195
rect 4435 8165 4440 8195
rect 4240 8160 4440 8165
rect 4480 8195 4680 8200
rect 4480 8165 4485 8195
rect 4515 8165 4645 8195
rect 4675 8165 4680 8195
rect 4480 8160 4680 8165
rect 4720 8195 5720 8200
rect 4720 8165 4725 8195
rect 4755 8165 4885 8195
rect 4915 8165 5045 8195
rect 5075 8165 5205 8195
rect 5235 8165 5365 8195
rect 5395 8165 5525 8195
rect 5555 8165 5685 8195
rect 5715 8165 5720 8195
rect 4720 8160 5720 8165
rect 5760 8195 5960 8200
rect 5760 8165 5765 8195
rect 5795 8165 5925 8195
rect 5955 8165 5960 8195
rect 5760 8160 5960 8165
rect 6000 8195 6200 8200
rect 6000 8165 6005 8195
rect 6035 8165 6165 8195
rect 6195 8165 6200 8195
rect 6000 8160 6200 8165
rect 4240 8115 4440 8120
rect 4240 8085 4245 8115
rect 4275 8085 4405 8115
rect 4435 8085 4440 8115
rect 4240 8080 4440 8085
rect 4480 8115 4680 8120
rect 4480 8085 4485 8115
rect 4515 8085 4645 8115
rect 4675 8085 4680 8115
rect 4480 8080 4680 8085
rect 4720 8115 5720 8120
rect 4720 8085 4725 8115
rect 4755 8085 4885 8115
rect 4915 8085 5045 8115
rect 5075 8085 5205 8115
rect 5235 8085 5365 8115
rect 5395 8085 5525 8115
rect 5555 8085 5685 8115
rect 5715 8085 5720 8115
rect 4720 8080 5720 8085
rect 5760 8115 5960 8120
rect 5760 8085 5765 8115
rect 5795 8085 5925 8115
rect 5955 8085 5960 8115
rect 5760 8080 5960 8085
rect 6000 8115 6200 8120
rect 6000 8085 6005 8115
rect 6035 8085 6165 8115
rect 6195 8085 6200 8115
rect 6000 8080 6200 8085
rect 4240 8035 4440 8040
rect 4240 8005 4245 8035
rect 4275 8005 4405 8035
rect 4435 8005 4440 8035
rect 4240 8000 4440 8005
rect 4480 8035 4680 8040
rect 4480 8005 4485 8035
rect 4515 8005 4645 8035
rect 4675 8005 4680 8035
rect 4480 8000 4680 8005
rect 4720 8035 5720 8040
rect 4720 8005 4725 8035
rect 4755 8005 4885 8035
rect 4915 8005 5045 8035
rect 5075 8005 5205 8035
rect 5235 8005 5365 8035
rect 5395 8005 5525 8035
rect 5555 8005 5685 8035
rect 5715 8005 5720 8035
rect 4720 8000 5720 8005
rect 5760 8035 5960 8040
rect 5760 8005 5765 8035
rect 5795 8005 5925 8035
rect 5955 8005 5960 8035
rect 5760 8000 5960 8005
rect 6000 8035 6200 8040
rect 6000 8005 6005 8035
rect 6035 8005 6165 8035
rect 6195 8005 6200 8035
rect 6000 8000 6200 8005
rect 4240 7955 4440 7960
rect 4240 7925 4245 7955
rect 4275 7925 4405 7955
rect 4435 7925 4440 7955
rect 4240 7920 4440 7925
rect 4480 7955 4680 7960
rect 4480 7925 4485 7955
rect 4515 7925 4645 7955
rect 4675 7925 4680 7955
rect 4480 7920 4680 7925
rect 4720 7955 5720 7960
rect 4720 7925 4725 7955
rect 4755 7925 4885 7955
rect 4915 7925 5045 7955
rect 5075 7925 5205 7955
rect 5235 7925 5365 7955
rect 5395 7925 5525 7955
rect 5555 7925 5685 7955
rect 5715 7925 5720 7955
rect 4720 7920 5720 7925
rect 5760 7955 5960 7960
rect 5760 7925 5765 7955
rect 5795 7925 5925 7955
rect 5955 7925 5960 7955
rect 5760 7920 5960 7925
rect 6000 7955 6200 7960
rect 6000 7925 6005 7955
rect 6035 7925 6165 7955
rect 6195 7925 6200 7955
rect 6000 7920 6200 7925
rect 4240 7875 4440 7880
rect 4240 7845 4245 7875
rect 4275 7845 4405 7875
rect 4435 7845 4440 7875
rect 4240 7840 4440 7845
rect 4480 7875 4680 7880
rect 4480 7845 4485 7875
rect 4515 7845 4645 7875
rect 4675 7845 4680 7875
rect 4480 7840 4680 7845
rect 4720 7875 5720 7880
rect 4720 7845 4725 7875
rect 4755 7845 4885 7875
rect 4915 7845 5045 7875
rect 5075 7845 5205 7875
rect 5235 7845 5365 7875
rect 5395 7845 5525 7875
rect 5555 7845 5685 7875
rect 5715 7845 5720 7875
rect 4720 7840 5720 7845
rect 5760 7875 5960 7880
rect 5760 7845 5765 7875
rect 5795 7845 5925 7875
rect 5955 7845 5960 7875
rect 5760 7840 5960 7845
rect 6000 7875 6200 7880
rect 6000 7845 6005 7875
rect 6035 7845 6165 7875
rect 6195 7845 6200 7875
rect 6000 7840 6200 7845
rect 4240 7795 4440 7800
rect 4240 7765 4245 7795
rect 4275 7765 4405 7795
rect 4435 7765 4440 7795
rect 4240 7760 4440 7765
rect 4480 7795 4680 7800
rect 4480 7765 4485 7795
rect 4515 7765 4645 7795
rect 4675 7765 4680 7795
rect 4480 7760 4680 7765
rect 4720 7795 5720 7800
rect 4720 7765 4725 7795
rect 4755 7765 4885 7795
rect 4915 7765 5045 7795
rect 5075 7765 5205 7795
rect 5235 7765 5365 7795
rect 5395 7765 5525 7795
rect 5555 7765 5685 7795
rect 5715 7765 5720 7795
rect 4720 7760 5720 7765
rect 5760 7795 5960 7800
rect 5760 7765 5765 7795
rect 5795 7765 5925 7795
rect 5955 7765 5960 7795
rect 5760 7760 5960 7765
rect 6000 7795 6200 7800
rect 6000 7765 6005 7795
rect 6035 7765 6165 7795
rect 6195 7765 6200 7795
rect 6000 7760 6200 7765
rect 4240 7715 4440 7720
rect 4240 7685 4245 7715
rect 4275 7685 4405 7715
rect 4435 7685 4440 7715
rect 4240 7680 4440 7685
rect 4480 7715 4680 7720
rect 4480 7685 4485 7715
rect 4515 7685 4645 7715
rect 4675 7685 4680 7715
rect 4480 7680 4680 7685
rect 4720 7715 5720 7720
rect 4720 7685 4725 7715
rect 4755 7685 4885 7715
rect 4915 7685 5045 7715
rect 5075 7685 5205 7715
rect 5235 7685 5365 7715
rect 5395 7685 5525 7715
rect 5555 7685 5685 7715
rect 5715 7685 5720 7715
rect 4720 7680 5720 7685
rect 5760 7715 5960 7720
rect 5760 7685 5765 7715
rect 5795 7685 5925 7715
rect 5955 7685 5960 7715
rect 5760 7680 5960 7685
rect 6000 7715 6200 7720
rect 6000 7685 6005 7715
rect 6035 7685 6165 7715
rect 6195 7685 6200 7715
rect 6000 7680 6200 7685
rect 4240 7635 4440 7640
rect 4240 7605 4245 7635
rect 4275 7605 4405 7635
rect 4435 7605 4440 7635
rect 4240 7600 4440 7605
rect 4480 7635 4680 7640
rect 4480 7605 4485 7635
rect 4515 7605 4645 7635
rect 4675 7605 4680 7635
rect 4480 7600 4680 7605
rect 4720 7635 5720 7640
rect 4720 7605 4725 7635
rect 4755 7605 4885 7635
rect 4915 7605 5045 7635
rect 5075 7605 5205 7635
rect 5235 7605 5365 7635
rect 5395 7605 5525 7635
rect 5555 7605 5685 7635
rect 5715 7605 5720 7635
rect 4720 7600 5720 7605
rect 5760 7635 5960 7640
rect 5760 7605 5765 7635
rect 5795 7605 5925 7635
rect 5955 7605 5960 7635
rect 5760 7600 5960 7605
rect 6000 7635 6200 7640
rect 6000 7605 6005 7635
rect 6035 7605 6165 7635
rect 6195 7605 6200 7635
rect 6000 7600 6200 7605
rect 4240 7555 4440 7560
rect 4240 7525 4245 7555
rect 4275 7525 4405 7555
rect 4435 7525 4440 7555
rect 4240 7520 4440 7525
rect 4480 7555 4680 7560
rect 4480 7525 4485 7555
rect 4515 7525 4645 7555
rect 4675 7525 4680 7555
rect 4480 7520 4680 7525
rect 4720 7555 5720 7560
rect 4720 7525 4725 7555
rect 4755 7525 4885 7555
rect 4915 7525 5045 7555
rect 5075 7525 5205 7555
rect 5235 7525 5365 7555
rect 5395 7525 5525 7555
rect 5555 7525 5685 7555
rect 5715 7525 5720 7555
rect 4720 7520 5720 7525
rect 5760 7555 5960 7560
rect 5760 7525 5765 7555
rect 5795 7525 5925 7555
rect 5955 7525 5960 7555
rect 5760 7520 5960 7525
rect 6000 7555 6200 7560
rect 6000 7525 6005 7555
rect 6035 7525 6165 7555
rect 6195 7525 6200 7555
rect 6000 7520 6200 7525
rect 4240 7475 4440 7480
rect 4240 7445 4245 7475
rect 4275 7445 4405 7475
rect 4435 7445 4440 7475
rect 4240 7440 4440 7445
rect 4480 7475 4680 7480
rect 4480 7445 4485 7475
rect 4515 7445 4645 7475
rect 4675 7445 4680 7475
rect 4480 7440 4680 7445
rect 4720 7475 5720 7480
rect 4720 7445 4725 7475
rect 4755 7445 4885 7475
rect 4915 7445 5045 7475
rect 5075 7445 5205 7475
rect 5235 7445 5365 7475
rect 5395 7445 5525 7475
rect 5555 7445 5685 7475
rect 5715 7445 5720 7475
rect 4720 7440 5720 7445
rect 5760 7475 5960 7480
rect 5760 7445 5765 7475
rect 5795 7445 5925 7475
rect 5955 7445 5960 7475
rect 5760 7440 5960 7445
rect 6000 7475 6200 7480
rect 6000 7445 6005 7475
rect 6035 7445 6165 7475
rect 6195 7445 6200 7475
rect 6000 7440 6200 7445
rect 4240 7395 4440 7400
rect 4240 7365 4245 7395
rect 4275 7365 4405 7395
rect 4435 7365 4440 7395
rect 4240 7360 4440 7365
rect 4480 7395 4680 7400
rect 4480 7365 4485 7395
rect 4515 7365 4645 7395
rect 4675 7365 4680 7395
rect 4480 7360 4680 7365
rect 4720 7395 5720 7400
rect 4720 7365 4725 7395
rect 4755 7365 4885 7395
rect 4915 7365 5045 7395
rect 5075 7365 5205 7395
rect 5235 7365 5365 7395
rect 5395 7365 5525 7395
rect 5555 7365 5685 7395
rect 5715 7365 5720 7395
rect 4720 7360 5720 7365
rect 5760 7395 5960 7400
rect 5760 7365 5765 7395
rect 5795 7365 5925 7395
rect 5955 7365 5960 7395
rect 5760 7360 5960 7365
rect 6000 7395 6200 7400
rect 6000 7365 6005 7395
rect 6035 7365 6165 7395
rect 6195 7365 6200 7395
rect 6000 7360 6200 7365
rect 4240 7315 4440 7320
rect 4240 7285 4245 7315
rect 4275 7285 4405 7315
rect 4435 7285 4440 7315
rect 4240 7280 4440 7285
rect 4480 7315 4680 7320
rect 4480 7285 4485 7315
rect 4515 7285 4645 7315
rect 4675 7285 4680 7315
rect 4480 7280 4680 7285
rect 4720 7315 5720 7320
rect 4720 7285 4725 7315
rect 4755 7285 4885 7315
rect 4915 7285 5045 7315
rect 5075 7285 5205 7315
rect 5235 7285 5365 7315
rect 5395 7285 5525 7315
rect 5555 7285 5685 7315
rect 5715 7285 5720 7315
rect 4720 7280 5720 7285
rect 5760 7315 5960 7320
rect 5760 7285 5765 7315
rect 5795 7285 5925 7315
rect 5955 7285 5960 7315
rect 5760 7280 5960 7285
rect 6000 7315 6200 7320
rect 6000 7285 6005 7315
rect 6035 7285 6165 7315
rect 6195 7285 6200 7315
rect 6000 7280 6200 7285
rect 4240 7235 4440 7240
rect 4240 7205 4245 7235
rect 4275 7205 4405 7235
rect 4435 7205 4440 7235
rect 4240 7200 4440 7205
rect 4480 7235 4680 7240
rect 4480 7205 4485 7235
rect 4515 7205 4645 7235
rect 4675 7205 4680 7235
rect 4480 7200 4680 7205
rect 4720 7235 5720 7240
rect 4720 7205 4725 7235
rect 4755 7205 4885 7235
rect 4915 7205 5045 7235
rect 5075 7205 5205 7235
rect 5235 7205 5365 7235
rect 5395 7205 5525 7235
rect 5555 7205 5685 7235
rect 5715 7205 5720 7235
rect 4720 7200 5720 7205
rect 5760 7235 5960 7240
rect 5760 7205 5765 7235
rect 5795 7205 5925 7235
rect 5955 7205 5960 7235
rect 5760 7200 5960 7205
rect 6000 7235 6200 7240
rect 6000 7205 6005 7235
rect 6035 7205 6165 7235
rect 6195 7205 6200 7235
rect 6000 7200 6200 7205
rect 4240 7155 4440 7160
rect 4240 7125 4245 7155
rect 4275 7125 4405 7155
rect 4435 7125 4440 7155
rect 4240 7120 4440 7125
rect 4480 7155 4680 7160
rect 4480 7125 4485 7155
rect 4515 7125 4645 7155
rect 4675 7125 4680 7155
rect 4480 7120 4680 7125
rect 4720 7155 5720 7160
rect 4720 7125 4725 7155
rect 4755 7125 4885 7155
rect 4915 7125 5045 7155
rect 5075 7125 5205 7155
rect 5235 7125 5365 7155
rect 5395 7125 5525 7155
rect 5555 7125 5685 7155
rect 5715 7125 5720 7155
rect 4720 7120 5720 7125
rect 5760 7155 5960 7160
rect 5760 7125 5765 7155
rect 5795 7125 5925 7155
rect 5955 7125 5960 7155
rect 5760 7120 5960 7125
rect 6000 7155 6200 7160
rect 6000 7125 6005 7155
rect 6035 7125 6165 7155
rect 6195 7125 6200 7155
rect 6000 7120 6200 7125
rect 4240 7075 4440 7080
rect 4240 7045 4245 7075
rect 4275 7045 4405 7075
rect 4435 7045 4440 7075
rect 4240 7040 4440 7045
rect 4480 7075 4680 7080
rect 4480 7045 4485 7075
rect 4515 7045 4645 7075
rect 4675 7045 4680 7075
rect 4480 7040 4680 7045
rect 4720 7075 5720 7080
rect 4720 7045 4725 7075
rect 4755 7045 4885 7075
rect 4915 7045 5045 7075
rect 5075 7045 5205 7075
rect 5235 7045 5365 7075
rect 5395 7045 5525 7075
rect 5555 7045 5685 7075
rect 5715 7045 5720 7075
rect 4720 7040 5720 7045
rect 5760 7075 5960 7080
rect 5760 7045 5765 7075
rect 5795 7045 5925 7075
rect 5955 7045 5960 7075
rect 5760 7040 5960 7045
rect 6000 7075 6200 7080
rect 6000 7045 6005 7075
rect 6035 7045 6165 7075
rect 6195 7045 6200 7075
rect 6000 7040 6200 7045
rect 4240 6995 4440 7000
rect 4240 6965 4245 6995
rect 4275 6965 4405 6995
rect 4435 6965 4440 6995
rect 4240 6960 4440 6965
rect 4480 6995 4680 7000
rect 4480 6965 4485 6995
rect 4515 6965 4645 6995
rect 4675 6965 4680 6995
rect 4480 6960 4680 6965
rect 4720 6995 5720 7000
rect 4720 6965 4725 6995
rect 4755 6965 4885 6995
rect 4915 6965 5045 6995
rect 5075 6965 5205 6995
rect 5235 6965 5365 6995
rect 5395 6965 5525 6995
rect 5555 6965 5685 6995
rect 5715 6965 5720 6995
rect 4720 6960 5720 6965
rect 5760 6995 5960 7000
rect 5760 6965 5765 6995
rect 5795 6965 5925 6995
rect 5955 6965 5960 6995
rect 5760 6960 5960 6965
rect 6000 6995 6200 7000
rect 6000 6965 6005 6995
rect 6035 6965 6165 6995
rect 6195 6965 6200 6995
rect 6000 6960 6200 6965
rect 0 6915 10440 6920
rect 0 6885 4565 6915
rect 4595 6885 10440 6915
rect 0 6880 10440 6885
rect 4240 6835 4440 6840
rect 4240 6805 4245 6835
rect 4275 6805 4405 6835
rect 4435 6805 4440 6835
rect 4240 6800 4440 6805
rect 4480 6835 4680 6840
rect 4480 6805 4485 6835
rect 4515 6805 4645 6835
rect 4675 6805 4680 6835
rect 4480 6800 4680 6805
rect 4720 6835 5720 6840
rect 4720 6805 4725 6835
rect 4755 6805 4885 6835
rect 4915 6805 5045 6835
rect 5075 6805 5205 6835
rect 5235 6805 5365 6835
rect 5395 6805 5525 6835
rect 5555 6805 5685 6835
rect 5715 6805 5720 6835
rect 4720 6800 5720 6805
rect 5760 6835 5960 6840
rect 5760 6805 5765 6835
rect 5795 6805 5925 6835
rect 5955 6805 5960 6835
rect 5760 6800 5960 6805
rect 6000 6835 6200 6840
rect 6000 6805 6005 6835
rect 6035 6805 6165 6835
rect 6195 6805 6200 6835
rect 6000 6800 6200 6805
rect 4240 6755 4440 6760
rect 4240 6725 4245 6755
rect 4275 6725 4405 6755
rect 4435 6725 4440 6755
rect 4240 6720 4440 6725
rect 4480 6755 4680 6760
rect 4480 6725 4485 6755
rect 4515 6725 4645 6755
rect 4675 6725 4680 6755
rect 4480 6720 4680 6725
rect 4720 6755 5720 6760
rect 4720 6725 4725 6755
rect 4755 6725 4885 6755
rect 4915 6725 5045 6755
rect 5075 6725 5205 6755
rect 5235 6725 5365 6755
rect 5395 6725 5525 6755
rect 5555 6725 5685 6755
rect 5715 6725 5720 6755
rect 4720 6720 5720 6725
rect 5760 6755 5960 6760
rect 5760 6725 5765 6755
rect 5795 6725 5925 6755
rect 5955 6725 5960 6755
rect 5760 6720 5960 6725
rect 6000 6755 6200 6760
rect 6000 6725 6005 6755
rect 6035 6725 6165 6755
rect 6195 6725 6200 6755
rect 6000 6720 6200 6725
rect 4240 6675 4440 6680
rect 4240 6645 4245 6675
rect 4275 6645 4405 6675
rect 4435 6645 4440 6675
rect 4240 6640 4440 6645
rect 4480 6675 4680 6680
rect 4480 6645 4485 6675
rect 4515 6645 4645 6675
rect 4675 6645 4680 6675
rect 4480 6640 4680 6645
rect 4720 6675 5720 6680
rect 4720 6645 4725 6675
rect 4755 6645 4885 6675
rect 4915 6645 5045 6675
rect 5075 6645 5205 6675
rect 5235 6645 5365 6675
rect 5395 6645 5525 6675
rect 5555 6645 5685 6675
rect 5715 6645 5720 6675
rect 4720 6640 5720 6645
rect 5760 6675 5960 6680
rect 5760 6645 5765 6675
rect 5795 6645 5925 6675
rect 5955 6645 5960 6675
rect 5760 6640 5960 6645
rect 6000 6675 6200 6680
rect 6000 6645 6005 6675
rect 6035 6645 6165 6675
rect 6195 6645 6200 6675
rect 6000 6640 6200 6645
rect 4240 6595 4440 6600
rect 4240 6565 4245 6595
rect 4275 6565 4405 6595
rect 4435 6565 4440 6595
rect 4240 6560 4440 6565
rect 4480 6595 4680 6600
rect 4480 6565 4485 6595
rect 4515 6565 4645 6595
rect 4675 6565 4680 6595
rect 4480 6560 4680 6565
rect 4720 6595 5720 6600
rect 4720 6565 4725 6595
rect 4755 6565 4885 6595
rect 4915 6565 5045 6595
rect 5075 6565 5205 6595
rect 5235 6565 5365 6595
rect 5395 6565 5525 6595
rect 5555 6565 5685 6595
rect 5715 6565 5720 6595
rect 4720 6560 5720 6565
rect 5760 6595 5960 6600
rect 5760 6565 5765 6595
rect 5795 6565 5925 6595
rect 5955 6565 5960 6595
rect 5760 6560 5960 6565
rect 6000 6595 6200 6600
rect 6000 6565 6005 6595
rect 6035 6565 6165 6595
rect 6195 6565 6200 6595
rect 6000 6560 6200 6565
rect 4240 6515 4440 6520
rect 4240 6485 4245 6515
rect 4275 6485 4405 6515
rect 4435 6485 4440 6515
rect 4240 6480 4440 6485
rect 4480 6515 4680 6520
rect 4480 6485 4485 6515
rect 4515 6485 4645 6515
rect 4675 6485 4680 6515
rect 4480 6480 4680 6485
rect 4720 6515 5720 6520
rect 4720 6485 4725 6515
rect 4755 6485 4885 6515
rect 4915 6485 5045 6515
rect 5075 6485 5205 6515
rect 5235 6485 5365 6515
rect 5395 6485 5525 6515
rect 5555 6485 5685 6515
rect 5715 6485 5720 6515
rect 4720 6480 5720 6485
rect 5760 6515 5960 6520
rect 5760 6485 5765 6515
rect 5795 6485 5925 6515
rect 5955 6485 5960 6515
rect 5760 6480 5960 6485
rect 6000 6515 6200 6520
rect 6000 6485 6005 6515
rect 6035 6485 6165 6515
rect 6195 6485 6200 6515
rect 6000 6480 6200 6485
rect 4240 6435 4440 6440
rect 4240 6405 4245 6435
rect 4275 6405 4405 6435
rect 4435 6405 4440 6435
rect 4240 6400 4440 6405
rect 4480 6435 4680 6440
rect 4480 6405 4485 6435
rect 4515 6405 4645 6435
rect 4675 6405 4680 6435
rect 4480 6400 4680 6405
rect 4720 6435 5720 6440
rect 4720 6405 4725 6435
rect 4755 6405 4885 6435
rect 4915 6405 5045 6435
rect 5075 6405 5205 6435
rect 5235 6405 5365 6435
rect 5395 6405 5525 6435
rect 5555 6405 5685 6435
rect 5715 6405 5720 6435
rect 4720 6400 5720 6405
rect 5760 6435 5960 6440
rect 5760 6405 5765 6435
rect 5795 6405 5925 6435
rect 5955 6405 5960 6435
rect 5760 6400 5960 6405
rect 6000 6435 6200 6440
rect 6000 6405 6005 6435
rect 6035 6405 6165 6435
rect 6195 6405 6200 6435
rect 6000 6400 6200 6405
rect 4240 6355 4440 6360
rect 4240 6325 4245 6355
rect 4275 6325 4405 6355
rect 4435 6325 4440 6355
rect 4240 6320 4440 6325
rect 4480 6355 4680 6360
rect 4480 6325 4485 6355
rect 4515 6325 4645 6355
rect 4675 6325 4680 6355
rect 4480 6320 4680 6325
rect 4720 6355 5720 6360
rect 4720 6325 4725 6355
rect 4755 6325 4885 6355
rect 4915 6325 5045 6355
rect 5075 6325 5205 6355
rect 5235 6325 5365 6355
rect 5395 6325 5525 6355
rect 5555 6325 5685 6355
rect 5715 6325 5720 6355
rect 4720 6320 5720 6325
rect 5760 6355 5960 6360
rect 5760 6325 5765 6355
rect 5795 6325 5925 6355
rect 5955 6325 5960 6355
rect 5760 6320 5960 6325
rect 6000 6355 6200 6360
rect 6000 6325 6005 6355
rect 6035 6325 6165 6355
rect 6195 6325 6200 6355
rect 6000 6320 6200 6325
rect 4240 6275 4440 6280
rect 4240 6245 4245 6275
rect 4275 6245 4405 6275
rect 4435 6245 4440 6275
rect 4240 6240 4440 6245
rect 4480 6275 4680 6280
rect 4480 6245 4485 6275
rect 4515 6245 4645 6275
rect 4675 6245 4680 6275
rect 4480 6240 4680 6245
rect 4720 6275 5720 6280
rect 4720 6245 4725 6275
rect 4755 6245 4885 6275
rect 4915 6245 5045 6275
rect 5075 6245 5205 6275
rect 5235 6245 5365 6275
rect 5395 6245 5525 6275
rect 5555 6245 5685 6275
rect 5715 6245 5720 6275
rect 4720 6240 5720 6245
rect 5760 6275 5960 6280
rect 5760 6245 5765 6275
rect 5795 6245 5925 6275
rect 5955 6245 5960 6275
rect 5760 6240 5960 6245
rect 6000 6275 6200 6280
rect 6000 6245 6005 6275
rect 6035 6245 6165 6275
rect 6195 6245 6200 6275
rect 6000 6240 6200 6245
rect 0 6155 4840 6160
rect 0 6125 4805 6155
rect 4835 6125 4840 6155
rect 0 6120 4840 6125
rect 5600 6155 10440 6160
rect 5600 6125 5605 6155
rect 5635 6125 10440 6155
rect 5600 6120 10440 6125
rect 0 5995 5000 6000
rect 0 5965 4965 5995
rect 4995 5965 5000 5995
rect 0 5960 5000 5965
rect 5440 5995 10440 6000
rect 5440 5965 5445 5995
rect 5475 5965 10440 5995
rect 5440 5960 10440 5965
rect 4240 5875 4440 5880
rect 4240 5845 4245 5875
rect 4275 5845 4405 5875
rect 4435 5845 4440 5875
rect 4240 5840 4440 5845
rect 4480 5875 4680 5880
rect 4480 5845 4485 5875
rect 4515 5845 4645 5875
rect 4675 5845 4680 5875
rect 4480 5840 4680 5845
rect 4720 5875 5720 5880
rect 4720 5845 4725 5875
rect 4755 5845 4885 5875
rect 4915 5845 5045 5875
rect 5075 5845 5205 5875
rect 5235 5845 5365 5875
rect 5395 5845 5525 5875
rect 5555 5845 5685 5875
rect 5715 5845 5720 5875
rect 4720 5840 5720 5845
rect 5760 5875 5960 5880
rect 5760 5845 5765 5875
rect 5795 5845 5925 5875
rect 5955 5845 5960 5875
rect 5760 5840 5960 5845
rect 6000 5875 6200 5880
rect 6000 5845 6005 5875
rect 6035 5845 6165 5875
rect 6195 5845 6200 5875
rect 6000 5840 6200 5845
rect 4240 5795 4440 5800
rect 4240 5765 4245 5795
rect 4275 5765 4405 5795
rect 4435 5765 4440 5795
rect 4240 5760 4440 5765
rect 4480 5795 4680 5800
rect 4480 5765 4485 5795
rect 4515 5765 4645 5795
rect 4675 5765 4680 5795
rect 4480 5760 4680 5765
rect 4720 5795 5720 5800
rect 4720 5765 4725 5795
rect 4755 5765 4885 5795
rect 4915 5765 5045 5795
rect 5075 5765 5205 5795
rect 5235 5765 5365 5795
rect 5395 5765 5525 5795
rect 5555 5765 5685 5795
rect 5715 5765 5720 5795
rect 4720 5760 5720 5765
rect 5760 5795 5960 5800
rect 5760 5765 5765 5795
rect 5795 5765 5925 5795
rect 5955 5765 5960 5795
rect 5760 5760 5960 5765
rect 6000 5795 6200 5800
rect 6000 5765 6005 5795
rect 6035 5765 6165 5795
rect 6195 5765 6200 5795
rect 6000 5760 6200 5765
rect 4240 5715 4440 5720
rect 4240 5685 4245 5715
rect 4275 5685 4405 5715
rect 4435 5685 4440 5715
rect 4240 5680 4440 5685
rect 4480 5715 4680 5720
rect 4480 5685 4485 5715
rect 4515 5685 4645 5715
rect 4675 5685 4680 5715
rect 4480 5680 4680 5685
rect 4720 5715 5720 5720
rect 4720 5685 4725 5715
rect 4755 5685 4885 5715
rect 4915 5685 5045 5715
rect 5075 5685 5205 5715
rect 5235 5685 5365 5715
rect 5395 5685 5525 5715
rect 5555 5685 5685 5715
rect 5715 5685 5720 5715
rect 4720 5680 5720 5685
rect 5760 5715 5960 5720
rect 5760 5685 5765 5715
rect 5795 5685 5925 5715
rect 5955 5685 5960 5715
rect 5760 5680 5960 5685
rect 6000 5715 6200 5720
rect 6000 5685 6005 5715
rect 6035 5685 6165 5715
rect 6195 5685 6200 5715
rect 6000 5680 6200 5685
rect 4240 5635 4440 5640
rect 4240 5605 4245 5635
rect 4275 5605 4405 5635
rect 4435 5605 4440 5635
rect 4240 5600 4440 5605
rect 4480 5635 4680 5640
rect 4480 5605 4485 5635
rect 4515 5605 4645 5635
rect 4675 5605 4680 5635
rect 4480 5600 4680 5605
rect 4720 5635 5720 5640
rect 4720 5605 4725 5635
rect 4755 5605 4885 5635
rect 4915 5605 5045 5635
rect 5075 5605 5205 5635
rect 5235 5605 5365 5635
rect 5395 5605 5525 5635
rect 5555 5605 5685 5635
rect 5715 5605 5720 5635
rect 4720 5600 5720 5605
rect 5760 5635 5960 5640
rect 5760 5605 5765 5635
rect 5795 5605 5925 5635
rect 5955 5605 5960 5635
rect 5760 5600 5960 5605
rect 6000 5635 6200 5640
rect 6000 5605 6005 5635
rect 6035 5605 6165 5635
rect 6195 5605 6200 5635
rect 6000 5600 6200 5605
rect 4240 5555 4440 5560
rect 4240 5525 4245 5555
rect 4275 5525 4405 5555
rect 4435 5525 4440 5555
rect 4240 5520 4440 5525
rect 4480 5555 4680 5560
rect 4480 5525 4485 5555
rect 4515 5525 4645 5555
rect 4675 5525 4680 5555
rect 4480 5520 4680 5525
rect 4720 5555 5720 5560
rect 4720 5525 4725 5555
rect 4755 5525 4885 5555
rect 4915 5525 5045 5555
rect 5075 5525 5205 5555
rect 5235 5525 5365 5555
rect 5395 5525 5525 5555
rect 5555 5525 5685 5555
rect 5715 5525 5720 5555
rect 4720 5520 5720 5525
rect 5760 5555 5960 5560
rect 5760 5525 5765 5555
rect 5795 5525 5925 5555
rect 5955 5525 5960 5555
rect 5760 5520 5960 5525
rect 6000 5555 6200 5560
rect 6000 5525 6005 5555
rect 6035 5525 6165 5555
rect 6195 5525 6200 5555
rect 6000 5520 6200 5525
rect 4240 5475 4440 5480
rect 4240 5445 4245 5475
rect 4275 5445 4405 5475
rect 4435 5445 4440 5475
rect 4240 5440 4440 5445
rect 4480 5475 4680 5480
rect 4480 5445 4485 5475
rect 4515 5445 4645 5475
rect 4675 5445 4680 5475
rect 4480 5440 4680 5445
rect 4720 5475 5720 5480
rect 4720 5445 4725 5475
rect 4755 5445 4885 5475
rect 4915 5445 5045 5475
rect 5075 5445 5205 5475
rect 5235 5445 5365 5475
rect 5395 5445 5525 5475
rect 5555 5445 5685 5475
rect 5715 5445 5720 5475
rect 4720 5440 5720 5445
rect 5760 5475 5960 5480
rect 5760 5445 5765 5475
rect 5795 5445 5925 5475
rect 5955 5445 5960 5475
rect 5760 5440 5960 5445
rect 6000 5475 6200 5480
rect 6000 5445 6005 5475
rect 6035 5445 6165 5475
rect 6195 5445 6200 5475
rect 6000 5440 6200 5445
rect 4240 5395 4440 5400
rect 4240 5365 4245 5395
rect 4275 5365 4405 5395
rect 4435 5365 4440 5395
rect 4240 5360 4440 5365
rect 4480 5395 4680 5400
rect 4480 5365 4485 5395
rect 4515 5365 4645 5395
rect 4675 5365 4680 5395
rect 4480 5360 4680 5365
rect 4720 5395 5720 5400
rect 4720 5365 4725 5395
rect 4755 5365 4885 5395
rect 4915 5365 5045 5395
rect 5075 5365 5205 5395
rect 5235 5365 5365 5395
rect 5395 5365 5525 5395
rect 5555 5365 5685 5395
rect 5715 5365 5720 5395
rect 4720 5360 5720 5365
rect 5760 5395 5960 5400
rect 5760 5365 5765 5395
rect 5795 5365 5925 5395
rect 5955 5365 5960 5395
rect 5760 5360 5960 5365
rect 6000 5395 6200 5400
rect 6000 5365 6005 5395
rect 6035 5365 6165 5395
rect 6195 5365 6200 5395
rect 6000 5360 6200 5365
rect 4240 5315 4440 5320
rect 4240 5285 4245 5315
rect 4275 5285 4405 5315
rect 4435 5285 4440 5315
rect 4240 5280 4440 5285
rect 4480 5315 4680 5320
rect 4480 5285 4485 5315
rect 4515 5285 4645 5315
rect 4675 5285 4680 5315
rect 4480 5280 4680 5285
rect 4720 5315 5720 5320
rect 4720 5285 4725 5315
rect 4755 5285 4885 5315
rect 4915 5285 5045 5315
rect 5075 5285 5205 5315
rect 5235 5285 5365 5315
rect 5395 5285 5525 5315
rect 5555 5285 5685 5315
rect 5715 5285 5720 5315
rect 4720 5280 5720 5285
rect 5760 5315 5960 5320
rect 5760 5285 5765 5315
rect 5795 5285 5925 5315
rect 5955 5285 5960 5315
rect 5760 5280 5960 5285
rect 6000 5315 6200 5320
rect 6000 5285 6005 5315
rect 6035 5285 6165 5315
rect 6195 5285 6200 5315
rect 6000 5280 6200 5285
rect 4240 5235 4440 5240
rect 4240 5205 4245 5235
rect 4275 5205 4405 5235
rect 4435 5205 4440 5235
rect 4240 5200 4440 5205
rect 4480 5235 4680 5240
rect 4480 5205 4485 5235
rect 4515 5205 4645 5235
rect 4675 5205 4680 5235
rect 4480 5200 4680 5205
rect 4720 5235 5720 5240
rect 4720 5205 4725 5235
rect 4755 5205 4885 5235
rect 4915 5205 5045 5235
rect 5075 5205 5205 5235
rect 5235 5205 5365 5235
rect 5395 5205 5525 5235
rect 5555 5205 5685 5235
rect 5715 5205 5720 5235
rect 4720 5200 5720 5205
rect 5760 5235 5960 5240
rect 5760 5205 5765 5235
rect 5795 5205 5925 5235
rect 5955 5205 5960 5235
rect 5760 5200 5960 5205
rect 6000 5235 6200 5240
rect 6000 5205 6005 5235
rect 6035 5205 6165 5235
rect 6195 5205 6200 5235
rect 6000 5200 6200 5205
rect 4240 5155 4440 5160
rect 4240 5125 4245 5155
rect 4275 5125 4405 5155
rect 4435 5125 4440 5155
rect 4240 5120 4440 5125
rect 4480 5155 4680 5160
rect 4480 5125 4485 5155
rect 4515 5125 4645 5155
rect 4675 5125 4680 5155
rect 4480 5120 4680 5125
rect 4720 5155 5720 5160
rect 4720 5125 4725 5155
rect 4755 5125 4885 5155
rect 4915 5125 5045 5155
rect 5075 5125 5205 5155
rect 5235 5125 5365 5155
rect 5395 5125 5525 5155
rect 5555 5125 5685 5155
rect 5715 5125 5720 5155
rect 4720 5120 5720 5125
rect 5760 5155 5960 5160
rect 5760 5125 5765 5155
rect 5795 5125 5925 5155
rect 5955 5125 5960 5155
rect 5760 5120 5960 5125
rect 6000 5155 6200 5160
rect 6000 5125 6005 5155
rect 6035 5125 6165 5155
rect 6195 5125 6200 5155
rect 6000 5120 6200 5125
rect 4240 5075 4440 5080
rect 4240 5045 4245 5075
rect 4275 5045 4405 5075
rect 4435 5045 4440 5075
rect 4240 5040 4440 5045
rect 4480 5075 4680 5080
rect 4480 5045 4485 5075
rect 4515 5045 4645 5075
rect 4675 5045 4680 5075
rect 4480 5040 4680 5045
rect 4720 5075 5720 5080
rect 4720 5045 4725 5075
rect 4755 5045 4885 5075
rect 4915 5045 5045 5075
rect 5075 5045 5205 5075
rect 5235 5045 5365 5075
rect 5395 5045 5525 5075
rect 5555 5045 5685 5075
rect 5715 5045 5720 5075
rect 4720 5040 5720 5045
rect 5760 5075 5960 5080
rect 5760 5045 5765 5075
rect 5795 5045 5925 5075
rect 5955 5045 5960 5075
rect 5760 5040 5960 5045
rect 6000 5075 6200 5080
rect 6000 5045 6005 5075
rect 6035 5045 6165 5075
rect 6195 5045 6200 5075
rect 6000 5040 6200 5045
rect 4240 4995 4440 5000
rect 4240 4965 4245 4995
rect 4275 4965 4405 4995
rect 4435 4965 4440 4995
rect 4240 4960 4440 4965
rect 4480 4995 4680 5000
rect 4480 4965 4485 4995
rect 4515 4965 4645 4995
rect 4675 4965 4680 4995
rect 4480 4960 4680 4965
rect 4720 4995 5720 5000
rect 4720 4965 4725 4995
rect 4755 4965 4885 4995
rect 4915 4965 5045 4995
rect 5075 4965 5205 4995
rect 5235 4965 5365 4995
rect 5395 4965 5525 4995
rect 5555 4965 5685 4995
rect 5715 4965 5720 4995
rect 4720 4960 5720 4965
rect 5760 4995 5960 5000
rect 5760 4965 5765 4995
rect 5795 4965 5925 4995
rect 5955 4965 5960 4995
rect 5760 4960 5960 4965
rect 6000 4995 6200 5000
rect 6000 4965 6005 4995
rect 6035 4965 6165 4995
rect 6195 4965 6200 4995
rect 6000 4960 6200 4965
rect 4240 4915 4440 4920
rect 4240 4885 4245 4915
rect 4275 4885 4405 4915
rect 4435 4885 4440 4915
rect 4240 4880 4440 4885
rect 4480 4915 4680 4920
rect 4480 4885 4485 4915
rect 4515 4885 4645 4915
rect 4675 4885 4680 4915
rect 4480 4880 4680 4885
rect 4720 4915 5720 4920
rect 4720 4885 4725 4915
rect 4755 4885 4885 4915
rect 4915 4885 5045 4915
rect 5075 4885 5205 4915
rect 5235 4885 5365 4915
rect 5395 4885 5525 4915
rect 5555 4885 5685 4915
rect 5715 4885 5720 4915
rect 4720 4880 5720 4885
rect 5760 4915 5960 4920
rect 5760 4885 5765 4915
rect 5795 4885 5925 4915
rect 5955 4885 5960 4915
rect 5760 4880 5960 4885
rect 6000 4915 6200 4920
rect 6000 4885 6005 4915
rect 6035 4885 6165 4915
rect 6195 4885 6200 4915
rect 6000 4880 6200 4885
rect 0 4835 10440 4840
rect 0 4805 5845 4835
rect 5875 4805 10440 4835
rect 0 4800 10440 4805
rect 4240 4755 4440 4760
rect 4240 4725 4245 4755
rect 4275 4725 4405 4755
rect 4435 4725 4440 4755
rect 4240 4720 4440 4725
rect 4480 4755 4680 4760
rect 4480 4725 4485 4755
rect 4515 4725 4645 4755
rect 4675 4725 4680 4755
rect 4480 4720 4680 4725
rect 4720 4755 5720 4760
rect 4720 4725 4725 4755
rect 4755 4725 4885 4755
rect 4915 4725 5045 4755
rect 5075 4725 5205 4755
rect 5235 4725 5365 4755
rect 5395 4725 5525 4755
rect 5555 4725 5685 4755
rect 5715 4725 5720 4755
rect 4720 4720 5720 4725
rect 5760 4755 5960 4760
rect 5760 4725 5765 4755
rect 5795 4725 5925 4755
rect 5955 4725 5960 4755
rect 5760 4720 5960 4725
rect 6000 4755 6200 4760
rect 6000 4725 6005 4755
rect 6035 4725 6165 4755
rect 6195 4725 6200 4755
rect 6000 4720 6200 4725
rect 4240 4675 4440 4680
rect 4240 4645 4245 4675
rect 4275 4645 4405 4675
rect 4435 4645 4440 4675
rect 4240 4640 4440 4645
rect 4480 4675 4680 4680
rect 4480 4645 4485 4675
rect 4515 4645 4645 4675
rect 4675 4645 4680 4675
rect 4480 4640 4680 4645
rect 4720 4675 5720 4680
rect 4720 4645 4725 4675
rect 4755 4645 4885 4675
rect 4915 4645 5045 4675
rect 5075 4645 5205 4675
rect 5235 4645 5365 4675
rect 5395 4645 5525 4675
rect 5555 4645 5685 4675
rect 5715 4645 5720 4675
rect 4720 4640 5720 4645
rect 5760 4675 5960 4680
rect 5760 4645 5765 4675
rect 5795 4645 5925 4675
rect 5955 4645 5960 4675
rect 5760 4640 5960 4645
rect 6000 4675 6200 4680
rect 6000 4645 6005 4675
rect 6035 4645 6165 4675
rect 6195 4645 6200 4675
rect 6000 4640 6200 4645
rect 0 4595 10440 4600
rect 0 4565 6085 4595
rect 6115 4565 10440 4595
rect 0 4560 10440 4565
rect 4240 4515 4440 4520
rect 4240 4485 4245 4515
rect 4275 4485 4405 4515
rect 4435 4485 4440 4515
rect 4240 4480 4440 4485
rect 4480 4515 4680 4520
rect 4480 4485 4485 4515
rect 4515 4485 4645 4515
rect 4675 4485 4680 4515
rect 4480 4480 4680 4485
rect 4720 4515 5720 4520
rect 4720 4485 4725 4515
rect 4755 4485 4885 4515
rect 4915 4485 5045 4515
rect 5075 4485 5205 4515
rect 5235 4485 5365 4515
rect 5395 4485 5525 4515
rect 5555 4485 5685 4515
rect 5715 4485 5720 4515
rect 4720 4480 5720 4485
rect 5760 4515 5960 4520
rect 5760 4485 5765 4515
rect 5795 4485 5925 4515
rect 5955 4485 5960 4515
rect 5760 4480 5960 4485
rect 6000 4515 6200 4520
rect 6000 4485 6005 4515
rect 6035 4485 6165 4515
rect 6195 4485 6200 4515
rect 6000 4480 6200 4485
rect 4240 4435 4440 4440
rect 4240 4405 4245 4435
rect 4275 4405 4405 4435
rect 4435 4405 4440 4435
rect 4240 4400 4440 4405
rect 4480 4435 4680 4440
rect 4480 4405 4485 4435
rect 4515 4405 4645 4435
rect 4675 4405 4680 4435
rect 4480 4400 4680 4405
rect 4720 4435 5720 4440
rect 4720 4405 4725 4435
rect 4755 4405 4885 4435
rect 4915 4405 5045 4435
rect 5075 4405 5205 4435
rect 5235 4405 5365 4435
rect 5395 4405 5525 4435
rect 5555 4405 5685 4435
rect 5715 4405 5720 4435
rect 4720 4400 5720 4405
rect 5760 4435 5960 4440
rect 5760 4405 5765 4435
rect 5795 4405 5925 4435
rect 5955 4405 5960 4435
rect 5760 4400 5960 4405
rect 6000 4435 6200 4440
rect 6000 4405 6005 4435
rect 6035 4405 6165 4435
rect 6195 4405 6200 4435
rect 6000 4400 6200 4405
rect 4240 4355 4440 4360
rect 4240 4325 4245 4355
rect 4275 4325 4405 4355
rect 4435 4325 4440 4355
rect 4240 4320 4440 4325
rect 4480 4355 4680 4360
rect 4480 4325 4485 4355
rect 4515 4325 4645 4355
rect 4675 4325 4680 4355
rect 4480 4320 4680 4325
rect 4720 4355 5720 4360
rect 4720 4325 4725 4355
rect 4755 4325 4885 4355
rect 4915 4325 5045 4355
rect 5075 4325 5205 4355
rect 5235 4325 5365 4355
rect 5395 4325 5525 4355
rect 5555 4325 5685 4355
rect 5715 4325 5720 4355
rect 4720 4320 5720 4325
rect 5760 4355 5960 4360
rect 5760 4325 5765 4355
rect 5795 4325 5925 4355
rect 5955 4325 5960 4355
rect 5760 4320 5960 4325
rect 6000 4355 6200 4360
rect 6000 4325 6005 4355
rect 6035 4325 6165 4355
rect 6195 4325 6200 4355
rect 6000 4320 6200 4325
rect 4240 4275 4440 4280
rect 4240 4245 4245 4275
rect 4275 4245 4405 4275
rect 4435 4245 4440 4275
rect 4240 4240 4440 4245
rect 4480 4275 4680 4280
rect 4480 4245 4485 4275
rect 4515 4245 4645 4275
rect 4675 4245 4680 4275
rect 4480 4240 4680 4245
rect 4720 4275 5720 4280
rect 4720 4245 4725 4275
rect 4755 4245 4885 4275
rect 4915 4245 5045 4275
rect 5075 4245 5205 4275
rect 5235 4245 5365 4275
rect 5395 4245 5525 4275
rect 5555 4245 5685 4275
rect 5715 4245 5720 4275
rect 4720 4240 5720 4245
rect 5760 4275 5960 4280
rect 5760 4245 5765 4275
rect 5795 4245 5925 4275
rect 5955 4245 5960 4275
rect 5760 4240 5960 4245
rect 6000 4275 6200 4280
rect 6000 4245 6005 4275
rect 6035 4245 6165 4275
rect 6195 4245 6200 4275
rect 6000 4240 6200 4245
rect 4240 4195 4440 4200
rect 4240 4165 4245 4195
rect 4275 4165 4405 4195
rect 4435 4165 4440 4195
rect 4240 4160 4440 4165
rect 4480 4195 4680 4200
rect 4480 4165 4485 4195
rect 4515 4165 4645 4195
rect 4675 4165 4680 4195
rect 4480 4160 4680 4165
rect 4720 4195 5720 4200
rect 4720 4165 4725 4195
rect 4755 4165 4885 4195
rect 4915 4165 5045 4195
rect 5075 4165 5205 4195
rect 5235 4165 5365 4195
rect 5395 4165 5525 4195
rect 5555 4165 5685 4195
rect 5715 4165 5720 4195
rect 4720 4160 5720 4165
rect 5760 4195 5960 4200
rect 5760 4165 5765 4195
rect 5795 4165 5925 4195
rect 5955 4165 5960 4195
rect 5760 4160 5960 4165
rect 6000 4195 6200 4200
rect 6000 4165 6005 4195
rect 6035 4165 6165 4195
rect 6195 4165 6200 4195
rect 6000 4160 6200 4165
rect 4240 4115 4440 4120
rect 4240 4085 4245 4115
rect 4275 4085 4405 4115
rect 4435 4085 4440 4115
rect 4240 4080 4440 4085
rect 4480 4115 4680 4120
rect 4480 4085 4485 4115
rect 4515 4085 4645 4115
rect 4675 4085 4680 4115
rect 4480 4080 4680 4085
rect 4720 4115 5720 4120
rect 4720 4085 4725 4115
rect 4755 4085 4885 4115
rect 4915 4085 5045 4115
rect 5075 4085 5205 4115
rect 5235 4085 5365 4115
rect 5395 4085 5525 4115
rect 5555 4085 5685 4115
rect 5715 4085 5720 4115
rect 4720 4080 5720 4085
rect 5760 4115 5960 4120
rect 5760 4085 5765 4115
rect 5795 4085 5925 4115
rect 5955 4085 5960 4115
rect 5760 4080 5960 4085
rect 6000 4115 6200 4120
rect 6000 4085 6005 4115
rect 6035 4085 6165 4115
rect 6195 4085 6200 4115
rect 6000 4080 6200 4085
rect 4240 4035 4440 4040
rect 4240 4005 4245 4035
rect 4275 4005 4405 4035
rect 4435 4005 4440 4035
rect 4240 4000 4440 4005
rect 4480 4035 4680 4040
rect 4480 4005 4485 4035
rect 4515 4005 4645 4035
rect 4675 4005 4680 4035
rect 4480 4000 4680 4005
rect 4720 4035 5720 4040
rect 4720 4005 4725 4035
rect 4755 4005 4885 4035
rect 4915 4005 5045 4035
rect 5075 4005 5205 4035
rect 5235 4005 5365 4035
rect 5395 4005 5525 4035
rect 5555 4005 5685 4035
rect 5715 4005 5720 4035
rect 4720 4000 5720 4005
rect 5760 4035 5960 4040
rect 5760 4005 5765 4035
rect 5795 4005 5925 4035
rect 5955 4005 5960 4035
rect 5760 4000 5960 4005
rect 6000 4035 6200 4040
rect 6000 4005 6005 4035
rect 6035 4005 6165 4035
rect 6195 4005 6200 4035
rect 6000 4000 6200 4005
rect 4240 3955 4440 3960
rect 4240 3925 4245 3955
rect 4275 3925 4405 3955
rect 4435 3925 4440 3955
rect 4240 3920 4440 3925
rect 4480 3955 4680 3960
rect 4480 3925 4485 3955
rect 4515 3925 4645 3955
rect 4675 3925 4680 3955
rect 4480 3920 4680 3925
rect 4720 3955 5720 3960
rect 4720 3925 4725 3955
rect 4755 3925 4885 3955
rect 4915 3925 5045 3955
rect 5075 3925 5205 3955
rect 5235 3925 5365 3955
rect 5395 3925 5525 3955
rect 5555 3925 5685 3955
rect 5715 3925 5720 3955
rect 4720 3920 5720 3925
rect 5760 3955 5960 3960
rect 5760 3925 5765 3955
rect 5795 3925 5925 3955
rect 5955 3925 5960 3955
rect 5760 3920 5960 3925
rect 6000 3955 6200 3960
rect 6000 3925 6005 3955
rect 6035 3925 6165 3955
rect 6195 3925 6200 3955
rect 6000 3920 6200 3925
rect 4240 3875 4440 3880
rect 4240 3845 4245 3875
rect 4275 3845 4405 3875
rect 4435 3845 4440 3875
rect 4240 3840 4440 3845
rect 4480 3875 4680 3880
rect 4480 3845 4485 3875
rect 4515 3845 4645 3875
rect 4675 3845 4680 3875
rect 4480 3840 4680 3845
rect 4720 3875 5720 3880
rect 4720 3845 4725 3875
rect 4755 3845 4885 3875
rect 4915 3845 5045 3875
rect 5075 3845 5205 3875
rect 5235 3845 5365 3875
rect 5395 3845 5525 3875
rect 5555 3845 5685 3875
rect 5715 3845 5720 3875
rect 4720 3840 5720 3845
rect 5760 3875 5960 3880
rect 5760 3845 5765 3875
rect 5795 3845 5925 3875
rect 5955 3845 5960 3875
rect 5760 3840 5960 3845
rect 6000 3875 6200 3880
rect 6000 3845 6005 3875
rect 6035 3845 6165 3875
rect 6195 3845 6200 3875
rect 6000 3840 6200 3845
rect 0 3795 10440 3800
rect 0 3765 4325 3795
rect 4355 3765 10440 3795
rect 0 3760 10440 3765
rect 4240 3715 4440 3720
rect 4240 3685 4245 3715
rect 4275 3685 4405 3715
rect 4435 3685 4440 3715
rect 4240 3680 4440 3685
rect 4480 3715 4680 3720
rect 4480 3685 4485 3715
rect 4515 3685 4645 3715
rect 4675 3685 4680 3715
rect 4480 3680 4680 3685
rect 4720 3715 5720 3720
rect 4720 3685 4725 3715
rect 4755 3685 4885 3715
rect 4915 3685 5045 3715
rect 5075 3685 5205 3715
rect 5235 3685 5365 3715
rect 5395 3685 5525 3715
rect 5555 3685 5685 3715
rect 5715 3685 5720 3715
rect 4720 3680 5720 3685
rect 5760 3715 5960 3720
rect 5760 3685 5765 3715
rect 5795 3685 5925 3715
rect 5955 3685 5960 3715
rect 5760 3680 5960 3685
rect 6000 3715 6200 3720
rect 6000 3685 6005 3715
rect 6035 3685 6165 3715
rect 6195 3685 6200 3715
rect 6000 3680 6200 3685
rect 4240 3635 4440 3640
rect 4240 3605 4245 3635
rect 4275 3605 4405 3635
rect 4435 3605 4440 3635
rect 4240 3600 4440 3605
rect 4480 3635 4680 3640
rect 4480 3605 4485 3635
rect 4515 3605 4645 3635
rect 4675 3605 4680 3635
rect 4480 3600 4680 3605
rect 4720 3635 5720 3640
rect 4720 3605 4725 3635
rect 4755 3605 4885 3635
rect 4915 3605 5045 3635
rect 5075 3605 5205 3635
rect 5235 3605 5365 3635
rect 5395 3605 5525 3635
rect 5555 3605 5685 3635
rect 5715 3605 5720 3635
rect 4720 3600 5720 3605
rect 5760 3635 5960 3640
rect 5760 3605 5765 3635
rect 5795 3605 5925 3635
rect 5955 3605 5960 3635
rect 5760 3600 5960 3605
rect 6000 3635 6200 3640
rect 6000 3605 6005 3635
rect 6035 3605 6165 3635
rect 6195 3605 6200 3635
rect 6000 3600 6200 3605
rect 0 3555 10440 3560
rect 0 3525 4565 3555
rect 4595 3525 10440 3555
rect 0 3520 10440 3525
rect 4240 3475 4440 3480
rect 4240 3445 4245 3475
rect 4275 3445 4405 3475
rect 4435 3445 4440 3475
rect 4240 3440 4440 3445
rect 4480 3475 4680 3480
rect 4480 3445 4485 3475
rect 4515 3445 4645 3475
rect 4675 3445 4680 3475
rect 4480 3440 4680 3445
rect 4720 3475 5720 3480
rect 4720 3445 4725 3475
rect 4755 3445 4885 3475
rect 4915 3445 5045 3475
rect 5075 3445 5205 3475
rect 5235 3445 5365 3475
rect 5395 3445 5525 3475
rect 5555 3445 5685 3475
rect 5715 3445 5720 3475
rect 4720 3440 5720 3445
rect 5760 3475 5960 3480
rect 5760 3445 5765 3475
rect 5795 3445 5925 3475
rect 5955 3445 5960 3475
rect 5760 3440 5960 3445
rect 6000 3475 6200 3480
rect 6000 3445 6005 3475
rect 6035 3445 6165 3475
rect 6195 3445 6200 3475
rect 6000 3440 6200 3445
rect 4240 3395 4440 3400
rect 4240 3365 4245 3395
rect 4275 3365 4405 3395
rect 4435 3365 4440 3395
rect 4240 3360 4440 3365
rect 4480 3395 4680 3400
rect 4480 3365 4485 3395
rect 4515 3365 4645 3395
rect 4675 3365 4680 3395
rect 4480 3360 4680 3365
rect 4720 3395 5720 3400
rect 4720 3365 4725 3395
rect 4755 3365 4885 3395
rect 4915 3365 5045 3395
rect 5075 3365 5205 3395
rect 5235 3365 5365 3395
rect 5395 3365 5525 3395
rect 5555 3365 5685 3395
rect 5715 3365 5720 3395
rect 4720 3360 5720 3365
rect 5760 3395 5960 3400
rect 5760 3365 5765 3395
rect 5795 3365 5925 3395
rect 5955 3365 5960 3395
rect 5760 3360 5960 3365
rect 6000 3395 6200 3400
rect 6000 3365 6005 3395
rect 6035 3365 6165 3395
rect 6195 3365 6200 3395
rect 6000 3360 6200 3365
rect 0 3315 10440 3320
rect 0 3285 5845 3315
rect 5875 3285 10440 3315
rect 0 3280 10440 3285
rect 4240 3235 4440 3240
rect 4240 3205 4245 3235
rect 4275 3205 4405 3235
rect 4435 3205 4440 3235
rect 4240 3200 4440 3205
rect 4480 3235 4680 3240
rect 4480 3205 4485 3235
rect 4515 3205 4645 3235
rect 4675 3205 4680 3235
rect 4480 3200 4680 3205
rect 4720 3235 5720 3240
rect 4720 3205 4725 3235
rect 4755 3205 4885 3235
rect 4915 3205 5045 3235
rect 5075 3205 5205 3235
rect 5235 3205 5365 3235
rect 5395 3205 5525 3235
rect 5555 3205 5685 3235
rect 5715 3205 5720 3235
rect 4720 3200 5720 3205
rect 5760 3235 5960 3240
rect 5760 3205 5765 3235
rect 5795 3205 5925 3235
rect 5955 3205 5960 3235
rect 5760 3200 5960 3205
rect 6000 3235 6200 3240
rect 6000 3205 6005 3235
rect 6035 3205 6165 3235
rect 6195 3205 6200 3235
rect 6000 3200 6200 3205
rect 4240 3155 4440 3160
rect 4240 3125 4245 3155
rect 4275 3125 4405 3155
rect 4435 3125 4440 3155
rect 4240 3120 4440 3125
rect 4480 3155 4680 3160
rect 4480 3125 4485 3155
rect 4515 3125 4645 3155
rect 4675 3125 4680 3155
rect 4480 3120 4680 3125
rect 4720 3155 5720 3160
rect 4720 3125 4725 3155
rect 4755 3125 4885 3155
rect 4915 3125 5045 3155
rect 5075 3125 5205 3155
rect 5235 3125 5365 3155
rect 5395 3125 5525 3155
rect 5555 3125 5685 3155
rect 5715 3125 5720 3155
rect 4720 3120 5720 3125
rect 5760 3155 5960 3160
rect 5760 3125 5765 3155
rect 5795 3125 5925 3155
rect 5955 3125 5960 3155
rect 5760 3120 5960 3125
rect 6000 3155 6200 3160
rect 6000 3125 6005 3155
rect 6035 3125 6165 3155
rect 6195 3125 6200 3155
rect 6000 3120 6200 3125
rect 4240 3075 4440 3080
rect 4240 3045 4245 3075
rect 4275 3045 4405 3075
rect 4435 3045 4440 3075
rect 4240 3040 4440 3045
rect 4480 3075 4680 3080
rect 4480 3045 4485 3075
rect 4515 3045 4645 3075
rect 4675 3045 4680 3075
rect 4480 3040 4680 3045
rect 4720 3075 5720 3080
rect 4720 3045 4725 3075
rect 4755 3045 4885 3075
rect 4915 3045 5045 3075
rect 5075 3045 5205 3075
rect 5235 3045 5365 3075
rect 5395 3045 5525 3075
rect 5555 3045 5685 3075
rect 5715 3045 5720 3075
rect 4720 3040 5720 3045
rect 5760 3075 5960 3080
rect 5760 3045 5765 3075
rect 5795 3045 5925 3075
rect 5955 3045 5960 3075
rect 5760 3040 5960 3045
rect 6000 3075 6200 3080
rect 6000 3045 6005 3075
rect 6035 3045 6165 3075
rect 6195 3045 6200 3075
rect 6000 3040 6200 3045
rect 4240 2995 4440 3000
rect 4240 2965 4245 2995
rect 4275 2965 4405 2995
rect 4435 2965 4440 2995
rect 4240 2960 4440 2965
rect 4480 2995 4680 3000
rect 4480 2965 4485 2995
rect 4515 2965 4645 2995
rect 4675 2965 4680 2995
rect 4480 2960 4680 2965
rect 4720 2995 5720 3000
rect 4720 2965 4725 2995
rect 4755 2965 4885 2995
rect 4915 2965 5045 2995
rect 5075 2965 5205 2995
rect 5235 2965 5365 2995
rect 5395 2965 5525 2995
rect 5555 2965 5685 2995
rect 5715 2965 5720 2995
rect 4720 2960 5720 2965
rect 5760 2995 5960 3000
rect 5760 2965 5765 2995
rect 5795 2965 5925 2995
rect 5955 2965 5960 2995
rect 5760 2960 5960 2965
rect 6000 2995 6200 3000
rect 6000 2965 6005 2995
rect 6035 2965 6165 2995
rect 6195 2965 6200 2995
rect 6000 2960 6200 2965
rect 4240 2915 4440 2920
rect 4240 2885 4245 2915
rect 4275 2885 4405 2915
rect 4435 2885 4440 2915
rect 4240 2880 4440 2885
rect 4480 2915 4680 2920
rect 4480 2885 4485 2915
rect 4515 2885 4645 2915
rect 4675 2885 4680 2915
rect 4480 2880 4680 2885
rect 4720 2915 5720 2920
rect 4720 2885 4725 2915
rect 4755 2885 4885 2915
rect 4915 2885 5045 2915
rect 5075 2885 5205 2915
rect 5235 2885 5365 2915
rect 5395 2885 5525 2915
rect 5555 2885 5685 2915
rect 5715 2885 5720 2915
rect 4720 2880 5720 2885
rect 5760 2915 5960 2920
rect 5760 2885 5765 2915
rect 5795 2885 5925 2915
rect 5955 2885 5960 2915
rect 5760 2880 5960 2885
rect 6000 2915 6200 2920
rect 6000 2885 6005 2915
rect 6035 2885 6165 2915
rect 6195 2885 6200 2915
rect 6000 2880 6200 2885
rect 4240 2835 4440 2840
rect 4240 2805 4245 2835
rect 4275 2805 4405 2835
rect 4435 2805 4440 2835
rect 4240 2800 4440 2805
rect 4480 2835 4680 2840
rect 4480 2805 4485 2835
rect 4515 2805 4645 2835
rect 4675 2805 4680 2835
rect 4480 2800 4680 2805
rect 4720 2835 5720 2840
rect 4720 2805 4725 2835
rect 4755 2805 4885 2835
rect 4915 2805 5045 2835
rect 5075 2805 5205 2835
rect 5235 2805 5365 2835
rect 5395 2805 5525 2835
rect 5555 2805 5685 2835
rect 5715 2805 5720 2835
rect 4720 2800 5720 2805
rect 5760 2835 5960 2840
rect 5760 2805 5765 2835
rect 5795 2805 5925 2835
rect 5955 2805 5960 2835
rect 5760 2800 5960 2805
rect 6000 2835 6200 2840
rect 6000 2805 6005 2835
rect 6035 2805 6165 2835
rect 6195 2805 6200 2835
rect 6000 2800 6200 2805
rect 4240 2755 4440 2760
rect 4240 2725 4245 2755
rect 4275 2725 4405 2755
rect 4435 2725 4440 2755
rect 4240 2720 4440 2725
rect 4480 2755 4680 2760
rect 4480 2725 4485 2755
rect 4515 2725 4645 2755
rect 4675 2725 4680 2755
rect 4480 2720 4680 2725
rect 4720 2755 5720 2760
rect 4720 2725 4725 2755
rect 4755 2725 4885 2755
rect 4915 2725 5045 2755
rect 5075 2725 5205 2755
rect 5235 2725 5365 2755
rect 5395 2725 5525 2755
rect 5555 2725 5685 2755
rect 5715 2725 5720 2755
rect 4720 2720 5720 2725
rect 5760 2755 5960 2760
rect 5760 2725 5765 2755
rect 5795 2725 5925 2755
rect 5955 2725 5960 2755
rect 5760 2720 5960 2725
rect 6000 2755 6200 2760
rect 6000 2725 6005 2755
rect 6035 2725 6165 2755
rect 6195 2725 6200 2755
rect 6000 2720 6200 2725
rect 4240 2675 4440 2680
rect 4240 2645 4245 2675
rect 4275 2645 4405 2675
rect 4435 2645 4440 2675
rect 4240 2640 4440 2645
rect 4480 2675 4680 2680
rect 4480 2645 4485 2675
rect 4515 2645 4645 2675
rect 4675 2645 4680 2675
rect 4480 2640 4680 2645
rect 4720 2675 5720 2680
rect 4720 2645 4725 2675
rect 4755 2645 4885 2675
rect 4915 2645 5045 2675
rect 5075 2645 5205 2675
rect 5235 2645 5365 2675
rect 5395 2645 5525 2675
rect 5555 2645 5685 2675
rect 5715 2645 5720 2675
rect 4720 2640 5720 2645
rect 5760 2675 5960 2680
rect 5760 2645 5765 2675
rect 5795 2645 5925 2675
rect 5955 2645 5960 2675
rect 5760 2640 5960 2645
rect 6000 2675 6200 2680
rect 6000 2645 6005 2675
rect 6035 2645 6165 2675
rect 6195 2645 6200 2675
rect 6000 2640 6200 2645
rect 4240 2595 4440 2600
rect 4240 2565 4245 2595
rect 4275 2565 4405 2595
rect 4435 2565 4440 2595
rect 4240 2560 4440 2565
rect 4480 2595 4680 2600
rect 4480 2565 4485 2595
rect 4515 2565 4645 2595
rect 4675 2565 4680 2595
rect 4480 2560 4680 2565
rect 4720 2595 5720 2600
rect 4720 2565 4725 2595
rect 4755 2565 4885 2595
rect 4915 2565 5045 2595
rect 5075 2565 5205 2595
rect 5235 2565 5365 2595
rect 5395 2565 5525 2595
rect 5555 2565 5685 2595
rect 5715 2565 5720 2595
rect 4720 2560 5720 2565
rect 5760 2595 5960 2600
rect 5760 2565 5765 2595
rect 5795 2565 5925 2595
rect 5955 2565 5960 2595
rect 5760 2560 5960 2565
rect 6000 2595 6200 2600
rect 6000 2565 6005 2595
rect 6035 2565 6165 2595
rect 6195 2565 6200 2595
rect 6000 2560 6200 2565
rect 4240 2515 4440 2520
rect 4240 2485 4245 2515
rect 4275 2485 4405 2515
rect 4435 2485 4440 2515
rect 4240 2480 4440 2485
rect 4480 2515 4680 2520
rect 4480 2485 4485 2515
rect 4515 2485 4645 2515
rect 4675 2485 4680 2515
rect 4480 2480 4680 2485
rect 4720 2515 5720 2520
rect 4720 2485 4725 2515
rect 4755 2485 4885 2515
rect 4915 2485 5045 2515
rect 5075 2485 5205 2515
rect 5235 2485 5365 2515
rect 5395 2485 5525 2515
rect 5555 2485 5685 2515
rect 5715 2485 5720 2515
rect 4720 2480 5720 2485
rect 5760 2515 5960 2520
rect 5760 2485 5765 2515
rect 5795 2485 5925 2515
rect 5955 2485 5960 2515
rect 5760 2480 5960 2485
rect 6000 2515 6200 2520
rect 6000 2485 6005 2515
rect 6035 2485 6165 2515
rect 6195 2485 6200 2515
rect 6000 2480 6200 2485
rect 4240 2435 4440 2440
rect 4240 2405 4245 2435
rect 4275 2405 4405 2435
rect 4435 2405 4440 2435
rect 4240 2400 4440 2405
rect 4480 2435 4680 2440
rect 4480 2405 4485 2435
rect 4515 2405 4645 2435
rect 4675 2405 4680 2435
rect 4480 2400 4680 2405
rect 4720 2435 5720 2440
rect 4720 2405 4725 2435
rect 4755 2405 4885 2435
rect 4915 2405 5045 2435
rect 5075 2405 5205 2435
rect 5235 2405 5365 2435
rect 5395 2405 5525 2435
rect 5555 2405 5685 2435
rect 5715 2405 5720 2435
rect 4720 2400 5720 2405
rect 5760 2435 5960 2440
rect 5760 2405 5765 2435
rect 5795 2405 5925 2435
rect 5955 2405 5960 2435
rect 5760 2400 5960 2405
rect 6000 2435 6200 2440
rect 6000 2405 6005 2435
rect 6035 2405 6165 2435
rect 6195 2405 6200 2435
rect 6000 2400 6200 2405
rect 4240 2355 4440 2360
rect 4240 2325 4245 2355
rect 4275 2325 4405 2355
rect 4435 2325 4440 2355
rect 4240 2320 4440 2325
rect 4480 2355 4680 2360
rect 4480 2325 4485 2355
rect 4515 2325 4645 2355
rect 4675 2325 4680 2355
rect 4480 2320 4680 2325
rect 4720 2355 5720 2360
rect 4720 2325 4725 2355
rect 4755 2325 4885 2355
rect 4915 2325 5045 2355
rect 5075 2325 5205 2355
rect 5235 2325 5365 2355
rect 5395 2325 5525 2355
rect 5555 2325 5685 2355
rect 5715 2325 5720 2355
rect 4720 2320 5720 2325
rect 5760 2355 5960 2360
rect 5760 2325 5765 2355
rect 5795 2325 5925 2355
rect 5955 2325 5960 2355
rect 5760 2320 5960 2325
rect 6000 2355 6200 2360
rect 6000 2325 6005 2355
rect 6035 2325 6165 2355
rect 6195 2325 6200 2355
rect 6000 2320 6200 2325
rect 4240 2275 4440 2280
rect 4240 2245 4245 2275
rect 4275 2245 4405 2275
rect 4435 2245 4440 2275
rect 4240 2240 4440 2245
rect 4480 2275 4680 2280
rect 4480 2245 4485 2275
rect 4515 2245 4645 2275
rect 4675 2245 4680 2275
rect 4480 2240 4680 2245
rect 4720 2275 5720 2280
rect 4720 2245 4725 2275
rect 4755 2245 4885 2275
rect 4915 2245 5045 2275
rect 5075 2245 5205 2275
rect 5235 2245 5365 2275
rect 5395 2245 5525 2275
rect 5555 2245 5685 2275
rect 5715 2245 5720 2275
rect 4720 2240 5720 2245
rect 5760 2275 5960 2280
rect 5760 2245 5765 2275
rect 5795 2245 5925 2275
rect 5955 2245 5960 2275
rect 5760 2240 5960 2245
rect 6000 2275 6200 2280
rect 6000 2245 6005 2275
rect 6035 2245 6165 2275
rect 6195 2245 6200 2275
rect 6000 2240 6200 2245
rect 4240 2195 4440 2200
rect 4240 2165 4245 2195
rect 4275 2165 4405 2195
rect 4435 2165 4440 2195
rect 4240 2160 4440 2165
rect 4480 2195 4680 2200
rect 4480 2165 4485 2195
rect 4515 2165 4645 2195
rect 4675 2165 4680 2195
rect 4480 2160 4680 2165
rect 4720 2195 5720 2200
rect 4720 2165 4725 2195
rect 4755 2165 4885 2195
rect 4915 2165 5045 2195
rect 5075 2165 5205 2195
rect 5235 2165 5365 2195
rect 5395 2165 5525 2195
rect 5555 2165 5685 2195
rect 5715 2165 5720 2195
rect 4720 2160 5720 2165
rect 5760 2195 5960 2200
rect 5760 2165 5765 2195
rect 5795 2165 5925 2195
rect 5955 2165 5960 2195
rect 5760 2160 5960 2165
rect 6000 2195 6200 2200
rect 6000 2165 6005 2195
rect 6035 2165 6165 2195
rect 6195 2165 6200 2195
rect 6000 2160 6200 2165
rect 4240 2115 4440 2120
rect 4240 2085 4245 2115
rect 4275 2085 4405 2115
rect 4435 2085 4440 2115
rect 4240 2080 4440 2085
rect 4480 2115 4680 2120
rect 4480 2085 4485 2115
rect 4515 2085 4645 2115
rect 4675 2085 4680 2115
rect 4480 2080 4680 2085
rect 4720 2115 5720 2120
rect 4720 2085 4725 2115
rect 4755 2085 4885 2115
rect 4915 2085 5045 2115
rect 5075 2085 5205 2115
rect 5235 2085 5365 2115
rect 5395 2085 5525 2115
rect 5555 2085 5685 2115
rect 5715 2085 5720 2115
rect 4720 2080 5720 2085
rect 5760 2115 5960 2120
rect 5760 2085 5765 2115
rect 5795 2085 5925 2115
rect 5955 2085 5960 2115
rect 5760 2080 5960 2085
rect 6000 2115 6200 2120
rect 6000 2085 6005 2115
rect 6035 2085 6165 2115
rect 6195 2085 6200 2115
rect 6000 2080 6200 2085
rect 4240 2035 4440 2040
rect 4240 2005 4245 2035
rect 4275 2005 4405 2035
rect 4435 2005 4440 2035
rect 4240 2000 4440 2005
rect 4480 2035 4680 2040
rect 4480 2005 4485 2035
rect 4515 2005 4645 2035
rect 4675 2005 4680 2035
rect 4480 2000 4680 2005
rect 4720 2035 5720 2040
rect 4720 2005 4725 2035
rect 4755 2005 4885 2035
rect 4915 2005 5045 2035
rect 5075 2005 5205 2035
rect 5235 2005 5365 2035
rect 5395 2005 5525 2035
rect 5555 2005 5685 2035
rect 5715 2005 5720 2035
rect 4720 2000 5720 2005
rect 5760 2035 5960 2040
rect 5760 2005 5765 2035
rect 5795 2005 5925 2035
rect 5955 2005 5960 2035
rect 5760 2000 5960 2005
rect 6000 2035 6200 2040
rect 6000 2005 6005 2035
rect 6035 2005 6165 2035
rect 6195 2005 6200 2035
rect 6000 2000 6200 2005
rect 4240 1955 4440 1960
rect 4240 1925 4245 1955
rect 4275 1925 4405 1955
rect 4435 1925 4440 1955
rect 4240 1920 4440 1925
rect 4480 1955 4680 1960
rect 4480 1925 4485 1955
rect 4515 1925 4645 1955
rect 4675 1925 4680 1955
rect 4480 1920 4680 1925
rect 4720 1955 5720 1960
rect 4720 1925 4725 1955
rect 4755 1925 4885 1955
rect 4915 1925 5045 1955
rect 5075 1925 5205 1955
rect 5235 1925 5365 1955
rect 5395 1925 5525 1955
rect 5555 1925 5685 1955
rect 5715 1925 5720 1955
rect 4720 1920 5720 1925
rect 5760 1955 5960 1960
rect 5760 1925 5765 1955
rect 5795 1925 5925 1955
rect 5955 1925 5960 1955
rect 5760 1920 5960 1925
rect 6000 1955 6200 1960
rect 6000 1925 6005 1955
rect 6035 1925 6165 1955
rect 6195 1925 6200 1955
rect 6000 1920 6200 1925
rect 0 1835 10440 1840
rect 0 1805 4565 1835
rect 4595 1805 10440 1835
rect 0 1800 10440 1805
rect 4240 1715 4440 1720
rect 4240 1685 4245 1715
rect 4275 1685 4405 1715
rect 4435 1685 4440 1715
rect 4240 1680 4440 1685
rect 4480 1715 4680 1720
rect 4480 1685 4485 1715
rect 4515 1685 4645 1715
rect 4675 1685 4680 1715
rect 4480 1680 4680 1685
rect 4720 1715 5720 1720
rect 4720 1685 4725 1715
rect 4755 1685 4885 1715
rect 4915 1685 5045 1715
rect 5075 1685 5205 1715
rect 5235 1685 5365 1715
rect 5395 1685 5525 1715
rect 5555 1685 5685 1715
rect 5715 1685 5720 1715
rect 4720 1680 5720 1685
rect 5760 1715 5960 1720
rect 5760 1685 5765 1715
rect 5795 1685 5925 1715
rect 5955 1685 5960 1715
rect 5760 1680 5960 1685
rect 6000 1715 6200 1720
rect 6000 1685 6005 1715
rect 6035 1685 6165 1715
rect 6195 1685 6200 1715
rect 6000 1680 6200 1685
rect 4240 1635 4440 1640
rect 4240 1605 4245 1635
rect 4275 1605 4405 1635
rect 4435 1605 4440 1635
rect 4240 1600 4440 1605
rect 4480 1635 4680 1640
rect 4480 1605 4485 1635
rect 4515 1605 4645 1635
rect 4675 1605 4680 1635
rect 4480 1600 4680 1605
rect 4720 1635 5720 1640
rect 4720 1605 4725 1635
rect 4755 1605 4885 1635
rect 4915 1605 5045 1635
rect 5075 1605 5205 1635
rect 5235 1605 5365 1635
rect 5395 1605 5525 1635
rect 5555 1605 5685 1635
rect 5715 1605 5720 1635
rect 4720 1600 5720 1605
rect 5760 1635 5960 1640
rect 5760 1605 5765 1635
rect 5795 1605 5925 1635
rect 5955 1605 5960 1635
rect 5760 1600 5960 1605
rect 6000 1635 6200 1640
rect 6000 1605 6005 1635
rect 6035 1605 6165 1635
rect 6195 1605 6200 1635
rect 6000 1600 6200 1605
rect 4240 1555 4440 1560
rect 4240 1525 4245 1555
rect 4275 1525 4405 1555
rect 4435 1525 4440 1555
rect 4240 1520 4440 1525
rect 4480 1555 4680 1560
rect 4480 1525 4485 1555
rect 4515 1525 4645 1555
rect 4675 1525 4680 1555
rect 4480 1520 4680 1525
rect 4720 1555 5720 1560
rect 4720 1525 4725 1555
rect 4755 1525 4885 1555
rect 4915 1525 5045 1555
rect 5075 1525 5205 1555
rect 5235 1525 5365 1555
rect 5395 1525 5525 1555
rect 5555 1525 5685 1555
rect 5715 1525 5720 1555
rect 4720 1520 5720 1525
rect 5760 1555 5960 1560
rect 5760 1525 5765 1555
rect 5795 1525 5925 1555
rect 5955 1525 5960 1555
rect 5760 1520 5960 1525
rect 6000 1555 6200 1560
rect 6000 1525 6005 1555
rect 6035 1525 6165 1555
rect 6195 1525 6200 1555
rect 6000 1520 6200 1525
rect 4240 1475 4440 1480
rect 4240 1445 4245 1475
rect 4275 1445 4405 1475
rect 4435 1445 4440 1475
rect 4240 1440 4440 1445
rect 4480 1475 4680 1480
rect 4480 1445 4485 1475
rect 4515 1445 4645 1475
rect 4675 1445 4680 1475
rect 4480 1440 4680 1445
rect 4720 1475 5720 1480
rect 4720 1445 4725 1475
rect 4755 1445 4885 1475
rect 4915 1445 5045 1475
rect 5075 1445 5205 1475
rect 5235 1445 5365 1475
rect 5395 1445 5525 1475
rect 5555 1445 5685 1475
rect 5715 1445 5720 1475
rect 4720 1440 5720 1445
rect 5760 1475 5960 1480
rect 5760 1445 5765 1475
rect 5795 1445 5925 1475
rect 5955 1445 5960 1475
rect 5760 1440 5960 1445
rect 6000 1475 6200 1480
rect 6000 1445 6005 1475
rect 6035 1445 6165 1475
rect 6195 1445 6200 1475
rect 6000 1440 6200 1445
rect 4240 1395 4440 1400
rect 4240 1365 4245 1395
rect 4275 1365 4405 1395
rect 4435 1365 4440 1395
rect 4240 1360 4440 1365
rect 4480 1395 4680 1400
rect 4480 1365 4485 1395
rect 4515 1365 4645 1395
rect 4675 1365 4680 1395
rect 4480 1360 4680 1365
rect 4720 1395 5720 1400
rect 4720 1365 4725 1395
rect 4755 1365 4885 1395
rect 4915 1365 5045 1395
rect 5075 1365 5205 1395
rect 5235 1365 5365 1395
rect 5395 1365 5525 1395
rect 5555 1365 5685 1395
rect 5715 1365 5720 1395
rect 4720 1360 5720 1365
rect 5760 1395 5960 1400
rect 5760 1365 5765 1395
rect 5795 1365 5925 1395
rect 5955 1365 5960 1395
rect 5760 1360 5960 1365
rect 6000 1395 6200 1400
rect 6000 1365 6005 1395
rect 6035 1365 6165 1395
rect 6195 1365 6200 1395
rect 6000 1360 6200 1365
rect 4240 1315 4440 1320
rect 4240 1285 4245 1315
rect 4275 1285 4405 1315
rect 4435 1285 4440 1315
rect 4240 1280 4440 1285
rect 4480 1315 4680 1320
rect 4480 1285 4485 1315
rect 4515 1285 4645 1315
rect 4675 1285 4680 1315
rect 4480 1280 4680 1285
rect 4720 1315 5720 1320
rect 4720 1285 4725 1315
rect 4755 1285 4885 1315
rect 4915 1285 5045 1315
rect 5075 1285 5205 1315
rect 5235 1285 5365 1315
rect 5395 1285 5525 1315
rect 5555 1285 5685 1315
rect 5715 1285 5720 1315
rect 4720 1280 5720 1285
rect 5760 1315 5960 1320
rect 5760 1285 5765 1315
rect 5795 1285 5925 1315
rect 5955 1285 5960 1315
rect 5760 1280 5960 1285
rect 6000 1315 6200 1320
rect 6000 1285 6005 1315
rect 6035 1285 6165 1315
rect 6195 1285 6200 1315
rect 6000 1280 6200 1285
rect 4240 1235 4440 1240
rect 4240 1205 4245 1235
rect 4275 1205 4405 1235
rect 4435 1205 4440 1235
rect 4240 1200 4440 1205
rect 4480 1235 4680 1240
rect 4480 1205 4485 1235
rect 4515 1205 4645 1235
rect 4675 1205 4680 1235
rect 4480 1200 4680 1205
rect 4720 1235 5720 1240
rect 4720 1205 4725 1235
rect 4755 1205 4885 1235
rect 4915 1205 5045 1235
rect 5075 1205 5205 1235
rect 5235 1205 5365 1235
rect 5395 1205 5525 1235
rect 5555 1205 5685 1235
rect 5715 1205 5720 1235
rect 4720 1200 5720 1205
rect 5760 1235 5960 1240
rect 5760 1205 5765 1235
rect 5795 1205 5925 1235
rect 5955 1205 5960 1235
rect 5760 1200 5960 1205
rect 6000 1235 6200 1240
rect 6000 1205 6005 1235
rect 6035 1205 6165 1235
rect 6195 1205 6200 1235
rect 6000 1200 6200 1205
rect 4240 1155 4440 1160
rect 4240 1125 4245 1155
rect 4275 1125 4405 1155
rect 4435 1125 4440 1155
rect 4240 1120 4440 1125
rect 4480 1155 4680 1160
rect 4480 1125 4485 1155
rect 4515 1125 4645 1155
rect 4675 1125 4680 1155
rect 4480 1120 4680 1125
rect 4720 1155 5720 1160
rect 4720 1125 4725 1155
rect 4755 1125 4885 1155
rect 4915 1125 5045 1155
rect 5075 1125 5205 1155
rect 5235 1125 5365 1155
rect 5395 1125 5525 1155
rect 5555 1125 5685 1155
rect 5715 1125 5720 1155
rect 4720 1120 5720 1125
rect 5760 1155 5960 1160
rect 5760 1125 5765 1155
rect 5795 1125 5925 1155
rect 5955 1125 5960 1155
rect 5760 1120 5960 1125
rect 6000 1155 6200 1160
rect 6000 1125 6005 1155
rect 6035 1125 6165 1155
rect 6195 1125 6200 1155
rect 6000 1120 6200 1125
rect 4240 1075 4440 1080
rect 4240 1045 4245 1075
rect 4275 1045 4405 1075
rect 4435 1045 4440 1075
rect 4240 1040 4440 1045
rect 4480 1075 4680 1080
rect 4480 1045 4485 1075
rect 4515 1045 4645 1075
rect 4675 1045 4680 1075
rect 4480 1040 4680 1045
rect 4720 1075 5720 1080
rect 4720 1045 4725 1075
rect 4755 1045 4885 1075
rect 4915 1045 5045 1075
rect 5075 1045 5205 1075
rect 5235 1045 5365 1075
rect 5395 1045 5525 1075
rect 5555 1045 5685 1075
rect 5715 1045 5720 1075
rect 4720 1040 5720 1045
rect 5760 1075 5960 1080
rect 5760 1045 5765 1075
rect 5795 1045 5925 1075
rect 5955 1045 5960 1075
rect 5760 1040 5960 1045
rect 6000 1075 6200 1080
rect 6000 1045 6005 1075
rect 6035 1045 6165 1075
rect 6195 1045 6200 1075
rect 6000 1040 6200 1045
rect 4240 995 4440 1000
rect 4240 965 4245 995
rect 4275 965 4405 995
rect 4435 965 4440 995
rect 4240 960 4440 965
rect 4480 995 4680 1000
rect 4480 965 4485 995
rect 4515 965 4645 995
rect 4675 965 4680 995
rect 4480 960 4680 965
rect 4720 995 5720 1000
rect 4720 965 4725 995
rect 4755 965 4885 995
rect 4915 965 5045 995
rect 5075 965 5205 995
rect 5235 965 5365 995
rect 5395 965 5525 995
rect 5555 965 5685 995
rect 5715 965 5720 995
rect 4720 960 5720 965
rect 5760 995 5960 1000
rect 5760 965 5765 995
rect 5795 965 5925 995
rect 5955 965 5960 995
rect 5760 960 5960 965
rect 6000 995 6200 1000
rect 6000 965 6005 995
rect 6035 965 6165 995
rect 6195 965 6200 995
rect 6000 960 6200 965
rect 0 915 10440 920
rect 0 885 6085 915
rect 6115 885 10440 915
rect 0 880 10440 885
rect 4240 835 4440 840
rect 4240 805 4245 835
rect 4275 805 4405 835
rect 4435 805 4440 835
rect 4240 800 4440 805
rect 4480 835 4680 840
rect 4480 805 4485 835
rect 4515 805 4645 835
rect 4675 805 4680 835
rect 4480 800 4680 805
rect 4720 835 5720 840
rect 4720 805 4725 835
rect 4755 805 4885 835
rect 4915 805 5045 835
rect 5075 805 5205 835
rect 5235 805 5365 835
rect 5395 805 5525 835
rect 5555 805 5685 835
rect 5715 805 5720 835
rect 4720 800 5720 805
rect 5760 835 5960 840
rect 5760 805 5765 835
rect 5795 805 5925 835
rect 5955 805 5960 835
rect 5760 800 5960 805
rect 6000 835 6200 840
rect 6000 805 6005 835
rect 6035 805 6165 835
rect 6195 805 6200 835
rect 6000 800 6200 805
rect 4240 755 4440 760
rect 4240 725 4245 755
rect 4275 725 4405 755
rect 4435 725 4440 755
rect 4240 720 4440 725
rect 4480 755 4680 760
rect 4480 725 4485 755
rect 4515 725 4645 755
rect 4675 725 4680 755
rect 4480 720 4680 725
rect 4720 755 5720 760
rect 4720 725 4725 755
rect 4755 725 4885 755
rect 4915 725 5045 755
rect 5075 725 5205 755
rect 5235 725 5365 755
rect 5395 725 5525 755
rect 5555 725 5685 755
rect 5715 725 5720 755
rect 4720 720 5720 725
rect 5760 755 5960 760
rect 5760 725 5765 755
rect 5795 725 5925 755
rect 5955 725 5960 755
rect 5760 720 5960 725
rect 6000 755 6200 760
rect 6000 725 6005 755
rect 6035 725 6165 755
rect 6195 725 6200 755
rect 6000 720 6200 725
rect 4240 675 4440 680
rect 4240 645 4245 675
rect 4275 645 4405 675
rect 4435 645 4440 675
rect 4240 640 4440 645
rect 4480 675 4680 680
rect 4480 645 4485 675
rect 4515 645 4645 675
rect 4675 645 4680 675
rect 4480 640 4680 645
rect 4720 675 5720 680
rect 4720 645 4725 675
rect 4755 645 4885 675
rect 4915 645 5045 675
rect 5075 645 5205 675
rect 5235 645 5365 675
rect 5395 645 5525 675
rect 5555 645 5685 675
rect 5715 645 5720 675
rect 4720 640 5720 645
rect 5760 675 5960 680
rect 5760 645 5765 675
rect 5795 645 5925 675
rect 5955 645 5960 675
rect 5760 640 5960 645
rect 6000 675 6200 680
rect 6000 645 6005 675
rect 6035 645 6165 675
rect 6195 645 6200 675
rect 6000 640 6200 645
rect 4240 595 4440 600
rect 4240 565 4245 595
rect 4275 565 4405 595
rect 4435 565 4440 595
rect 4240 560 4440 565
rect 4480 595 4680 600
rect 4480 565 4485 595
rect 4515 565 4645 595
rect 4675 565 4680 595
rect 4480 560 4680 565
rect 4720 595 5720 600
rect 4720 565 4725 595
rect 4755 565 4885 595
rect 4915 565 5045 595
rect 5075 565 5205 595
rect 5235 565 5365 595
rect 5395 565 5525 595
rect 5555 565 5685 595
rect 5715 565 5720 595
rect 4720 560 5720 565
rect 5760 595 5960 600
rect 5760 565 5765 595
rect 5795 565 5925 595
rect 5955 565 5960 595
rect 5760 560 5960 565
rect 6000 595 6200 600
rect 6000 565 6005 595
rect 6035 565 6165 595
rect 6195 565 6200 595
rect 6000 560 6200 565
rect 4240 515 4440 520
rect 4240 485 4245 515
rect 4275 485 4405 515
rect 4435 485 4440 515
rect 4240 480 4440 485
rect 4480 515 4680 520
rect 4480 485 4485 515
rect 4515 485 4645 515
rect 4675 485 4680 515
rect 4480 480 4680 485
rect 4720 515 5720 520
rect 4720 485 4725 515
rect 4755 485 4885 515
rect 4915 485 5045 515
rect 5075 485 5205 515
rect 5235 485 5365 515
rect 5395 485 5525 515
rect 5555 485 5685 515
rect 5715 485 5720 515
rect 4720 480 5720 485
rect 5760 515 5960 520
rect 5760 485 5765 515
rect 5795 485 5925 515
rect 5955 485 5960 515
rect 5760 480 5960 485
rect 6000 515 6200 520
rect 6000 485 6005 515
rect 6035 485 6165 515
rect 6195 485 6200 515
rect 6000 480 6200 485
rect 0 395 10440 400
rect 0 365 4325 395
rect 4355 365 10440 395
rect 0 360 10440 365
rect 4240 275 4440 280
rect 4240 245 4245 275
rect 4275 245 4405 275
rect 4435 245 4440 275
rect 4240 240 4440 245
rect 4480 275 4680 280
rect 4480 245 4485 275
rect 4515 245 4645 275
rect 4675 245 4680 275
rect 4480 240 4680 245
rect 4720 275 5720 280
rect 4720 245 4725 275
rect 4755 245 4885 275
rect 4915 245 5045 275
rect 5075 245 5205 275
rect 5235 245 5365 275
rect 5395 245 5525 275
rect 5555 245 5685 275
rect 5715 245 5720 275
rect 4720 240 5720 245
rect 5760 275 5960 280
rect 5760 245 5765 275
rect 5795 245 5925 275
rect 5955 245 5960 275
rect 5760 240 5960 245
rect 6000 275 6200 280
rect 6000 245 6005 275
rect 6035 245 6165 275
rect 6195 245 6200 275
rect 6000 240 6200 245
rect 4240 195 4440 200
rect 4240 165 4245 195
rect 4275 165 4405 195
rect 4435 165 4440 195
rect 4240 160 4440 165
rect 4480 195 4680 200
rect 4480 165 4485 195
rect 4515 165 4645 195
rect 4675 165 4680 195
rect 4480 160 4680 165
rect 4720 195 5720 200
rect 4720 165 4725 195
rect 4755 165 4885 195
rect 4915 165 5045 195
rect 5075 165 5205 195
rect 5235 165 5365 195
rect 5395 165 5525 195
rect 5555 165 5685 195
rect 5715 165 5720 195
rect 4720 160 5720 165
rect 5760 195 5960 200
rect 5760 165 5765 195
rect 5795 165 5925 195
rect 5955 165 5960 195
rect 5760 160 5960 165
rect 6000 195 6200 200
rect 6000 165 6005 195
rect 6035 165 6165 195
rect 6195 165 6200 195
rect 6000 160 6200 165
rect 4240 115 4440 120
rect 4240 85 4245 115
rect 4275 85 4405 115
rect 4435 85 4440 115
rect 4240 80 4440 85
rect 4480 115 4680 120
rect 4480 85 4485 115
rect 4515 85 4645 115
rect 4675 85 4680 115
rect 4480 80 4680 85
rect 4720 115 5720 120
rect 4720 85 4725 115
rect 4755 85 4885 115
rect 4915 85 5045 115
rect 5075 85 5205 115
rect 5235 85 5365 115
rect 5395 85 5525 115
rect 5555 85 5685 115
rect 5715 85 5720 115
rect 4720 80 5720 85
rect 5760 115 5960 120
rect 5760 85 5765 115
rect 5795 85 5925 115
rect 5955 85 5960 115
rect 5760 80 5960 85
rect 6000 115 6200 120
rect 6000 85 6005 115
rect 6035 85 6165 115
rect 6195 85 6200 115
rect 6000 80 6200 85
rect 4240 35 4440 40
rect 4240 5 4245 35
rect 4275 5 4405 35
rect 4435 5 4440 35
rect 4240 0 4440 5
rect 4480 35 4680 40
rect 4480 5 4485 35
rect 4515 5 4645 35
rect 4675 5 4680 35
rect 4480 0 4680 5
rect 4720 35 5720 40
rect 4720 5 4725 35
rect 4755 5 4885 35
rect 4915 5 5045 35
rect 5075 5 5205 35
rect 5235 5 5365 35
rect 5395 5 5525 35
rect 5555 5 5685 35
rect 5715 5 5720 35
rect 4720 0 5720 5
rect 5760 35 5960 40
rect 5760 5 5765 35
rect 5795 5 5925 35
rect 5955 5 5960 35
rect 5760 0 5960 5
rect 6000 35 6200 40
rect 6000 5 6005 35
rect 6035 5 6165 35
rect 6195 5 6200 35
rect 6000 0 6200 5
<< via2 >>
rect 4245 15685 4275 15715
rect 4405 15685 4435 15715
rect 4485 15685 4515 15715
rect 4645 15685 4675 15715
rect 4725 15685 4755 15715
rect 4885 15685 4915 15715
rect 5045 15685 5075 15715
rect 5205 15685 5235 15715
rect 5365 15685 5395 15715
rect 5525 15685 5555 15715
rect 5685 15685 5715 15715
rect 5765 15685 5795 15715
rect 5925 15685 5955 15715
rect 6005 15685 6035 15715
rect 6165 15685 6195 15715
rect 4245 15605 4275 15635
rect 4405 15605 4435 15635
rect 4485 15605 4515 15635
rect 4645 15605 4675 15635
rect 4725 15605 4755 15635
rect 4885 15605 4915 15635
rect 5045 15605 5075 15635
rect 5205 15605 5235 15635
rect 5365 15605 5395 15635
rect 5525 15605 5555 15635
rect 5685 15605 5715 15635
rect 5765 15605 5795 15635
rect 5925 15605 5955 15635
rect 6005 15605 6035 15635
rect 6165 15605 6195 15635
rect 4245 15525 4275 15555
rect 4405 15525 4435 15555
rect 4485 15525 4515 15555
rect 4645 15525 4675 15555
rect 4725 15525 4755 15555
rect 4885 15525 4915 15555
rect 5045 15525 5075 15555
rect 5205 15525 5235 15555
rect 5365 15525 5395 15555
rect 5525 15525 5555 15555
rect 5685 15525 5715 15555
rect 5765 15525 5795 15555
rect 5925 15525 5955 15555
rect 6005 15525 6035 15555
rect 6165 15525 6195 15555
rect 4245 15445 4275 15475
rect 4405 15445 4435 15475
rect 4485 15445 4515 15475
rect 4645 15445 4675 15475
rect 4725 15445 4755 15475
rect 4885 15445 4915 15475
rect 5045 15445 5075 15475
rect 5205 15445 5235 15475
rect 5365 15445 5395 15475
rect 5525 15445 5555 15475
rect 5685 15445 5715 15475
rect 5765 15445 5795 15475
rect 5925 15445 5955 15475
rect 6005 15445 6035 15475
rect 6165 15445 6195 15475
rect 4245 15365 4275 15395
rect 4405 15365 4435 15395
rect 4485 15365 4515 15395
rect 4645 15365 4675 15395
rect 4725 15365 4755 15395
rect 4885 15365 4915 15395
rect 5045 15365 5075 15395
rect 5205 15365 5235 15395
rect 5365 15365 5395 15395
rect 5525 15365 5555 15395
rect 5685 15365 5715 15395
rect 5765 15365 5795 15395
rect 5925 15365 5955 15395
rect 6005 15365 6035 15395
rect 6165 15365 6195 15395
rect 4245 15285 4275 15315
rect 4405 15285 4435 15315
rect 4485 15285 4515 15315
rect 4645 15285 4675 15315
rect 4725 15285 4755 15315
rect 4885 15285 4915 15315
rect 5045 15285 5075 15315
rect 5205 15285 5235 15315
rect 5365 15285 5395 15315
rect 5525 15285 5555 15315
rect 5685 15285 5715 15315
rect 5765 15285 5795 15315
rect 5925 15285 5955 15315
rect 6005 15285 6035 15315
rect 6165 15285 6195 15315
rect 4245 15205 4275 15235
rect 4405 15205 4435 15235
rect 4485 15205 4515 15235
rect 4645 15205 4675 15235
rect 4725 15205 4755 15235
rect 4885 15205 4915 15235
rect 5045 15205 5075 15235
rect 5205 15205 5235 15235
rect 5365 15205 5395 15235
rect 5525 15205 5555 15235
rect 5685 15205 5715 15235
rect 5765 15205 5795 15235
rect 5925 15205 5955 15235
rect 6005 15205 6035 15235
rect 6165 15205 6195 15235
rect 4245 15125 4275 15155
rect 4405 15125 4435 15155
rect 4485 15125 4515 15155
rect 4645 15125 4675 15155
rect 4725 15125 4755 15155
rect 4885 15125 4915 15155
rect 5045 15125 5075 15155
rect 5205 15125 5235 15155
rect 5365 15125 5395 15155
rect 5525 15125 5555 15155
rect 5685 15125 5715 15155
rect 5765 15125 5795 15155
rect 5925 15125 5955 15155
rect 6005 15125 6035 15155
rect 6165 15125 6195 15155
rect 4565 15045 4595 15075
rect 4245 14965 4275 14995
rect 4405 14965 4435 14995
rect 4485 14965 4515 14995
rect 4645 14965 4675 14995
rect 4725 14965 4755 14995
rect 4885 14965 4915 14995
rect 5045 14965 5075 14995
rect 5205 14965 5235 14995
rect 5365 14965 5395 14995
rect 5525 14965 5555 14995
rect 5685 14965 5715 14995
rect 5765 14965 5795 14995
rect 5925 14965 5955 14995
rect 6005 14965 6035 14995
rect 6165 14965 6195 14995
rect 4245 14885 4275 14915
rect 4405 14885 4435 14915
rect 4485 14885 4515 14915
rect 4645 14885 4675 14915
rect 4725 14885 4755 14915
rect 4885 14885 4915 14915
rect 5045 14885 5075 14915
rect 5205 14885 5235 14915
rect 5365 14885 5395 14915
rect 5525 14885 5555 14915
rect 5685 14885 5715 14915
rect 5765 14885 5795 14915
rect 5925 14885 5955 14915
rect 6005 14885 6035 14915
rect 6165 14885 6195 14915
rect 4245 14805 4275 14835
rect 4405 14805 4435 14835
rect 4485 14805 4515 14835
rect 4645 14805 4675 14835
rect 4725 14805 4755 14835
rect 4885 14805 4915 14835
rect 5045 14805 5075 14835
rect 5205 14805 5235 14835
rect 5365 14805 5395 14835
rect 5525 14805 5555 14835
rect 5685 14805 5715 14835
rect 5765 14805 5795 14835
rect 5925 14805 5955 14835
rect 6005 14805 6035 14835
rect 6165 14805 6195 14835
rect 4245 14725 4275 14755
rect 4405 14725 4435 14755
rect 4485 14725 4515 14755
rect 4645 14725 4675 14755
rect 4725 14725 4755 14755
rect 4885 14725 4915 14755
rect 5045 14725 5075 14755
rect 5205 14725 5235 14755
rect 5365 14725 5395 14755
rect 5525 14725 5555 14755
rect 5685 14725 5715 14755
rect 5765 14725 5795 14755
rect 5925 14725 5955 14755
rect 6005 14725 6035 14755
rect 6165 14725 6195 14755
rect 4245 14645 4275 14675
rect 4405 14645 4435 14675
rect 4485 14645 4515 14675
rect 4645 14645 4675 14675
rect 4725 14645 4755 14675
rect 4885 14645 4915 14675
rect 5045 14645 5075 14675
rect 5205 14645 5235 14675
rect 5365 14645 5395 14675
rect 5525 14645 5555 14675
rect 5685 14645 5715 14675
rect 5765 14645 5795 14675
rect 5925 14645 5955 14675
rect 6005 14645 6035 14675
rect 6165 14645 6195 14675
rect 4245 14565 4275 14595
rect 4405 14565 4435 14595
rect 4485 14565 4515 14595
rect 4645 14565 4675 14595
rect 4725 14565 4755 14595
rect 4885 14565 4915 14595
rect 5045 14565 5075 14595
rect 5205 14565 5235 14595
rect 5365 14565 5395 14595
rect 5525 14565 5555 14595
rect 5685 14565 5715 14595
rect 5765 14565 5795 14595
rect 5925 14565 5955 14595
rect 6005 14565 6035 14595
rect 6165 14565 6195 14595
rect 4245 14485 4275 14515
rect 4405 14485 4435 14515
rect 4485 14485 4515 14515
rect 4645 14485 4675 14515
rect 4725 14485 4755 14515
rect 4885 14485 4915 14515
rect 5045 14485 5075 14515
rect 5205 14485 5235 14515
rect 5365 14485 5395 14515
rect 5525 14485 5555 14515
rect 5685 14485 5715 14515
rect 5765 14485 5795 14515
rect 5925 14485 5955 14515
rect 6005 14485 6035 14515
rect 6165 14485 6195 14515
rect 4245 14405 4275 14435
rect 4405 14405 4435 14435
rect 4485 14405 4515 14435
rect 4645 14405 4675 14435
rect 4725 14405 4755 14435
rect 4885 14405 4915 14435
rect 5045 14405 5075 14435
rect 5205 14405 5235 14435
rect 5365 14405 5395 14435
rect 5525 14405 5555 14435
rect 5685 14405 5715 14435
rect 5765 14405 5795 14435
rect 5925 14405 5955 14435
rect 6005 14405 6035 14435
rect 6165 14405 6195 14435
rect 5285 14285 5315 14315
rect 4965 14125 4995 14155
rect 5445 14125 5475 14155
rect 4245 14005 4275 14035
rect 4405 14005 4435 14035
rect 4485 14005 4515 14035
rect 4645 14005 4675 14035
rect 4725 14005 4755 14035
rect 4885 14005 4915 14035
rect 5045 14005 5075 14035
rect 5205 14005 5235 14035
rect 5365 14005 5395 14035
rect 5525 14005 5555 14035
rect 5685 14005 5715 14035
rect 5765 14005 5795 14035
rect 5925 14005 5955 14035
rect 6005 14005 6035 14035
rect 6165 14005 6195 14035
rect 4245 13925 4275 13955
rect 4405 13925 4435 13955
rect 4485 13925 4515 13955
rect 4645 13925 4675 13955
rect 4725 13925 4755 13955
rect 4885 13925 4915 13955
rect 5045 13925 5075 13955
rect 5205 13925 5235 13955
rect 5365 13925 5395 13955
rect 5525 13925 5555 13955
rect 5685 13925 5715 13955
rect 5765 13925 5795 13955
rect 5925 13925 5955 13955
rect 6005 13925 6035 13955
rect 6165 13925 6195 13955
rect 4245 13845 4275 13875
rect 4405 13845 4435 13875
rect 4485 13845 4515 13875
rect 4645 13845 4675 13875
rect 4725 13845 4755 13875
rect 4885 13845 4915 13875
rect 5045 13845 5075 13875
rect 5205 13845 5235 13875
rect 5365 13845 5395 13875
rect 5525 13845 5555 13875
rect 5685 13845 5715 13875
rect 5765 13845 5795 13875
rect 5925 13845 5955 13875
rect 6005 13845 6035 13875
rect 6165 13845 6195 13875
rect 4245 13765 4275 13795
rect 4405 13765 4435 13795
rect 4485 13765 4515 13795
rect 4645 13765 4675 13795
rect 4725 13765 4755 13795
rect 4885 13765 4915 13795
rect 5045 13765 5075 13795
rect 5205 13765 5235 13795
rect 5365 13765 5395 13795
rect 5525 13765 5555 13795
rect 5685 13765 5715 13795
rect 5765 13765 5795 13795
rect 5925 13765 5955 13795
rect 6005 13765 6035 13795
rect 6165 13765 6195 13795
rect 4245 13685 4275 13715
rect 4405 13685 4435 13715
rect 4485 13685 4515 13715
rect 4645 13685 4675 13715
rect 4725 13685 4755 13715
rect 4885 13685 4915 13715
rect 5045 13685 5075 13715
rect 5205 13685 5235 13715
rect 5365 13685 5395 13715
rect 5525 13685 5555 13715
rect 5685 13685 5715 13715
rect 5765 13685 5795 13715
rect 5925 13685 5955 13715
rect 6005 13685 6035 13715
rect 6165 13685 6195 13715
rect 4245 13605 4275 13635
rect 4405 13605 4435 13635
rect 4485 13605 4515 13635
rect 4645 13605 4675 13635
rect 4725 13605 4755 13635
rect 4885 13605 4915 13635
rect 5045 13605 5075 13635
rect 5205 13605 5235 13635
rect 5365 13605 5395 13635
rect 5525 13605 5555 13635
rect 5685 13605 5715 13635
rect 5765 13605 5795 13635
rect 5925 13605 5955 13635
rect 6005 13605 6035 13635
rect 6165 13605 6195 13635
rect 4245 13525 4275 13555
rect 4405 13525 4435 13555
rect 4485 13525 4515 13555
rect 4645 13525 4675 13555
rect 4725 13525 4755 13555
rect 4885 13525 4915 13555
rect 5045 13525 5075 13555
rect 5205 13525 5235 13555
rect 5365 13525 5395 13555
rect 5525 13525 5555 13555
rect 5685 13525 5715 13555
rect 5765 13525 5795 13555
rect 5925 13525 5955 13555
rect 6005 13525 6035 13555
rect 6165 13525 6195 13555
rect 4245 13445 4275 13475
rect 4405 13445 4435 13475
rect 4485 13445 4515 13475
rect 4645 13445 4675 13475
rect 4725 13445 4755 13475
rect 4885 13445 4915 13475
rect 5045 13445 5075 13475
rect 5205 13445 5235 13475
rect 5365 13445 5395 13475
rect 5525 13445 5555 13475
rect 5685 13445 5715 13475
rect 5765 13445 5795 13475
rect 5925 13445 5955 13475
rect 6005 13445 6035 13475
rect 6165 13445 6195 13475
rect 5285 13325 5315 13355
rect 5125 13165 5155 13195
rect 5285 13165 5315 13195
rect 4245 13045 4275 13075
rect 4405 13045 4435 13075
rect 4485 13045 4515 13075
rect 4645 13045 4675 13075
rect 4725 13045 4755 13075
rect 4885 13045 4915 13075
rect 5045 13045 5075 13075
rect 5205 13045 5235 13075
rect 5365 13045 5395 13075
rect 5525 13045 5555 13075
rect 5685 13045 5715 13075
rect 5765 13045 5795 13075
rect 5925 13045 5955 13075
rect 6005 13045 6035 13075
rect 6165 13045 6195 13075
rect 4245 12965 4275 12995
rect 4405 12965 4435 12995
rect 4485 12965 4515 12995
rect 4645 12965 4675 12995
rect 4725 12965 4755 12995
rect 4885 12965 4915 12995
rect 5045 12965 5075 12995
rect 5205 12965 5235 12995
rect 5365 12965 5395 12995
rect 5525 12965 5555 12995
rect 5685 12965 5715 12995
rect 5765 12965 5795 12995
rect 5925 12965 5955 12995
rect 6005 12965 6035 12995
rect 6165 12965 6195 12995
rect 4245 12885 4275 12915
rect 4405 12885 4435 12915
rect 4485 12885 4515 12915
rect 4645 12885 4675 12915
rect 4725 12885 4755 12915
rect 4885 12885 4915 12915
rect 5045 12885 5075 12915
rect 5205 12885 5235 12915
rect 5365 12885 5395 12915
rect 5525 12885 5555 12915
rect 5685 12885 5715 12915
rect 5765 12885 5795 12915
rect 5925 12885 5955 12915
rect 6005 12885 6035 12915
rect 6165 12885 6195 12915
rect 4245 12805 4275 12835
rect 4405 12805 4435 12835
rect 4485 12805 4515 12835
rect 4645 12805 4675 12835
rect 4725 12805 4755 12835
rect 4885 12805 4915 12835
rect 5045 12805 5075 12835
rect 5205 12805 5235 12835
rect 5365 12805 5395 12835
rect 5525 12805 5555 12835
rect 5685 12805 5715 12835
rect 5765 12805 5795 12835
rect 5925 12805 5955 12835
rect 6005 12805 6035 12835
rect 6165 12805 6195 12835
rect 4245 12725 4275 12755
rect 4405 12725 4435 12755
rect 4485 12725 4515 12755
rect 4645 12725 4675 12755
rect 4725 12725 4755 12755
rect 4885 12725 4915 12755
rect 5045 12725 5075 12755
rect 5205 12725 5235 12755
rect 5365 12725 5395 12755
rect 5525 12725 5555 12755
rect 5685 12725 5715 12755
rect 5765 12725 5795 12755
rect 5925 12725 5955 12755
rect 6005 12725 6035 12755
rect 6165 12725 6195 12755
rect 4245 12645 4275 12675
rect 4405 12645 4435 12675
rect 4485 12645 4515 12675
rect 4645 12645 4675 12675
rect 4725 12645 4755 12675
rect 4885 12645 4915 12675
rect 5045 12645 5075 12675
rect 5205 12645 5235 12675
rect 5365 12645 5395 12675
rect 5525 12645 5555 12675
rect 5685 12645 5715 12675
rect 5765 12645 5795 12675
rect 5925 12645 5955 12675
rect 6005 12645 6035 12675
rect 6165 12645 6195 12675
rect 4245 12565 4275 12595
rect 4405 12565 4435 12595
rect 4485 12565 4515 12595
rect 4645 12565 4675 12595
rect 4725 12565 4755 12595
rect 4885 12565 4915 12595
rect 5045 12565 5075 12595
rect 5205 12565 5235 12595
rect 5365 12565 5395 12595
rect 5525 12565 5555 12595
rect 5685 12565 5715 12595
rect 5765 12565 5795 12595
rect 5925 12565 5955 12595
rect 6005 12565 6035 12595
rect 6165 12565 6195 12595
rect 4245 12485 4275 12515
rect 4405 12485 4435 12515
rect 4485 12485 4515 12515
rect 4645 12485 4675 12515
rect 4725 12485 4755 12515
rect 4885 12485 4915 12515
rect 5045 12485 5075 12515
rect 5205 12485 5235 12515
rect 5365 12485 5395 12515
rect 5525 12485 5555 12515
rect 5685 12485 5715 12515
rect 5765 12485 5795 12515
rect 5925 12485 5955 12515
rect 6005 12485 6035 12515
rect 6165 12485 6195 12515
rect 4565 12405 4595 12435
rect 4245 12325 4275 12355
rect 4405 12325 4435 12355
rect 4485 12325 4515 12355
rect 4645 12325 4675 12355
rect 4725 12325 4755 12355
rect 4885 12325 4915 12355
rect 5045 12325 5075 12355
rect 5205 12325 5235 12355
rect 5365 12325 5395 12355
rect 5525 12325 5555 12355
rect 5685 12325 5715 12355
rect 5765 12325 5795 12355
rect 5925 12325 5955 12355
rect 6005 12325 6035 12355
rect 6165 12325 6195 12355
rect 4245 12245 4275 12275
rect 4405 12245 4435 12275
rect 4485 12245 4515 12275
rect 4645 12245 4675 12275
rect 4725 12245 4755 12275
rect 4885 12245 4915 12275
rect 5045 12245 5075 12275
rect 5205 12245 5235 12275
rect 5365 12245 5395 12275
rect 5525 12245 5555 12275
rect 5685 12245 5715 12275
rect 5765 12245 5795 12275
rect 5925 12245 5955 12275
rect 6005 12245 6035 12275
rect 6165 12245 6195 12275
rect 4245 12165 4275 12195
rect 4405 12165 4435 12195
rect 4485 12165 4515 12195
rect 4645 12165 4675 12195
rect 4725 12165 4755 12195
rect 4885 12165 4915 12195
rect 5045 12165 5075 12195
rect 5205 12165 5235 12195
rect 5365 12165 5395 12195
rect 5525 12165 5555 12195
rect 5685 12165 5715 12195
rect 5765 12165 5795 12195
rect 5925 12165 5955 12195
rect 6005 12165 6035 12195
rect 6165 12165 6195 12195
rect 4245 12085 4275 12115
rect 4405 12085 4435 12115
rect 4485 12085 4515 12115
rect 4645 12085 4675 12115
rect 4725 12085 4755 12115
rect 4885 12085 4915 12115
rect 5045 12085 5075 12115
rect 5205 12085 5235 12115
rect 5365 12085 5395 12115
rect 5525 12085 5555 12115
rect 5685 12085 5715 12115
rect 5765 12085 5795 12115
rect 5925 12085 5955 12115
rect 6005 12085 6035 12115
rect 6165 12085 6195 12115
rect 4245 12005 4275 12035
rect 4405 12005 4435 12035
rect 4485 12005 4515 12035
rect 4645 12005 4675 12035
rect 4725 12005 4755 12035
rect 4885 12005 4915 12035
rect 5045 12005 5075 12035
rect 5205 12005 5235 12035
rect 5365 12005 5395 12035
rect 5525 12005 5555 12035
rect 5685 12005 5715 12035
rect 5765 12005 5795 12035
rect 5925 12005 5955 12035
rect 6005 12005 6035 12035
rect 6165 12005 6195 12035
rect 4245 11925 4275 11955
rect 4405 11925 4435 11955
rect 4485 11925 4515 11955
rect 4645 11925 4675 11955
rect 4725 11925 4755 11955
rect 4885 11925 4915 11955
rect 5045 11925 5075 11955
rect 5205 11925 5235 11955
rect 5365 11925 5395 11955
rect 5525 11925 5555 11955
rect 5685 11925 5715 11955
rect 5765 11925 5795 11955
rect 5925 11925 5955 11955
rect 6005 11925 6035 11955
rect 6165 11925 6195 11955
rect 4245 11845 4275 11875
rect 4405 11845 4435 11875
rect 4485 11845 4515 11875
rect 4645 11845 4675 11875
rect 4725 11845 4755 11875
rect 4885 11845 4915 11875
rect 5045 11845 5075 11875
rect 5205 11845 5235 11875
rect 5365 11845 5395 11875
rect 5525 11845 5555 11875
rect 5685 11845 5715 11875
rect 5765 11845 5795 11875
rect 5925 11845 5955 11875
rect 6005 11845 6035 11875
rect 6165 11845 6195 11875
rect 4245 11765 4275 11795
rect 4405 11765 4435 11795
rect 4485 11765 4515 11795
rect 4645 11765 4675 11795
rect 4725 11765 4755 11795
rect 4885 11765 4915 11795
rect 5045 11765 5075 11795
rect 5205 11765 5235 11795
rect 5365 11765 5395 11795
rect 5525 11765 5555 11795
rect 5685 11765 5715 11795
rect 5765 11765 5795 11795
rect 5925 11765 5955 11795
rect 6005 11765 6035 11795
rect 6165 11765 6195 11795
rect 4245 11685 4275 11715
rect 4405 11685 4435 11715
rect 4485 11685 4515 11715
rect 4645 11685 4675 11715
rect 4725 11685 4755 11715
rect 4885 11685 4915 11715
rect 5045 11685 5075 11715
rect 5205 11685 5235 11715
rect 5365 11685 5395 11715
rect 5525 11685 5555 11715
rect 5685 11685 5715 11715
rect 5765 11685 5795 11715
rect 5925 11685 5955 11715
rect 6005 11685 6035 11715
rect 6165 11685 6195 11715
rect 4245 11605 4275 11635
rect 4405 11605 4435 11635
rect 4485 11605 4515 11635
rect 4645 11605 4675 11635
rect 4725 11605 4755 11635
rect 4885 11605 4915 11635
rect 5045 11605 5075 11635
rect 5205 11605 5235 11635
rect 5365 11605 5395 11635
rect 5525 11605 5555 11635
rect 5685 11605 5715 11635
rect 5765 11605 5795 11635
rect 5925 11605 5955 11635
rect 6005 11605 6035 11635
rect 6165 11605 6195 11635
rect 4245 11525 4275 11555
rect 4405 11525 4435 11555
rect 4485 11525 4515 11555
rect 4645 11525 4675 11555
rect 4725 11525 4755 11555
rect 4885 11525 4915 11555
rect 5045 11525 5075 11555
rect 5205 11525 5235 11555
rect 5365 11525 5395 11555
rect 5525 11525 5555 11555
rect 5685 11525 5715 11555
rect 5765 11525 5795 11555
rect 5925 11525 5955 11555
rect 6005 11525 6035 11555
rect 6165 11525 6195 11555
rect 4245 11445 4275 11475
rect 4405 11445 4435 11475
rect 4485 11445 4515 11475
rect 4645 11445 4675 11475
rect 4725 11445 4755 11475
rect 4885 11445 4915 11475
rect 5045 11445 5075 11475
rect 5205 11445 5235 11475
rect 5365 11445 5395 11475
rect 5525 11445 5555 11475
rect 5685 11445 5715 11475
rect 5765 11445 5795 11475
rect 5925 11445 5955 11475
rect 6005 11445 6035 11475
rect 6165 11445 6195 11475
rect 4245 11365 4275 11395
rect 4405 11365 4435 11395
rect 4485 11365 4515 11395
rect 4645 11365 4675 11395
rect 4725 11365 4755 11395
rect 4885 11365 4915 11395
rect 5045 11365 5075 11395
rect 5205 11365 5235 11395
rect 5365 11365 5395 11395
rect 5525 11365 5555 11395
rect 5685 11365 5715 11395
rect 5765 11365 5795 11395
rect 5925 11365 5955 11395
rect 6005 11365 6035 11395
rect 6165 11365 6195 11395
rect 4245 11285 4275 11315
rect 4405 11285 4435 11315
rect 4485 11285 4515 11315
rect 4645 11285 4675 11315
rect 4725 11285 4755 11315
rect 4885 11285 4915 11315
rect 5045 11285 5075 11315
rect 5205 11285 5235 11315
rect 5365 11285 5395 11315
rect 5525 11285 5555 11315
rect 5685 11285 5715 11315
rect 5765 11285 5795 11315
rect 5925 11285 5955 11315
rect 6005 11285 6035 11315
rect 6165 11285 6195 11315
rect 4245 11205 4275 11235
rect 4405 11205 4435 11235
rect 4485 11205 4515 11235
rect 4645 11205 4675 11235
rect 4725 11205 4755 11235
rect 4885 11205 4915 11235
rect 5045 11205 5075 11235
rect 5205 11205 5235 11235
rect 5365 11205 5395 11235
rect 5525 11205 5555 11235
rect 5685 11205 5715 11235
rect 5765 11205 5795 11235
rect 5925 11205 5955 11235
rect 6005 11205 6035 11235
rect 6165 11205 6195 11235
rect 4245 11125 4275 11155
rect 4405 11125 4435 11155
rect 4485 11125 4515 11155
rect 4645 11125 4675 11155
rect 4725 11125 4755 11155
rect 4885 11125 4915 11155
rect 5045 11125 5075 11155
rect 5205 11125 5235 11155
rect 5365 11125 5395 11155
rect 5525 11125 5555 11155
rect 5685 11125 5715 11155
rect 5765 11125 5795 11155
rect 5925 11125 5955 11155
rect 6005 11125 6035 11155
rect 6165 11125 6195 11155
rect 4245 11045 4275 11075
rect 4405 11045 4435 11075
rect 4485 11045 4515 11075
rect 4645 11045 4675 11075
rect 4725 11045 4755 11075
rect 4885 11045 4915 11075
rect 5045 11045 5075 11075
rect 5205 11045 5235 11075
rect 5365 11045 5395 11075
rect 5525 11045 5555 11075
rect 5685 11045 5715 11075
rect 5765 11045 5795 11075
rect 5925 11045 5955 11075
rect 6005 11045 6035 11075
rect 6165 11045 6195 11075
rect 4565 10965 4595 10995
rect 4245 10885 4275 10915
rect 4405 10885 4435 10915
rect 4485 10885 4515 10915
rect 4645 10885 4675 10915
rect 4725 10885 4755 10915
rect 4885 10885 4915 10915
rect 5045 10885 5075 10915
rect 5205 10885 5235 10915
rect 5365 10885 5395 10915
rect 5525 10885 5555 10915
rect 5685 10885 5715 10915
rect 5765 10885 5795 10915
rect 5925 10885 5955 10915
rect 6005 10885 6035 10915
rect 6165 10885 6195 10915
rect 4245 10805 4275 10835
rect 4405 10805 4435 10835
rect 4485 10805 4515 10835
rect 4645 10805 4675 10835
rect 4725 10805 4755 10835
rect 4885 10805 4915 10835
rect 5045 10805 5075 10835
rect 5205 10805 5235 10835
rect 5365 10805 5395 10835
rect 5525 10805 5555 10835
rect 5685 10805 5715 10835
rect 5765 10805 5795 10835
rect 5925 10805 5955 10835
rect 6005 10805 6035 10835
rect 6165 10805 6195 10835
rect 4245 10725 4275 10755
rect 4405 10725 4435 10755
rect 4485 10725 4515 10755
rect 4645 10725 4675 10755
rect 4725 10725 4755 10755
rect 4885 10725 4915 10755
rect 5045 10725 5075 10755
rect 5205 10725 5235 10755
rect 5365 10725 5395 10755
rect 5525 10725 5555 10755
rect 5685 10725 5715 10755
rect 5765 10725 5795 10755
rect 5925 10725 5955 10755
rect 6005 10725 6035 10755
rect 6165 10725 6195 10755
rect 4245 10645 4275 10675
rect 4405 10645 4435 10675
rect 4485 10645 4515 10675
rect 4645 10645 4675 10675
rect 4725 10645 4755 10675
rect 4885 10645 4915 10675
rect 5045 10645 5075 10675
rect 5205 10645 5235 10675
rect 5365 10645 5395 10675
rect 5525 10645 5555 10675
rect 5685 10645 5715 10675
rect 5765 10645 5795 10675
rect 5925 10645 5955 10675
rect 6005 10645 6035 10675
rect 6165 10645 6195 10675
rect 4245 10565 4275 10595
rect 4405 10565 4435 10595
rect 4485 10565 4515 10595
rect 4645 10565 4675 10595
rect 4725 10565 4755 10595
rect 4885 10565 4915 10595
rect 5045 10565 5075 10595
rect 5205 10565 5235 10595
rect 5365 10565 5395 10595
rect 5525 10565 5555 10595
rect 5685 10565 5715 10595
rect 5765 10565 5795 10595
rect 5925 10565 5955 10595
rect 6005 10565 6035 10595
rect 6165 10565 6195 10595
rect 4245 10485 4275 10515
rect 4405 10485 4435 10515
rect 4485 10485 4515 10515
rect 4645 10485 4675 10515
rect 4725 10485 4755 10515
rect 4885 10485 4915 10515
rect 5045 10485 5075 10515
rect 5205 10485 5235 10515
rect 5365 10485 5395 10515
rect 5525 10485 5555 10515
rect 5685 10485 5715 10515
rect 5765 10485 5795 10515
rect 5925 10485 5955 10515
rect 6005 10485 6035 10515
rect 6165 10485 6195 10515
rect 4245 10405 4275 10435
rect 4405 10405 4435 10435
rect 4485 10405 4515 10435
rect 4645 10405 4675 10435
rect 4725 10405 4755 10435
rect 4885 10405 4915 10435
rect 5045 10405 5075 10435
rect 5205 10405 5235 10435
rect 5365 10405 5395 10435
rect 5525 10405 5555 10435
rect 5685 10405 5715 10435
rect 5765 10405 5795 10435
rect 5925 10405 5955 10435
rect 6005 10405 6035 10435
rect 6165 10405 6195 10435
rect 4245 10325 4275 10355
rect 4405 10325 4435 10355
rect 4485 10325 4515 10355
rect 4645 10325 4675 10355
rect 4725 10325 4755 10355
rect 4885 10325 4915 10355
rect 5045 10325 5075 10355
rect 5205 10325 5235 10355
rect 5365 10325 5395 10355
rect 5525 10325 5555 10355
rect 5685 10325 5715 10355
rect 5765 10325 5795 10355
rect 5925 10325 5955 10355
rect 6005 10325 6035 10355
rect 6165 10325 6195 10355
rect 5125 10205 5155 10235
rect 5125 10045 5155 10075
rect 4245 9925 4275 9955
rect 4405 9925 4435 9955
rect 4485 9925 4515 9955
rect 4645 9925 4675 9955
rect 4725 9925 4755 9955
rect 4885 9925 4915 9955
rect 5045 9925 5075 9955
rect 5205 9925 5235 9955
rect 5365 9925 5395 9955
rect 5525 9925 5555 9955
rect 5685 9925 5715 9955
rect 5765 9925 5795 9955
rect 5925 9925 5955 9955
rect 6005 9925 6035 9955
rect 6165 9925 6195 9955
rect 4245 9845 4275 9875
rect 4405 9845 4435 9875
rect 4485 9845 4515 9875
rect 4645 9845 4675 9875
rect 4725 9845 4755 9875
rect 4885 9845 4915 9875
rect 5045 9845 5075 9875
rect 5205 9845 5235 9875
rect 5365 9845 5395 9875
rect 5525 9845 5555 9875
rect 5685 9845 5715 9875
rect 5765 9845 5795 9875
rect 5925 9845 5955 9875
rect 6005 9845 6035 9875
rect 6165 9845 6195 9875
rect 4245 9765 4275 9795
rect 4405 9765 4435 9795
rect 4485 9765 4515 9795
rect 4645 9765 4675 9795
rect 4725 9765 4755 9795
rect 4885 9765 4915 9795
rect 5045 9765 5075 9795
rect 5205 9765 5235 9795
rect 5365 9765 5395 9795
rect 5525 9765 5555 9795
rect 5685 9765 5715 9795
rect 5765 9765 5795 9795
rect 5925 9765 5955 9795
rect 6005 9765 6035 9795
rect 6165 9765 6195 9795
rect 4245 9685 4275 9715
rect 4405 9685 4435 9715
rect 4485 9685 4515 9715
rect 4645 9685 4675 9715
rect 4725 9685 4755 9715
rect 4885 9685 4915 9715
rect 5045 9685 5075 9715
rect 5205 9685 5235 9715
rect 5365 9685 5395 9715
rect 5525 9685 5555 9715
rect 5685 9685 5715 9715
rect 5765 9685 5795 9715
rect 5925 9685 5955 9715
rect 6005 9685 6035 9715
rect 6165 9685 6195 9715
rect 4245 9605 4275 9635
rect 4405 9605 4435 9635
rect 4485 9605 4515 9635
rect 4645 9605 4675 9635
rect 4725 9605 4755 9635
rect 4885 9605 4915 9635
rect 5045 9605 5075 9635
rect 5205 9605 5235 9635
rect 5365 9605 5395 9635
rect 5525 9605 5555 9635
rect 5685 9605 5715 9635
rect 5765 9605 5795 9635
rect 5925 9605 5955 9635
rect 6005 9605 6035 9635
rect 6165 9605 6195 9635
rect 4245 9525 4275 9555
rect 4405 9525 4435 9555
rect 4485 9525 4515 9555
rect 4645 9525 4675 9555
rect 4725 9525 4755 9555
rect 4885 9525 4915 9555
rect 5045 9525 5075 9555
rect 5205 9525 5235 9555
rect 5365 9525 5395 9555
rect 5525 9525 5555 9555
rect 5685 9525 5715 9555
rect 5765 9525 5795 9555
rect 5925 9525 5955 9555
rect 6005 9525 6035 9555
rect 6165 9525 6195 9555
rect 4245 9445 4275 9475
rect 4405 9445 4435 9475
rect 4485 9445 4515 9475
rect 4645 9445 4675 9475
rect 4725 9445 4755 9475
rect 4885 9445 4915 9475
rect 5045 9445 5075 9475
rect 5205 9445 5235 9475
rect 5365 9445 5395 9475
rect 5525 9445 5555 9475
rect 5685 9445 5715 9475
rect 5765 9445 5795 9475
rect 5925 9445 5955 9475
rect 6005 9445 6035 9475
rect 6165 9445 6195 9475
rect 4245 9365 4275 9395
rect 4405 9365 4435 9395
rect 4485 9365 4515 9395
rect 4645 9365 4675 9395
rect 4725 9365 4755 9395
rect 4885 9365 4915 9395
rect 5045 9365 5075 9395
rect 5205 9365 5235 9395
rect 5365 9365 5395 9395
rect 5525 9365 5555 9395
rect 5685 9365 5715 9395
rect 5765 9365 5795 9395
rect 5925 9365 5955 9395
rect 6005 9365 6035 9395
rect 6165 9365 6195 9395
rect 5125 9245 5155 9275
rect 4965 9085 4995 9115
rect 5445 9085 5475 9115
rect 4245 8965 4275 8995
rect 4405 8965 4435 8995
rect 4485 8965 4515 8995
rect 4645 8965 4675 8995
rect 4725 8965 4755 8995
rect 4885 8965 4915 8995
rect 5045 8965 5075 8995
rect 5205 8965 5235 8995
rect 5365 8965 5395 8995
rect 5525 8965 5555 8995
rect 5685 8965 5715 8995
rect 5765 8965 5795 8995
rect 5925 8965 5955 8995
rect 6005 8965 6035 8995
rect 6165 8965 6195 8995
rect 4245 8885 4275 8915
rect 4405 8885 4435 8915
rect 4485 8885 4515 8915
rect 4645 8885 4675 8915
rect 4725 8885 4755 8915
rect 4885 8885 4915 8915
rect 5045 8885 5075 8915
rect 5205 8885 5235 8915
rect 5365 8885 5395 8915
rect 5525 8885 5555 8915
rect 5685 8885 5715 8915
rect 5765 8885 5795 8915
rect 5925 8885 5955 8915
rect 6005 8885 6035 8915
rect 6165 8885 6195 8915
rect 4245 8805 4275 8835
rect 4405 8805 4435 8835
rect 4485 8805 4515 8835
rect 4645 8805 4675 8835
rect 4725 8805 4755 8835
rect 4885 8805 4915 8835
rect 5045 8805 5075 8835
rect 5205 8805 5235 8835
rect 5365 8805 5395 8835
rect 5525 8805 5555 8835
rect 5685 8805 5715 8835
rect 5765 8805 5795 8835
rect 5925 8805 5955 8835
rect 6005 8805 6035 8835
rect 6165 8805 6195 8835
rect 4245 8725 4275 8755
rect 4405 8725 4435 8755
rect 4485 8725 4515 8755
rect 4645 8725 4675 8755
rect 4725 8725 4755 8755
rect 4885 8725 4915 8755
rect 5045 8725 5075 8755
rect 5205 8725 5235 8755
rect 5365 8725 5395 8755
rect 5525 8725 5555 8755
rect 5685 8725 5715 8755
rect 5765 8725 5795 8755
rect 5925 8725 5955 8755
rect 6005 8725 6035 8755
rect 6165 8725 6195 8755
rect 4245 8645 4275 8675
rect 4405 8645 4435 8675
rect 4485 8645 4515 8675
rect 4645 8645 4675 8675
rect 4725 8645 4755 8675
rect 4885 8645 4915 8675
rect 5045 8645 5075 8675
rect 5205 8645 5235 8675
rect 5365 8645 5395 8675
rect 5525 8645 5555 8675
rect 5685 8645 5715 8675
rect 5765 8645 5795 8675
rect 5925 8645 5955 8675
rect 6005 8645 6035 8675
rect 6165 8645 6195 8675
rect 4245 8565 4275 8595
rect 4405 8565 4435 8595
rect 4485 8565 4515 8595
rect 4645 8565 4675 8595
rect 4725 8565 4755 8595
rect 4885 8565 4915 8595
rect 5045 8565 5075 8595
rect 5205 8565 5235 8595
rect 5365 8565 5395 8595
rect 5525 8565 5555 8595
rect 5685 8565 5715 8595
rect 5765 8565 5795 8595
rect 5925 8565 5955 8595
rect 6005 8565 6035 8595
rect 6165 8565 6195 8595
rect 4245 8485 4275 8515
rect 4405 8485 4435 8515
rect 4485 8485 4515 8515
rect 4645 8485 4675 8515
rect 4725 8485 4755 8515
rect 4885 8485 4915 8515
rect 5045 8485 5075 8515
rect 5205 8485 5235 8515
rect 5365 8485 5395 8515
rect 5525 8485 5555 8515
rect 5685 8485 5715 8515
rect 5765 8485 5795 8515
rect 5925 8485 5955 8515
rect 6005 8485 6035 8515
rect 6165 8485 6195 8515
rect 4245 8405 4275 8435
rect 4405 8405 4435 8435
rect 4485 8405 4515 8435
rect 4645 8405 4675 8435
rect 4725 8405 4755 8435
rect 4885 8405 4915 8435
rect 5045 8405 5075 8435
rect 5205 8405 5235 8435
rect 5365 8405 5395 8435
rect 5525 8405 5555 8435
rect 5685 8405 5715 8435
rect 5765 8405 5795 8435
rect 5925 8405 5955 8435
rect 6005 8405 6035 8435
rect 6165 8405 6195 8435
rect 4565 8325 4595 8355
rect 4245 8245 4275 8275
rect 4405 8245 4435 8275
rect 4485 8245 4515 8275
rect 4645 8245 4675 8275
rect 4725 8245 4755 8275
rect 4885 8245 4915 8275
rect 5045 8245 5075 8275
rect 5205 8245 5235 8275
rect 5365 8245 5395 8275
rect 5525 8245 5555 8275
rect 5685 8245 5715 8275
rect 5765 8245 5795 8275
rect 5925 8245 5955 8275
rect 6005 8245 6035 8275
rect 6165 8245 6195 8275
rect 4245 8165 4275 8195
rect 4405 8165 4435 8195
rect 4485 8165 4515 8195
rect 4645 8165 4675 8195
rect 4725 8165 4755 8195
rect 4885 8165 4915 8195
rect 5045 8165 5075 8195
rect 5205 8165 5235 8195
rect 5365 8165 5395 8195
rect 5525 8165 5555 8195
rect 5685 8165 5715 8195
rect 5765 8165 5795 8195
rect 5925 8165 5955 8195
rect 6005 8165 6035 8195
rect 6165 8165 6195 8195
rect 4245 8085 4275 8115
rect 4405 8085 4435 8115
rect 4485 8085 4515 8115
rect 4645 8085 4675 8115
rect 4725 8085 4755 8115
rect 4885 8085 4915 8115
rect 5045 8085 5075 8115
rect 5205 8085 5235 8115
rect 5365 8085 5395 8115
rect 5525 8085 5555 8115
rect 5685 8085 5715 8115
rect 5765 8085 5795 8115
rect 5925 8085 5955 8115
rect 6005 8085 6035 8115
rect 6165 8085 6195 8115
rect 4245 8005 4275 8035
rect 4405 8005 4435 8035
rect 4485 8005 4515 8035
rect 4645 8005 4675 8035
rect 4725 8005 4755 8035
rect 4885 8005 4915 8035
rect 5045 8005 5075 8035
rect 5205 8005 5235 8035
rect 5365 8005 5395 8035
rect 5525 8005 5555 8035
rect 5685 8005 5715 8035
rect 5765 8005 5795 8035
rect 5925 8005 5955 8035
rect 6005 8005 6035 8035
rect 6165 8005 6195 8035
rect 4245 7925 4275 7955
rect 4405 7925 4435 7955
rect 4485 7925 4515 7955
rect 4645 7925 4675 7955
rect 4725 7925 4755 7955
rect 4885 7925 4915 7955
rect 5045 7925 5075 7955
rect 5205 7925 5235 7955
rect 5365 7925 5395 7955
rect 5525 7925 5555 7955
rect 5685 7925 5715 7955
rect 5765 7925 5795 7955
rect 5925 7925 5955 7955
rect 6005 7925 6035 7955
rect 6165 7925 6195 7955
rect 4245 7845 4275 7875
rect 4405 7845 4435 7875
rect 4485 7845 4515 7875
rect 4645 7845 4675 7875
rect 4725 7845 4755 7875
rect 4885 7845 4915 7875
rect 5045 7845 5075 7875
rect 5205 7845 5235 7875
rect 5365 7845 5395 7875
rect 5525 7845 5555 7875
rect 5685 7845 5715 7875
rect 5765 7845 5795 7875
rect 5925 7845 5955 7875
rect 6005 7845 6035 7875
rect 6165 7845 6195 7875
rect 4245 7765 4275 7795
rect 4405 7765 4435 7795
rect 4485 7765 4515 7795
rect 4645 7765 4675 7795
rect 4725 7765 4755 7795
rect 4885 7765 4915 7795
rect 5045 7765 5075 7795
rect 5205 7765 5235 7795
rect 5365 7765 5395 7795
rect 5525 7765 5555 7795
rect 5685 7765 5715 7795
rect 5765 7765 5795 7795
rect 5925 7765 5955 7795
rect 6005 7765 6035 7795
rect 6165 7765 6195 7795
rect 4245 7685 4275 7715
rect 4405 7685 4435 7715
rect 4485 7685 4515 7715
rect 4645 7685 4675 7715
rect 4725 7685 4755 7715
rect 4885 7685 4915 7715
rect 5045 7685 5075 7715
rect 5205 7685 5235 7715
rect 5365 7685 5395 7715
rect 5525 7685 5555 7715
rect 5685 7685 5715 7715
rect 5765 7685 5795 7715
rect 5925 7685 5955 7715
rect 6005 7685 6035 7715
rect 6165 7685 6195 7715
rect 4245 7605 4275 7635
rect 4405 7605 4435 7635
rect 4485 7605 4515 7635
rect 4645 7605 4675 7635
rect 4725 7605 4755 7635
rect 4885 7605 4915 7635
rect 5045 7605 5075 7635
rect 5205 7605 5235 7635
rect 5365 7605 5395 7635
rect 5525 7605 5555 7635
rect 5685 7605 5715 7635
rect 5765 7605 5795 7635
rect 5925 7605 5955 7635
rect 6005 7605 6035 7635
rect 6165 7605 6195 7635
rect 4245 7525 4275 7555
rect 4405 7525 4435 7555
rect 4485 7525 4515 7555
rect 4645 7525 4675 7555
rect 4725 7525 4755 7555
rect 4885 7525 4915 7555
rect 5045 7525 5075 7555
rect 5205 7525 5235 7555
rect 5365 7525 5395 7555
rect 5525 7525 5555 7555
rect 5685 7525 5715 7555
rect 5765 7525 5795 7555
rect 5925 7525 5955 7555
rect 6005 7525 6035 7555
rect 6165 7525 6195 7555
rect 4245 7445 4275 7475
rect 4405 7445 4435 7475
rect 4485 7445 4515 7475
rect 4645 7445 4675 7475
rect 4725 7445 4755 7475
rect 4885 7445 4915 7475
rect 5045 7445 5075 7475
rect 5205 7445 5235 7475
rect 5365 7445 5395 7475
rect 5525 7445 5555 7475
rect 5685 7445 5715 7475
rect 5765 7445 5795 7475
rect 5925 7445 5955 7475
rect 6005 7445 6035 7475
rect 6165 7445 6195 7475
rect 4245 7365 4275 7395
rect 4405 7365 4435 7395
rect 4485 7365 4515 7395
rect 4645 7365 4675 7395
rect 4725 7365 4755 7395
rect 4885 7365 4915 7395
rect 5045 7365 5075 7395
rect 5205 7365 5235 7395
rect 5365 7365 5395 7395
rect 5525 7365 5555 7395
rect 5685 7365 5715 7395
rect 5765 7365 5795 7395
rect 5925 7365 5955 7395
rect 6005 7365 6035 7395
rect 6165 7365 6195 7395
rect 4245 7285 4275 7315
rect 4405 7285 4435 7315
rect 4485 7285 4515 7315
rect 4645 7285 4675 7315
rect 4725 7285 4755 7315
rect 4885 7285 4915 7315
rect 5045 7285 5075 7315
rect 5205 7285 5235 7315
rect 5365 7285 5395 7315
rect 5525 7285 5555 7315
rect 5685 7285 5715 7315
rect 5765 7285 5795 7315
rect 5925 7285 5955 7315
rect 6005 7285 6035 7315
rect 6165 7285 6195 7315
rect 4245 7205 4275 7235
rect 4405 7205 4435 7235
rect 4485 7205 4515 7235
rect 4645 7205 4675 7235
rect 4725 7205 4755 7235
rect 4885 7205 4915 7235
rect 5045 7205 5075 7235
rect 5205 7205 5235 7235
rect 5365 7205 5395 7235
rect 5525 7205 5555 7235
rect 5685 7205 5715 7235
rect 5765 7205 5795 7235
rect 5925 7205 5955 7235
rect 6005 7205 6035 7235
rect 6165 7205 6195 7235
rect 4245 7125 4275 7155
rect 4405 7125 4435 7155
rect 4485 7125 4515 7155
rect 4645 7125 4675 7155
rect 4725 7125 4755 7155
rect 4885 7125 4915 7155
rect 5045 7125 5075 7155
rect 5205 7125 5235 7155
rect 5365 7125 5395 7155
rect 5525 7125 5555 7155
rect 5685 7125 5715 7155
rect 5765 7125 5795 7155
rect 5925 7125 5955 7155
rect 6005 7125 6035 7155
rect 6165 7125 6195 7155
rect 4245 7045 4275 7075
rect 4405 7045 4435 7075
rect 4485 7045 4515 7075
rect 4645 7045 4675 7075
rect 4725 7045 4755 7075
rect 4885 7045 4915 7075
rect 5045 7045 5075 7075
rect 5205 7045 5235 7075
rect 5365 7045 5395 7075
rect 5525 7045 5555 7075
rect 5685 7045 5715 7075
rect 5765 7045 5795 7075
rect 5925 7045 5955 7075
rect 6005 7045 6035 7075
rect 6165 7045 6195 7075
rect 4245 6965 4275 6995
rect 4405 6965 4435 6995
rect 4485 6965 4515 6995
rect 4645 6965 4675 6995
rect 4725 6965 4755 6995
rect 4885 6965 4915 6995
rect 5045 6965 5075 6995
rect 5205 6965 5235 6995
rect 5365 6965 5395 6995
rect 5525 6965 5555 6995
rect 5685 6965 5715 6995
rect 5765 6965 5795 6995
rect 5925 6965 5955 6995
rect 6005 6965 6035 6995
rect 6165 6965 6195 6995
rect 4565 6885 4595 6915
rect 4245 6805 4275 6835
rect 4405 6805 4435 6835
rect 4485 6805 4515 6835
rect 4645 6805 4675 6835
rect 4725 6805 4755 6835
rect 4885 6805 4915 6835
rect 5045 6805 5075 6835
rect 5205 6805 5235 6835
rect 5365 6805 5395 6835
rect 5525 6805 5555 6835
rect 5685 6805 5715 6835
rect 5765 6805 5795 6835
rect 5925 6805 5955 6835
rect 6005 6805 6035 6835
rect 6165 6805 6195 6835
rect 4245 6725 4275 6755
rect 4405 6725 4435 6755
rect 4485 6725 4515 6755
rect 4645 6725 4675 6755
rect 4725 6725 4755 6755
rect 4885 6725 4915 6755
rect 5045 6725 5075 6755
rect 5205 6725 5235 6755
rect 5365 6725 5395 6755
rect 5525 6725 5555 6755
rect 5685 6725 5715 6755
rect 5765 6725 5795 6755
rect 5925 6725 5955 6755
rect 6005 6725 6035 6755
rect 6165 6725 6195 6755
rect 4245 6645 4275 6675
rect 4405 6645 4435 6675
rect 4485 6645 4515 6675
rect 4645 6645 4675 6675
rect 4725 6645 4755 6675
rect 4885 6645 4915 6675
rect 5045 6645 5075 6675
rect 5205 6645 5235 6675
rect 5365 6645 5395 6675
rect 5525 6645 5555 6675
rect 5685 6645 5715 6675
rect 5765 6645 5795 6675
rect 5925 6645 5955 6675
rect 6005 6645 6035 6675
rect 6165 6645 6195 6675
rect 4245 6565 4275 6595
rect 4405 6565 4435 6595
rect 4485 6565 4515 6595
rect 4645 6565 4675 6595
rect 4725 6565 4755 6595
rect 4885 6565 4915 6595
rect 5045 6565 5075 6595
rect 5205 6565 5235 6595
rect 5365 6565 5395 6595
rect 5525 6565 5555 6595
rect 5685 6565 5715 6595
rect 5765 6565 5795 6595
rect 5925 6565 5955 6595
rect 6005 6565 6035 6595
rect 6165 6565 6195 6595
rect 4245 6485 4275 6515
rect 4405 6485 4435 6515
rect 4485 6485 4515 6515
rect 4645 6485 4675 6515
rect 4725 6485 4755 6515
rect 4885 6485 4915 6515
rect 5045 6485 5075 6515
rect 5205 6485 5235 6515
rect 5365 6485 5395 6515
rect 5525 6485 5555 6515
rect 5685 6485 5715 6515
rect 5765 6485 5795 6515
rect 5925 6485 5955 6515
rect 6005 6485 6035 6515
rect 6165 6485 6195 6515
rect 4245 6405 4275 6435
rect 4405 6405 4435 6435
rect 4485 6405 4515 6435
rect 4645 6405 4675 6435
rect 4725 6405 4755 6435
rect 4885 6405 4915 6435
rect 5045 6405 5075 6435
rect 5205 6405 5235 6435
rect 5365 6405 5395 6435
rect 5525 6405 5555 6435
rect 5685 6405 5715 6435
rect 5765 6405 5795 6435
rect 5925 6405 5955 6435
rect 6005 6405 6035 6435
rect 6165 6405 6195 6435
rect 4245 6325 4275 6355
rect 4405 6325 4435 6355
rect 4485 6325 4515 6355
rect 4645 6325 4675 6355
rect 4725 6325 4755 6355
rect 4885 6325 4915 6355
rect 5045 6325 5075 6355
rect 5205 6325 5235 6355
rect 5365 6325 5395 6355
rect 5525 6325 5555 6355
rect 5685 6325 5715 6355
rect 5765 6325 5795 6355
rect 5925 6325 5955 6355
rect 6005 6325 6035 6355
rect 6165 6325 6195 6355
rect 4245 6245 4275 6275
rect 4405 6245 4435 6275
rect 4485 6245 4515 6275
rect 4645 6245 4675 6275
rect 4725 6245 4755 6275
rect 4885 6245 4915 6275
rect 5045 6245 5075 6275
rect 5205 6245 5235 6275
rect 5365 6245 5395 6275
rect 5525 6245 5555 6275
rect 5685 6245 5715 6275
rect 5765 6245 5795 6275
rect 5925 6245 5955 6275
rect 6005 6245 6035 6275
rect 6165 6245 6195 6275
rect 4805 6125 4835 6155
rect 5605 6125 5635 6155
rect 4965 5965 4995 5995
rect 5445 5965 5475 5995
rect 4245 5845 4275 5875
rect 4405 5845 4435 5875
rect 4485 5845 4515 5875
rect 4645 5845 4675 5875
rect 4725 5845 4755 5875
rect 4885 5845 4915 5875
rect 5045 5845 5075 5875
rect 5205 5845 5235 5875
rect 5365 5845 5395 5875
rect 5525 5845 5555 5875
rect 5685 5845 5715 5875
rect 5765 5845 5795 5875
rect 5925 5845 5955 5875
rect 6005 5845 6035 5875
rect 6165 5845 6195 5875
rect 4245 5765 4275 5795
rect 4405 5765 4435 5795
rect 4485 5765 4515 5795
rect 4645 5765 4675 5795
rect 4725 5765 4755 5795
rect 4885 5765 4915 5795
rect 5045 5765 5075 5795
rect 5205 5765 5235 5795
rect 5365 5765 5395 5795
rect 5525 5765 5555 5795
rect 5685 5765 5715 5795
rect 5765 5765 5795 5795
rect 5925 5765 5955 5795
rect 6005 5765 6035 5795
rect 6165 5765 6195 5795
rect 4245 5685 4275 5715
rect 4405 5685 4435 5715
rect 4485 5685 4515 5715
rect 4645 5685 4675 5715
rect 4725 5685 4755 5715
rect 4885 5685 4915 5715
rect 5045 5685 5075 5715
rect 5205 5685 5235 5715
rect 5365 5685 5395 5715
rect 5525 5685 5555 5715
rect 5685 5685 5715 5715
rect 5765 5685 5795 5715
rect 5925 5685 5955 5715
rect 6005 5685 6035 5715
rect 6165 5685 6195 5715
rect 4245 5605 4275 5635
rect 4405 5605 4435 5635
rect 4485 5605 4515 5635
rect 4645 5605 4675 5635
rect 4725 5605 4755 5635
rect 4885 5605 4915 5635
rect 5045 5605 5075 5635
rect 5205 5605 5235 5635
rect 5365 5605 5395 5635
rect 5525 5605 5555 5635
rect 5685 5605 5715 5635
rect 5765 5605 5795 5635
rect 5925 5605 5955 5635
rect 6005 5605 6035 5635
rect 6165 5605 6195 5635
rect 4245 5525 4275 5555
rect 4405 5525 4435 5555
rect 4485 5525 4515 5555
rect 4645 5525 4675 5555
rect 4725 5525 4755 5555
rect 4885 5525 4915 5555
rect 5045 5525 5075 5555
rect 5205 5525 5235 5555
rect 5365 5525 5395 5555
rect 5525 5525 5555 5555
rect 5685 5525 5715 5555
rect 5765 5525 5795 5555
rect 5925 5525 5955 5555
rect 6005 5525 6035 5555
rect 6165 5525 6195 5555
rect 4245 5445 4275 5475
rect 4405 5445 4435 5475
rect 4485 5445 4515 5475
rect 4645 5445 4675 5475
rect 4725 5445 4755 5475
rect 4885 5445 4915 5475
rect 5045 5445 5075 5475
rect 5205 5445 5235 5475
rect 5365 5445 5395 5475
rect 5525 5445 5555 5475
rect 5685 5445 5715 5475
rect 5765 5445 5795 5475
rect 5925 5445 5955 5475
rect 6005 5445 6035 5475
rect 6165 5445 6195 5475
rect 4245 5365 4275 5395
rect 4405 5365 4435 5395
rect 4485 5365 4515 5395
rect 4645 5365 4675 5395
rect 4725 5365 4755 5395
rect 4885 5365 4915 5395
rect 5045 5365 5075 5395
rect 5205 5365 5235 5395
rect 5365 5365 5395 5395
rect 5525 5365 5555 5395
rect 5685 5365 5715 5395
rect 5765 5365 5795 5395
rect 5925 5365 5955 5395
rect 6005 5365 6035 5395
rect 6165 5365 6195 5395
rect 4245 5285 4275 5315
rect 4405 5285 4435 5315
rect 4485 5285 4515 5315
rect 4645 5285 4675 5315
rect 4725 5285 4755 5315
rect 4885 5285 4915 5315
rect 5045 5285 5075 5315
rect 5205 5285 5235 5315
rect 5365 5285 5395 5315
rect 5525 5285 5555 5315
rect 5685 5285 5715 5315
rect 5765 5285 5795 5315
rect 5925 5285 5955 5315
rect 6005 5285 6035 5315
rect 6165 5285 6195 5315
rect 4245 5205 4275 5235
rect 4405 5205 4435 5235
rect 4485 5205 4515 5235
rect 4645 5205 4675 5235
rect 4725 5205 4755 5235
rect 4885 5205 4915 5235
rect 5045 5205 5075 5235
rect 5205 5205 5235 5235
rect 5365 5205 5395 5235
rect 5525 5205 5555 5235
rect 5685 5205 5715 5235
rect 5765 5205 5795 5235
rect 5925 5205 5955 5235
rect 6005 5205 6035 5235
rect 6165 5205 6195 5235
rect 4245 5125 4275 5155
rect 4405 5125 4435 5155
rect 4485 5125 4515 5155
rect 4645 5125 4675 5155
rect 4725 5125 4755 5155
rect 4885 5125 4915 5155
rect 5045 5125 5075 5155
rect 5205 5125 5235 5155
rect 5365 5125 5395 5155
rect 5525 5125 5555 5155
rect 5685 5125 5715 5155
rect 5765 5125 5795 5155
rect 5925 5125 5955 5155
rect 6005 5125 6035 5155
rect 6165 5125 6195 5155
rect 4245 5045 4275 5075
rect 4405 5045 4435 5075
rect 4485 5045 4515 5075
rect 4645 5045 4675 5075
rect 4725 5045 4755 5075
rect 4885 5045 4915 5075
rect 5045 5045 5075 5075
rect 5205 5045 5235 5075
rect 5365 5045 5395 5075
rect 5525 5045 5555 5075
rect 5685 5045 5715 5075
rect 5765 5045 5795 5075
rect 5925 5045 5955 5075
rect 6005 5045 6035 5075
rect 6165 5045 6195 5075
rect 4245 4965 4275 4995
rect 4405 4965 4435 4995
rect 4485 4965 4515 4995
rect 4645 4965 4675 4995
rect 4725 4965 4755 4995
rect 4885 4965 4915 4995
rect 5045 4965 5075 4995
rect 5205 4965 5235 4995
rect 5365 4965 5395 4995
rect 5525 4965 5555 4995
rect 5685 4965 5715 4995
rect 5765 4965 5795 4995
rect 5925 4965 5955 4995
rect 6005 4965 6035 4995
rect 6165 4965 6195 4995
rect 4245 4885 4275 4915
rect 4405 4885 4435 4915
rect 4485 4885 4515 4915
rect 4645 4885 4675 4915
rect 4725 4885 4755 4915
rect 4885 4885 4915 4915
rect 5045 4885 5075 4915
rect 5205 4885 5235 4915
rect 5365 4885 5395 4915
rect 5525 4885 5555 4915
rect 5685 4885 5715 4915
rect 5765 4885 5795 4915
rect 5925 4885 5955 4915
rect 6005 4885 6035 4915
rect 6165 4885 6195 4915
rect 5845 4805 5875 4835
rect 4245 4725 4275 4755
rect 4405 4725 4435 4755
rect 4485 4725 4515 4755
rect 4645 4725 4675 4755
rect 4725 4725 4755 4755
rect 4885 4725 4915 4755
rect 5045 4725 5075 4755
rect 5205 4725 5235 4755
rect 5365 4725 5395 4755
rect 5525 4725 5555 4755
rect 5685 4725 5715 4755
rect 5765 4725 5795 4755
rect 5925 4725 5955 4755
rect 6005 4725 6035 4755
rect 6165 4725 6195 4755
rect 4245 4645 4275 4675
rect 4405 4645 4435 4675
rect 4485 4645 4515 4675
rect 4645 4645 4675 4675
rect 4725 4645 4755 4675
rect 4885 4645 4915 4675
rect 5045 4645 5075 4675
rect 5205 4645 5235 4675
rect 5365 4645 5395 4675
rect 5525 4645 5555 4675
rect 5685 4645 5715 4675
rect 5765 4645 5795 4675
rect 5925 4645 5955 4675
rect 6005 4645 6035 4675
rect 6165 4645 6195 4675
rect 6085 4565 6115 4595
rect 4245 4485 4275 4515
rect 4405 4485 4435 4515
rect 4485 4485 4515 4515
rect 4645 4485 4675 4515
rect 4725 4485 4755 4515
rect 4885 4485 4915 4515
rect 5045 4485 5075 4515
rect 5205 4485 5235 4515
rect 5365 4485 5395 4515
rect 5525 4485 5555 4515
rect 5685 4485 5715 4515
rect 5765 4485 5795 4515
rect 5925 4485 5955 4515
rect 6005 4485 6035 4515
rect 6165 4485 6195 4515
rect 4245 4405 4275 4435
rect 4405 4405 4435 4435
rect 4485 4405 4515 4435
rect 4645 4405 4675 4435
rect 4725 4405 4755 4435
rect 4885 4405 4915 4435
rect 5045 4405 5075 4435
rect 5205 4405 5235 4435
rect 5365 4405 5395 4435
rect 5525 4405 5555 4435
rect 5685 4405 5715 4435
rect 5765 4405 5795 4435
rect 5925 4405 5955 4435
rect 6005 4405 6035 4435
rect 6165 4405 6195 4435
rect 4245 4325 4275 4355
rect 4405 4325 4435 4355
rect 4485 4325 4515 4355
rect 4645 4325 4675 4355
rect 4725 4325 4755 4355
rect 4885 4325 4915 4355
rect 5045 4325 5075 4355
rect 5205 4325 5235 4355
rect 5365 4325 5395 4355
rect 5525 4325 5555 4355
rect 5685 4325 5715 4355
rect 5765 4325 5795 4355
rect 5925 4325 5955 4355
rect 6005 4325 6035 4355
rect 6165 4325 6195 4355
rect 4245 4245 4275 4275
rect 4405 4245 4435 4275
rect 4485 4245 4515 4275
rect 4645 4245 4675 4275
rect 4725 4245 4755 4275
rect 4885 4245 4915 4275
rect 5045 4245 5075 4275
rect 5205 4245 5235 4275
rect 5365 4245 5395 4275
rect 5525 4245 5555 4275
rect 5685 4245 5715 4275
rect 5765 4245 5795 4275
rect 5925 4245 5955 4275
rect 6005 4245 6035 4275
rect 6165 4245 6195 4275
rect 4245 4165 4275 4195
rect 4405 4165 4435 4195
rect 4485 4165 4515 4195
rect 4645 4165 4675 4195
rect 4725 4165 4755 4195
rect 4885 4165 4915 4195
rect 5045 4165 5075 4195
rect 5205 4165 5235 4195
rect 5365 4165 5395 4195
rect 5525 4165 5555 4195
rect 5685 4165 5715 4195
rect 5765 4165 5795 4195
rect 5925 4165 5955 4195
rect 6005 4165 6035 4195
rect 6165 4165 6195 4195
rect 4245 4085 4275 4115
rect 4405 4085 4435 4115
rect 4485 4085 4515 4115
rect 4645 4085 4675 4115
rect 4725 4085 4755 4115
rect 4885 4085 4915 4115
rect 5045 4085 5075 4115
rect 5205 4085 5235 4115
rect 5365 4085 5395 4115
rect 5525 4085 5555 4115
rect 5685 4085 5715 4115
rect 5765 4085 5795 4115
rect 5925 4085 5955 4115
rect 6005 4085 6035 4115
rect 6165 4085 6195 4115
rect 4245 4005 4275 4035
rect 4405 4005 4435 4035
rect 4485 4005 4515 4035
rect 4645 4005 4675 4035
rect 4725 4005 4755 4035
rect 4885 4005 4915 4035
rect 5045 4005 5075 4035
rect 5205 4005 5235 4035
rect 5365 4005 5395 4035
rect 5525 4005 5555 4035
rect 5685 4005 5715 4035
rect 5765 4005 5795 4035
rect 5925 4005 5955 4035
rect 6005 4005 6035 4035
rect 6165 4005 6195 4035
rect 4245 3925 4275 3955
rect 4405 3925 4435 3955
rect 4485 3925 4515 3955
rect 4645 3925 4675 3955
rect 4725 3925 4755 3955
rect 4885 3925 4915 3955
rect 5045 3925 5075 3955
rect 5205 3925 5235 3955
rect 5365 3925 5395 3955
rect 5525 3925 5555 3955
rect 5685 3925 5715 3955
rect 5765 3925 5795 3955
rect 5925 3925 5955 3955
rect 6005 3925 6035 3955
rect 6165 3925 6195 3955
rect 4245 3845 4275 3875
rect 4405 3845 4435 3875
rect 4485 3845 4515 3875
rect 4645 3845 4675 3875
rect 4725 3845 4755 3875
rect 4885 3845 4915 3875
rect 5045 3845 5075 3875
rect 5205 3845 5235 3875
rect 5365 3845 5395 3875
rect 5525 3845 5555 3875
rect 5685 3845 5715 3875
rect 5765 3845 5795 3875
rect 5925 3845 5955 3875
rect 6005 3845 6035 3875
rect 6165 3845 6195 3875
rect 4325 3765 4355 3795
rect 4245 3685 4275 3715
rect 4405 3685 4435 3715
rect 4485 3685 4515 3715
rect 4645 3685 4675 3715
rect 4725 3685 4755 3715
rect 4885 3685 4915 3715
rect 5045 3685 5075 3715
rect 5205 3685 5235 3715
rect 5365 3685 5395 3715
rect 5525 3685 5555 3715
rect 5685 3685 5715 3715
rect 5765 3685 5795 3715
rect 5925 3685 5955 3715
rect 6005 3685 6035 3715
rect 6165 3685 6195 3715
rect 4245 3605 4275 3635
rect 4405 3605 4435 3635
rect 4485 3605 4515 3635
rect 4645 3605 4675 3635
rect 4725 3605 4755 3635
rect 4885 3605 4915 3635
rect 5045 3605 5075 3635
rect 5205 3605 5235 3635
rect 5365 3605 5395 3635
rect 5525 3605 5555 3635
rect 5685 3605 5715 3635
rect 5765 3605 5795 3635
rect 5925 3605 5955 3635
rect 6005 3605 6035 3635
rect 6165 3605 6195 3635
rect 4565 3525 4595 3555
rect 4245 3445 4275 3475
rect 4405 3445 4435 3475
rect 4485 3445 4515 3475
rect 4645 3445 4675 3475
rect 4725 3445 4755 3475
rect 4885 3445 4915 3475
rect 5045 3445 5075 3475
rect 5205 3445 5235 3475
rect 5365 3445 5395 3475
rect 5525 3445 5555 3475
rect 5685 3445 5715 3475
rect 5765 3445 5795 3475
rect 5925 3445 5955 3475
rect 6005 3445 6035 3475
rect 6165 3445 6195 3475
rect 4245 3365 4275 3395
rect 4405 3365 4435 3395
rect 4485 3365 4515 3395
rect 4645 3365 4675 3395
rect 4725 3365 4755 3395
rect 4885 3365 4915 3395
rect 5045 3365 5075 3395
rect 5205 3365 5235 3395
rect 5365 3365 5395 3395
rect 5525 3365 5555 3395
rect 5685 3365 5715 3395
rect 5765 3365 5795 3395
rect 5925 3365 5955 3395
rect 6005 3365 6035 3395
rect 6165 3365 6195 3395
rect 5845 3285 5875 3315
rect 4245 3205 4275 3235
rect 4405 3205 4435 3235
rect 4485 3205 4515 3235
rect 4645 3205 4675 3235
rect 4725 3205 4755 3235
rect 4885 3205 4915 3235
rect 5045 3205 5075 3235
rect 5205 3205 5235 3235
rect 5365 3205 5395 3235
rect 5525 3205 5555 3235
rect 5685 3205 5715 3235
rect 5765 3205 5795 3235
rect 5925 3205 5955 3235
rect 6005 3205 6035 3235
rect 6165 3205 6195 3235
rect 4245 3125 4275 3155
rect 4405 3125 4435 3155
rect 4485 3125 4515 3155
rect 4645 3125 4675 3155
rect 4725 3125 4755 3155
rect 4885 3125 4915 3155
rect 5045 3125 5075 3155
rect 5205 3125 5235 3155
rect 5365 3125 5395 3155
rect 5525 3125 5555 3155
rect 5685 3125 5715 3155
rect 5765 3125 5795 3155
rect 5925 3125 5955 3155
rect 6005 3125 6035 3155
rect 6165 3125 6195 3155
rect 4245 3045 4275 3075
rect 4405 3045 4435 3075
rect 4485 3045 4515 3075
rect 4645 3045 4675 3075
rect 4725 3045 4755 3075
rect 4885 3045 4915 3075
rect 5045 3045 5075 3075
rect 5205 3045 5235 3075
rect 5365 3045 5395 3075
rect 5525 3045 5555 3075
rect 5685 3045 5715 3075
rect 5765 3045 5795 3075
rect 5925 3045 5955 3075
rect 6005 3045 6035 3075
rect 6165 3045 6195 3075
rect 4245 2965 4275 2995
rect 4405 2965 4435 2995
rect 4485 2965 4515 2995
rect 4645 2965 4675 2995
rect 4725 2965 4755 2995
rect 4885 2965 4915 2995
rect 5045 2965 5075 2995
rect 5205 2965 5235 2995
rect 5365 2965 5395 2995
rect 5525 2965 5555 2995
rect 5685 2965 5715 2995
rect 5765 2965 5795 2995
rect 5925 2965 5955 2995
rect 6005 2965 6035 2995
rect 6165 2965 6195 2995
rect 4245 2885 4275 2915
rect 4405 2885 4435 2915
rect 4485 2885 4515 2915
rect 4645 2885 4675 2915
rect 4725 2885 4755 2915
rect 4885 2885 4915 2915
rect 5045 2885 5075 2915
rect 5205 2885 5235 2915
rect 5365 2885 5395 2915
rect 5525 2885 5555 2915
rect 5685 2885 5715 2915
rect 5765 2885 5795 2915
rect 5925 2885 5955 2915
rect 6005 2885 6035 2915
rect 6165 2885 6195 2915
rect 4245 2805 4275 2835
rect 4405 2805 4435 2835
rect 4485 2805 4515 2835
rect 4645 2805 4675 2835
rect 4725 2805 4755 2835
rect 4885 2805 4915 2835
rect 5045 2805 5075 2835
rect 5205 2805 5235 2835
rect 5365 2805 5395 2835
rect 5525 2805 5555 2835
rect 5685 2805 5715 2835
rect 5765 2805 5795 2835
rect 5925 2805 5955 2835
rect 6005 2805 6035 2835
rect 6165 2805 6195 2835
rect 4245 2725 4275 2755
rect 4405 2725 4435 2755
rect 4485 2725 4515 2755
rect 4645 2725 4675 2755
rect 4725 2725 4755 2755
rect 4885 2725 4915 2755
rect 5045 2725 5075 2755
rect 5205 2725 5235 2755
rect 5365 2725 5395 2755
rect 5525 2725 5555 2755
rect 5685 2725 5715 2755
rect 5765 2725 5795 2755
rect 5925 2725 5955 2755
rect 6005 2725 6035 2755
rect 6165 2725 6195 2755
rect 4245 2645 4275 2675
rect 4405 2645 4435 2675
rect 4485 2645 4515 2675
rect 4645 2645 4675 2675
rect 4725 2645 4755 2675
rect 4885 2645 4915 2675
rect 5045 2645 5075 2675
rect 5205 2645 5235 2675
rect 5365 2645 5395 2675
rect 5525 2645 5555 2675
rect 5685 2645 5715 2675
rect 5765 2645 5795 2675
rect 5925 2645 5955 2675
rect 6005 2645 6035 2675
rect 6165 2645 6195 2675
rect 4245 2565 4275 2595
rect 4405 2565 4435 2595
rect 4485 2565 4515 2595
rect 4645 2565 4675 2595
rect 4725 2565 4755 2595
rect 4885 2565 4915 2595
rect 5045 2565 5075 2595
rect 5205 2565 5235 2595
rect 5365 2565 5395 2595
rect 5525 2565 5555 2595
rect 5685 2565 5715 2595
rect 5765 2565 5795 2595
rect 5925 2565 5955 2595
rect 6005 2565 6035 2595
rect 6165 2565 6195 2595
rect 4245 2485 4275 2515
rect 4405 2485 4435 2515
rect 4485 2485 4515 2515
rect 4645 2485 4675 2515
rect 4725 2485 4755 2515
rect 4885 2485 4915 2515
rect 5045 2485 5075 2515
rect 5205 2485 5235 2515
rect 5365 2485 5395 2515
rect 5525 2485 5555 2515
rect 5685 2485 5715 2515
rect 5765 2485 5795 2515
rect 5925 2485 5955 2515
rect 6005 2485 6035 2515
rect 6165 2485 6195 2515
rect 4245 2405 4275 2435
rect 4405 2405 4435 2435
rect 4485 2405 4515 2435
rect 4645 2405 4675 2435
rect 4725 2405 4755 2435
rect 4885 2405 4915 2435
rect 5045 2405 5075 2435
rect 5205 2405 5235 2435
rect 5365 2405 5395 2435
rect 5525 2405 5555 2435
rect 5685 2405 5715 2435
rect 5765 2405 5795 2435
rect 5925 2405 5955 2435
rect 6005 2405 6035 2435
rect 6165 2405 6195 2435
rect 4245 2325 4275 2355
rect 4405 2325 4435 2355
rect 4485 2325 4515 2355
rect 4645 2325 4675 2355
rect 4725 2325 4755 2355
rect 4885 2325 4915 2355
rect 5045 2325 5075 2355
rect 5205 2325 5235 2355
rect 5365 2325 5395 2355
rect 5525 2325 5555 2355
rect 5685 2325 5715 2355
rect 5765 2325 5795 2355
rect 5925 2325 5955 2355
rect 6005 2325 6035 2355
rect 6165 2325 6195 2355
rect 4245 2245 4275 2275
rect 4405 2245 4435 2275
rect 4485 2245 4515 2275
rect 4645 2245 4675 2275
rect 4725 2245 4755 2275
rect 4885 2245 4915 2275
rect 5045 2245 5075 2275
rect 5205 2245 5235 2275
rect 5365 2245 5395 2275
rect 5525 2245 5555 2275
rect 5685 2245 5715 2275
rect 5765 2245 5795 2275
rect 5925 2245 5955 2275
rect 6005 2245 6035 2275
rect 6165 2245 6195 2275
rect 4245 2165 4275 2195
rect 4405 2165 4435 2195
rect 4485 2165 4515 2195
rect 4645 2165 4675 2195
rect 4725 2165 4755 2195
rect 4885 2165 4915 2195
rect 5045 2165 5075 2195
rect 5205 2165 5235 2195
rect 5365 2165 5395 2195
rect 5525 2165 5555 2195
rect 5685 2165 5715 2195
rect 5765 2165 5795 2195
rect 5925 2165 5955 2195
rect 6005 2165 6035 2195
rect 6165 2165 6195 2195
rect 4245 2085 4275 2115
rect 4405 2085 4435 2115
rect 4485 2085 4515 2115
rect 4645 2085 4675 2115
rect 4725 2085 4755 2115
rect 4885 2085 4915 2115
rect 5045 2085 5075 2115
rect 5205 2085 5235 2115
rect 5365 2085 5395 2115
rect 5525 2085 5555 2115
rect 5685 2085 5715 2115
rect 5765 2085 5795 2115
rect 5925 2085 5955 2115
rect 6005 2085 6035 2115
rect 6165 2085 6195 2115
rect 4245 2005 4275 2035
rect 4405 2005 4435 2035
rect 4485 2005 4515 2035
rect 4645 2005 4675 2035
rect 4725 2005 4755 2035
rect 4885 2005 4915 2035
rect 5045 2005 5075 2035
rect 5205 2005 5235 2035
rect 5365 2005 5395 2035
rect 5525 2005 5555 2035
rect 5685 2005 5715 2035
rect 5765 2005 5795 2035
rect 5925 2005 5955 2035
rect 6005 2005 6035 2035
rect 6165 2005 6195 2035
rect 4245 1925 4275 1955
rect 4405 1925 4435 1955
rect 4485 1925 4515 1955
rect 4645 1925 4675 1955
rect 4725 1925 4755 1955
rect 4885 1925 4915 1955
rect 5045 1925 5075 1955
rect 5205 1925 5235 1955
rect 5365 1925 5395 1955
rect 5525 1925 5555 1955
rect 5685 1925 5715 1955
rect 5765 1925 5795 1955
rect 5925 1925 5955 1955
rect 6005 1925 6035 1955
rect 6165 1925 6195 1955
rect 4565 1805 4595 1835
rect 4245 1685 4275 1715
rect 4405 1685 4435 1715
rect 4485 1685 4515 1715
rect 4645 1685 4675 1715
rect 4725 1685 4755 1715
rect 4885 1685 4915 1715
rect 5045 1685 5075 1715
rect 5205 1685 5235 1715
rect 5365 1685 5395 1715
rect 5525 1685 5555 1715
rect 5685 1685 5715 1715
rect 5765 1685 5795 1715
rect 5925 1685 5955 1715
rect 6005 1685 6035 1715
rect 6165 1685 6195 1715
rect 4245 1605 4275 1635
rect 4405 1605 4435 1635
rect 4485 1605 4515 1635
rect 4645 1605 4675 1635
rect 4725 1605 4755 1635
rect 4885 1605 4915 1635
rect 5045 1605 5075 1635
rect 5205 1605 5235 1635
rect 5365 1605 5395 1635
rect 5525 1605 5555 1635
rect 5685 1605 5715 1635
rect 5765 1605 5795 1635
rect 5925 1605 5955 1635
rect 6005 1605 6035 1635
rect 6165 1605 6195 1635
rect 4245 1525 4275 1555
rect 4405 1525 4435 1555
rect 4485 1525 4515 1555
rect 4645 1525 4675 1555
rect 4725 1525 4755 1555
rect 4885 1525 4915 1555
rect 5045 1525 5075 1555
rect 5205 1525 5235 1555
rect 5365 1525 5395 1555
rect 5525 1525 5555 1555
rect 5685 1525 5715 1555
rect 5765 1525 5795 1555
rect 5925 1525 5955 1555
rect 6005 1525 6035 1555
rect 6165 1525 6195 1555
rect 4245 1445 4275 1475
rect 4405 1445 4435 1475
rect 4485 1445 4515 1475
rect 4645 1445 4675 1475
rect 4725 1445 4755 1475
rect 4885 1445 4915 1475
rect 5045 1445 5075 1475
rect 5205 1445 5235 1475
rect 5365 1445 5395 1475
rect 5525 1445 5555 1475
rect 5685 1445 5715 1475
rect 5765 1445 5795 1475
rect 5925 1445 5955 1475
rect 6005 1445 6035 1475
rect 6165 1445 6195 1475
rect 4245 1365 4275 1395
rect 4405 1365 4435 1395
rect 4485 1365 4515 1395
rect 4645 1365 4675 1395
rect 4725 1365 4755 1395
rect 4885 1365 4915 1395
rect 5045 1365 5075 1395
rect 5205 1365 5235 1395
rect 5365 1365 5395 1395
rect 5525 1365 5555 1395
rect 5685 1365 5715 1395
rect 5765 1365 5795 1395
rect 5925 1365 5955 1395
rect 6005 1365 6035 1395
rect 6165 1365 6195 1395
rect 4245 1285 4275 1315
rect 4405 1285 4435 1315
rect 4485 1285 4515 1315
rect 4645 1285 4675 1315
rect 4725 1285 4755 1315
rect 4885 1285 4915 1315
rect 5045 1285 5075 1315
rect 5205 1285 5235 1315
rect 5365 1285 5395 1315
rect 5525 1285 5555 1315
rect 5685 1285 5715 1315
rect 5765 1285 5795 1315
rect 5925 1285 5955 1315
rect 6005 1285 6035 1315
rect 6165 1285 6195 1315
rect 4245 1205 4275 1235
rect 4405 1205 4435 1235
rect 4485 1205 4515 1235
rect 4645 1205 4675 1235
rect 4725 1205 4755 1235
rect 4885 1205 4915 1235
rect 5045 1205 5075 1235
rect 5205 1205 5235 1235
rect 5365 1205 5395 1235
rect 5525 1205 5555 1235
rect 5685 1205 5715 1235
rect 5765 1205 5795 1235
rect 5925 1205 5955 1235
rect 6005 1205 6035 1235
rect 6165 1205 6195 1235
rect 4245 1125 4275 1155
rect 4405 1125 4435 1155
rect 4485 1125 4515 1155
rect 4645 1125 4675 1155
rect 4725 1125 4755 1155
rect 4885 1125 4915 1155
rect 5045 1125 5075 1155
rect 5205 1125 5235 1155
rect 5365 1125 5395 1155
rect 5525 1125 5555 1155
rect 5685 1125 5715 1155
rect 5765 1125 5795 1155
rect 5925 1125 5955 1155
rect 6005 1125 6035 1155
rect 6165 1125 6195 1155
rect 4245 1045 4275 1075
rect 4405 1045 4435 1075
rect 4485 1045 4515 1075
rect 4645 1045 4675 1075
rect 4725 1045 4755 1075
rect 4885 1045 4915 1075
rect 5045 1045 5075 1075
rect 5205 1045 5235 1075
rect 5365 1045 5395 1075
rect 5525 1045 5555 1075
rect 5685 1045 5715 1075
rect 5765 1045 5795 1075
rect 5925 1045 5955 1075
rect 6005 1045 6035 1075
rect 6165 1045 6195 1075
rect 4245 965 4275 995
rect 4405 965 4435 995
rect 4485 965 4515 995
rect 4645 965 4675 995
rect 4725 965 4755 995
rect 4885 965 4915 995
rect 5045 965 5075 995
rect 5205 965 5235 995
rect 5365 965 5395 995
rect 5525 965 5555 995
rect 5685 965 5715 995
rect 5765 965 5795 995
rect 5925 965 5955 995
rect 6005 965 6035 995
rect 6165 965 6195 995
rect 6085 885 6115 915
rect 4245 805 4275 835
rect 4405 805 4435 835
rect 4485 805 4515 835
rect 4645 805 4675 835
rect 4725 805 4755 835
rect 4885 805 4915 835
rect 5045 805 5075 835
rect 5205 805 5235 835
rect 5365 805 5395 835
rect 5525 805 5555 835
rect 5685 805 5715 835
rect 5765 805 5795 835
rect 5925 805 5955 835
rect 6005 805 6035 835
rect 6165 805 6195 835
rect 4245 725 4275 755
rect 4405 725 4435 755
rect 4485 725 4515 755
rect 4645 725 4675 755
rect 4725 725 4755 755
rect 4885 725 4915 755
rect 5045 725 5075 755
rect 5205 725 5235 755
rect 5365 725 5395 755
rect 5525 725 5555 755
rect 5685 725 5715 755
rect 5765 725 5795 755
rect 5925 725 5955 755
rect 6005 725 6035 755
rect 6165 725 6195 755
rect 4245 645 4275 675
rect 4405 645 4435 675
rect 4485 645 4515 675
rect 4645 645 4675 675
rect 4725 645 4755 675
rect 4885 645 4915 675
rect 5045 645 5075 675
rect 5205 645 5235 675
rect 5365 645 5395 675
rect 5525 645 5555 675
rect 5685 645 5715 675
rect 5765 645 5795 675
rect 5925 645 5955 675
rect 6005 645 6035 675
rect 6165 645 6195 675
rect 4245 565 4275 595
rect 4405 565 4435 595
rect 4485 565 4515 595
rect 4645 565 4675 595
rect 4725 565 4755 595
rect 4885 565 4915 595
rect 5045 565 5075 595
rect 5205 565 5235 595
rect 5365 565 5395 595
rect 5525 565 5555 595
rect 5685 565 5715 595
rect 5765 565 5795 595
rect 5925 565 5955 595
rect 6005 565 6035 595
rect 6165 565 6195 595
rect 4245 485 4275 515
rect 4405 485 4435 515
rect 4485 485 4515 515
rect 4645 485 4675 515
rect 4725 485 4755 515
rect 4885 485 4915 515
rect 5045 485 5075 515
rect 5205 485 5235 515
rect 5365 485 5395 515
rect 5525 485 5555 515
rect 5685 485 5715 515
rect 5765 485 5795 515
rect 5925 485 5955 515
rect 6005 485 6035 515
rect 6165 485 6195 515
rect 4325 365 4355 395
rect 4245 245 4275 275
rect 4405 245 4435 275
rect 4485 245 4515 275
rect 4645 245 4675 275
rect 4725 245 4755 275
rect 4885 245 4915 275
rect 5045 245 5075 275
rect 5205 245 5235 275
rect 5365 245 5395 275
rect 5525 245 5555 275
rect 5685 245 5715 275
rect 5765 245 5795 275
rect 5925 245 5955 275
rect 6005 245 6035 275
rect 6165 245 6195 275
rect 4245 165 4275 195
rect 4405 165 4435 195
rect 4485 165 4515 195
rect 4645 165 4675 195
rect 4725 165 4755 195
rect 4885 165 4915 195
rect 5045 165 5075 195
rect 5205 165 5235 195
rect 5365 165 5395 195
rect 5525 165 5555 195
rect 5685 165 5715 195
rect 5765 165 5795 195
rect 5925 165 5955 195
rect 6005 165 6035 195
rect 6165 165 6195 195
rect 4245 85 4275 115
rect 4405 85 4435 115
rect 4485 85 4515 115
rect 4645 85 4675 115
rect 4725 85 4755 115
rect 4885 85 4915 115
rect 5045 85 5075 115
rect 5205 85 5235 115
rect 5365 85 5395 115
rect 5525 85 5555 115
rect 5685 85 5715 115
rect 5765 85 5795 115
rect 5925 85 5955 115
rect 6005 85 6035 115
rect 6165 85 6195 115
rect 4245 5 4275 35
rect 4405 5 4435 35
rect 4485 5 4515 35
rect 4645 5 4675 35
rect 4725 5 4755 35
rect 4885 5 4915 35
rect 5045 5 5075 35
rect 5205 5 5235 35
rect 5365 5 5395 35
rect 5525 5 5555 35
rect 5685 5 5715 35
rect 5765 5 5795 35
rect 5925 5 5955 35
rect 6005 5 6035 35
rect 6165 5 6195 35
<< metal3 >>
rect 4240 15716 4280 15760
rect 4240 15684 4244 15716
rect 4276 15684 4280 15716
rect 4240 15636 4280 15684
rect 4240 15604 4244 15636
rect 4276 15604 4280 15636
rect 4240 15556 4280 15604
rect 4240 15524 4244 15556
rect 4276 15524 4280 15556
rect 4240 15476 4280 15524
rect 4240 15444 4244 15476
rect 4276 15444 4280 15476
rect 4240 15396 4280 15444
rect 4240 15364 4244 15396
rect 4276 15364 4280 15396
rect 4240 15316 4280 15364
rect 4240 15284 4244 15316
rect 4276 15284 4280 15316
rect 4240 15236 4280 15284
rect 4240 15204 4244 15236
rect 4276 15204 4280 15236
rect 4240 15156 4280 15204
rect 4240 15124 4244 15156
rect 4276 15124 4280 15156
rect 4240 15076 4280 15124
rect 4240 15044 4244 15076
rect 4276 15044 4280 15076
rect 4240 14996 4280 15044
rect 4240 14964 4244 14996
rect 4276 14964 4280 14996
rect 4240 14916 4280 14964
rect 4240 14884 4244 14916
rect 4276 14884 4280 14916
rect 4240 14836 4280 14884
rect 4240 14804 4244 14836
rect 4276 14804 4280 14836
rect 4240 14756 4280 14804
rect 4240 14724 4244 14756
rect 4276 14724 4280 14756
rect 4240 14676 4280 14724
rect 4240 14644 4244 14676
rect 4276 14644 4280 14676
rect 4240 14596 4280 14644
rect 4240 14564 4244 14596
rect 4276 14564 4280 14596
rect 4240 14516 4280 14564
rect 4240 14484 4244 14516
rect 4276 14484 4280 14516
rect 4240 14436 4280 14484
rect 4240 14404 4244 14436
rect 4276 14404 4280 14436
rect 4240 14356 4280 14404
rect 4240 14324 4244 14356
rect 4276 14324 4280 14356
rect 4240 14276 4280 14324
rect 4240 14244 4244 14276
rect 4276 14244 4280 14276
rect 4240 14196 4280 14244
rect 4240 14164 4244 14196
rect 4276 14164 4280 14196
rect 4240 14116 4280 14164
rect 4240 14084 4244 14116
rect 4276 14084 4280 14116
rect 4240 14036 4280 14084
rect 4240 14004 4244 14036
rect 4276 14004 4280 14036
rect 4240 13956 4280 14004
rect 4240 13924 4244 13956
rect 4276 13924 4280 13956
rect 4240 13876 4280 13924
rect 4240 13844 4244 13876
rect 4276 13844 4280 13876
rect 4240 13796 4280 13844
rect 4240 13764 4244 13796
rect 4276 13764 4280 13796
rect 4240 13716 4280 13764
rect 4240 13684 4244 13716
rect 4276 13684 4280 13716
rect 4240 13636 4280 13684
rect 4240 13604 4244 13636
rect 4276 13604 4280 13636
rect 4240 13556 4280 13604
rect 4240 13524 4244 13556
rect 4276 13524 4280 13556
rect 4240 13476 4280 13524
rect 4240 13444 4244 13476
rect 4276 13444 4280 13476
rect 4240 13396 4280 13444
rect 4240 13364 4244 13396
rect 4276 13364 4280 13396
rect 4240 13316 4280 13364
rect 4240 13284 4244 13316
rect 4276 13284 4280 13316
rect 4240 13236 4280 13284
rect 4240 13204 4244 13236
rect 4276 13204 4280 13236
rect 4240 13156 4280 13204
rect 4240 13124 4244 13156
rect 4276 13124 4280 13156
rect 4240 13076 4280 13124
rect 4240 13044 4244 13076
rect 4276 13044 4280 13076
rect 4240 12996 4280 13044
rect 4240 12964 4244 12996
rect 4276 12964 4280 12996
rect 4240 12916 4280 12964
rect 4240 12884 4244 12916
rect 4276 12884 4280 12916
rect 4240 12836 4280 12884
rect 4240 12804 4244 12836
rect 4276 12804 4280 12836
rect 4240 12756 4280 12804
rect 4240 12724 4244 12756
rect 4276 12724 4280 12756
rect 4240 12676 4280 12724
rect 4240 12644 4244 12676
rect 4276 12644 4280 12676
rect 4240 12596 4280 12644
rect 4240 12564 4244 12596
rect 4276 12564 4280 12596
rect 4240 12516 4280 12564
rect 4240 12484 4244 12516
rect 4276 12484 4280 12516
rect 4240 12436 4280 12484
rect 4240 12404 4244 12436
rect 4276 12404 4280 12436
rect 4240 12356 4280 12404
rect 4240 12324 4244 12356
rect 4276 12324 4280 12356
rect 4240 12276 4280 12324
rect 4240 12244 4244 12276
rect 4276 12244 4280 12276
rect 4240 12196 4280 12244
rect 4240 12164 4244 12196
rect 4276 12164 4280 12196
rect 4240 12116 4280 12164
rect 4240 12084 4244 12116
rect 4276 12084 4280 12116
rect 4240 12036 4280 12084
rect 4240 12004 4244 12036
rect 4276 12004 4280 12036
rect 4240 11956 4280 12004
rect 4240 11924 4244 11956
rect 4276 11924 4280 11956
rect 4240 11876 4280 11924
rect 4240 11844 4244 11876
rect 4276 11844 4280 11876
rect 4240 11796 4280 11844
rect 4240 11764 4244 11796
rect 4276 11764 4280 11796
rect 4240 11716 4280 11764
rect 4240 11684 4244 11716
rect 4276 11684 4280 11716
rect 4240 11636 4280 11684
rect 4240 11604 4244 11636
rect 4276 11604 4280 11636
rect 4240 11556 4280 11604
rect 4240 11524 4244 11556
rect 4276 11524 4280 11556
rect 4240 11476 4280 11524
rect 4240 11444 4244 11476
rect 4276 11444 4280 11476
rect 4240 11396 4280 11444
rect 4240 11364 4244 11396
rect 4276 11364 4280 11396
rect 4240 11316 4280 11364
rect 4240 11284 4244 11316
rect 4276 11284 4280 11316
rect 4240 11236 4280 11284
rect 4240 11204 4244 11236
rect 4276 11204 4280 11236
rect 4240 11156 4280 11204
rect 4240 11124 4244 11156
rect 4276 11124 4280 11156
rect 4240 11076 4280 11124
rect 4240 11044 4244 11076
rect 4276 11044 4280 11076
rect 4240 10996 4280 11044
rect 4240 10964 4244 10996
rect 4276 10964 4280 10996
rect 4240 10916 4280 10964
rect 4240 10884 4244 10916
rect 4276 10884 4280 10916
rect 4240 10836 4280 10884
rect 4240 10804 4244 10836
rect 4276 10804 4280 10836
rect 4240 10756 4280 10804
rect 4240 10724 4244 10756
rect 4276 10724 4280 10756
rect 4240 10676 4280 10724
rect 4240 10644 4244 10676
rect 4276 10644 4280 10676
rect 4240 10596 4280 10644
rect 4240 10564 4244 10596
rect 4276 10564 4280 10596
rect 4240 10516 4280 10564
rect 4240 10484 4244 10516
rect 4276 10484 4280 10516
rect 4240 10436 4280 10484
rect 4240 10404 4244 10436
rect 4276 10404 4280 10436
rect 4240 10356 4280 10404
rect 4240 10324 4244 10356
rect 4276 10324 4280 10356
rect 4240 10276 4280 10324
rect 4240 10244 4244 10276
rect 4276 10244 4280 10276
rect 4240 10196 4280 10244
rect 4240 10164 4244 10196
rect 4276 10164 4280 10196
rect 4240 10116 4280 10164
rect 4240 10084 4244 10116
rect 4276 10084 4280 10116
rect 4240 10036 4280 10084
rect 4240 10004 4244 10036
rect 4276 10004 4280 10036
rect 4240 9956 4280 10004
rect 4240 9924 4244 9956
rect 4276 9924 4280 9956
rect 4240 9876 4280 9924
rect 4240 9844 4244 9876
rect 4276 9844 4280 9876
rect 4240 9796 4280 9844
rect 4240 9764 4244 9796
rect 4276 9764 4280 9796
rect 4240 9716 4280 9764
rect 4240 9684 4244 9716
rect 4276 9684 4280 9716
rect 4240 9636 4280 9684
rect 4240 9604 4244 9636
rect 4276 9604 4280 9636
rect 4240 9556 4280 9604
rect 4240 9524 4244 9556
rect 4276 9524 4280 9556
rect 4240 9476 4280 9524
rect 4240 9444 4244 9476
rect 4276 9444 4280 9476
rect 4240 9396 4280 9444
rect 4240 9364 4244 9396
rect 4276 9364 4280 9396
rect 4240 9316 4280 9364
rect 4240 9284 4244 9316
rect 4276 9284 4280 9316
rect 4240 9236 4280 9284
rect 4240 9204 4244 9236
rect 4276 9204 4280 9236
rect 4240 9156 4280 9204
rect 4240 9124 4244 9156
rect 4276 9124 4280 9156
rect 4240 9076 4280 9124
rect 4240 9044 4244 9076
rect 4276 9044 4280 9076
rect 4240 8996 4280 9044
rect 4240 8964 4244 8996
rect 4276 8964 4280 8996
rect 4240 8916 4280 8964
rect 4240 8884 4244 8916
rect 4276 8884 4280 8916
rect 4240 8836 4280 8884
rect 4240 8804 4244 8836
rect 4276 8804 4280 8836
rect 4240 8756 4280 8804
rect 4240 8724 4244 8756
rect 4276 8724 4280 8756
rect 4240 8676 4280 8724
rect 4240 8644 4244 8676
rect 4276 8644 4280 8676
rect 4240 8596 4280 8644
rect 4240 8564 4244 8596
rect 4276 8564 4280 8596
rect 4240 8516 4280 8564
rect 4240 8484 4244 8516
rect 4276 8484 4280 8516
rect 4240 8436 4280 8484
rect 4240 8404 4244 8436
rect 4276 8404 4280 8436
rect 4240 8356 4280 8404
rect 4240 8324 4244 8356
rect 4276 8324 4280 8356
rect 4240 8276 4280 8324
rect 4240 8244 4244 8276
rect 4276 8244 4280 8276
rect 4240 8196 4280 8244
rect 4240 8164 4244 8196
rect 4276 8164 4280 8196
rect 4240 8116 4280 8164
rect 4240 8084 4244 8116
rect 4276 8084 4280 8116
rect 4240 8036 4280 8084
rect 4240 8004 4244 8036
rect 4276 8004 4280 8036
rect 4240 7956 4280 8004
rect 4240 7924 4244 7956
rect 4276 7924 4280 7956
rect 4240 7876 4280 7924
rect 4240 7844 4244 7876
rect 4276 7844 4280 7876
rect 4240 7796 4280 7844
rect 4240 7764 4244 7796
rect 4276 7764 4280 7796
rect 4240 7716 4280 7764
rect 4240 7684 4244 7716
rect 4276 7684 4280 7716
rect 4240 7636 4280 7684
rect 4240 7604 4244 7636
rect 4276 7604 4280 7636
rect 4240 7556 4280 7604
rect 4240 7524 4244 7556
rect 4276 7524 4280 7556
rect 4240 7476 4280 7524
rect 4240 7444 4244 7476
rect 4276 7444 4280 7476
rect 4240 7396 4280 7444
rect 4240 7364 4244 7396
rect 4276 7364 4280 7396
rect 4240 7316 4280 7364
rect 4240 7284 4244 7316
rect 4276 7284 4280 7316
rect 4240 7236 4280 7284
rect 4240 7204 4244 7236
rect 4276 7204 4280 7236
rect 4240 7156 4280 7204
rect 4240 7124 4244 7156
rect 4276 7124 4280 7156
rect 4240 7076 4280 7124
rect 4240 7044 4244 7076
rect 4276 7044 4280 7076
rect 4240 6996 4280 7044
rect 4240 6964 4244 6996
rect 4276 6964 4280 6996
rect 4240 6916 4280 6964
rect 4240 6884 4244 6916
rect 4276 6884 4280 6916
rect 4240 6836 4280 6884
rect 4240 6804 4244 6836
rect 4276 6804 4280 6836
rect 4240 6756 4280 6804
rect 4240 6724 4244 6756
rect 4276 6724 4280 6756
rect 4240 6676 4280 6724
rect 4240 6644 4244 6676
rect 4276 6644 4280 6676
rect 4240 6596 4280 6644
rect 4240 6564 4244 6596
rect 4276 6564 4280 6596
rect 4240 6516 4280 6564
rect 4240 6484 4244 6516
rect 4276 6484 4280 6516
rect 4240 6436 4280 6484
rect 4240 6404 4244 6436
rect 4276 6404 4280 6436
rect 4240 6356 4280 6404
rect 4240 6324 4244 6356
rect 4276 6324 4280 6356
rect 4240 6276 4280 6324
rect 4240 6244 4244 6276
rect 4276 6244 4280 6276
rect 4240 6196 4280 6244
rect 4240 6164 4244 6196
rect 4276 6164 4280 6196
rect 4240 6116 4280 6164
rect 4240 6084 4244 6116
rect 4276 6084 4280 6116
rect 4240 6036 4280 6084
rect 4240 6004 4244 6036
rect 4276 6004 4280 6036
rect 4240 5956 4280 6004
rect 4240 5924 4244 5956
rect 4276 5924 4280 5956
rect 4240 5876 4280 5924
rect 4240 5844 4244 5876
rect 4276 5844 4280 5876
rect 4240 5796 4280 5844
rect 4240 5764 4244 5796
rect 4276 5764 4280 5796
rect 4240 5716 4280 5764
rect 4240 5684 4244 5716
rect 4276 5684 4280 5716
rect 4240 5636 4280 5684
rect 4240 5604 4244 5636
rect 4276 5604 4280 5636
rect 4240 5556 4280 5604
rect 4240 5524 4244 5556
rect 4276 5524 4280 5556
rect 4240 5476 4280 5524
rect 4240 5444 4244 5476
rect 4276 5444 4280 5476
rect 4240 5396 4280 5444
rect 4240 5364 4244 5396
rect 4276 5364 4280 5396
rect 4240 5316 4280 5364
rect 4240 5284 4244 5316
rect 4276 5284 4280 5316
rect 4240 5236 4280 5284
rect 4240 5204 4244 5236
rect 4276 5204 4280 5236
rect 4240 5156 4280 5204
rect 4240 5124 4244 5156
rect 4276 5124 4280 5156
rect 4240 5076 4280 5124
rect 4240 5044 4244 5076
rect 4276 5044 4280 5076
rect 4240 4996 4280 5044
rect 4240 4964 4244 4996
rect 4276 4964 4280 4996
rect 4240 4916 4280 4964
rect 4240 4884 4244 4916
rect 4276 4884 4280 4916
rect 4240 4836 4280 4884
rect 4240 4804 4244 4836
rect 4276 4804 4280 4836
rect 4240 4756 4280 4804
rect 4240 4724 4244 4756
rect 4276 4724 4280 4756
rect 4240 4676 4280 4724
rect 4240 4644 4244 4676
rect 4276 4644 4280 4676
rect 4240 4596 4280 4644
rect 4240 4564 4244 4596
rect 4276 4564 4280 4596
rect 4240 4516 4280 4564
rect 4240 4484 4244 4516
rect 4276 4484 4280 4516
rect 4240 4436 4280 4484
rect 4240 4404 4244 4436
rect 4276 4404 4280 4436
rect 4240 4356 4280 4404
rect 4240 4324 4244 4356
rect 4276 4324 4280 4356
rect 4240 4276 4280 4324
rect 4240 4244 4244 4276
rect 4276 4244 4280 4276
rect 4240 4196 4280 4244
rect 4240 4164 4244 4196
rect 4276 4164 4280 4196
rect 4240 4116 4280 4164
rect 4240 4084 4244 4116
rect 4276 4084 4280 4116
rect 4240 4036 4280 4084
rect 4240 4004 4244 4036
rect 4276 4004 4280 4036
rect 4240 3956 4280 4004
rect 4240 3924 4244 3956
rect 4276 3924 4280 3956
rect 4240 3876 4280 3924
rect 4240 3844 4244 3876
rect 4276 3844 4280 3876
rect 4240 3796 4280 3844
rect 4240 3764 4244 3796
rect 4276 3764 4280 3796
rect 4240 3716 4280 3764
rect 4240 3684 4244 3716
rect 4276 3684 4280 3716
rect 4240 3636 4280 3684
rect 4240 3604 4244 3636
rect 4276 3604 4280 3636
rect 4240 3556 4280 3604
rect 4240 3524 4244 3556
rect 4276 3524 4280 3556
rect 4240 3476 4280 3524
rect 4240 3444 4244 3476
rect 4276 3444 4280 3476
rect 4240 3396 4280 3444
rect 4240 3364 4244 3396
rect 4276 3364 4280 3396
rect 4240 3316 4280 3364
rect 4240 3284 4244 3316
rect 4276 3284 4280 3316
rect 4240 3236 4280 3284
rect 4240 3204 4244 3236
rect 4276 3204 4280 3236
rect 4240 3156 4280 3204
rect 4240 3124 4244 3156
rect 4276 3124 4280 3156
rect 4240 3076 4280 3124
rect 4240 3044 4244 3076
rect 4276 3044 4280 3076
rect 4240 2996 4280 3044
rect 4240 2964 4244 2996
rect 4276 2964 4280 2996
rect 4240 2916 4280 2964
rect 4240 2884 4244 2916
rect 4276 2884 4280 2916
rect 4240 2836 4280 2884
rect 4240 2804 4244 2836
rect 4276 2804 4280 2836
rect 4240 2756 4280 2804
rect 4240 2724 4244 2756
rect 4276 2724 4280 2756
rect 4240 2676 4280 2724
rect 4240 2644 4244 2676
rect 4276 2644 4280 2676
rect 4240 2596 4280 2644
rect 4240 2564 4244 2596
rect 4276 2564 4280 2596
rect 4240 2516 4280 2564
rect 4240 2484 4244 2516
rect 4276 2484 4280 2516
rect 4240 2436 4280 2484
rect 4240 2404 4244 2436
rect 4276 2404 4280 2436
rect 4240 2356 4280 2404
rect 4240 2324 4244 2356
rect 4276 2324 4280 2356
rect 4240 2276 4280 2324
rect 4240 2244 4244 2276
rect 4276 2244 4280 2276
rect 4240 2196 4280 2244
rect 4240 2164 4244 2196
rect 4276 2164 4280 2196
rect 4240 2116 4280 2164
rect 4240 2084 4244 2116
rect 4276 2084 4280 2116
rect 4240 2036 4280 2084
rect 4240 2004 4244 2036
rect 4276 2004 4280 2036
rect 4240 1956 4280 2004
rect 4240 1924 4244 1956
rect 4276 1924 4280 1956
rect 4240 1876 4280 1924
rect 4240 1844 4244 1876
rect 4276 1844 4280 1876
rect 4240 1796 4280 1844
rect 4240 1764 4244 1796
rect 4276 1764 4280 1796
rect 4240 1716 4280 1764
rect 4240 1684 4244 1716
rect 4276 1684 4280 1716
rect 4240 1636 4280 1684
rect 4240 1604 4244 1636
rect 4276 1604 4280 1636
rect 4240 1556 4280 1604
rect 4240 1524 4244 1556
rect 4276 1524 4280 1556
rect 4240 1476 4280 1524
rect 4240 1444 4244 1476
rect 4276 1444 4280 1476
rect 4240 1396 4280 1444
rect 4240 1364 4244 1396
rect 4276 1364 4280 1396
rect 4240 1316 4280 1364
rect 4240 1284 4244 1316
rect 4276 1284 4280 1316
rect 4240 1236 4280 1284
rect 4240 1204 4244 1236
rect 4276 1204 4280 1236
rect 4240 1156 4280 1204
rect 4240 1124 4244 1156
rect 4276 1124 4280 1156
rect 4240 1076 4280 1124
rect 4240 1044 4244 1076
rect 4276 1044 4280 1076
rect 4240 996 4280 1044
rect 4240 964 4244 996
rect 4276 964 4280 996
rect 4240 916 4280 964
rect 4240 884 4244 916
rect 4276 884 4280 916
rect 4240 836 4280 884
rect 4240 804 4244 836
rect 4276 804 4280 836
rect 4240 756 4280 804
rect 4240 724 4244 756
rect 4276 724 4280 756
rect 4240 676 4280 724
rect 4240 644 4244 676
rect 4276 644 4280 676
rect 4240 596 4280 644
rect 4240 564 4244 596
rect 4276 564 4280 596
rect 4240 516 4280 564
rect 4240 484 4244 516
rect 4276 484 4280 516
rect 4240 436 4280 484
rect 4240 404 4244 436
rect 4276 404 4280 436
rect 4240 356 4280 404
rect 4240 324 4244 356
rect 4276 324 4280 356
rect 4240 276 4280 324
rect 4240 244 4244 276
rect 4276 244 4280 276
rect 4240 196 4280 244
rect 4240 164 4244 196
rect 4276 164 4280 196
rect 4240 116 4280 164
rect 4240 84 4244 116
rect 4276 84 4280 116
rect 4240 36 4280 84
rect 4240 4 4244 36
rect 4276 4 4280 36
rect 4240 -764 4280 4
rect 4320 3795 4360 15760
rect 4320 3765 4325 3795
rect 4355 3765 4360 3795
rect 4320 395 4360 3765
rect 4320 365 4325 395
rect 4355 365 4360 395
rect 4320 0 4360 365
rect 4400 15716 4440 15760
rect 4400 15684 4404 15716
rect 4436 15684 4440 15716
rect 4400 15636 4440 15684
rect 4400 15604 4404 15636
rect 4436 15604 4440 15636
rect 4400 15556 4440 15604
rect 4400 15524 4404 15556
rect 4436 15524 4440 15556
rect 4400 15476 4440 15524
rect 4400 15444 4404 15476
rect 4436 15444 4440 15476
rect 4400 15396 4440 15444
rect 4400 15364 4404 15396
rect 4436 15364 4440 15396
rect 4400 15316 4440 15364
rect 4400 15284 4404 15316
rect 4436 15284 4440 15316
rect 4400 15236 4440 15284
rect 4400 15204 4404 15236
rect 4436 15204 4440 15236
rect 4400 15156 4440 15204
rect 4400 15124 4404 15156
rect 4436 15124 4440 15156
rect 4400 15076 4440 15124
rect 4400 15044 4404 15076
rect 4436 15044 4440 15076
rect 4400 14996 4440 15044
rect 4400 14964 4404 14996
rect 4436 14964 4440 14996
rect 4400 14916 4440 14964
rect 4400 14884 4404 14916
rect 4436 14884 4440 14916
rect 4400 14836 4440 14884
rect 4400 14804 4404 14836
rect 4436 14804 4440 14836
rect 4400 14756 4440 14804
rect 4400 14724 4404 14756
rect 4436 14724 4440 14756
rect 4400 14676 4440 14724
rect 4400 14644 4404 14676
rect 4436 14644 4440 14676
rect 4400 14596 4440 14644
rect 4400 14564 4404 14596
rect 4436 14564 4440 14596
rect 4400 14516 4440 14564
rect 4400 14484 4404 14516
rect 4436 14484 4440 14516
rect 4400 14436 4440 14484
rect 4400 14404 4404 14436
rect 4436 14404 4440 14436
rect 4400 14356 4440 14404
rect 4400 14324 4404 14356
rect 4436 14324 4440 14356
rect 4400 14276 4440 14324
rect 4400 14244 4404 14276
rect 4436 14244 4440 14276
rect 4400 14196 4440 14244
rect 4400 14164 4404 14196
rect 4436 14164 4440 14196
rect 4400 14116 4440 14164
rect 4400 14084 4404 14116
rect 4436 14084 4440 14116
rect 4400 14036 4440 14084
rect 4400 14004 4404 14036
rect 4436 14004 4440 14036
rect 4400 13956 4440 14004
rect 4400 13924 4404 13956
rect 4436 13924 4440 13956
rect 4400 13876 4440 13924
rect 4400 13844 4404 13876
rect 4436 13844 4440 13876
rect 4400 13796 4440 13844
rect 4400 13764 4404 13796
rect 4436 13764 4440 13796
rect 4400 13716 4440 13764
rect 4400 13684 4404 13716
rect 4436 13684 4440 13716
rect 4400 13636 4440 13684
rect 4400 13604 4404 13636
rect 4436 13604 4440 13636
rect 4400 13556 4440 13604
rect 4400 13524 4404 13556
rect 4436 13524 4440 13556
rect 4400 13476 4440 13524
rect 4400 13444 4404 13476
rect 4436 13444 4440 13476
rect 4400 13396 4440 13444
rect 4400 13364 4404 13396
rect 4436 13364 4440 13396
rect 4400 13316 4440 13364
rect 4400 13284 4404 13316
rect 4436 13284 4440 13316
rect 4400 13236 4440 13284
rect 4400 13204 4404 13236
rect 4436 13204 4440 13236
rect 4400 13156 4440 13204
rect 4400 13124 4404 13156
rect 4436 13124 4440 13156
rect 4400 13076 4440 13124
rect 4400 13044 4404 13076
rect 4436 13044 4440 13076
rect 4400 12996 4440 13044
rect 4400 12964 4404 12996
rect 4436 12964 4440 12996
rect 4400 12916 4440 12964
rect 4400 12884 4404 12916
rect 4436 12884 4440 12916
rect 4400 12836 4440 12884
rect 4400 12804 4404 12836
rect 4436 12804 4440 12836
rect 4400 12756 4440 12804
rect 4400 12724 4404 12756
rect 4436 12724 4440 12756
rect 4400 12676 4440 12724
rect 4400 12644 4404 12676
rect 4436 12644 4440 12676
rect 4400 12596 4440 12644
rect 4400 12564 4404 12596
rect 4436 12564 4440 12596
rect 4400 12516 4440 12564
rect 4400 12484 4404 12516
rect 4436 12484 4440 12516
rect 4400 12436 4440 12484
rect 4400 12404 4404 12436
rect 4436 12404 4440 12436
rect 4400 12356 4440 12404
rect 4400 12324 4404 12356
rect 4436 12324 4440 12356
rect 4400 12276 4440 12324
rect 4400 12244 4404 12276
rect 4436 12244 4440 12276
rect 4400 12196 4440 12244
rect 4400 12164 4404 12196
rect 4436 12164 4440 12196
rect 4400 12116 4440 12164
rect 4400 12084 4404 12116
rect 4436 12084 4440 12116
rect 4400 12036 4440 12084
rect 4400 12004 4404 12036
rect 4436 12004 4440 12036
rect 4400 11956 4440 12004
rect 4400 11924 4404 11956
rect 4436 11924 4440 11956
rect 4400 11876 4440 11924
rect 4400 11844 4404 11876
rect 4436 11844 4440 11876
rect 4400 11796 4440 11844
rect 4400 11764 4404 11796
rect 4436 11764 4440 11796
rect 4400 11716 4440 11764
rect 4400 11684 4404 11716
rect 4436 11684 4440 11716
rect 4400 11636 4440 11684
rect 4400 11604 4404 11636
rect 4436 11604 4440 11636
rect 4400 11556 4440 11604
rect 4400 11524 4404 11556
rect 4436 11524 4440 11556
rect 4400 11476 4440 11524
rect 4400 11444 4404 11476
rect 4436 11444 4440 11476
rect 4400 11396 4440 11444
rect 4400 11364 4404 11396
rect 4436 11364 4440 11396
rect 4400 11316 4440 11364
rect 4400 11284 4404 11316
rect 4436 11284 4440 11316
rect 4400 11236 4440 11284
rect 4400 11204 4404 11236
rect 4436 11204 4440 11236
rect 4400 11156 4440 11204
rect 4400 11124 4404 11156
rect 4436 11124 4440 11156
rect 4400 11076 4440 11124
rect 4400 11044 4404 11076
rect 4436 11044 4440 11076
rect 4400 10996 4440 11044
rect 4400 10964 4404 10996
rect 4436 10964 4440 10996
rect 4400 10916 4440 10964
rect 4400 10884 4404 10916
rect 4436 10884 4440 10916
rect 4400 10836 4440 10884
rect 4400 10804 4404 10836
rect 4436 10804 4440 10836
rect 4400 10756 4440 10804
rect 4400 10724 4404 10756
rect 4436 10724 4440 10756
rect 4400 10676 4440 10724
rect 4400 10644 4404 10676
rect 4436 10644 4440 10676
rect 4400 10596 4440 10644
rect 4400 10564 4404 10596
rect 4436 10564 4440 10596
rect 4400 10516 4440 10564
rect 4400 10484 4404 10516
rect 4436 10484 4440 10516
rect 4400 10436 4440 10484
rect 4400 10404 4404 10436
rect 4436 10404 4440 10436
rect 4400 10356 4440 10404
rect 4400 10324 4404 10356
rect 4436 10324 4440 10356
rect 4400 10276 4440 10324
rect 4400 10244 4404 10276
rect 4436 10244 4440 10276
rect 4400 10196 4440 10244
rect 4400 10164 4404 10196
rect 4436 10164 4440 10196
rect 4400 10116 4440 10164
rect 4400 10084 4404 10116
rect 4436 10084 4440 10116
rect 4400 10036 4440 10084
rect 4400 10004 4404 10036
rect 4436 10004 4440 10036
rect 4400 9956 4440 10004
rect 4400 9924 4404 9956
rect 4436 9924 4440 9956
rect 4400 9876 4440 9924
rect 4400 9844 4404 9876
rect 4436 9844 4440 9876
rect 4400 9796 4440 9844
rect 4400 9764 4404 9796
rect 4436 9764 4440 9796
rect 4400 9716 4440 9764
rect 4400 9684 4404 9716
rect 4436 9684 4440 9716
rect 4400 9636 4440 9684
rect 4400 9604 4404 9636
rect 4436 9604 4440 9636
rect 4400 9556 4440 9604
rect 4400 9524 4404 9556
rect 4436 9524 4440 9556
rect 4400 9476 4440 9524
rect 4400 9444 4404 9476
rect 4436 9444 4440 9476
rect 4400 9396 4440 9444
rect 4400 9364 4404 9396
rect 4436 9364 4440 9396
rect 4400 9316 4440 9364
rect 4400 9284 4404 9316
rect 4436 9284 4440 9316
rect 4400 9236 4440 9284
rect 4400 9204 4404 9236
rect 4436 9204 4440 9236
rect 4400 9156 4440 9204
rect 4400 9124 4404 9156
rect 4436 9124 4440 9156
rect 4400 9076 4440 9124
rect 4400 9044 4404 9076
rect 4436 9044 4440 9076
rect 4400 8996 4440 9044
rect 4400 8964 4404 8996
rect 4436 8964 4440 8996
rect 4400 8916 4440 8964
rect 4400 8884 4404 8916
rect 4436 8884 4440 8916
rect 4400 8836 4440 8884
rect 4400 8804 4404 8836
rect 4436 8804 4440 8836
rect 4400 8756 4440 8804
rect 4400 8724 4404 8756
rect 4436 8724 4440 8756
rect 4400 8676 4440 8724
rect 4400 8644 4404 8676
rect 4436 8644 4440 8676
rect 4400 8596 4440 8644
rect 4400 8564 4404 8596
rect 4436 8564 4440 8596
rect 4400 8516 4440 8564
rect 4400 8484 4404 8516
rect 4436 8484 4440 8516
rect 4400 8436 4440 8484
rect 4400 8404 4404 8436
rect 4436 8404 4440 8436
rect 4400 8356 4440 8404
rect 4400 8324 4404 8356
rect 4436 8324 4440 8356
rect 4400 8276 4440 8324
rect 4400 8244 4404 8276
rect 4436 8244 4440 8276
rect 4400 8196 4440 8244
rect 4400 8164 4404 8196
rect 4436 8164 4440 8196
rect 4400 8116 4440 8164
rect 4400 8084 4404 8116
rect 4436 8084 4440 8116
rect 4400 8036 4440 8084
rect 4400 8004 4404 8036
rect 4436 8004 4440 8036
rect 4400 7956 4440 8004
rect 4400 7924 4404 7956
rect 4436 7924 4440 7956
rect 4400 7876 4440 7924
rect 4400 7844 4404 7876
rect 4436 7844 4440 7876
rect 4400 7796 4440 7844
rect 4400 7764 4404 7796
rect 4436 7764 4440 7796
rect 4400 7716 4440 7764
rect 4400 7684 4404 7716
rect 4436 7684 4440 7716
rect 4400 7636 4440 7684
rect 4400 7604 4404 7636
rect 4436 7604 4440 7636
rect 4400 7556 4440 7604
rect 4400 7524 4404 7556
rect 4436 7524 4440 7556
rect 4400 7476 4440 7524
rect 4400 7444 4404 7476
rect 4436 7444 4440 7476
rect 4400 7396 4440 7444
rect 4400 7364 4404 7396
rect 4436 7364 4440 7396
rect 4400 7316 4440 7364
rect 4400 7284 4404 7316
rect 4436 7284 4440 7316
rect 4400 7236 4440 7284
rect 4400 7204 4404 7236
rect 4436 7204 4440 7236
rect 4400 7156 4440 7204
rect 4400 7124 4404 7156
rect 4436 7124 4440 7156
rect 4400 7076 4440 7124
rect 4400 7044 4404 7076
rect 4436 7044 4440 7076
rect 4400 6996 4440 7044
rect 4400 6964 4404 6996
rect 4436 6964 4440 6996
rect 4400 6916 4440 6964
rect 4400 6884 4404 6916
rect 4436 6884 4440 6916
rect 4400 6836 4440 6884
rect 4400 6804 4404 6836
rect 4436 6804 4440 6836
rect 4400 6756 4440 6804
rect 4400 6724 4404 6756
rect 4436 6724 4440 6756
rect 4400 6676 4440 6724
rect 4400 6644 4404 6676
rect 4436 6644 4440 6676
rect 4400 6596 4440 6644
rect 4400 6564 4404 6596
rect 4436 6564 4440 6596
rect 4400 6516 4440 6564
rect 4400 6484 4404 6516
rect 4436 6484 4440 6516
rect 4400 6436 4440 6484
rect 4400 6404 4404 6436
rect 4436 6404 4440 6436
rect 4400 6356 4440 6404
rect 4400 6324 4404 6356
rect 4436 6324 4440 6356
rect 4400 6276 4440 6324
rect 4400 6244 4404 6276
rect 4436 6244 4440 6276
rect 4400 6196 4440 6244
rect 4400 6164 4404 6196
rect 4436 6164 4440 6196
rect 4400 6116 4440 6164
rect 4400 6084 4404 6116
rect 4436 6084 4440 6116
rect 4400 6036 4440 6084
rect 4400 6004 4404 6036
rect 4436 6004 4440 6036
rect 4400 5956 4440 6004
rect 4400 5924 4404 5956
rect 4436 5924 4440 5956
rect 4400 5876 4440 5924
rect 4400 5844 4404 5876
rect 4436 5844 4440 5876
rect 4400 5796 4440 5844
rect 4400 5764 4404 5796
rect 4436 5764 4440 5796
rect 4400 5716 4440 5764
rect 4400 5684 4404 5716
rect 4436 5684 4440 5716
rect 4400 5636 4440 5684
rect 4400 5604 4404 5636
rect 4436 5604 4440 5636
rect 4400 5556 4440 5604
rect 4400 5524 4404 5556
rect 4436 5524 4440 5556
rect 4400 5476 4440 5524
rect 4400 5444 4404 5476
rect 4436 5444 4440 5476
rect 4400 5396 4440 5444
rect 4400 5364 4404 5396
rect 4436 5364 4440 5396
rect 4400 5316 4440 5364
rect 4400 5284 4404 5316
rect 4436 5284 4440 5316
rect 4400 5236 4440 5284
rect 4400 5204 4404 5236
rect 4436 5204 4440 5236
rect 4400 5156 4440 5204
rect 4400 5124 4404 5156
rect 4436 5124 4440 5156
rect 4400 5076 4440 5124
rect 4400 5044 4404 5076
rect 4436 5044 4440 5076
rect 4400 4996 4440 5044
rect 4400 4964 4404 4996
rect 4436 4964 4440 4996
rect 4400 4916 4440 4964
rect 4400 4884 4404 4916
rect 4436 4884 4440 4916
rect 4400 4836 4440 4884
rect 4400 4804 4404 4836
rect 4436 4804 4440 4836
rect 4400 4756 4440 4804
rect 4400 4724 4404 4756
rect 4436 4724 4440 4756
rect 4400 4676 4440 4724
rect 4400 4644 4404 4676
rect 4436 4644 4440 4676
rect 4400 4596 4440 4644
rect 4400 4564 4404 4596
rect 4436 4564 4440 4596
rect 4400 4516 4440 4564
rect 4400 4484 4404 4516
rect 4436 4484 4440 4516
rect 4400 4436 4440 4484
rect 4400 4404 4404 4436
rect 4436 4404 4440 4436
rect 4400 4356 4440 4404
rect 4400 4324 4404 4356
rect 4436 4324 4440 4356
rect 4400 4276 4440 4324
rect 4400 4244 4404 4276
rect 4436 4244 4440 4276
rect 4400 4196 4440 4244
rect 4400 4164 4404 4196
rect 4436 4164 4440 4196
rect 4400 4116 4440 4164
rect 4400 4084 4404 4116
rect 4436 4084 4440 4116
rect 4400 4036 4440 4084
rect 4400 4004 4404 4036
rect 4436 4004 4440 4036
rect 4400 3956 4440 4004
rect 4400 3924 4404 3956
rect 4436 3924 4440 3956
rect 4400 3876 4440 3924
rect 4400 3844 4404 3876
rect 4436 3844 4440 3876
rect 4400 3796 4440 3844
rect 4400 3764 4404 3796
rect 4436 3764 4440 3796
rect 4400 3716 4440 3764
rect 4400 3684 4404 3716
rect 4436 3684 4440 3716
rect 4400 3636 4440 3684
rect 4400 3604 4404 3636
rect 4436 3604 4440 3636
rect 4400 3556 4440 3604
rect 4400 3524 4404 3556
rect 4436 3524 4440 3556
rect 4400 3476 4440 3524
rect 4400 3444 4404 3476
rect 4436 3444 4440 3476
rect 4400 3396 4440 3444
rect 4400 3364 4404 3396
rect 4436 3364 4440 3396
rect 4400 3316 4440 3364
rect 4400 3284 4404 3316
rect 4436 3284 4440 3316
rect 4400 3236 4440 3284
rect 4400 3204 4404 3236
rect 4436 3204 4440 3236
rect 4400 3156 4440 3204
rect 4400 3124 4404 3156
rect 4436 3124 4440 3156
rect 4400 3076 4440 3124
rect 4400 3044 4404 3076
rect 4436 3044 4440 3076
rect 4400 2996 4440 3044
rect 4400 2964 4404 2996
rect 4436 2964 4440 2996
rect 4400 2916 4440 2964
rect 4400 2884 4404 2916
rect 4436 2884 4440 2916
rect 4400 2836 4440 2884
rect 4400 2804 4404 2836
rect 4436 2804 4440 2836
rect 4400 2756 4440 2804
rect 4400 2724 4404 2756
rect 4436 2724 4440 2756
rect 4400 2676 4440 2724
rect 4400 2644 4404 2676
rect 4436 2644 4440 2676
rect 4400 2596 4440 2644
rect 4400 2564 4404 2596
rect 4436 2564 4440 2596
rect 4400 2516 4440 2564
rect 4400 2484 4404 2516
rect 4436 2484 4440 2516
rect 4400 2436 4440 2484
rect 4400 2404 4404 2436
rect 4436 2404 4440 2436
rect 4400 2356 4440 2404
rect 4400 2324 4404 2356
rect 4436 2324 4440 2356
rect 4400 2276 4440 2324
rect 4400 2244 4404 2276
rect 4436 2244 4440 2276
rect 4400 2196 4440 2244
rect 4400 2164 4404 2196
rect 4436 2164 4440 2196
rect 4400 2116 4440 2164
rect 4400 2084 4404 2116
rect 4436 2084 4440 2116
rect 4400 2036 4440 2084
rect 4400 2004 4404 2036
rect 4436 2004 4440 2036
rect 4400 1956 4440 2004
rect 4400 1924 4404 1956
rect 4436 1924 4440 1956
rect 4400 1876 4440 1924
rect 4400 1844 4404 1876
rect 4436 1844 4440 1876
rect 4400 1796 4440 1844
rect 4400 1764 4404 1796
rect 4436 1764 4440 1796
rect 4400 1716 4440 1764
rect 4400 1684 4404 1716
rect 4436 1684 4440 1716
rect 4400 1636 4440 1684
rect 4400 1604 4404 1636
rect 4436 1604 4440 1636
rect 4400 1556 4440 1604
rect 4400 1524 4404 1556
rect 4436 1524 4440 1556
rect 4400 1476 4440 1524
rect 4400 1444 4404 1476
rect 4436 1444 4440 1476
rect 4400 1396 4440 1444
rect 4400 1364 4404 1396
rect 4436 1364 4440 1396
rect 4400 1316 4440 1364
rect 4400 1284 4404 1316
rect 4436 1284 4440 1316
rect 4400 1236 4440 1284
rect 4400 1204 4404 1236
rect 4436 1204 4440 1236
rect 4400 1156 4440 1204
rect 4400 1124 4404 1156
rect 4436 1124 4440 1156
rect 4400 1076 4440 1124
rect 4400 1044 4404 1076
rect 4436 1044 4440 1076
rect 4400 996 4440 1044
rect 4400 964 4404 996
rect 4436 964 4440 996
rect 4400 916 4440 964
rect 4400 884 4404 916
rect 4436 884 4440 916
rect 4400 836 4440 884
rect 4400 804 4404 836
rect 4436 804 4440 836
rect 4400 756 4440 804
rect 4400 724 4404 756
rect 4436 724 4440 756
rect 4400 676 4440 724
rect 4400 644 4404 676
rect 4436 644 4440 676
rect 4400 596 4440 644
rect 4400 564 4404 596
rect 4436 564 4440 596
rect 4400 516 4440 564
rect 4400 484 4404 516
rect 4436 484 4440 516
rect 4400 436 4440 484
rect 4400 404 4404 436
rect 4436 404 4440 436
rect 4400 356 4440 404
rect 4400 324 4404 356
rect 4436 324 4440 356
rect 4400 276 4440 324
rect 4400 244 4404 276
rect 4436 244 4440 276
rect 4400 196 4440 244
rect 4400 164 4404 196
rect 4436 164 4440 196
rect 4400 116 4440 164
rect 4400 84 4404 116
rect 4436 84 4440 116
rect 4400 36 4440 84
rect 4400 4 4404 36
rect 4436 4 4440 36
rect 4240 -956 4244 -764
rect 4276 -956 4280 -764
rect 4240 -960 4280 -956
rect 4400 -764 4440 4
rect 4400 -956 4404 -764
rect 4436 -956 4440 -764
rect 4400 -960 4440 -956
rect 4480 15716 4520 15760
rect 4480 15684 4484 15716
rect 4516 15684 4520 15716
rect 4480 15636 4520 15684
rect 4480 15604 4484 15636
rect 4516 15604 4520 15636
rect 4480 15556 4520 15604
rect 4480 15524 4484 15556
rect 4516 15524 4520 15556
rect 4480 15476 4520 15524
rect 4480 15444 4484 15476
rect 4516 15444 4520 15476
rect 4480 15396 4520 15444
rect 4480 15364 4484 15396
rect 4516 15364 4520 15396
rect 4480 15316 4520 15364
rect 4480 15284 4484 15316
rect 4516 15284 4520 15316
rect 4480 15236 4520 15284
rect 4480 15204 4484 15236
rect 4516 15204 4520 15236
rect 4480 15156 4520 15204
rect 4480 15124 4484 15156
rect 4516 15124 4520 15156
rect 4480 15076 4520 15124
rect 4480 15044 4484 15076
rect 4516 15044 4520 15076
rect 4480 14996 4520 15044
rect 4480 14964 4484 14996
rect 4516 14964 4520 14996
rect 4480 14916 4520 14964
rect 4480 14884 4484 14916
rect 4516 14884 4520 14916
rect 4480 14836 4520 14884
rect 4480 14804 4484 14836
rect 4516 14804 4520 14836
rect 4480 14756 4520 14804
rect 4480 14724 4484 14756
rect 4516 14724 4520 14756
rect 4480 14676 4520 14724
rect 4480 14644 4484 14676
rect 4516 14644 4520 14676
rect 4480 14596 4520 14644
rect 4480 14564 4484 14596
rect 4516 14564 4520 14596
rect 4480 14516 4520 14564
rect 4480 14484 4484 14516
rect 4516 14484 4520 14516
rect 4480 14436 4520 14484
rect 4480 14404 4484 14436
rect 4516 14404 4520 14436
rect 4480 14356 4520 14404
rect 4480 14324 4484 14356
rect 4516 14324 4520 14356
rect 4480 14276 4520 14324
rect 4480 14244 4484 14276
rect 4516 14244 4520 14276
rect 4480 14196 4520 14244
rect 4480 14164 4484 14196
rect 4516 14164 4520 14196
rect 4480 14116 4520 14164
rect 4480 14084 4484 14116
rect 4516 14084 4520 14116
rect 4480 14036 4520 14084
rect 4480 14004 4484 14036
rect 4516 14004 4520 14036
rect 4480 13956 4520 14004
rect 4480 13924 4484 13956
rect 4516 13924 4520 13956
rect 4480 13876 4520 13924
rect 4480 13844 4484 13876
rect 4516 13844 4520 13876
rect 4480 13796 4520 13844
rect 4480 13764 4484 13796
rect 4516 13764 4520 13796
rect 4480 13716 4520 13764
rect 4480 13684 4484 13716
rect 4516 13684 4520 13716
rect 4480 13636 4520 13684
rect 4480 13604 4484 13636
rect 4516 13604 4520 13636
rect 4480 13556 4520 13604
rect 4480 13524 4484 13556
rect 4516 13524 4520 13556
rect 4480 13476 4520 13524
rect 4480 13444 4484 13476
rect 4516 13444 4520 13476
rect 4480 13396 4520 13444
rect 4480 13364 4484 13396
rect 4516 13364 4520 13396
rect 4480 13316 4520 13364
rect 4480 13284 4484 13316
rect 4516 13284 4520 13316
rect 4480 13236 4520 13284
rect 4480 13204 4484 13236
rect 4516 13204 4520 13236
rect 4480 13156 4520 13204
rect 4480 13124 4484 13156
rect 4516 13124 4520 13156
rect 4480 13076 4520 13124
rect 4480 13044 4484 13076
rect 4516 13044 4520 13076
rect 4480 12996 4520 13044
rect 4480 12964 4484 12996
rect 4516 12964 4520 12996
rect 4480 12916 4520 12964
rect 4480 12884 4484 12916
rect 4516 12884 4520 12916
rect 4480 12836 4520 12884
rect 4480 12804 4484 12836
rect 4516 12804 4520 12836
rect 4480 12756 4520 12804
rect 4480 12724 4484 12756
rect 4516 12724 4520 12756
rect 4480 12676 4520 12724
rect 4480 12644 4484 12676
rect 4516 12644 4520 12676
rect 4480 12596 4520 12644
rect 4480 12564 4484 12596
rect 4516 12564 4520 12596
rect 4480 12516 4520 12564
rect 4480 12484 4484 12516
rect 4516 12484 4520 12516
rect 4480 12436 4520 12484
rect 4480 12404 4484 12436
rect 4516 12404 4520 12436
rect 4480 12356 4520 12404
rect 4480 12324 4484 12356
rect 4516 12324 4520 12356
rect 4480 12276 4520 12324
rect 4480 12244 4484 12276
rect 4516 12244 4520 12276
rect 4480 12196 4520 12244
rect 4480 12164 4484 12196
rect 4516 12164 4520 12196
rect 4480 12116 4520 12164
rect 4480 12084 4484 12116
rect 4516 12084 4520 12116
rect 4480 12036 4520 12084
rect 4480 12004 4484 12036
rect 4516 12004 4520 12036
rect 4480 11956 4520 12004
rect 4480 11924 4484 11956
rect 4516 11924 4520 11956
rect 4480 11876 4520 11924
rect 4480 11844 4484 11876
rect 4516 11844 4520 11876
rect 4480 11796 4520 11844
rect 4480 11764 4484 11796
rect 4516 11764 4520 11796
rect 4480 11716 4520 11764
rect 4480 11684 4484 11716
rect 4516 11684 4520 11716
rect 4480 11636 4520 11684
rect 4480 11604 4484 11636
rect 4516 11604 4520 11636
rect 4480 11556 4520 11604
rect 4480 11524 4484 11556
rect 4516 11524 4520 11556
rect 4480 11476 4520 11524
rect 4480 11444 4484 11476
rect 4516 11444 4520 11476
rect 4480 11396 4520 11444
rect 4480 11364 4484 11396
rect 4516 11364 4520 11396
rect 4480 11316 4520 11364
rect 4480 11284 4484 11316
rect 4516 11284 4520 11316
rect 4480 11236 4520 11284
rect 4480 11204 4484 11236
rect 4516 11204 4520 11236
rect 4480 11156 4520 11204
rect 4480 11124 4484 11156
rect 4516 11124 4520 11156
rect 4480 11076 4520 11124
rect 4480 11044 4484 11076
rect 4516 11044 4520 11076
rect 4480 10996 4520 11044
rect 4480 10964 4484 10996
rect 4516 10964 4520 10996
rect 4480 10916 4520 10964
rect 4480 10884 4484 10916
rect 4516 10884 4520 10916
rect 4480 10836 4520 10884
rect 4480 10804 4484 10836
rect 4516 10804 4520 10836
rect 4480 10756 4520 10804
rect 4480 10724 4484 10756
rect 4516 10724 4520 10756
rect 4480 10676 4520 10724
rect 4480 10644 4484 10676
rect 4516 10644 4520 10676
rect 4480 10596 4520 10644
rect 4480 10564 4484 10596
rect 4516 10564 4520 10596
rect 4480 10516 4520 10564
rect 4480 10484 4484 10516
rect 4516 10484 4520 10516
rect 4480 10436 4520 10484
rect 4480 10404 4484 10436
rect 4516 10404 4520 10436
rect 4480 10356 4520 10404
rect 4480 10324 4484 10356
rect 4516 10324 4520 10356
rect 4480 10276 4520 10324
rect 4480 10244 4484 10276
rect 4516 10244 4520 10276
rect 4480 10196 4520 10244
rect 4480 10164 4484 10196
rect 4516 10164 4520 10196
rect 4480 10116 4520 10164
rect 4480 10084 4484 10116
rect 4516 10084 4520 10116
rect 4480 10036 4520 10084
rect 4480 10004 4484 10036
rect 4516 10004 4520 10036
rect 4480 9956 4520 10004
rect 4480 9924 4484 9956
rect 4516 9924 4520 9956
rect 4480 9876 4520 9924
rect 4480 9844 4484 9876
rect 4516 9844 4520 9876
rect 4480 9796 4520 9844
rect 4480 9764 4484 9796
rect 4516 9764 4520 9796
rect 4480 9716 4520 9764
rect 4480 9684 4484 9716
rect 4516 9684 4520 9716
rect 4480 9636 4520 9684
rect 4480 9604 4484 9636
rect 4516 9604 4520 9636
rect 4480 9556 4520 9604
rect 4480 9524 4484 9556
rect 4516 9524 4520 9556
rect 4480 9476 4520 9524
rect 4480 9444 4484 9476
rect 4516 9444 4520 9476
rect 4480 9396 4520 9444
rect 4480 9364 4484 9396
rect 4516 9364 4520 9396
rect 4480 9316 4520 9364
rect 4480 9284 4484 9316
rect 4516 9284 4520 9316
rect 4480 9236 4520 9284
rect 4480 9204 4484 9236
rect 4516 9204 4520 9236
rect 4480 9156 4520 9204
rect 4480 9124 4484 9156
rect 4516 9124 4520 9156
rect 4480 9076 4520 9124
rect 4480 9044 4484 9076
rect 4516 9044 4520 9076
rect 4480 8996 4520 9044
rect 4480 8964 4484 8996
rect 4516 8964 4520 8996
rect 4480 8916 4520 8964
rect 4480 8884 4484 8916
rect 4516 8884 4520 8916
rect 4480 8836 4520 8884
rect 4480 8804 4484 8836
rect 4516 8804 4520 8836
rect 4480 8756 4520 8804
rect 4480 8724 4484 8756
rect 4516 8724 4520 8756
rect 4480 8676 4520 8724
rect 4480 8644 4484 8676
rect 4516 8644 4520 8676
rect 4480 8596 4520 8644
rect 4480 8564 4484 8596
rect 4516 8564 4520 8596
rect 4480 8516 4520 8564
rect 4480 8484 4484 8516
rect 4516 8484 4520 8516
rect 4480 8436 4520 8484
rect 4480 8404 4484 8436
rect 4516 8404 4520 8436
rect 4480 8356 4520 8404
rect 4480 8324 4484 8356
rect 4516 8324 4520 8356
rect 4480 8276 4520 8324
rect 4480 8244 4484 8276
rect 4516 8244 4520 8276
rect 4480 8196 4520 8244
rect 4480 8164 4484 8196
rect 4516 8164 4520 8196
rect 4480 8116 4520 8164
rect 4480 8084 4484 8116
rect 4516 8084 4520 8116
rect 4480 8036 4520 8084
rect 4480 8004 4484 8036
rect 4516 8004 4520 8036
rect 4480 7956 4520 8004
rect 4480 7924 4484 7956
rect 4516 7924 4520 7956
rect 4480 7876 4520 7924
rect 4480 7844 4484 7876
rect 4516 7844 4520 7876
rect 4480 7796 4520 7844
rect 4480 7764 4484 7796
rect 4516 7764 4520 7796
rect 4480 7716 4520 7764
rect 4480 7684 4484 7716
rect 4516 7684 4520 7716
rect 4480 7636 4520 7684
rect 4480 7604 4484 7636
rect 4516 7604 4520 7636
rect 4480 7556 4520 7604
rect 4480 7524 4484 7556
rect 4516 7524 4520 7556
rect 4480 7476 4520 7524
rect 4480 7444 4484 7476
rect 4516 7444 4520 7476
rect 4480 7396 4520 7444
rect 4480 7364 4484 7396
rect 4516 7364 4520 7396
rect 4480 7316 4520 7364
rect 4480 7284 4484 7316
rect 4516 7284 4520 7316
rect 4480 7236 4520 7284
rect 4480 7204 4484 7236
rect 4516 7204 4520 7236
rect 4480 7156 4520 7204
rect 4480 7124 4484 7156
rect 4516 7124 4520 7156
rect 4480 7076 4520 7124
rect 4480 7044 4484 7076
rect 4516 7044 4520 7076
rect 4480 6996 4520 7044
rect 4480 6964 4484 6996
rect 4516 6964 4520 6996
rect 4480 6916 4520 6964
rect 4480 6884 4484 6916
rect 4516 6884 4520 6916
rect 4480 6836 4520 6884
rect 4480 6804 4484 6836
rect 4516 6804 4520 6836
rect 4480 6756 4520 6804
rect 4480 6724 4484 6756
rect 4516 6724 4520 6756
rect 4480 6676 4520 6724
rect 4480 6644 4484 6676
rect 4516 6644 4520 6676
rect 4480 6596 4520 6644
rect 4480 6564 4484 6596
rect 4516 6564 4520 6596
rect 4480 6516 4520 6564
rect 4480 6484 4484 6516
rect 4516 6484 4520 6516
rect 4480 6436 4520 6484
rect 4480 6404 4484 6436
rect 4516 6404 4520 6436
rect 4480 6356 4520 6404
rect 4480 6324 4484 6356
rect 4516 6324 4520 6356
rect 4480 6276 4520 6324
rect 4480 6244 4484 6276
rect 4516 6244 4520 6276
rect 4480 6196 4520 6244
rect 4480 6164 4484 6196
rect 4516 6164 4520 6196
rect 4480 6116 4520 6164
rect 4480 6084 4484 6116
rect 4516 6084 4520 6116
rect 4480 6036 4520 6084
rect 4480 6004 4484 6036
rect 4516 6004 4520 6036
rect 4480 5956 4520 6004
rect 4480 5924 4484 5956
rect 4516 5924 4520 5956
rect 4480 5876 4520 5924
rect 4480 5844 4484 5876
rect 4516 5844 4520 5876
rect 4480 5796 4520 5844
rect 4480 5764 4484 5796
rect 4516 5764 4520 5796
rect 4480 5716 4520 5764
rect 4480 5684 4484 5716
rect 4516 5684 4520 5716
rect 4480 5636 4520 5684
rect 4480 5604 4484 5636
rect 4516 5604 4520 5636
rect 4480 5556 4520 5604
rect 4480 5524 4484 5556
rect 4516 5524 4520 5556
rect 4480 5476 4520 5524
rect 4480 5444 4484 5476
rect 4516 5444 4520 5476
rect 4480 5396 4520 5444
rect 4480 5364 4484 5396
rect 4516 5364 4520 5396
rect 4480 5316 4520 5364
rect 4480 5284 4484 5316
rect 4516 5284 4520 5316
rect 4480 5236 4520 5284
rect 4480 5204 4484 5236
rect 4516 5204 4520 5236
rect 4480 5156 4520 5204
rect 4480 5124 4484 5156
rect 4516 5124 4520 5156
rect 4480 5076 4520 5124
rect 4480 5044 4484 5076
rect 4516 5044 4520 5076
rect 4480 4996 4520 5044
rect 4480 4964 4484 4996
rect 4516 4964 4520 4996
rect 4480 4916 4520 4964
rect 4480 4884 4484 4916
rect 4516 4884 4520 4916
rect 4480 4836 4520 4884
rect 4480 4804 4484 4836
rect 4516 4804 4520 4836
rect 4480 4756 4520 4804
rect 4480 4724 4484 4756
rect 4516 4724 4520 4756
rect 4480 4676 4520 4724
rect 4480 4644 4484 4676
rect 4516 4644 4520 4676
rect 4480 4596 4520 4644
rect 4480 4564 4484 4596
rect 4516 4564 4520 4596
rect 4480 4516 4520 4564
rect 4480 4484 4484 4516
rect 4516 4484 4520 4516
rect 4480 4436 4520 4484
rect 4480 4404 4484 4436
rect 4516 4404 4520 4436
rect 4480 4356 4520 4404
rect 4480 4324 4484 4356
rect 4516 4324 4520 4356
rect 4480 4276 4520 4324
rect 4480 4244 4484 4276
rect 4516 4244 4520 4276
rect 4480 4196 4520 4244
rect 4480 4164 4484 4196
rect 4516 4164 4520 4196
rect 4480 4116 4520 4164
rect 4480 4084 4484 4116
rect 4516 4084 4520 4116
rect 4480 4036 4520 4084
rect 4480 4004 4484 4036
rect 4516 4004 4520 4036
rect 4480 3956 4520 4004
rect 4480 3924 4484 3956
rect 4516 3924 4520 3956
rect 4480 3876 4520 3924
rect 4480 3844 4484 3876
rect 4516 3844 4520 3876
rect 4480 3796 4520 3844
rect 4480 3764 4484 3796
rect 4516 3764 4520 3796
rect 4480 3716 4520 3764
rect 4480 3684 4484 3716
rect 4516 3684 4520 3716
rect 4480 3636 4520 3684
rect 4480 3604 4484 3636
rect 4516 3604 4520 3636
rect 4480 3556 4520 3604
rect 4480 3524 4484 3556
rect 4516 3524 4520 3556
rect 4480 3476 4520 3524
rect 4480 3444 4484 3476
rect 4516 3444 4520 3476
rect 4480 3396 4520 3444
rect 4480 3364 4484 3396
rect 4516 3364 4520 3396
rect 4480 3316 4520 3364
rect 4480 3284 4484 3316
rect 4516 3284 4520 3316
rect 4480 3236 4520 3284
rect 4480 3204 4484 3236
rect 4516 3204 4520 3236
rect 4480 3156 4520 3204
rect 4480 3124 4484 3156
rect 4516 3124 4520 3156
rect 4480 3076 4520 3124
rect 4480 3044 4484 3076
rect 4516 3044 4520 3076
rect 4480 2996 4520 3044
rect 4480 2964 4484 2996
rect 4516 2964 4520 2996
rect 4480 2916 4520 2964
rect 4480 2884 4484 2916
rect 4516 2884 4520 2916
rect 4480 2836 4520 2884
rect 4480 2804 4484 2836
rect 4516 2804 4520 2836
rect 4480 2756 4520 2804
rect 4480 2724 4484 2756
rect 4516 2724 4520 2756
rect 4480 2676 4520 2724
rect 4480 2644 4484 2676
rect 4516 2644 4520 2676
rect 4480 2596 4520 2644
rect 4480 2564 4484 2596
rect 4516 2564 4520 2596
rect 4480 2516 4520 2564
rect 4480 2484 4484 2516
rect 4516 2484 4520 2516
rect 4480 2436 4520 2484
rect 4480 2404 4484 2436
rect 4516 2404 4520 2436
rect 4480 2356 4520 2404
rect 4480 2324 4484 2356
rect 4516 2324 4520 2356
rect 4480 2276 4520 2324
rect 4480 2244 4484 2276
rect 4516 2244 4520 2276
rect 4480 2196 4520 2244
rect 4480 2164 4484 2196
rect 4516 2164 4520 2196
rect 4480 2116 4520 2164
rect 4480 2084 4484 2116
rect 4516 2084 4520 2116
rect 4480 2036 4520 2084
rect 4480 2004 4484 2036
rect 4516 2004 4520 2036
rect 4480 1956 4520 2004
rect 4480 1924 4484 1956
rect 4516 1924 4520 1956
rect 4480 1876 4520 1924
rect 4480 1844 4484 1876
rect 4516 1844 4520 1876
rect 4480 1796 4520 1844
rect 4480 1764 4484 1796
rect 4516 1764 4520 1796
rect 4480 1716 4520 1764
rect 4480 1684 4484 1716
rect 4516 1684 4520 1716
rect 4480 1636 4520 1684
rect 4480 1604 4484 1636
rect 4516 1604 4520 1636
rect 4480 1556 4520 1604
rect 4480 1524 4484 1556
rect 4516 1524 4520 1556
rect 4480 1476 4520 1524
rect 4480 1444 4484 1476
rect 4516 1444 4520 1476
rect 4480 1396 4520 1444
rect 4480 1364 4484 1396
rect 4516 1364 4520 1396
rect 4480 1316 4520 1364
rect 4480 1284 4484 1316
rect 4516 1284 4520 1316
rect 4480 1236 4520 1284
rect 4480 1204 4484 1236
rect 4516 1204 4520 1236
rect 4480 1156 4520 1204
rect 4480 1124 4484 1156
rect 4516 1124 4520 1156
rect 4480 1076 4520 1124
rect 4480 1044 4484 1076
rect 4516 1044 4520 1076
rect 4480 996 4520 1044
rect 4480 964 4484 996
rect 4516 964 4520 996
rect 4480 916 4520 964
rect 4480 884 4484 916
rect 4516 884 4520 916
rect 4480 836 4520 884
rect 4480 804 4484 836
rect 4516 804 4520 836
rect 4480 756 4520 804
rect 4480 724 4484 756
rect 4516 724 4520 756
rect 4480 676 4520 724
rect 4480 644 4484 676
rect 4516 644 4520 676
rect 4480 596 4520 644
rect 4480 564 4484 596
rect 4516 564 4520 596
rect 4480 516 4520 564
rect 4480 484 4484 516
rect 4516 484 4520 516
rect 4480 436 4520 484
rect 4480 404 4484 436
rect 4516 404 4520 436
rect 4480 356 4520 404
rect 4480 324 4484 356
rect 4516 324 4520 356
rect 4480 276 4520 324
rect 4480 244 4484 276
rect 4516 244 4520 276
rect 4480 196 4520 244
rect 4480 164 4484 196
rect 4516 164 4520 196
rect 4480 116 4520 164
rect 4480 84 4484 116
rect 4516 84 4520 116
rect 4480 36 4520 84
rect 4480 4 4484 36
rect 4516 4 4520 36
rect 4480 -284 4520 4
rect 4480 -476 4484 -284
rect 4516 -476 4520 -284
rect 120 -1004 160 -1000
rect 120 -1036 124 -1004
rect 156 -1036 160 -1004
rect 120 -2284 160 -1036
rect 4480 -1004 4520 -476
rect 4480 -1036 4484 -1004
rect 4516 -1036 4520 -1004
rect 4480 -1040 4520 -1036
rect 4560 15075 4600 15760
rect 4560 15045 4565 15075
rect 4595 15045 4600 15075
rect 4560 12435 4600 15045
rect 4560 12405 4565 12435
rect 4595 12405 4600 12435
rect 4560 10995 4600 12405
rect 4560 10965 4565 10995
rect 4595 10965 4600 10995
rect 4560 8355 4600 10965
rect 4560 8325 4565 8355
rect 4595 8325 4600 8355
rect 4560 6915 4600 8325
rect 4560 6885 4565 6915
rect 4595 6885 4600 6915
rect 4560 3555 4600 6885
rect 4560 3525 4565 3555
rect 4595 3525 4600 3555
rect 4560 1835 4600 3525
rect 4560 1805 4565 1835
rect 4595 1805 4600 1835
rect 4560 -1080 4600 1805
rect 4640 15716 4680 15760
rect 4640 15684 4644 15716
rect 4676 15684 4680 15716
rect 4640 15636 4680 15684
rect 4640 15604 4644 15636
rect 4676 15604 4680 15636
rect 4640 15556 4680 15604
rect 4640 15524 4644 15556
rect 4676 15524 4680 15556
rect 4640 15476 4680 15524
rect 4640 15444 4644 15476
rect 4676 15444 4680 15476
rect 4640 15396 4680 15444
rect 4640 15364 4644 15396
rect 4676 15364 4680 15396
rect 4640 15316 4680 15364
rect 4640 15284 4644 15316
rect 4676 15284 4680 15316
rect 4640 15236 4680 15284
rect 4640 15204 4644 15236
rect 4676 15204 4680 15236
rect 4640 15156 4680 15204
rect 4640 15124 4644 15156
rect 4676 15124 4680 15156
rect 4640 15076 4680 15124
rect 4640 15044 4644 15076
rect 4676 15044 4680 15076
rect 4640 14996 4680 15044
rect 4640 14964 4644 14996
rect 4676 14964 4680 14996
rect 4640 14916 4680 14964
rect 4640 14884 4644 14916
rect 4676 14884 4680 14916
rect 4640 14836 4680 14884
rect 4640 14804 4644 14836
rect 4676 14804 4680 14836
rect 4640 14756 4680 14804
rect 4640 14724 4644 14756
rect 4676 14724 4680 14756
rect 4640 14676 4680 14724
rect 4640 14644 4644 14676
rect 4676 14644 4680 14676
rect 4640 14596 4680 14644
rect 4640 14564 4644 14596
rect 4676 14564 4680 14596
rect 4640 14516 4680 14564
rect 4640 14484 4644 14516
rect 4676 14484 4680 14516
rect 4640 14436 4680 14484
rect 4640 14404 4644 14436
rect 4676 14404 4680 14436
rect 4640 14356 4680 14404
rect 4640 14324 4644 14356
rect 4676 14324 4680 14356
rect 4640 14276 4680 14324
rect 4640 14244 4644 14276
rect 4676 14244 4680 14276
rect 4640 14196 4680 14244
rect 4640 14164 4644 14196
rect 4676 14164 4680 14196
rect 4640 14116 4680 14164
rect 4640 14084 4644 14116
rect 4676 14084 4680 14116
rect 4640 14036 4680 14084
rect 4640 14004 4644 14036
rect 4676 14004 4680 14036
rect 4640 13956 4680 14004
rect 4640 13924 4644 13956
rect 4676 13924 4680 13956
rect 4640 13876 4680 13924
rect 4640 13844 4644 13876
rect 4676 13844 4680 13876
rect 4640 13796 4680 13844
rect 4640 13764 4644 13796
rect 4676 13764 4680 13796
rect 4640 13716 4680 13764
rect 4640 13684 4644 13716
rect 4676 13684 4680 13716
rect 4640 13636 4680 13684
rect 4640 13604 4644 13636
rect 4676 13604 4680 13636
rect 4640 13556 4680 13604
rect 4640 13524 4644 13556
rect 4676 13524 4680 13556
rect 4640 13476 4680 13524
rect 4640 13444 4644 13476
rect 4676 13444 4680 13476
rect 4640 13396 4680 13444
rect 4640 13364 4644 13396
rect 4676 13364 4680 13396
rect 4640 13316 4680 13364
rect 4640 13284 4644 13316
rect 4676 13284 4680 13316
rect 4640 13236 4680 13284
rect 4640 13204 4644 13236
rect 4676 13204 4680 13236
rect 4640 13156 4680 13204
rect 4640 13124 4644 13156
rect 4676 13124 4680 13156
rect 4640 13076 4680 13124
rect 4640 13044 4644 13076
rect 4676 13044 4680 13076
rect 4640 12996 4680 13044
rect 4640 12964 4644 12996
rect 4676 12964 4680 12996
rect 4640 12916 4680 12964
rect 4640 12884 4644 12916
rect 4676 12884 4680 12916
rect 4640 12836 4680 12884
rect 4640 12804 4644 12836
rect 4676 12804 4680 12836
rect 4640 12756 4680 12804
rect 4640 12724 4644 12756
rect 4676 12724 4680 12756
rect 4640 12676 4680 12724
rect 4640 12644 4644 12676
rect 4676 12644 4680 12676
rect 4640 12596 4680 12644
rect 4640 12564 4644 12596
rect 4676 12564 4680 12596
rect 4640 12516 4680 12564
rect 4640 12484 4644 12516
rect 4676 12484 4680 12516
rect 4640 12436 4680 12484
rect 4640 12404 4644 12436
rect 4676 12404 4680 12436
rect 4640 12356 4680 12404
rect 4640 12324 4644 12356
rect 4676 12324 4680 12356
rect 4640 12276 4680 12324
rect 4640 12244 4644 12276
rect 4676 12244 4680 12276
rect 4640 12196 4680 12244
rect 4640 12164 4644 12196
rect 4676 12164 4680 12196
rect 4640 12116 4680 12164
rect 4640 12084 4644 12116
rect 4676 12084 4680 12116
rect 4640 12036 4680 12084
rect 4640 12004 4644 12036
rect 4676 12004 4680 12036
rect 4640 11956 4680 12004
rect 4640 11924 4644 11956
rect 4676 11924 4680 11956
rect 4640 11876 4680 11924
rect 4640 11844 4644 11876
rect 4676 11844 4680 11876
rect 4640 11796 4680 11844
rect 4640 11764 4644 11796
rect 4676 11764 4680 11796
rect 4640 11716 4680 11764
rect 4640 11684 4644 11716
rect 4676 11684 4680 11716
rect 4640 11636 4680 11684
rect 4640 11604 4644 11636
rect 4676 11604 4680 11636
rect 4640 11556 4680 11604
rect 4640 11524 4644 11556
rect 4676 11524 4680 11556
rect 4640 11476 4680 11524
rect 4640 11444 4644 11476
rect 4676 11444 4680 11476
rect 4640 11396 4680 11444
rect 4640 11364 4644 11396
rect 4676 11364 4680 11396
rect 4640 11316 4680 11364
rect 4640 11284 4644 11316
rect 4676 11284 4680 11316
rect 4640 11236 4680 11284
rect 4640 11204 4644 11236
rect 4676 11204 4680 11236
rect 4640 11156 4680 11204
rect 4640 11124 4644 11156
rect 4676 11124 4680 11156
rect 4640 11076 4680 11124
rect 4640 11044 4644 11076
rect 4676 11044 4680 11076
rect 4640 10996 4680 11044
rect 4640 10964 4644 10996
rect 4676 10964 4680 10996
rect 4640 10916 4680 10964
rect 4640 10884 4644 10916
rect 4676 10884 4680 10916
rect 4640 10836 4680 10884
rect 4640 10804 4644 10836
rect 4676 10804 4680 10836
rect 4640 10756 4680 10804
rect 4640 10724 4644 10756
rect 4676 10724 4680 10756
rect 4640 10676 4680 10724
rect 4640 10644 4644 10676
rect 4676 10644 4680 10676
rect 4640 10596 4680 10644
rect 4640 10564 4644 10596
rect 4676 10564 4680 10596
rect 4640 10516 4680 10564
rect 4640 10484 4644 10516
rect 4676 10484 4680 10516
rect 4640 10436 4680 10484
rect 4640 10404 4644 10436
rect 4676 10404 4680 10436
rect 4640 10356 4680 10404
rect 4640 10324 4644 10356
rect 4676 10324 4680 10356
rect 4640 10276 4680 10324
rect 4640 10244 4644 10276
rect 4676 10244 4680 10276
rect 4640 10196 4680 10244
rect 4640 10164 4644 10196
rect 4676 10164 4680 10196
rect 4640 10116 4680 10164
rect 4640 10084 4644 10116
rect 4676 10084 4680 10116
rect 4640 10036 4680 10084
rect 4640 10004 4644 10036
rect 4676 10004 4680 10036
rect 4640 9956 4680 10004
rect 4640 9924 4644 9956
rect 4676 9924 4680 9956
rect 4640 9876 4680 9924
rect 4640 9844 4644 9876
rect 4676 9844 4680 9876
rect 4640 9796 4680 9844
rect 4640 9764 4644 9796
rect 4676 9764 4680 9796
rect 4640 9716 4680 9764
rect 4640 9684 4644 9716
rect 4676 9684 4680 9716
rect 4640 9636 4680 9684
rect 4640 9604 4644 9636
rect 4676 9604 4680 9636
rect 4640 9556 4680 9604
rect 4640 9524 4644 9556
rect 4676 9524 4680 9556
rect 4640 9476 4680 9524
rect 4640 9444 4644 9476
rect 4676 9444 4680 9476
rect 4640 9396 4680 9444
rect 4640 9364 4644 9396
rect 4676 9364 4680 9396
rect 4640 9316 4680 9364
rect 4640 9284 4644 9316
rect 4676 9284 4680 9316
rect 4640 9236 4680 9284
rect 4640 9204 4644 9236
rect 4676 9204 4680 9236
rect 4640 9156 4680 9204
rect 4640 9124 4644 9156
rect 4676 9124 4680 9156
rect 4640 9076 4680 9124
rect 4640 9044 4644 9076
rect 4676 9044 4680 9076
rect 4640 8996 4680 9044
rect 4640 8964 4644 8996
rect 4676 8964 4680 8996
rect 4640 8916 4680 8964
rect 4640 8884 4644 8916
rect 4676 8884 4680 8916
rect 4640 8836 4680 8884
rect 4640 8804 4644 8836
rect 4676 8804 4680 8836
rect 4640 8756 4680 8804
rect 4640 8724 4644 8756
rect 4676 8724 4680 8756
rect 4640 8676 4680 8724
rect 4640 8644 4644 8676
rect 4676 8644 4680 8676
rect 4640 8596 4680 8644
rect 4640 8564 4644 8596
rect 4676 8564 4680 8596
rect 4640 8516 4680 8564
rect 4640 8484 4644 8516
rect 4676 8484 4680 8516
rect 4640 8436 4680 8484
rect 4640 8404 4644 8436
rect 4676 8404 4680 8436
rect 4640 8356 4680 8404
rect 4640 8324 4644 8356
rect 4676 8324 4680 8356
rect 4640 8276 4680 8324
rect 4640 8244 4644 8276
rect 4676 8244 4680 8276
rect 4640 8196 4680 8244
rect 4640 8164 4644 8196
rect 4676 8164 4680 8196
rect 4640 8116 4680 8164
rect 4640 8084 4644 8116
rect 4676 8084 4680 8116
rect 4640 8036 4680 8084
rect 4640 8004 4644 8036
rect 4676 8004 4680 8036
rect 4640 7956 4680 8004
rect 4640 7924 4644 7956
rect 4676 7924 4680 7956
rect 4640 7876 4680 7924
rect 4640 7844 4644 7876
rect 4676 7844 4680 7876
rect 4640 7796 4680 7844
rect 4640 7764 4644 7796
rect 4676 7764 4680 7796
rect 4640 7716 4680 7764
rect 4640 7684 4644 7716
rect 4676 7684 4680 7716
rect 4640 7636 4680 7684
rect 4640 7604 4644 7636
rect 4676 7604 4680 7636
rect 4640 7556 4680 7604
rect 4640 7524 4644 7556
rect 4676 7524 4680 7556
rect 4640 7476 4680 7524
rect 4640 7444 4644 7476
rect 4676 7444 4680 7476
rect 4640 7396 4680 7444
rect 4640 7364 4644 7396
rect 4676 7364 4680 7396
rect 4640 7316 4680 7364
rect 4640 7284 4644 7316
rect 4676 7284 4680 7316
rect 4640 7236 4680 7284
rect 4640 7204 4644 7236
rect 4676 7204 4680 7236
rect 4640 7156 4680 7204
rect 4640 7124 4644 7156
rect 4676 7124 4680 7156
rect 4640 7076 4680 7124
rect 4640 7044 4644 7076
rect 4676 7044 4680 7076
rect 4640 6996 4680 7044
rect 4640 6964 4644 6996
rect 4676 6964 4680 6996
rect 4640 6916 4680 6964
rect 4640 6884 4644 6916
rect 4676 6884 4680 6916
rect 4640 6836 4680 6884
rect 4640 6804 4644 6836
rect 4676 6804 4680 6836
rect 4640 6756 4680 6804
rect 4640 6724 4644 6756
rect 4676 6724 4680 6756
rect 4640 6676 4680 6724
rect 4640 6644 4644 6676
rect 4676 6644 4680 6676
rect 4640 6596 4680 6644
rect 4640 6564 4644 6596
rect 4676 6564 4680 6596
rect 4640 6516 4680 6564
rect 4640 6484 4644 6516
rect 4676 6484 4680 6516
rect 4640 6436 4680 6484
rect 4640 6404 4644 6436
rect 4676 6404 4680 6436
rect 4640 6356 4680 6404
rect 4640 6324 4644 6356
rect 4676 6324 4680 6356
rect 4640 6276 4680 6324
rect 4640 6244 4644 6276
rect 4676 6244 4680 6276
rect 4640 6196 4680 6244
rect 4640 6164 4644 6196
rect 4676 6164 4680 6196
rect 4640 6116 4680 6164
rect 4640 6084 4644 6116
rect 4676 6084 4680 6116
rect 4640 6036 4680 6084
rect 4640 6004 4644 6036
rect 4676 6004 4680 6036
rect 4640 5956 4680 6004
rect 4640 5924 4644 5956
rect 4676 5924 4680 5956
rect 4640 5876 4680 5924
rect 4640 5844 4644 5876
rect 4676 5844 4680 5876
rect 4640 5796 4680 5844
rect 4640 5764 4644 5796
rect 4676 5764 4680 5796
rect 4640 5716 4680 5764
rect 4640 5684 4644 5716
rect 4676 5684 4680 5716
rect 4640 5636 4680 5684
rect 4640 5604 4644 5636
rect 4676 5604 4680 5636
rect 4640 5556 4680 5604
rect 4640 5524 4644 5556
rect 4676 5524 4680 5556
rect 4640 5476 4680 5524
rect 4640 5444 4644 5476
rect 4676 5444 4680 5476
rect 4640 5396 4680 5444
rect 4640 5364 4644 5396
rect 4676 5364 4680 5396
rect 4640 5316 4680 5364
rect 4640 5284 4644 5316
rect 4676 5284 4680 5316
rect 4640 5236 4680 5284
rect 4640 5204 4644 5236
rect 4676 5204 4680 5236
rect 4640 5156 4680 5204
rect 4640 5124 4644 5156
rect 4676 5124 4680 5156
rect 4640 5076 4680 5124
rect 4640 5044 4644 5076
rect 4676 5044 4680 5076
rect 4640 4996 4680 5044
rect 4640 4964 4644 4996
rect 4676 4964 4680 4996
rect 4640 4916 4680 4964
rect 4640 4884 4644 4916
rect 4676 4884 4680 4916
rect 4640 4836 4680 4884
rect 4640 4804 4644 4836
rect 4676 4804 4680 4836
rect 4640 4756 4680 4804
rect 4640 4724 4644 4756
rect 4676 4724 4680 4756
rect 4640 4676 4680 4724
rect 4640 4644 4644 4676
rect 4676 4644 4680 4676
rect 4640 4596 4680 4644
rect 4640 4564 4644 4596
rect 4676 4564 4680 4596
rect 4640 4516 4680 4564
rect 4640 4484 4644 4516
rect 4676 4484 4680 4516
rect 4640 4436 4680 4484
rect 4640 4404 4644 4436
rect 4676 4404 4680 4436
rect 4640 4356 4680 4404
rect 4640 4324 4644 4356
rect 4676 4324 4680 4356
rect 4640 4276 4680 4324
rect 4640 4244 4644 4276
rect 4676 4244 4680 4276
rect 4640 4196 4680 4244
rect 4640 4164 4644 4196
rect 4676 4164 4680 4196
rect 4640 4116 4680 4164
rect 4640 4084 4644 4116
rect 4676 4084 4680 4116
rect 4640 4036 4680 4084
rect 4640 4004 4644 4036
rect 4676 4004 4680 4036
rect 4640 3956 4680 4004
rect 4640 3924 4644 3956
rect 4676 3924 4680 3956
rect 4640 3876 4680 3924
rect 4640 3844 4644 3876
rect 4676 3844 4680 3876
rect 4640 3796 4680 3844
rect 4640 3764 4644 3796
rect 4676 3764 4680 3796
rect 4640 3716 4680 3764
rect 4640 3684 4644 3716
rect 4676 3684 4680 3716
rect 4640 3636 4680 3684
rect 4640 3604 4644 3636
rect 4676 3604 4680 3636
rect 4640 3556 4680 3604
rect 4640 3524 4644 3556
rect 4676 3524 4680 3556
rect 4640 3476 4680 3524
rect 4640 3444 4644 3476
rect 4676 3444 4680 3476
rect 4640 3396 4680 3444
rect 4640 3364 4644 3396
rect 4676 3364 4680 3396
rect 4640 3316 4680 3364
rect 4640 3284 4644 3316
rect 4676 3284 4680 3316
rect 4640 3236 4680 3284
rect 4640 3204 4644 3236
rect 4676 3204 4680 3236
rect 4640 3156 4680 3204
rect 4640 3124 4644 3156
rect 4676 3124 4680 3156
rect 4640 3076 4680 3124
rect 4640 3044 4644 3076
rect 4676 3044 4680 3076
rect 4640 2996 4680 3044
rect 4640 2964 4644 2996
rect 4676 2964 4680 2996
rect 4640 2916 4680 2964
rect 4640 2884 4644 2916
rect 4676 2884 4680 2916
rect 4640 2836 4680 2884
rect 4640 2804 4644 2836
rect 4676 2804 4680 2836
rect 4640 2756 4680 2804
rect 4640 2724 4644 2756
rect 4676 2724 4680 2756
rect 4640 2676 4680 2724
rect 4640 2644 4644 2676
rect 4676 2644 4680 2676
rect 4640 2596 4680 2644
rect 4640 2564 4644 2596
rect 4676 2564 4680 2596
rect 4640 2516 4680 2564
rect 4640 2484 4644 2516
rect 4676 2484 4680 2516
rect 4640 2436 4680 2484
rect 4640 2404 4644 2436
rect 4676 2404 4680 2436
rect 4640 2356 4680 2404
rect 4640 2324 4644 2356
rect 4676 2324 4680 2356
rect 4640 2276 4680 2324
rect 4640 2244 4644 2276
rect 4676 2244 4680 2276
rect 4640 2196 4680 2244
rect 4640 2164 4644 2196
rect 4676 2164 4680 2196
rect 4640 2116 4680 2164
rect 4640 2084 4644 2116
rect 4676 2084 4680 2116
rect 4640 2036 4680 2084
rect 4640 2004 4644 2036
rect 4676 2004 4680 2036
rect 4640 1956 4680 2004
rect 4640 1924 4644 1956
rect 4676 1924 4680 1956
rect 4640 1876 4680 1924
rect 4640 1844 4644 1876
rect 4676 1844 4680 1876
rect 4640 1796 4680 1844
rect 4640 1764 4644 1796
rect 4676 1764 4680 1796
rect 4640 1716 4680 1764
rect 4640 1684 4644 1716
rect 4676 1684 4680 1716
rect 4640 1636 4680 1684
rect 4640 1604 4644 1636
rect 4676 1604 4680 1636
rect 4640 1556 4680 1604
rect 4640 1524 4644 1556
rect 4676 1524 4680 1556
rect 4640 1476 4680 1524
rect 4640 1444 4644 1476
rect 4676 1444 4680 1476
rect 4640 1396 4680 1444
rect 4640 1364 4644 1396
rect 4676 1364 4680 1396
rect 4640 1316 4680 1364
rect 4640 1284 4644 1316
rect 4676 1284 4680 1316
rect 4640 1236 4680 1284
rect 4640 1204 4644 1236
rect 4676 1204 4680 1236
rect 4640 1156 4680 1204
rect 4640 1124 4644 1156
rect 4676 1124 4680 1156
rect 4640 1076 4680 1124
rect 4640 1044 4644 1076
rect 4676 1044 4680 1076
rect 4640 996 4680 1044
rect 4640 964 4644 996
rect 4676 964 4680 996
rect 4640 916 4680 964
rect 4640 884 4644 916
rect 4676 884 4680 916
rect 4640 836 4680 884
rect 4640 804 4644 836
rect 4676 804 4680 836
rect 4640 756 4680 804
rect 4640 724 4644 756
rect 4676 724 4680 756
rect 4640 676 4680 724
rect 4640 644 4644 676
rect 4676 644 4680 676
rect 4640 596 4680 644
rect 4640 564 4644 596
rect 4676 564 4680 596
rect 4640 516 4680 564
rect 4640 484 4644 516
rect 4676 484 4680 516
rect 4640 436 4680 484
rect 4640 404 4644 436
rect 4676 404 4680 436
rect 4640 356 4680 404
rect 4640 324 4644 356
rect 4676 324 4680 356
rect 4640 276 4680 324
rect 4640 244 4644 276
rect 4676 244 4680 276
rect 4640 196 4680 244
rect 4640 164 4644 196
rect 4676 164 4680 196
rect 4640 116 4680 164
rect 4640 84 4644 116
rect 4676 84 4680 116
rect 4640 36 4680 84
rect 4640 4 4644 36
rect 4676 4 4680 36
rect 4640 -284 4680 4
rect 4640 -476 4644 -284
rect 4676 -476 4680 -284
rect 4640 -1004 4680 -476
rect 4720 15716 4760 15760
rect 4720 15684 4724 15716
rect 4756 15684 4760 15716
rect 4720 15636 4760 15684
rect 4720 15604 4724 15636
rect 4756 15604 4760 15636
rect 4720 15556 4760 15604
rect 4720 15524 4724 15556
rect 4756 15524 4760 15556
rect 4720 15476 4760 15524
rect 4720 15444 4724 15476
rect 4756 15444 4760 15476
rect 4720 15396 4760 15444
rect 4720 15364 4724 15396
rect 4756 15364 4760 15396
rect 4720 15316 4760 15364
rect 4720 15284 4724 15316
rect 4756 15284 4760 15316
rect 4720 15236 4760 15284
rect 4720 15204 4724 15236
rect 4756 15204 4760 15236
rect 4720 15156 4760 15204
rect 4720 15124 4724 15156
rect 4756 15124 4760 15156
rect 4720 15076 4760 15124
rect 4720 15044 4724 15076
rect 4756 15044 4760 15076
rect 4720 14996 4760 15044
rect 4720 14964 4724 14996
rect 4756 14964 4760 14996
rect 4720 14916 4760 14964
rect 4720 14884 4724 14916
rect 4756 14884 4760 14916
rect 4720 14836 4760 14884
rect 4720 14804 4724 14836
rect 4756 14804 4760 14836
rect 4720 14756 4760 14804
rect 4720 14724 4724 14756
rect 4756 14724 4760 14756
rect 4720 14676 4760 14724
rect 4720 14644 4724 14676
rect 4756 14644 4760 14676
rect 4720 14596 4760 14644
rect 4720 14564 4724 14596
rect 4756 14564 4760 14596
rect 4720 14516 4760 14564
rect 4720 14484 4724 14516
rect 4756 14484 4760 14516
rect 4720 14436 4760 14484
rect 4720 14404 4724 14436
rect 4756 14404 4760 14436
rect 4720 14356 4760 14404
rect 4720 14324 4724 14356
rect 4756 14324 4760 14356
rect 4720 14276 4760 14324
rect 4720 14244 4724 14276
rect 4756 14244 4760 14276
rect 4720 14196 4760 14244
rect 4720 14164 4724 14196
rect 4756 14164 4760 14196
rect 4720 14116 4760 14164
rect 4720 14084 4724 14116
rect 4756 14084 4760 14116
rect 4720 14036 4760 14084
rect 4720 14004 4724 14036
rect 4756 14004 4760 14036
rect 4720 13956 4760 14004
rect 4720 13924 4724 13956
rect 4756 13924 4760 13956
rect 4720 13876 4760 13924
rect 4720 13844 4724 13876
rect 4756 13844 4760 13876
rect 4720 13796 4760 13844
rect 4720 13764 4724 13796
rect 4756 13764 4760 13796
rect 4720 13716 4760 13764
rect 4720 13684 4724 13716
rect 4756 13684 4760 13716
rect 4720 13636 4760 13684
rect 4720 13604 4724 13636
rect 4756 13604 4760 13636
rect 4720 13556 4760 13604
rect 4720 13524 4724 13556
rect 4756 13524 4760 13556
rect 4720 13476 4760 13524
rect 4720 13444 4724 13476
rect 4756 13444 4760 13476
rect 4720 13396 4760 13444
rect 4720 13364 4724 13396
rect 4756 13364 4760 13396
rect 4720 13316 4760 13364
rect 4720 13284 4724 13316
rect 4756 13284 4760 13316
rect 4720 13236 4760 13284
rect 4720 13204 4724 13236
rect 4756 13204 4760 13236
rect 4720 13156 4760 13204
rect 4720 13124 4724 13156
rect 4756 13124 4760 13156
rect 4720 13076 4760 13124
rect 4720 13044 4724 13076
rect 4756 13044 4760 13076
rect 4720 12996 4760 13044
rect 4720 12964 4724 12996
rect 4756 12964 4760 12996
rect 4720 12916 4760 12964
rect 4720 12884 4724 12916
rect 4756 12884 4760 12916
rect 4720 12836 4760 12884
rect 4720 12804 4724 12836
rect 4756 12804 4760 12836
rect 4720 12756 4760 12804
rect 4720 12724 4724 12756
rect 4756 12724 4760 12756
rect 4720 12676 4760 12724
rect 4720 12644 4724 12676
rect 4756 12644 4760 12676
rect 4720 12596 4760 12644
rect 4720 12564 4724 12596
rect 4756 12564 4760 12596
rect 4720 12516 4760 12564
rect 4720 12484 4724 12516
rect 4756 12484 4760 12516
rect 4720 12436 4760 12484
rect 4720 12404 4724 12436
rect 4756 12404 4760 12436
rect 4720 12356 4760 12404
rect 4720 12324 4724 12356
rect 4756 12324 4760 12356
rect 4720 12276 4760 12324
rect 4720 12244 4724 12276
rect 4756 12244 4760 12276
rect 4720 12196 4760 12244
rect 4720 12164 4724 12196
rect 4756 12164 4760 12196
rect 4720 12116 4760 12164
rect 4720 12084 4724 12116
rect 4756 12084 4760 12116
rect 4720 12036 4760 12084
rect 4720 12004 4724 12036
rect 4756 12004 4760 12036
rect 4720 11956 4760 12004
rect 4720 11924 4724 11956
rect 4756 11924 4760 11956
rect 4720 11876 4760 11924
rect 4720 11844 4724 11876
rect 4756 11844 4760 11876
rect 4720 11796 4760 11844
rect 4720 11764 4724 11796
rect 4756 11764 4760 11796
rect 4720 11716 4760 11764
rect 4720 11684 4724 11716
rect 4756 11684 4760 11716
rect 4720 11636 4760 11684
rect 4720 11604 4724 11636
rect 4756 11604 4760 11636
rect 4720 11556 4760 11604
rect 4720 11524 4724 11556
rect 4756 11524 4760 11556
rect 4720 11476 4760 11524
rect 4720 11444 4724 11476
rect 4756 11444 4760 11476
rect 4720 11396 4760 11444
rect 4720 11364 4724 11396
rect 4756 11364 4760 11396
rect 4720 11316 4760 11364
rect 4720 11284 4724 11316
rect 4756 11284 4760 11316
rect 4720 11236 4760 11284
rect 4720 11204 4724 11236
rect 4756 11204 4760 11236
rect 4720 11156 4760 11204
rect 4720 11124 4724 11156
rect 4756 11124 4760 11156
rect 4720 11076 4760 11124
rect 4720 11044 4724 11076
rect 4756 11044 4760 11076
rect 4720 10996 4760 11044
rect 4720 10964 4724 10996
rect 4756 10964 4760 10996
rect 4720 10916 4760 10964
rect 4720 10884 4724 10916
rect 4756 10884 4760 10916
rect 4720 10836 4760 10884
rect 4720 10804 4724 10836
rect 4756 10804 4760 10836
rect 4720 10756 4760 10804
rect 4720 10724 4724 10756
rect 4756 10724 4760 10756
rect 4720 10676 4760 10724
rect 4720 10644 4724 10676
rect 4756 10644 4760 10676
rect 4720 10596 4760 10644
rect 4720 10564 4724 10596
rect 4756 10564 4760 10596
rect 4720 10516 4760 10564
rect 4720 10484 4724 10516
rect 4756 10484 4760 10516
rect 4720 10436 4760 10484
rect 4720 10404 4724 10436
rect 4756 10404 4760 10436
rect 4720 10356 4760 10404
rect 4720 10324 4724 10356
rect 4756 10324 4760 10356
rect 4720 10276 4760 10324
rect 4720 10244 4724 10276
rect 4756 10244 4760 10276
rect 4720 10196 4760 10244
rect 4720 10164 4724 10196
rect 4756 10164 4760 10196
rect 4720 10116 4760 10164
rect 4720 10084 4724 10116
rect 4756 10084 4760 10116
rect 4720 10036 4760 10084
rect 4720 10004 4724 10036
rect 4756 10004 4760 10036
rect 4720 9956 4760 10004
rect 4720 9924 4724 9956
rect 4756 9924 4760 9956
rect 4720 9876 4760 9924
rect 4720 9844 4724 9876
rect 4756 9844 4760 9876
rect 4720 9796 4760 9844
rect 4720 9764 4724 9796
rect 4756 9764 4760 9796
rect 4720 9716 4760 9764
rect 4720 9684 4724 9716
rect 4756 9684 4760 9716
rect 4720 9636 4760 9684
rect 4720 9604 4724 9636
rect 4756 9604 4760 9636
rect 4720 9556 4760 9604
rect 4720 9524 4724 9556
rect 4756 9524 4760 9556
rect 4720 9476 4760 9524
rect 4720 9444 4724 9476
rect 4756 9444 4760 9476
rect 4720 9396 4760 9444
rect 4720 9364 4724 9396
rect 4756 9364 4760 9396
rect 4720 9316 4760 9364
rect 4720 9284 4724 9316
rect 4756 9284 4760 9316
rect 4720 9236 4760 9284
rect 4720 9204 4724 9236
rect 4756 9204 4760 9236
rect 4720 9156 4760 9204
rect 4720 9124 4724 9156
rect 4756 9124 4760 9156
rect 4720 9076 4760 9124
rect 4720 9044 4724 9076
rect 4756 9044 4760 9076
rect 4720 8996 4760 9044
rect 4720 8964 4724 8996
rect 4756 8964 4760 8996
rect 4720 8916 4760 8964
rect 4720 8884 4724 8916
rect 4756 8884 4760 8916
rect 4720 8836 4760 8884
rect 4720 8804 4724 8836
rect 4756 8804 4760 8836
rect 4720 8756 4760 8804
rect 4720 8724 4724 8756
rect 4756 8724 4760 8756
rect 4720 8676 4760 8724
rect 4720 8644 4724 8676
rect 4756 8644 4760 8676
rect 4720 8596 4760 8644
rect 4720 8564 4724 8596
rect 4756 8564 4760 8596
rect 4720 8516 4760 8564
rect 4720 8484 4724 8516
rect 4756 8484 4760 8516
rect 4720 8436 4760 8484
rect 4720 8404 4724 8436
rect 4756 8404 4760 8436
rect 4720 8356 4760 8404
rect 4720 8324 4724 8356
rect 4756 8324 4760 8356
rect 4720 8276 4760 8324
rect 4720 8244 4724 8276
rect 4756 8244 4760 8276
rect 4720 8196 4760 8244
rect 4720 8164 4724 8196
rect 4756 8164 4760 8196
rect 4720 8116 4760 8164
rect 4720 8084 4724 8116
rect 4756 8084 4760 8116
rect 4720 8036 4760 8084
rect 4720 8004 4724 8036
rect 4756 8004 4760 8036
rect 4720 7956 4760 8004
rect 4720 7924 4724 7956
rect 4756 7924 4760 7956
rect 4720 7876 4760 7924
rect 4720 7844 4724 7876
rect 4756 7844 4760 7876
rect 4720 7796 4760 7844
rect 4720 7764 4724 7796
rect 4756 7764 4760 7796
rect 4720 7716 4760 7764
rect 4720 7684 4724 7716
rect 4756 7684 4760 7716
rect 4720 7636 4760 7684
rect 4720 7604 4724 7636
rect 4756 7604 4760 7636
rect 4720 7556 4760 7604
rect 4720 7524 4724 7556
rect 4756 7524 4760 7556
rect 4720 7476 4760 7524
rect 4720 7444 4724 7476
rect 4756 7444 4760 7476
rect 4720 7396 4760 7444
rect 4720 7364 4724 7396
rect 4756 7364 4760 7396
rect 4720 7316 4760 7364
rect 4720 7284 4724 7316
rect 4756 7284 4760 7316
rect 4720 7236 4760 7284
rect 4720 7204 4724 7236
rect 4756 7204 4760 7236
rect 4720 7156 4760 7204
rect 4720 7124 4724 7156
rect 4756 7124 4760 7156
rect 4720 7076 4760 7124
rect 4720 7044 4724 7076
rect 4756 7044 4760 7076
rect 4720 6996 4760 7044
rect 4720 6964 4724 6996
rect 4756 6964 4760 6996
rect 4720 6916 4760 6964
rect 4720 6884 4724 6916
rect 4756 6884 4760 6916
rect 4720 6836 4760 6884
rect 4720 6804 4724 6836
rect 4756 6804 4760 6836
rect 4720 6756 4760 6804
rect 4720 6724 4724 6756
rect 4756 6724 4760 6756
rect 4720 6676 4760 6724
rect 4720 6644 4724 6676
rect 4756 6644 4760 6676
rect 4720 6596 4760 6644
rect 4720 6564 4724 6596
rect 4756 6564 4760 6596
rect 4720 6516 4760 6564
rect 4720 6484 4724 6516
rect 4756 6484 4760 6516
rect 4720 6436 4760 6484
rect 4720 6404 4724 6436
rect 4756 6404 4760 6436
rect 4720 6356 4760 6404
rect 4720 6324 4724 6356
rect 4756 6324 4760 6356
rect 4720 6276 4760 6324
rect 4720 6244 4724 6276
rect 4756 6244 4760 6276
rect 4720 6196 4760 6244
rect 4720 6164 4724 6196
rect 4756 6164 4760 6196
rect 4720 6116 4760 6164
rect 4720 6084 4724 6116
rect 4756 6084 4760 6116
rect 4720 6036 4760 6084
rect 4720 6004 4724 6036
rect 4756 6004 4760 6036
rect 4720 5956 4760 6004
rect 4720 5924 4724 5956
rect 4756 5924 4760 5956
rect 4720 5876 4760 5924
rect 4720 5844 4724 5876
rect 4756 5844 4760 5876
rect 4720 5796 4760 5844
rect 4720 5764 4724 5796
rect 4756 5764 4760 5796
rect 4720 5716 4760 5764
rect 4720 5684 4724 5716
rect 4756 5684 4760 5716
rect 4720 5636 4760 5684
rect 4720 5604 4724 5636
rect 4756 5604 4760 5636
rect 4720 5556 4760 5604
rect 4720 5524 4724 5556
rect 4756 5524 4760 5556
rect 4720 5476 4760 5524
rect 4720 5444 4724 5476
rect 4756 5444 4760 5476
rect 4720 5396 4760 5444
rect 4720 5364 4724 5396
rect 4756 5364 4760 5396
rect 4720 5316 4760 5364
rect 4720 5284 4724 5316
rect 4756 5284 4760 5316
rect 4720 5236 4760 5284
rect 4720 5204 4724 5236
rect 4756 5204 4760 5236
rect 4720 5156 4760 5204
rect 4720 5124 4724 5156
rect 4756 5124 4760 5156
rect 4720 5076 4760 5124
rect 4720 5044 4724 5076
rect 4756 5044 4760 5076
rect 4720 4996 4760 5044
rect 4720 4964 4724 4996
rect 4756 4964 4760 4996
rect 4720 4916 4760 4964
rect 4720 4884 4724 4916
rect 4756 4884 4760 4916
rect 4720 4836 4760 4884
rect 4720 4804 4724 4836
rect 4756 4804 4760 4836
rect 4720 4756 4760 4804
rect 4720 4724 4724 4756
rect 4756 4724 4760 4756
rect 4720 4676 4760 4724
rect 4720 4644 4724 4676
rect 4756 4644 4760 4676
rect 4720 4596 4760 4644
rect 4720 4564 4724 4596
rect 4756 4564 4760 4596
rect 4720 4516 4760 4564
rect 4720 4484 4724 4516
rect 4756 4484 4760 4516
rect 4720 4436 4760 4484
rect 4720 4404 4724 4436
rect 4756 4404 4760 4436
rect 4720 4356 4760 4404
rect 4720 4324 4724 4356
rect 4756 4324 4760 4356
rect 4720 4276 4760 4324
rect 4720 4244 4724 4276
rect 4756 4244 4760 4276
rect 4720 4196 4760 4244
rect 4720 4164 4724 4196
rect 4756 4164 4760 4196
rect 4720 4116 4760 4164
rect 4720 4084 4724 4116
rect 4756 4084 4760 4116
rect 4720 4036 4760 4084
rect 4720 4004 4724 4036
rect 4756 4004 4760 4036
rect 4720 3956 4760 4004
rect 4720 3924 4724 3956
rect 4756 3924 4760 3956
rect 4720 3876 4760 3924
rect 4720 3844 4724 3876
rect 4756 3844 4760 3876
rect 4720 3796 4760 3844
rect 4720 3764 4724 3796
rect 4756 3764 4760 3796
rect 4720 3716 4760 3764
rect 4720 3684 4724 3716
rect 4756 3684 4760 3716
rect 4720 3636 4760 3684
rect 4720 3604 4724 3636
rect 4756 3604 4760 3636
rect 4720 3556 4760 3604
rect 4720 3524 4724 3556
rect 4756 3524 4760 3556
rect 4720 3476 4760 3524
rect 4720 3444 4724 3476
rect 4756 3444 4760 3476
rect 4720 3396 4760 3444
rect 4720 3364 4724 3396
rect 4756 3364 4760 3396
rect 4720 3316 4760 3364
rect 4720 3284 4724 3316
rect 4756 3284 4760 3316
rect 4720 3236 4760 3284
rect 4720 3204 4724 3236
rect 4756 3204 4760 3236
rect 4720 3156 4760 3204
rect 4720 3124 4724 3156
rect 4756 3124 4760 3156
rect 4720 3076 4760 3124
rect 4720 3044 4724 3076
rect 4756 3044 4760 3076
rect 4720 2996 4760 3044
rect 4720 2964 4724 2996
rect 4756 2964 4760 2996
rect 4720 2916 4760 2964
rect 4720 2884 4724 2916
rect 4756 2884 4760 2916
rect 4720 2836 4760 2884
rect 4720 2804 4724 2836
rect 4756 2804 4760 2836
rect 4720 2756 4760 2804
rect 4720 2724 4724 2756
rect 4756 2724 4760 2756
rect 4720 2676 4760 2724
rect 4720 2644 4724 2676
rect 4756 2644 4760 2676
rect 4720 2596 4760 2644
rect 4720 2564 4724 2596
rect 4756 2564 4760 2596
rect 4720 2516 4760 2564
rect 4720 2484 4724 2516
rect 4756 2484 4760 2516
rect 4720 2436 4760 2484
rect 4720 2404 4724 2436
rect 4756 2404 4760 2436
rect 4720 2356 4760 2404
rect 4720 2324 4724 2356
rect 4756 2324 4760 2356
rect 4720 2276 4760 2324
rect 4720 2244 4724 2276
rect 4756 2244 4760 2276
rect 4720 2196 4760 2244
rect 4720 2164 4724 2196
rect 4756 2164 4760 2196
rect 4720 2116 4760 2164
rect 4720 2084 4724 2116
rect 4756 2084 4760 2116
rect 4720 2036 4760 2084
rect 4720 2004 4724 2036
rect 4756 2004 4760 2036
rect 4720 1956 4760 2004
rect 4720 1924 4724 1956
rect 4756 1924 4760 1956
rect 4720 1876 4760 1924
rect 4720 1844 4724 1876
rect 4756 1844 4760 1876
rect 4720 1796 4760 1844
rect 4720 1764 4724 1796
rect 4756 1764 4760 1796
rect 4720 1716 4760 1764
rect 4720 1684 4724 1716
rect 4756 1684 4760 1716
rect 4720 1636 4760 1684
rect 4720 1604 4724 1636
rect 4756 1604 4760 1636
rect 4720 1556 4760 1604
rect 4720 1524 4724 1556
rect 4756 1524 4760 1556
rect 4720 1476 4760 1524
rect 4720 1444 4724 1476
rect 4756 1444 4760 1476
rect 4720 1396 4760 1444
rect 4720 1364 4724 1396
rect 4756 1364 4760 1396
rect 4720 1316 4760 1364
rect 4720 1284 4724 1316
rect 4756 1284 4760 1316
rect 4720 1236 4760 1284
rect 4720 1204 4724 1236
rect 4756 1204 4760 1236
rect 4720 1156 4760 1204
rect 4720 1124 4724 1156
rect 4756 1124 4760 1156
rect 4720 1076 4760 1124
rect 4720 1044 4724 1076
rect 4756 1044 4760 1076
rect 4720 996 4760 1044
rect 4720 964 4724 996
rect 4756 964 4760 996
rect 4720 916 4760 964
rect 4720 884 4724 916
rect 4756 884 4760 916
rect 4720 836 4760 884
rect 4720 804 4724 836
rect 4756 804 4760 836
rect 4720 756 4760 804
rect 4720 724 4724 756
rect 4756 724 4760 756
rect 4720 676 4760 724
rect 4720 644 4724 676
rect 4756 644 4760 676
rect 4720 596 4760 644
rect 4720 564 4724 596
rect 4756 564 4760 596
rect 4720 516 4760 564
rect 4720 484 4724 516
rect 4756 484 4760 516
rect 4720 436 4760 484
rect 4720 404 4724 436
rect 4756 404 4760 436
rect 4720 356 4760 404
rect 4720 324 4724 356
rect 4756 324 4760 356
rect 4720 276 4760 324
rect 4720 244 4724 276
rect 4756 244 4760 276
rect 4720 196 4760 244
rect 4720 164 4724 196
rect 4756 164 4760 196
rect 4720 116 4760 164
rect 4720 84 4724 116
rect 4756 84 4760 116
rect 4720 36 4760 84
rect 4720 4 4724 36
rect 4756 4 4760 36
rect 4720 -524 4760 4
rect 4800 6155 4840 15760
rect 4800 6125 4805 6155
rect 4835 6125 4840 6155
rect 4800 0 4840 6125
rect 4880 15716 4920 15760
rect 4880 15684 4884 15716
rect 4916 15684 4920 15716
rect 4880 15636 4920 15684
rect 4880 15604 4884 15636
rect 4916 15604 4920 15636
rect 4880 15556 4920 15604
rect 4880 15524 4884 15556
rect 4916 15524 4920 15556
rect 4880 15476 4920 15524
rect 4880 15444 4884 15476
rect 4916 15444 4920 15476
rect 4880 15396 4920 15444
rect 4880 15364 4884 15396
rect 4916 15364 4920 15396
rect 4880 15316 4920 15364
rect 4880 15284 4884 15316
rect 4916 15284 4920 15316
rect 4880 15236 4920 15284
rect 4880 15204 4884 15236
rect 4916 15204 4920 15236
rect 4880 15156 4920 15204
rect 4880 15124 4884 15156
rect 4916 15124 4920 15156
rect 4880 15076 4920 15124
rect 4880 15044 4884 15076
rect 4916 15044 4920 15076
rect 4880 14996 4920 15044
rect 4880 14964 4884 14996
rect 4916 14964 4920 14996
rect 4880 14916 4920 14964
rect 4880 14884 4884 14916
rect 4916 14884 4920 14916
rect 4880 14836 4920 14884
rect 4880 14804 4884 14836
rect 4916 14804 4920 14836
rect 4880 14756 4920 14804
rect 4880 14724 4884 14756
rect 4916 14724 4920 14756
rect 4880 14676 4920 14724
rect 4880 14644 4884 14676
rect 4916 14644 4920 14676
rect 4880 14596 4920 14644
rect 4880 14564 4884 14596
rect 4916 14564 4920 14596
rect 4880 14516 4920 14564
rect 4880 14484 4884 14516
rect 4916 14484 4920 14516
rect 4880 14436 4920 14484
rect 4880 14404 4884 14436
rect 4916 14404 4920 14436
rect 4880 14356 4920 14404
rect 4880 14324 4884 14356
rect 4916 14324 4920 14356
rect 4880 14276 4920 14324
rect 4880 14244 4884 14276
rect 4916 14244 4920 14276
rect 4880 14196 4920 14244
rect 4880 14164 4884 14196
rect 4916 14164 4920 14196
rect 4880 14116 4920 14164
rect 4880 14084 4884 14116
rect 4916 14084 4920 14116
rect 4880 14036 4920 14084
rect 4880 14004 4884 14036
rect 4916 14004 4920 14036
rect 4880 13956 4920 14004
rect 4880 13924 4884 13956
rect 4916 13924 4920 13956
rect 4880 13876 4920 13924
rect 4880 13844 4884 13876
rect 4916 13844 4920 13876
rect 4880 13796 4920 13844
rect 4880 13764 4884 13796
rect 4916 13764 4920 13796
rect 4880 13716 4920 13764
rect 4880 13684 4884 13716
rect 4916 13684 4920 13716
rect 4880 13636 4920 13684
rect 4880 13604 4884 13636
rect 4916 13604 4920 13636
rect 4880 13556 4920 13604
rect 4880 13524 4884 13556
rect 4916 13524 4920 13556
rect 4880 13476 4920 13524
rect 4880 13444 4884 13476
rect 4916 13444 4920 13476
rect 4880 13396 4920 13444
rect 4880 13364 4884 13396
rect 4916 13364 4920 13396
rect 4880 13316 4920 13364
rect 4880 13284 4884 13316
rect 4916 13284 4920 13316
rect 4880 13236 4920 13284
rect 4880 13204 4884 13236
rect 4916 13204 4920 13236
rect 4880 13156 4920 13204
rect 4880 13124 4884 13156
rect 4916 13124 4920 13156
rect 4880 13076 4920 13124
rect 4880 13044 4884 13076
rect 4916 13044 4920 13076
rect 4880 12996 4920 13044
rect 4880 12964 4884 12996
rect 4916 12964 4920 12996
rect 4880 12916 4920 12964
rect 4880 12884 4884 12916
rect 4916 12884 4920 12916
rect 4880 12836 4920 12884
rect 4880 12804 4884 12836
rect 4916 12804 4920 12836
rect 4880 12756 4920 12804
rect 4880 12724 4884 12756
rect 4916 12724 4920 12756
rect 4880 12676 4920 12724
rect 4880 12644 4884 12676
rect 4916 12644 4920 12676
rect 4880 12596 4920 12644
rect 4880 12564 4884 12596
rect 4916 12564 4920 12596
rect 4880 12516 4920 12564
rect 4880 12484 4884 12516
rect 4916 12484 4920 12516
rect 4880 12436 4920 12484
rect 4880 12404 4884 12436
rect 4916 12404 4920 12436
rect 4880 12356 4920 12404
rect 4880 12324 4884 12356
rect 4916 12324 4920 12356
rect 4880 12276 4920 12324
rect 4880 12244 4884 12276
rect 4916 12244 4920 12276
rect 4880 12196 4920 12244
rect 4880 12164 4884 12196
rect 4916 12164 4920 12196
rect 4880 12116 4920 12164
rect 4880 12084 4884 12116
rect 4916 12084 4920 12116
rect 4880 12036 4920 12084
rect 4880 12004 4884 12036
rect 4916 12004 4920 12036
rect 4880 11956 4920 12004
rect 4880 11924 4884 11956
rect 4916 11924 4920 11956
rect 4880 11876 4920 11924
rect 4880 11844 4884 11876
rect 4916 11844 4920 11876
rect 4880 11796 4920 11844
rect 4880 11764 4884 11796
rect 4916 11764 4920 11796
rect 4880 11716 4920 11764
rect 4880 11684 4884 11716
rect 4916 11684 4920 11716
rect 4880 11636 4920 11684
rect 4880 11604 4884 11636
rect 4916 11604 4920 11636
rect 4880 11556 4920 11604
rect 4880 11524 4884 11556
rect 4916 11524 4920 11556
rect 4880 11476 4920 11524
rect 4880 11444 4884 11476
rect 4916 11444 4920 11476
rect 4880 11396 4920 11444
rect 4880 11364 4884 11396
rect 4916 11364 4920 11396
rect 4880 11316 4920 11364
rect 4880 11284 4884 11316
rect 4916 11284 4920 11316
rect 4880 11236 4920 11284
rect 4880 11204 4884 11236
rect 4916 11204 4920 11236
rect 4880 11156 4920 11204
rect 4880 11124 4884 11156
rect 4916 11124 4920 11156
rect 4880 11076 4920 11124
rect 4880 11044 4884 11076
rect 4916 11044 4920 11076
rect 4880 10996 4920 11044
rect 4880 10964 4884 10996
rect 4916 10964 4920 10996
rect 4880 10916 4920 10964
rect 4880 10884 4884 10916
rect 4916 10884 4920 10916
rect 4880 10836 4920 10884
rect 4880 10804 4884 10836
rect 4916 10804 4920 10836
rect 4880 10756 4920 10804
rect 4880 10724 4884 10756
rect 4916 10724 4920 10756
rect 4880 10676 4920 10724
rect 4880 10644 4884 10676
rect 4916 10644 4920 10676
rect 4880 10596 4920 10644
rect 4880 10564 4884 10596
rect 4916 10564 4920 10596
rect 4880 10516 4920 10564
rect 4880 10484 4884 10516
rect 4916 10484 4920 10516
rect 4880 10436 4920 10484
rect 4880 10404 4884 10436
rect 4916 10404 4920 10436
rect 4880 10356 4920 10404
rect 4880 10324 4884 10356
rect 4916 10324 4920 10356
rect 4880 10276 4920 10324
rect 4880 10244 4884 10276
rect 4916 10244 4920 10276
rect 4880 10196 4920 10244
rect 4880 10164 4884 10196
rect 4916 10164 4920 10196
rect 4880 10116 4920 10164
rect 4880 10084 4884 10116
rect 4916 10084 4920 10116
rect 4880 10036 4920 10084
rect 4880 10004 4884 10036
rect 4916 10004 4920 10036
rect 4880 9956 4920 10004
rect 4880 9924 4884 9956
rect 4916 9924 4920 9956
rect 4880 9876 4920 9924
rect 4880 9844 4884 9876
rect 4916 9844 4920 9876
rect 4880 9796 4920 9844
rect 4880 9764 4884 9796
rect 4916 9764 4920 9796
rect 4880 9716 4920 9764
rect 4880 9684 4884 9716
rect 4916 9684 4920 9716
rect 4880 9636 4920 9684
rect 4880 9604 4884 9636
rect 4916 9604 4920 9636
rect 4880 9556 4920 9604
rect 4880 9524 4884 9556
rect 4916 9524 4920 9556
rect 4880 9476 4920 9524
rect 4880 9444 4884 9476
rect 4916 9444 4920 9476
rect 4880 9396 4920 9444
rect 4880 9364 4884 9396
rect 4916 9364 4920 9396
rect 4880 9316 4920 9364
rect 4880 9284 4884 9316
rect 4916 9284 4920 9316
rect 4880 9236 4920 9284
rect 4880 9204 4884 9236
rect 4916 9204 4920 9236
rect 4880 9156 4920 9204
rect 4880 9124 4884 9156
rect 4916 9124 4920 9156
rect 4880 9076 4920 9124
rect 4880 9044 4884 9076
rect 4916 9044 4920 9076
rect 4880 8996 4920 9044
rect 4880 8964 4884 8996
rect 4916 8964 4920 8996
rect 4880 8916 4920 8964
rect 4880 8884 4884 8916
rect 4916 8884 4920 8916
rect 4880 8836 4920 8884
rect 4880 8804 4884 8836
rect 4916 8804 4920 8836
rect 4880 8756 4920 8804
rect 4880 8724 4884 8756
rect 4916 8724 4920 8756
rect 4880 8676 4920 8724
rect 4880 8644 4884 8676
rect 4916 8644 4920 8676
rect 4880 8596 4920 8644
rect 4880 8564 4884 8596
rect 4916 8564 4920 8596
rect 4880 8516 4920 8564
rect 4880 8484 4884 8516
rect 4916 8484 4920 8516
rect 4880 8436 4920 8484
rect 4880 8404 4884 8436
rect 4916 8404 4920 8436
rect 4880 8356 4920 8404
rect 4880 8324 4884 8356
rect 4916 8324 4920 8356
rect 4880 8276 4920 8324
rect 4880 8244 4884 8276
rect 4916 8244 4920 8276
rect 4880 8196 4920 8244
rect 4880 8164 4884 8196
rect 4916 8164 4920 8196
rect 4880 8116 4920 8164
rect 4880 8084 4884 8116
rect 4916 8084 4920 8116
rect 4880 8036 4920 8084
rect 4880 8004 4884 8036
rect 4916 8004 4920 8036
rect 4880 7956 4920 8004
rect 4880 7924 4884 7956
rect 4916 7924 4920 7956
rect 4880 7876 4920 7924
rect 4880 7844 4884 7876
rect 4916 7844 4920 7876
rect 4880 7796 4920 7844
rect 4880 7764 4884 7796
rect 4916 7764 4920 7796
rect 4880 7716 4920 7764
rect 4880 7684 4884 7716
rect 4916 7684 4920 7716
rect 4880 7636 4920 7684
rect 4880 7604 4884 7636
rect 4916 7604 4920 7636
rect 4880 7556 4920 7604
rect 4880 7524 4884 7556
rect 4916 7524 4920 7556
rect 4880 7476 4920 7524
rect 4880 7444 4884 7476
rect 4916 7444 4920 7476
rect 4880 7396 4920 7444
rect 4880 7364 4884 7396
rect 4916 7364 4920 7396
rect 4880 7316 4920 7364
rect 4880 7284 4884 7316
rect 4916 7284 4920 7316
rect 4880 7236 4920 7284
rect 4880 7204 4884 7236
rect 4916 7204 4920 7236
rect 4880 7156 4920 7204
rect 4880 7124 4884 7156
rect 4916 7124 4920 7156
rect 4880 7076 4920 7124
rect 4880 7044 4884 7076
rect 4916 7044 4920 7076
rect 4880 6996 4920 7044
rect 4880 6964 4884 6996
rect 4916 6964 4920 6996
rect 4880 6916 4920 6964
rect 4880 6884 4884 6916
rect 4916 6884 4920 6916
rect 4880 6836 4920 6884
rect 4880 6804 4884 6836
rect 4916 6804 4920 6836
rect 4880 6756 4920 6804
rect 4880 6724 4884 6756
rect 4916 6724 4920 6756
rect 4880 6676 4920 6724
rect 4880 6644 4884 6676
rect 4916 6644 4920 6676
rect 4880 6596 4920 6644
rect 4880 6564 4884 6596
rect 4916 6564 4920 6596
rect 4880 6516 4920 6564
rect 4880 6484 4884 6516
rect 4916 6484 4920 6516
rect 4880 6436 4920 6484
rect 4880 6404 4884 6436
rect 4916 6404 4920 6436
rect 4880 6356 4920 6404
rect 4880 6324 4884 6356
rect 4916 6324 4920 6356
rect 4880 6276 4920 6324
rect 4880 6244 4884 6276
rect 4916 6244 4920 6276
rect 4880 6196 4920 6244
rect 4880 6164 4884 6196
rect 4916 6164 4920 6196
rect 4880 6116 4920 6164
rect 4880 6084 4884 6116
rect 4916 6084 4920 6116
rect 4880 6036 4920 6084
rect 4880 6004 4884 6036
rect 4916 6004 4920 6036
rect 4880 5956 4920 6004
rect 4880 5924 4884 5956
rect 4916 5924 4920 5956
rect 4880 5876 4920 5924
rect 4880 5844 4884 5876
rect 4916 5844 4920 5876
rect 4880 5796 4920 5844
rect 4880 5764 4884 5796
rect 4916 5764 4920 5796
rect 4880 5716 4920 5764
rect 4880 5684 4884 5716
rect 4916 5684 4920 5716
rect 4880 5636 4920 5684
rect 4880 5604 4884 5636
rect 4916 5604 4920 5636
rect 4880 5556 4920 5604
rect 4880 5524 4884 5556
rect 4916 5524 4920 5556
rect 4880 5476 4920 5524
rect 4880 5444 4884 5476
rect 4916 5444 4920 5476
rect 4880 5396 4920 5444
rect 4880 5364 4884 5396
rect 4916 5364 4920 5396
rect 4880 5316 4920 5364
rect 4880 5284 4884 5316
rect 4916 5284 4920 5316
rect 4880 5236 4920 5284
rect 4880 5204 4884 5236
rect 4916 5204 4920 5236
rect 4880 5156 4920 5204
rect 4880 5124 4884 5156
rect 4916 5124 4920 5156
rect 4880 5076 4920 5124
rect 4880 5044 4884 5076
rect 4916 5044 4920 5076
rect 4880 4996 4920 5044
rect 4880 4964 4884 4996
rect 4916 4964 4920 4996
rect 4880 4916 4920 4964
rect 4880 4884 4884 4916
rect 4916 4884 4920 4916
rect 4880 4836 4920 4884
rect 4880 4804 4884 4836
rect 4916 4804 4920 4836
rect 4880 4756 4920 4804
rect 4880 4724 4884 4756
rect 4916 4724 4920 4756
rect 4880 4676 4920 4724
rect 4880 4644 4884 4676
rect 4916 4644 4920 4676
rect 4880 4596 4920 4644
rect 4880 4564 4884 4596
rect 4916 4564 4920 4596
rect 4880 4516 4920 4564
rect 4880 4484 4884 4516
rect 4916 4484 4920 4516
rect 4880 4436 4920 4484
rect 4880 4404 4884 4436
rect 4916 4404 4920 4436
rect 4880 4356 4920 4404
rect 4880 4324 4884 4356
rect 4916 4324 4920 4356
rect 4880 4276 4920 4324
rect 4880 4244 4884 4276
rect 4916 4244 4920 4276
rect 4880 4196 4920 4244
rect 4880 4164 4884 4196
rect 4916 4164 4920 4196
rect 4880 4116 4920 4164
rect 4880 4084 4884 4116
rect 4916 4084 4920 4116
rect 4880 4036 4920 4084
rect 4880 4004 4884 4036
rect 4916 4004 4920 4036
rect 4880 3956 4920 4004
rect 4880 3924 4884 3956
rect 4916 3924 4920 3956
rect 4880 3876 4920 3924
rect 4880 3844 4884 3876
rect 4916 3844 4920 3876
rect 4880 3796 4920 3844
rect 4880 3764 4884 3796
rect 4916 3764 4920 3796
rect 4880 3716 4920 3764
rect 4880 3684 4884 3716
rect 4916 3684 4920 3716
rect 4880 3636 4920 3684
rect 4880 3604 4884 3636
rect 4916 3604 4920 3636
rect 4880 3556 4920 3604
rect 4880 3524 4884 3556
rect 4916 3524 4920 3556
rect 4880 3476 4920 3524
rect 4880 3444 4884 3476
rect 4916 3444 4920 3476
rect 4880 3396 4920 3444
rect 4880 3364 4884 3396
rect 4916 3364 4920 3396
rect 4880 3316 4920 3364
rect 4880 3284 4884 3316
rect 4916 3284 4920 3316
rect 4880 3236 4920 3284
rect 4880 3204 4884 3236
rect 4916 3204 4920 3236
rect 4880 3156 4920 3204
rect 4880 3124 4884 3156
rect 4916 3124 4920 3156
rect 4880 3076 4920 3124
rect 4880 3044 4884 3076
rect 4916 3044 4920 3076
rect 4880 2996 4920 3044
rect 4880 2964 4884 2996
rect 4916 2964 4920 2996
rect 4880 2916 4920 2964
rect 4880 2884 4884 2916
rect 4916 2884 4920 2916
rect 4880 2836 4920 2884
rect 4880 2804 4884 2836
rect 4916 2804 4920 2836
rect 4880 2756 4920 2804
rect 4880 2724 4884 2756
rect 4916 2724 4920 2756
rect 4880 2676 4920 2724
rect 4880 2644 4884 2676
rect 4916 2644 4920 2676
rect 4880 2596 4920 2644
rect 4880 2564 4884 2596
rect 4916 2564 4920 2596
rect 4880 2516 4920 2564
rect 4880 2484 4884 2516
rect 4916 2484 4920 2516
rect 4880 2436 4920 2484
rect 4880 2404 4884 2436
rect 4916 2404 4920 2436
rect 4880 2356 4920 2404
rect 4880 2324 4884 2356
rect 4916 2324 4920 2356
rect 4880 2276 4920 2324
rect 4880 2244 4884 2276
rect 4916 2244 4920 2276
rect 4880 2196 4920 2244
rect 4880 2164 4884 2196
rect 4916 2164 4920 2196
rect 4880 2116 4920 2164
rect 4880 2084 4884 2116
rect 4916 2084 4920 2116
rect 4880 2036 4920 2084
rect 4880 2004 4884 2036
rect 4916 2004 4920 2036
rect 4880 1956 4920 2004
rect 4880 1924 4884 1956
rect 4916 1924 4920 1956
rect 4880 1876 4920 1924
rect 4880 1844 4884 1876
rect 4916 1844 4920 1876
rect 4880 1796 4920 1844
rect 4880 1764 4884 1796
rect 4916 1764 4920 1796
rect 4880 1716 4920 1764
rect 4880 1684 4884 1716
rect 4916 1684 4920 1716
rect 4880 1636 4920 1684
rect 4880 1604 4884 1636
rect 4916 1604 4920 1636
rect 4880 1556 4920 1604
rect 4880 1524 4884 1556
rect 4916 1524 4920 1556
rect 4880 1476 4920 1524
rect 4880 1444 4884 1476
rect 4916 1444 4920 1476
rect 4880 1396 4920 1444
rect 4880 1364 4884 1396
rect 4916 1364 4920 1396
rect 4880 1316 4920 1364
rect 4880 1284 4884 1316
rect 4916 1284 4920 1316
rect 4880 1236 4920 1284
rect 4880 1204 4884 1236
rect 4916 1204 4920 1236
rect 4880 1156 4920 1204
rect 4880 1124 4884 1156
rect 4916 1124 4920 1156
rect 4880 1076 4920 1124
rect 4880 1044 4884 1076
rect 4916 1044 4920 1076
rect 4880 996 4920 1044
rect 4880 964 4884 996
rect 4916 964 4920 996
rect 4880 916 4920 964
rect 4880 884 4884 916
rect 4916 884 4920 916
rect 4880 836 4920 884
rect 4880 804 4884 836
rect 4916 804 4920 836
rect 4880 756 4920 804
rect 4880 724 4884 756
rect 4916 724 4920 756
rect 4880 676 4920 724
rect 4880 644 4884 676
rect 4916 644 4920 676
rect 4880 596 4920 644
rect 4880 564 4884 596
rect 4916 564 4920 596
rect 4880 516 4920 564
rect 4880 484 4884 516
rect 4916 484 4920 516
rect 4880 436 4920 484
rect 4880 404 4884 436
rect 4916 404 4920 436
rect 4880 356 4920 404
rect 4880 324 4884 356
rect 4916 324 4920 356
rect 4880 276 4920 324
rect 4880 244 4884 276
rect 4916 244 4920 276
rect 4880 196 4920 244
rect 4880 164 4884 196
rect 4916 164 4920 196
rect 4880 116 4920 164
rect 4880 84 4884 116
rect 4916 84 4920 116
rect 4880 36 4920 84
rect 4880 4 4884 36
rect 4916 4 4920 36
rect 4720 -716 4724 -524
rect 4756 -716 4760 -524
rect 4720 -960 4760 -716
rect 4880 -524 4920 4
rect 4960 14155 5000 15760
rect 4960 14125 4965 14155
rect 4995 14125 5000 14155
rect 4960 9115 5000 14125
rect 4960 9085 4965 9115
rect 4995 9085 5000 9115
rect 4960 5995 5000 9085
rect 4960 5965 4965 5995
rect 4995 5965 5000 5995
rect 4960 0 5000 5965
rect 5040 15716 5080 15760
rect 5040 15684 5044 15716
rect 5076 15684 5080 15716
rect 5040 15636 5080 15684
rect 5040 15604 5044 15636
rect 5076 15604 5080 15636
rect 5040 15556 5080 15604
rect 5040 15524 5044 15556
rect 5076 15524 5080 15556
rect 5040 15476 5080 15524
rect 5040 15444 5044 15476
rect 5076 15444 5080 15476
rect 5040 15396 5080 15444
rect 5040 15364 5044 15396
rect 5076 15364 5080 15396
rect 5040 15316 5080 15364
rect 5040 15284 5044 15316
rect 5076 15284 5080 15316
rect 5040 15236 5080 15284
rect 5040 15204 5044 15236
rect 5076 15204 5080 15236
rect 5040 15156 5080 15204
rect 5040 15124 5044 15156
rect 5076 15124 5080 15156
rect 5040 15076 5080 15124
rect 5040 15044 5044 15076
rect 5076 15044 5080 15076
rect 5040 14996 5080 15044
rect 5040 14964 5044 14996
rect 5076 14964 5080 14996
rect 5040 14916 5080 14964
rect 5040 14884 5044 14916
rect 5076 14884 5080 14916
rect 5040 14836 5080 14884
rect 5040 14804 5044 14836
rect 5076 14804 5080 14836
rect 5040 14756 5080 14804
rect 5040 14724 5044 14756
rect 5076 14724 5080 14756
rect 5040 14676 5080 14724
rect 5040 14644 5044 14676
rect 5076 14644 5080 14676
rect 5040 14596 5080 14644
rect 5040 14564 5044 14596
rect 5076 14564 5080 14596
rect 5040 14516 5080 14564
rect 5040 14484 5044 14516
rect 5076 14484 5080 14516
rect 5040 14436 5080 14484
rect 5040 14404 5044 14436
rect 5076 14404 5080 14436
rect 5040 14356 5080 14404
rect 5040 14324 5044 14356
rect 5076 14324 5080 14356
rect 5040 14276 5080 14324
rect 5040 14244 5044 14276
rect 5076 14244 5080 14276
rect 5040 14196 5080 14244
rect 5040 14164 5044 14196
rect 5076 14164 5080 14196
rect 5040 14116 5080 14164
rect 5040 14084 5044 14116
rect 5076 14084 5080 14116
rect 5040 14036 5080 14084
rect 5040 14004 5044 14036
rect 5076 14004 5080 14036
rect 5040 13956 5080 14004
rect 5040 13924 5044 13956
rect 5076 13924 5080 13956
rect 5040 13876 5080 13924
rect 5040 13844 5044 13876
rect 5076 13844 5080 13876
rect 5040 13796 5080 13844
rect 5040 13764 5044 13796
rect 5076 13764 5080 13796
rect 5040 13716 5080 13764
rect 5040 13684 5044 13716
rect 5076 13684 5080 13716
rect 5040 13636 5080 13684
rect 5040 13604 5044 13636
rect 5076 13604 5080 13636
rect 5040 13556 5080 13604
rect 5040 13524 5044 13556
rect 5076 13524 5080 13556
rect 5040 13476 5080 13524
rect 5040 13444 5044 13476
rect 5076 13444 5080 13476
rect 5040 13396 5080 13444
rect 5040 13364 5044 13396
rect 5076 13364 5080 13396
rect 5040 13316 5080 13364
rect 5040 13284 5044 13316
rect 5076 13284 5080 13316
rect 5040 13236 5080 13284
rect 5040 13204 5044 13236
rect 5076 13204 5080 13236
rect 5040 13156 5080 13204
rect 5040 13124 5044 13156
rect 5076 13124 5080 13156
rect 5040 13076 5080 13124
rect 5040 13044 5044 13076
rect 5076 13044 5080 13076
rect 5040 12996 5080 13044
rect 5040 12964 5044 12996
rect 5076 12964 5080 12996
rect 5040 12916 5080 12964
rect 5040 12884 5044 12916
rect 5076 12884 5080 12916
rect 5040 12836 5080 12884
rect 5040 12804 5044 12836
rect 5076 12804 5080 12836
rect 5040 12756 5080 12804
rect 5040 12724 5044 12756
rect 5076 12724 5080 12756
rect 5040 12676 5080 12724
rect 5040 12644 5044 12676
rect 5076 12644 5080 12676
rect 5040 12596 5080 12644
rect 5040 12564 5044 12596
rect 5076 12564 5080 12596
rect 5040 12516 5080 12564
rect 5040 12484 5044 12516
rect 5076 12484 5080 12516
rect 5040 12436 5080 12484
rect 5040 12404 5044 12436
rect 5076 12404 5080 12436
rect 5040 12356 5080 12404
rect 5040 12324 5044 12356
rect 5076 12324 5080 12356
rect 5040 12276 5080 12324
rect 5040 12244 5044 12276
rect 5076 12244 5080 12276
rect 5040 12196 5080 12244
rect 5040 12164 5044 12196
rect 5076 12164 5080 12196
rect 5040 12116 5080 12164
rect 5040 12084 5044 12116
rect 5076 12084 5080 12116
rect 5040 12036 5080 12084
rect 5040 12004 5044 12036
rect 5076 12004 5080 12036
rect 5040 11956 5080 12004
rect 5040 11924 5044 11956
rect 5076 11924 5080 11956
rect 5040 11876 5080 11924
rect 5040 11844 5044 11876
rect 5076 11844 5080 11876
rect 5040 11796 5080 11844
rect 5040 11764 5044 11796
rect 5076 11764 5080 11796
rect 5040 11716 5080 11764
rect 5040 11684 5044 11716
rect 5076 11684 5080 11716
rect 5040 11636 5080 11684
rect 5040 11604 5044 11636
rect 5076 11604 5080 11636
rect 5040 11556 5080 11604
rect 5040 11524 5044 11556
rect 5076 11524 5080 11556
rect 5040 11476 5080 11524
rect 5040 11444 5044 11476
rect 5076 11444 5080 11476
rect 5040 11396 5080 11444
rect 5040 11364 5044 11396
rect 5076 11364 5080 11396
rect 5040 11316 5080 11364
rect 5040 11284 5044 11316
rect 5076 11284 5080 11316
rect 5040 11236 5080 11284
rect 5040 11204 5044 11236
rect 5076 11204 5080 11236
rect 5040 11156 5080 11204
rect 5040 11124 5044 11156
rect 5076 11124 5080 11156
rect 5040 11076 5080 11124
rect 5040 11044 5044 11076
rect 5076 11044 5080 11076
rect 5040 10996 5080 11044
rect 5040 10964 5044 10996
rect 5076 10964 5080 10996
rect 5040 10916 5080 10964
rect 5040 10884 5044 10916
rect 5076 10884 5080 10916
rect 5040 10836 5080 10884
rect 5040 10804 5044 10836
rect 5076 10804 5080 10836
rect 5040 10756 5080 10804
rect 5040 10724 5044 10756
rect 5076 10724 5080 10756
rect 5040 10676 5080 10724
rect 5040 10644 5044 10676
rect 5076 10644 5080 10676
rect 5040 10596 5080 10644
rect 5040 10564 5044 10596
rect 5076 10564 5080 10596
rect 5040 10516 5080 10564
rect 5040 10484 5044 10516
rect 5076 10484 5080 10516
rect 5040 10436 5080 10484
rect 5040 10404 5044 10436
rect 5076 10404 5080 10436
rect 5040 10356 5080 10404
rect 5040 10324 5044 10356
rect 5076 10324 5080 10356
rect 5040 10276 5080 10324
rect 5040 10244 5044 10276
rect 5076 10244 5080 10276
rect 5040 10196 5080 10244
rect 5040 10164 5044 10196
rect 5076 10164 5080 10196
rect 5040 10116 5080 10164
rect 5040 10084 5044 10116
rect 5076 10084 5080 10116
rect 5040 10036 5080 10084
rect 5040 10004 5044 10036
rect 5076 10004 5080 10036
rect 5040 9956 5080 10004
rect 5040 9924 5044 9956
rect 5076 9924 5080 9956
rect 5040 9876 5080 9924
rect 5040 9844 5044 9876
rect 5076 9844 5080 9876
rect 5040 9796 5080 9844
rect 5040 9764 5044 9796
rect 5076 9764 5080 9796
rect 5040 9716 5080 9764
rect 5040 9684 5044 9716
rect 5076 9684 5080 9716
rect 5040 9636 5080 9684
rect 5040 9604 5044 9636
rect 5076 9604 5080 9636
rect 5040 9556 5080 9604
rect 5040 9524 5044 9556
rect 5076 9524 5080 9556
rect 5040 9476 5080 9524
rect 5040 9444 5044 9476
rect 5076 9444 5080 9476
rect 5040 9396 5080 9444
rect 5040 9364 5044 9396
rect 5076 9364 5080 9396
rect 5040 9316 5080 9364
rect 5040 9284 5044 9316
rect 5076 9284 5080 9316
rect 5040 9236 5080 9284
rect 5040 9204 5044 9236
rect 5076 9204 5080 9236
rect 5040 9156 5080 9204
rect 5040 9124 5044 9156
rect 5076 9124 5080 9156
rect 5040 9076 5080 9124
rect 5040 9044 5044 9076
rect 5076 9044 5080 9076
rect 5040 8996 5080 9044
rect 5040 8964 5044 8996
rect 5076 8964 5080 8996
rect 5040 8916 5080 8964
rect 5040 8884 5044 8916
rect 5076 8884 5080 8916
rect 5040 8836 5080 8884
rect 5040 8804 5044 8836
rect 5076 8804 5080 8836
rect 5040 8756 5080 8804
rect 5040 8724 5044 8756
rect 5076 8724 5080 8756
rect 5040 8676 5080 8724
rect 5040 8644 5044 8676
rect 5076 8644 5080 8676
rect 5040 8596 5080 8644
rect 5040 8564 5044 8596
rect 5076 8564 5080 8596
rect 5040 8516 5080 8564
rect 5040 8484 5044 8516
rect 5076 8484 5080 8516
rect 5040 8436 5080 8484
rect 5040 8404 5044 8436
rect 5076 8404 5080 8436
rect 5040 8356 5080 8404
rect 5040 8324 5044 8356
rect 5076 8324 5080 8356
rect 5040 8276 5080 8324
rect 5040 8244 5044 8276
rect 5076 8244 5080 8276
rect 5040 8196 5080 8244
rect 5040 8164 5044 8196
rect 5076 8164 5080 8196
rect 5040 8116 5080 8164
rect 5040 8084 5044 8116
rect 5076 8084 5080 8116
rect 5040 8036 5080 8084
rect 5040 8004 5044 8036
rect 5076 8004 5080 8036
rect 5040 7956 5080 8004
rect 5040 7924 5044 7956
rect 5076 7924 5080 7956
rect 5040 7876 5080 7924
rect 5040 7844 5044 7876
rect 5076 7844 5080 7876
rect 5040 7796 5080 7844
rect 5040 7764 5044 7796
rect 5076 7764 5080 7796
rect 5040 7716 5080 7764
rect 5040 7684 5044 7716
rect 5076 7684 5080 7716
rect 5040 7636 5080 7684
rect 5040 7604 5044 7636
rect 5076 7604 5080 7636
rect 5040 7556 5080 7604
rect 5040 7524 5044 7556
rect 5076 7524 5080 7556
rect 5040 7476 5080 7524
rect 5040 7444 5044 7476
rect 5076 7444 5080 7476
rect 5040 7396 5080 7444
rect 5040 7364 5044 7396
rect 5076 7364 5080 7396
rect 5040 7316 5080 7364
rect 5040 7284 5044 7316
rect 5076 7284 5080 7316
rect 5040 7236 5080 7284
rect 5040 7204 5044 7236
rect 5076 7204 5080 7236
rect 5040 7156 5080 7204
rect 5040 7124 5044 7156
rect 5076 7124 5080 7156
rect 5040 7076 5080 7124
rect 5040 7044 5044 7076
rect 5076 7044 5080 7076
rect 5040 6996 5080 7044
rect 5040 6964 5044 6996
rect 5076 6964 5080 6996
rect 5040 6916 5080 6964
rect 5040 6884 5044 6916
rect 5076 6884 5080 6916
rect 5040 6836 5080 6884
rect 5040 6804 5044 6836
rect 5076 6804 5080 6836
rect 5040 6756 5080 6804
rect 5040 6724 5044 6756
rect 5076 6724 5080 6756
rect 5040 6676 5080 6724
rect 5040 6644 5044 6676
rect 5076 6644 5080 6676
rect 5040 6596 5080 6644
rect 5040 6564 5044 6596
rect 5076 6564 5080 6596
rect 5040 6516 5080 6564
rect 5040 6484 5044 6516
rect 5076 6484 5080 6516
rect 5040 6436 5080 6484
rect 5040 6404 5044 6436
rect 5076 6404 5080 6436
rect 5040 6356 5080 6404
rect 5040 6324 5044 6356
rect 5076 6324 5080 6356
rect 5040 6276 5080 6324
rect 5040 6244 5044 6276
rect 5076 6244 5080 6276
rect 5040 6196 5080 6244
rect 5040 6164 5044 6196
rect 5076 6164 5080 6196
rect 5040 6116 5080 6164
rect 5040 6084 5044 6116
rect 5076 6084 5080 6116
rect 5040 6036 5080 6084
rect 5040 6004 5044 6036
rect 5076 6004 5080 6036
rect 5040 5956 5080 6004
rect 5040 5924 5044 5956
rect 5076 5924 5080 5956
rect 5040 5876 5080 5924
rect 5040 5844 5044 5876
rect 5076 5844 5080 5876
rect 5040 5796 5080 5844
rect 5040 5764 5044 5796
rect 5076 5764 5080 5796
rect 5040 5716 5080 5764
rect 5040 5684 5044 5716
rect 5076 5684 5080 5716
rect 5040 5636 5080 5684
rect 5040 5604 5044 5636
rect 5076 5604 5080 5636
rect 5040 5556 5080 5604
rect 5040 5524 5044 5556
rect 5076 5524 5080 5556
rect 5040 5476 5080 5524
rect 5040 5444 5044 5476
rect 5076 5444 5080 5476
rect 5040 5396 5080 5444
rect 5040 5364 5044 5396
rect 5076 5364 5080 5396
rect 5040 5316 5080 5364
rect 5040 5284 5044 5316
rect 5076 5284 5080 5316
rect 5040 5236 5080 5284
rect 5040 5204 5044 5236
rect 5076 5204 5080 5236
rect 5040 5156 5080 5204
rect 5040 5124 5044 5156
rect 5076 5124 5080 5156
rect 5040 5076 5080 5124
rect 5040 5044 5044 5076
rect 5076 5044 5080 5076
rect 5040 4996 5080 5044
rect 5040 4964 5044 4996
rect 5076 4964 5080 4996
rect 5040 4916 5080 4964
rect 5040 4884 5044 4916
rect 5076 4884 5080 4916
rect 5040 4836 5080 4884
rect 5040 4804 5044 4836
rect 5076 4804 5080 4836
rect 5040 4756 5080 4804
rect 5040 4724 5044 4756
rect 5076 4724 5080 4756
rect 5040 4676 5080 4724
rect 5040 4644 5044 4676
rect 5076 4644 5080 4676
rect 5040 4596 5080 4644
rect 5040 4564 5044 4596
rect 5076 4564 5080 4596
rect 5040 4516 5080 4564
rect 5040 4484 5044 4516
rect 5076 4484 5080 4516
rect 5040 4436 5080 4484
rect 5040 4404 5044 4436
rect 5076 4404 5080 4436
rect 5040 4356 5080 4404
rect 5040 4324 5044 4356
rect 5076 4324 5080 4356
rect 5040 4276 5080 4324
rect 5040 4244 5044 4276
rect 5076 4244 5080 4276
rect 5040 4196 5080 4244
rect 5040 4164 5044 4196
rect 5076 4164 5080 4196
rect 5040 4116 5080 4164
rect 5040 4084 5044 4116
rect 5076 4084 5080 4116
rect 5040 4036 5080 4084
rect 5040 4004 5044 4036
rect 5076 4004 5080 4036
rect 5040 3956 5080 4004
rect 5040 3924 5044 3956
rect 5076 3924 5080 3956
rect 5040 3876 5080 3924
rect 5040 3844 5044 3876
rect 5076 3844 5080 3876
rect 5040 3796 5080 3844
rect 5040 3764 5044 3796
rect 5076 3764 5080 3796
rect 5040 3716 5080 3764
rect 5040 3684 5044 3716
rect 5076 3684 5080 3716
rect 5040 3636 5080 3684
rect 5040 3604 5044 3636
rect 5076 3604 5080 3636
rect 5040 3556 5080 3604
rect 5040 3524 5044 3556
rect 5076 3524 5080 3556
rect 5040 3476 5080 3524
rect 5040 3444 5044 3476
rect 5076 3444 5080 3476
rect 5040 3396 5080 3444
rect 5040 3364 5044 3396
rect 5076 3364 5080 3396
rect 5040 3316 5080 3364
rect 5040 3284 5044 3316
rect 5076 3284 5080 3316
rect 5040 3236 5080 3284
rect 5040 3204 5044 3236
rect 5076 3204 5080 3236
rect 5040 3156 5080 3204
rect 5040 3124 5044 3156
rect 5076 3124 5080 3156
rect 5040 3076 5080 3124
rect 5040 3044 5044 3076
rect 5076 3044 5080 3076
rect 5040 2996 5080 3044
rect 5040 2964 5044 2996
rect 5076 2964 5080 2996
rect 5040 2916 5080 2964
rect 5040 2884 5044 2916
rect 5076 2884 5080 2916
rect 5040 2836 5080 2884
rect 5040 2804 5044 2836
rect 5076 2804 5080 2836
rect 5040 2756 5080 2804
rect 5040 2724 5044 2756
rect 5076 2724 5080 2756
rect 5040 2676 5080 2724
rect 5040 2644 5044 2676
rect 5076 2644 5080 2676
rect 5040 2596 5080 2644
rect 5040 2564 5044 2596
rect 5076 2564 5080 2596
rect 5040 2516 5080 2564
rect 5040 2484 5044 2516
rect 5076 2484 5080 2516
rect 5040 2436 5080 2484
rect 5040 2404 5044 2436
rect 5076 2404 5080 2436
rect 5040 2356 5080 2404
rect 5040 2324 5044 2356
rect 5076 2324 5080 2356
rect 5040 2276 5080 2324
rect 5040 2244 5044 2276
rect 5076 2244 5080 2276
rect 5040 2196 5080 2244
rect 5040 2164 5044 2196
rect 5076 2164 5080 2196
rect 5040 2116 5080 2164
rect 5040 2084 5044 2116
rect 5076 2084 5080 2116
rect 5040 2036 5080 2084
rect 5040 2004 5044 2036
rect 5076 2004 5080 2036
rect 5040 1956 5080 2004
rect 5040 1924 5044 1956
rect 5076 1924 5080 1956
rect 5040 1876 5080 1924
rect 5040 1844 5044 1876
rect 5076 1844 5080 1876
rect 5040 1796 5080 1844
rect 5040 1764 5044 1796
rect 5076 1764 5080 1796
rect 5040 1716 5080 1764
rect 5040 1684 5044 1716
rect 5076 1684 5080 1716
rect 5040 1636 5080 1684
rect 5040 1604 5044 1636
rect 5076 1604 5080 1636
rect 5040 1556 5080 1604
rect 5040 1524 5044 1556
rect 5076 1524 5080 1556
rect 5040 1476 5080 1524
rect 5040 1444 5044 1476
rect 5076 1444 5080 1476
rect 5040 1396 5080 1444
rect 5040 1364 5044 1396
rect 5076 1364 5080 1396
rect 5040 1316 5080 1364
rect 5040 1284 5044 1316
rect 5076 1284 5080 1316
rect 5040 1236 5080 1284
rect 5040 1204 5044 1236
rect 5076 1204 5080 1236
rect 5040 1156 5080 1204
rect 5040 1124 5044 1156
rect 5076 1124 5080 1156
rect 5040 1076 5080 1124
rect 5040 1044 5044 1076
rect 5076 1044 5080 1076
rect 5040 996 5080 1044
rect 5040 964 5044 996
rect 5076 964 5080 996
rect 5040 916 5080 964
rect 5040 884 5044 916
rect 5076 884 5080 916
rect 5040 836 5080 884
rect 5040 804 5044 836
rect 5076 804 5080 836
rect 5040 756 5080 804
rect 5040 724 5044 756
rect 5076 724 5080 756
rect 5040 676 5080 724
rect 5040 644 5044 676
rect 5076 644 5080 676
rect 5040 596 5080 644
rect 5040 564 5044 596
rect 5076 564 5080 596
rect 5040 516 5080 564
rect 5040 484 5044 516
rect 5076 484 5080 516
rect 5040 436 5080 484
rect 5040 404 5044 436
rect 5076 404 5080 436
rect 5040 356 5080 404
rect 5040 324 5044 356
rect 5076 324 5080 356
rect 5040 276 5080 324
rect 5040 244 5044 276
rect 5076 244 5080 276
rect 5040 196 5080 244
rect 5040 164 5044 196
rect 5076 164 5080 196
rect 5040 116 5080 164
rect 5040 84 5044 116
rect 5076 84 5080 116
rect 5040 36 5080 84
rect 5040 4 5044 36
rect 5076 4 5080 36
rect 4880 -716 4884 -524
rect 4916 -716 4920 -524
rect 4880 -960 4920 -716
rect 5040 -524 5080 4
rect 5120 13195 5160 15760
rect 5120 13165 5125 13195
rect 5155 13165 5160 13195
rect 5120 10235 5160 13165
rect 5120 10205 5125 10235
rect 5155 10205 5160 10235
rect 5120 10075 5160 10205
rect 5120 10045 5125 10075
rect 5155 10045 5160 10075
rect 5120 9275 5160 10045
rect 5120 9245 5125 9275
rect 5155 9245 5160 9275
rect 5120 0 5160 9245
rect 5200 15716 5240 15760
rect 5200 15684 5204 15716
rect 5236 15684 5240 15716
rect 5200 15636 5240 15684
rect 5200 15604 5204 15636
rect 5236 15604 5240 15636
rect 5200 15556 5240 15604
rect 5200 15524 5204 15556
rect 5236 15524 5240 15556
rect 5200 15476 5240 15524
rect 5200 15444 5204 15476
rect 5236 15444 5240 15476
rect 5200 15396 5240 15444
rect 5200 15364 5204 15396
rect 5236 15364 5240 15396
rect 5200 15316 5240 15364
rect 5200 15284 5204 15316
rect 5236 15284 5240 15316
rect 5200 15236 5240 15284
rect 5200 15204 5204 15236
rect 5236 15204 5240 15236
rect 5200 15156 5240 15204
rect 5200 15124 5204 15156
rect 5236 15124 5240 15156
rect 5200 15076 5240 15124
rect 5200 15044 5204 15076
rect 5236 15044 5240 15076
rect 5200 14996 5240 15044
rect 5200 14964 5204 14996
rect 5236 14964 5240 14996
rect 5200 14916 5240 14964
rect 5200 14884 5204 14916
rect 5236 14884 5240 14916
rect 5200 14836 5240 14884
rect 5200 14804 5204 14836
rect 5236 14804 5240 14836
rect 5200 14756 5240 14804
rect 5200 14724 5204 14756
rect 5236 14724 5240 14756
rect 5200 14676 5240 14724
rect 5200 14644 5204 14676
rect 5236 14644 5240 14676
rect 5200 14596 5240 14644
rect 5200 14564 5204 14596
rect 5236 14564 5240 14596
rect 5200 14516 5240 14564
rect 5200 14484 5204 14516
rect 5236 14484 5240 14516
rect 5200 14436 5240 14484
rect 5200 14404 5204 14436
rect 5236 14404 5240 14436
rect 5200 14356 5240 14404
rect 5200 14324 5204 14356
rect 5236 14324 5240 14356
rect 5200 14276 5240 14324
rect 5200 14244 5204 14276
rect 5236 14244 5240 14276
rect 5200 14196 5240 14244
rect 5200 14164 5204 14196
rect 5236 14164 5240 14196
rect 5200 14116 5240 14164
rect 5200 14084 5204 14116
rect 5236 14084 5240 14116
rect 5200 14036 5240 14084
rect 5200 14004 5204 14036
rect 5236 14004 5240 14036
rect 5200 13956 5240 14004
rect 5200 13924 5204 13956
rect 5236 13924 5240 13956
rect 5200 13876 5240 13924
rect 5200 13844 5204 13876
rect 5236 13844 5240 13876
rect 5200 13796 5240 13844
rect 5200 13764 5204 13796
rect 5236 13764 5240 13796
rect 5200 13716 5240 13764
rect 5200 13684 5204 13716
rect 5236 13684 5240 13716
rect 5200 13636 5240 13684
rect 5200 13604 5204 13636
rect 5236 13604 5240 13636
rect 5200 13556 5240 13604
rect 5200 13524 5204 13556
rect 5236 13524 5240 13556
rect 5200 13476 5240 13524
rect 5200 13444 5204 13476
rect 5236 13444 5240 13476
rect 5200 13396 5240 13444
rect 5200 13364 5204 13396
rect 5236 13364 5240 13396
rect 5200 13316 5240 13364
rect 5200 13284 5204 13316
rect 5236 13284 5240 13316
rect 5200 13236 5240 13284
rect 5200 13204 5204 13236
rect 5236 13204 5240 13236
rect 5200 13156 5240 13204
rect 5200 13124 5204 13156
rect 5236 13124 5240 13156
rect 5200 13076 5240 13124
rect 5200 13044 5204 13076
rect 5236 13044 5240 13076
rect 5200 12996 5240 13044
rect 5200 12964 5204 12996
rect 5236 12964 5240 12996
rect 5200 12916 5240 12964
rect 5200 12884 5204 12916
rect 5236 12884 5240 12916
rect 5200 12836 5240 12884
rect 5200 12804 5204 12836
rect 5236 12804 5240 12836
rect 5200 12756 5240 12804
rect 5200 12724 5204 12756
rect 5236 12724 5240 12756
rect 5200 12676 5240 12724
rect 5200 12644 5204 12676
rect 5236 12644 5240 12676
rect 5200 12596 5240 12644
rect 5200 12564 5204 12596
rect 5236 12564 5240 12596
rect 5200 12516 5240 12564
rect 5200 12484 5204 12516
rect 5236 12484 5240 12516
rect 5200 12436 5240 12484
rect 5200 12404 5204 12436
rect 5236 12404 5240 12436
rect 5200 12356 5240 12404
rect 5200 12324 5204 12356
rect 5236 12324 5240 12356
rect 5200 12276 5240 12324
rect 5200 12244 5204 12276
rect 5236 12244 5240 12276
rect 5200 12196 5240 12244
rect 5200 12164 5204 12196
rect 5236 12164 5240 12196
rect 5200 12116 5240 12164
rect 5200 12084 5204 12116
rect 5236 12084 5240 12116
rect 5200 12036 5240 12084
rect 5200 12004 5204 12036
rect 5236 12004 5240 12036
rect 5200 11956 5240 12004
rect 5200 11924 5204 11956
rect 5236 11924 5240 11956
rect 5200 11876 5240 11924
rect 5200 11844 5204 11876
rect 5236 11844 5240 11876
rect 5200 11796 5240 11844
rect 5200 11764 5204 11796
rect 5236 11764 5240 11796
rect 5200 11716 5240 11764
rect 5200 11684 5204 11716
rect 5236 11684 5240 11716
rect 5200 11636 5240 11684
rect 5200 11604 5204 11636
rect 5236 11604 5240 11636
rect 5200 11556 5240 11604
rect 5200 11524 5204 11556
rect 5236 11524 5240 11556
rect 5200 11476 5240 11524
rect 5200 11444 5204 11476
rect 5236 11444 5240 11476
rect 5200 11396 5240 11444
rect 5200 11364 5204 11396
rect 5236 11364 5240 11396
rect 5200 11316 5240 11364
rect 5200 11284 5204 11316
rect 5236 11284 5240 11316
rect 5200 11236 5240 11284
rect 5200 11204 5204 11236
rect 5236 11204 5240 11236
rect 5200 11156 5240 11204
rect 5200 11124 5204 11156
rect 5236 11124 5240 11156
rect 5200 11076 5240 11124
rect 5200 11044 5204 11076
rect 5236 11044 5240 11076
rect 5200 10996 5240 11044
rect 5200 10964 5204 10996
rect 5236 10964 5240 10996
rect 5200 10916 5240 10964
rect 5200 10884 5204 10916
rect 5236 10884 5240 10916
rect 5200 10836 5240 10884
rect 5200 10804 5204 10836
rect 5236 10804 5240 10836
rect 5200 10756 5240 10804
rect 5200 10724 5204 10756
rect 5236 10724 5240 10756
rect 5200 10676 5240 10724
rect 5200 10644 5204 10676
rect 5236 10644 5240 10676
rect 5200 10596 5240 10644
rect 5200 10564 5204 10596
rect 5236 10564 5240 10596
rect 5200 10516 5240 10564
rect 5200 10484 5204 10516
rect 5236 10484 5240 10516
rect 5200 10436 5240 10484
rect 5200 10404 5204 10436
rect 5236 10404 5240 10436
rect 5200 10356 5240 10404
rect 5200 10324 5204 10356
rect 5236 10324 5240 10356
rect 5200 10276 5240 10324
rect 5200 10244 5204 10276
rect 5236 10244 5240 10276
rect 5200 10196 5240 10244
rect 5200 10164 5204 10196
rect 5236 10164 5240 10196
rect 5200 10116 5240 10164
rect 5200 10084 5204 10116
rect 5236 10084 5240 10116
rect 5200 10036 5240 10084
rect 5200 10004 5204 10036
rect 5236 10004 5240 10036
rect 5200 9956 5240 10004
rect 5200 9924 5204 9956
rect 5236 9924 5240 9956
rect 5200 9876 5240 9924
rect 5200 9844 5204 9876
rect 5236 9844 5240 9876
rect 5200 9796 5240 9844
rect 5200 9764 5204 9796
rect 5236 9764 5240 9796
rect 5200 9716 5240 9764
rect 5200 9684 5204 9716
rect 5236 9684 5240 9716
rect 5200 9636 5240 9684
rect 5200 9604 5204 9636
rect 5236 9604 5240 9636
rect 5200 9556 5240 9604
rect 5200 9524 5204 9556
rect 5236 9524 5240 9556
rect 5200 9476 5240 9524
rect 5200 9444 5204 9476
rect 5236 9444 5240 9476
rect 5200 9396 5240 9444
rect 5200 9364 5204 9396
rect 5236 9364 5240 9396
rect 5200 9316 5240 9364
rect 5200 9284 5204 9316
rect 5236 9284 5240 9316
rect 5200 9236 5240 9284
rect 5200 9204 5204 9236
rect 5236 9204 5240 9236
rect 5200 9156 5240 9204
rect 5200 9124 5204 9156
rect 5236 9124 5240 9156
rect 5200 9076 5240 9124
rect 5200 9044 5204 9076
rect 5236 9044 5240 9076
rect 5200 8996 5240 9044
rect 5200 8964 5204 8996
rect 5236 8964 5240 8996
rect 5200 8916 5240 8964
rect 5200 8884 5204 8916
rect 5236 8884 5240 8916
rect 5200 8836 5240 8884
rect 5200 8804 5204 8836
rect 5236 8804 5240 8836
rect 5200 8756 5240 8804
rect 5200 8724 5204 8756
rect 5236 8724 5240 8756
rect 5200 8676 5240 8724
rect 5200 8644 5204 8676
rect 5236 8644 5240 8676
rect 5200 8596 5240 8644
rect 5200 8564 5204 8596
rect 5236 8564 5240 8596
rect 5200 8516 5240 8564
rect 5200 8484 5204 8516
rect 5236 8484 5240 8516
rect 5200 8436 5240 8484
rect 5200 8404 5204 8436
rect 5236 8404 5240 8436
rect 5200 8356 5240 8404
rect 5200 8324 5204 8356
rect 5236 8324 5240 8356
rect 5200 8276 5240 8324
rect 5200 8244 5204 8276
rect 5236 8244 5240 8276
rect 5200 8196 5240 8244
rect 5200 8164 5204 8196
rect 5236 8164 5240 8196
rect 5200 8116 5240 8164
rect 5200 8084 5204 8116
rect 5236 8084 5240 8116
rect 5200 8036 5240 8084
rect 5200 8004 5204 8036
rect 5236 8004 5240 8036
rect 5200 7956 5240 8004
rect 5200 7924 5204 7956
rect 5236 7924 5240 7956
rect 5200 7876 5240 7924
rect 5200 7844 5204 7876
rect 5236 7844 5240 7876
rect 5200 7796 5240 7844
rect 5200 7764 5204 7796
rect 5236 7764 5240 7796
rect 5200 7716 5240 7764
rect 5200 7684 5204 7716
rect 5236 7684 5240 7716
rect 5200 7636 5240 7684
rect 5200 7604 5204 7636
rect 5236 7604 5240 7636
rect 5200 7556 5240 7604
rect 5200 7524 5204 7556
rect 5236 7524 5240 7556
rect 5200 7476 5240 7524
rect 5200 7444 5204 7476
rect 5236 7444 5240 7476
rect 5200 7396 5240 7444
rect 5200 7364 5204 7396
rect 5236 7364 5240 7396
rect 5200 7316 5240 7364
rect 5200 7284 5204 7316
rect 5236 7284 5240 7316
rect 5200 7236 5240 7284
rect 5200 7204 5204 7236
rect 5236 7204 5240 7236
rect 5200 7156 5240 7204
rect 5200 7124 5204 7156
rect 5236 7124 5240 7156
rect 5200 7076 5240 7124
rect 5200 7044 5204 7076
rect 5236 7044 5240 7076
rect 5200 6996 5240 7044
rect 5200 6964 5204 6996
rect 5236 6964 5240 6996
rect 5200 6916 5240 6964
rect 5200 6884 5204 6916
rect 5236 6884 5240 6916
rect 5200 6836 5240 6884
rect 5200 6804 5204 6836
rect 5236 6804 5240 6836
rect 5200 6756 5240 6804
rect 5200 6724 5204 6756
rect 5236 6724 5240 6756
rect 5200 6676 5240 6724
rect 5200 6644 5204 6676
rect 5236 6644 5240 6676
rect 5200 6596 5240 6644
rect 5200 6564 5204 6596
rect 5236 6564 5240 6596
rect 5200 6516 5240 6564
rect 5200 6484 5204 6516
rect 5236 6484 5240 6516
rect 5200 6436 5240 6484
rect 5200 6404 5204 6436
rect 5236 6404 5240 6436
rect 5200 6356 5240 6404
rect 5200 6324 5204 6356
rect 5236 6324 5240 6356
rect 5200 6276 5240 6324
rect 5200 6244 5204 6276
rect 5236 6244 5240 6276
rect 5200 6196 5240 6244
rect 5200 6164 5204 6196
rect 5236 6164 5240 6196
rect 5200 6116 5240 6164
rect 5200 6084 5204 6116
rect 5236 6084 5240 6116
rect 5200 6036 5240 6084
rect 5200 6004 5204 6036
rect 5236 6004 5240 6036
rect 5200 5956 5240 6004
rect 5200 5924 5204 5956
rect 5236 5924 5240 5956
rect 5200 5876 5240 5924
rect 5200 5844 5204 5876
rect 5236 5844 5240 5876
rect 5200 5796 5240 5844
rect 5200 5764 5204 5796
rect 5236 5764 5240 5796
rect 5200 5716 5240 5764
rect 5200 5684 5204 5716
rect 5236 5684 5240 5716
rect 5200 5636 5240 5684
rect 5200 5604 5204 5636
rect 5236 5604 5240 5636
rect 5200 5556 5240 5604
rect 5200 5524 5204 5556
rect 5236 5524 5240 5556
rect 5200 5476 5240 5524
rect 5200 5444 5204 5476
rect 5236 5444 5240 5476
rect 5200 5396 5240 5444
rect 5200 5364 5204 5396
rect 5236 5364 5240 5396
rect 5200 5316 5240 5364
rect 5200 5284 5204 5316
rect 5236 5284 5240 5316
rect 5200 5236 5240 5284
rect 5200 5204 5204 5236
rect 5236 5204 5240 5236
rect 5200 5156 5240 5204
rect 5200 5124 5204 5156
rect 5236 5124 5240 5156
rect 5200 5076 5240 5124
rect 5200 5044 5204 5076
rect 5236 5044 5240 5076
rect 5200 4996 5240 5044
rect 5200 4964 5204 4996
rect 5236 4964 5240 4996
rect 5200 4916 5240 4964
rect 5200 4884 5204 4916
rect 5236 4884 5240 4916
rect 5200 4836 5240 4884
rect 5200 4804 5204 4836
rect 5236 4804 5240 4836
rect 5200 4756 5240 4804
rect 5200 4724 5204 4756
rect 5236 4724 5240 4756
rect 5200 4676 5240 4724
rect 5200 4644 5204 4676
rect 5236 4644 5240 4676
rect 5200 4596 5240 4644
rect 5200 4564 5204 4596
rect 5236 4564 5240 4596
rect 5200 4516 5240 4564
rect 5200 4484 5204 4516
rect 5236 4484 5240 4516
rect 5200 4436 5240 4484
rect 5200 4404 5204 4436
rect 5236 4404 5240 4436
rect 5200 4356 5240 4404
rect 5200 4324 5204 4356
rect 5236 4324 5240 4356
rect 5200 4276 5240 4324
rect 5200 4244 5204 4276
rect 5236 4244 5240 4276
rect 5200 4196 5240 4244
rect 5200 4164 5204 4196
rect 5236 4164 5240 4196
rect 5200 4116 5240 4164
rect 5200 4084 5204 4116
rect 5236 4084 5240 4116
rect 5200 4036 5240 4084
rect 5200 4004 5204 4036
rect 5236 4004 5240 4036
rect 5200 3956 5240 4004
rect 5200 3924 5204 3956
rect 5236 3924 5240 3956
rect 5200 3876 5240 3924
rect 5200 3844 5204 3876
rect 5236 3844 5240 3876
rect 5200 3796 5240 3844
rect 5200 3764 5204 3796
rect 5236 3764 5240 3796
rect 5200 3716 5240 3764
rect 5200 3684 5204 3716
rect 5236 3684 5240 3716
rect 5200 3636 5240 3684
rect 5200 3604 5204 3636
rect 5236 3604 5240 3636
rect 5200 3556 5240 3604
rect 5200 3524 5204 3556
rect 5236 3524 5240 3556
rect 5200 3476 5240 3524
rect 5200 3444 5204 3476
rect 5236 3444 5240 3476
rect 5200 3396 5240 3444
rect 5200 3364 5204 3396
rect 5236 3364 5240 3396
rect 5200 3316 5240 3364
rect 5200 3284 5204 3316
rect 5236 3284 5240 3316
rect 5200 3236 5240 3284
rect 5200 3204 5204 3236
rect 5236 3204 5240 3236
rect 5200 3156 5240 3204
rect 5200 3124 5204 3156
rect 5236 3124 5240 3156
rect 5200 3076 5240 3124
rect 5200 3044 5204 3076
rect 5236 3044 5240 3076
rect 5200 2996 5240 3044
rect 5200 2964 5204 2996
rect 5236 2964 5240 2996
rect 5200 2916 5240 2964
rect 5200 2884 5204 2916
rect 5236 2884 5240 2916
rect 5200 2836 5240 2884
rect 5200 2804 5204 2836
rect 5236 2804 5240 2836
rect 5200 2756 5240 2804
rect 5200 2724 5204 2756
rect 5236 2724 5240 2756
rect 5200 2676 5240 2724
rect 5200 2644 5204 2676
rect 5236 2644 5240 2676
rect 5200 2596 5240 2644
rect 5200 2564 5204 2596
rect 5236 2564 5240 2596
rect 5200 2516 5240 2564
rect 5200 2484 5204 2516
rect 5236 2484 5240 2516
rect 5200 2436 5240 2484
rect 5200 2404 5204 2436
rect 5236 2404 5240 2436
rect 5200 2356 5240 2404
rect 5200 2324 5204 2356
rect 5236 2324 5240 2356
rect 5200 2276 5240 2324
rect 5200 2244 5204 2276
rect 5236 2244 5240 2276
rect 5200 2196 5240 2244
rect 5200 2164 5204 2196
rect 5236 2164 5240 2196
rect 5200 2116 5240 2164
rect 5200 2084 5204 2116
rect 5236 2084 5240 2116
rect 5200 2036 5240 2084
rect 5200 2004 5204 2036
rect 5236 2004 5240 2036
rect 5200 1956 5240 2004
rect 5200 1924 5204 1956
rect 5236 1924 5240 1956
rect 5200 1876 5240 1924
rect 5200 1844 5204 1876
rect 5236 1844 5240 1876
rect 5200 1796 5240 1844
rect 5200 1764 5204 1796
rect 5236 1764 5240 1796
rect 5200 1716 5240 1764
rect 5200 1684 5204 1716
rect 5236 1684 5240 1716
rect 5200 1636 5240 1684
rect 5200 1604 5204 1636
rect 5236 1604 5240 1636
rect 5200 1556 5240 1604
rect 5200 1524 5204 1556
rect 5236 1524 5240 1556
rect 5200 1476 5240 1524
rect 5200 1444 5204 1476
rect 5236 1444 5240 1476
rect 5200 1396 5240 1444
rect 5200 1364 5204 1396
rect 5236 1364 5240 1396
rect 5200 1316 5240 1364
rect 5200 1284 5204 1316
rect 5236 1284 5240 1316
rect 5200 1236 5240 1284
rect 5200 1204 5204 1236
rect 5236 1204 5240 1236
rect 5200 1156 5240 1204
rect 5200 1124 5204 1156
rect 5236 1124 5240 1156
rect 5200 1076 5240 1124
rect 5200 1044 5204 1076
rect 5236 1044 5240 1076
rect 5200 996 5240 1044
rect 5200 964 5204 996
rect 5236 964 5240 996
rect 5200 916 5240 964
rect 5200 884 5204 916
rect 5236 884 5240 916
rect 5200 836 5240 884
rect 5200 804 5204 836
rect 5236 804 5240 836
rect 5200 756 5240 804
rect 5200 724 5204 756
rect 5236 724 5240 756
rect 5200 676 5240 724
rect 5200 644 5204 676
rect 5236 644 5240 676
rect 5200 596 5240 644
rect 5200 564 5204 596
rect 5236 564 5240 596
rect 5200 516 5240 564
rect 5200 484 5204 516
rect 5236 484 5240 516
rect 5200 436 5240 484
rect 5200 404 5204 436
rect 5236 404 5240 436
rect 5200 356 5240 404
rect 5200 324 5204 356
rect 5236 324 5240 356
rect 5200 276 5240 324
rect 5200 244 5204 276
rect 5236 244 5240 276
rect 5200 196 5240 244
rect 5200 164 5204 196
rect 5236 164 5240 196
rect 5200 116 5240 164
rect 5200 84 5204 116
rect 5236 84 5240 116
rect 5200 36 5240 84
rect 5200 4 5204 36
rect 5236 4 5240 36
rect 5040 -716 5044 -524
rect 5076 -716 5080 -524
rect 5040 -960 5080 -716
rect 5200 -524 5240 4
rect 5280 14315 5320 15760
rect 5280 14285 5285 14315
rect 5315 14285 5320 14315
rect 5280 13355 5320 14285
rect 5280 13325 5285 13355
rect 5315 13325 5320 13355
rect 5280 13195 5320 13325
rect 5280 13165 5285 13195
rect 5315 13165 5320 13195
rect 5280 0 5320 13165
rect 5360 15716 5400 15760
rect 5360 15684 5364 15716
rect 5396 15684 5400 15716
rect 5360 15636 5400 15684
rect 5360 15604 5364 15636
rect 5396 15604 5400 15636
rect 5360 15556 5400 15604
rect 5360 15524 5364 15556
rect 5396 15524 5400 15556
rect 5360 15476 5400 15524
rect 5360 15444 5364 15476
rect 5396 15444 5400 15476
rect 5360 15396 5400 15444
rect 5360 15364 5364 15396
rect 5396 15364 5400 15396
rect 5360 15316 5400 15364
rect 5360 15284 5364 15316
rect 5396 15284 5400 15316
rect 5360 15236 5400 15284
rect 5360 15204 5364 15236
rect 5396 15204 5400 15236
rect 5360 15156 5400 15204
rect 5360 15124 5364 15156
rect 5396 15124 5400 15156
rect 5360 15076 5400 15124
rect 5360 15044 5364 15076
rect 5396 15044 5400 15076
rect 5360 14996 5400 15044
rect 5360 14964 5364 14996
rect 5396 14964 5400 14996
rect 5360 14916 5400 14964
rect 5360 14884 5364 14916
rect 5396 14884 5400 14916
rect 5360 14836 5400 14884
rect 5360 14804 5364 14836
rect 5396 14804 5400 14836
rect 5360 14756 5400 14804
rect 5360 14724 5364 14756
rect 5396 14724 5400 14756
rect 5360 14676 5400 14724
rect 5360 14644 5364 14676
rect 5396 14644 5400 14676
rect 5360 14596 5400 14644
rect 5360 14564 5364 14596
rect 5396 14564 5400 14596
rect 5360 14516 5400 14564
rect 5360 14484 5364 14516
rect 5396 14484 5400 14516
rect 5360 14436 5400 14484
rect 5360 14404 5364 14436
rect 5396 14404 5400 14436
rect 5360 14356 5400 14404
rect 5360 14324 5364 14356
rect 5396 14324 5400 14356
rect 5360 14276 5400 14324
rect 5360 14244 5364 14276
rect 5396 14244 5400 14276
rect 5360 14196 5400 14244
rect 5360 14164 5364 14196
rect 5396 14164 5400 14196
rect 5360 14116 5400 14164
rect 5360 14084 5364 14116
rect 5396 14084 5400 14116
rect 5360 14036 5400 14084
rect 5360 14004 5364 14036
rect 5396 14004 5400 14036
rect 5360 13956 5400 14004
rect 5360 13924 5364 13956
rect 5396 13924 5400 13956
rect 5360 13876 5400 13924
rect 5360 13844 5364 13876
rect 5396 13844 5400 13876
rect 5360 13796 5400 13844
rect 5360 13764 5364 13796
rect 5396 13764 5400 13796
rect 5360 13716 5400 13764
rect 5360 13684 5364 13716
rect 5396 13684 5400 13716
rect 5360 13636 5400 13684
rect 5360 13604 5364 13636
rect 5396 13604 5400 13636
rect 5360 13556 5400 13604
rect 5360 13524 5364 13556
rect 5396 13524 5400 13556
rect 5360 13476 5400 13524
rect 5360 13444 5364 13476
rect 5396 13444 5400 13476
rect 5360 13396 5400 13444
rect 5360 13364 5364 13396
rect 5396 13364 5400 13396
rect 5360 13316 5400 13364
rect 5360 13284 5364 13316
rect 5396 13284 5400 13316
rect 5360 13236 5400 13284
rect 5360 13204 5364 13236
rect 5396 13204 5400 13236
rect 5360 13156 5400 13204
rect 5360 13124 5364 13156
rect 5396 13124 5400 13156
rect 5360 13076 5400 13124
rect 5360 13044 5364 13076
rect 5396 13044 5400 13076
rect 5360 12996 5400 13044
rect 5360 12964 5364 12996
rect 5396 12964 5400 12996
rect 5360 12916 5400 12964
rect 5360 12884 5364 12916
rect 5396 12884 5400 12916
rect 5360 12836 5400 12884
rect 5360 12804 5364 12836
rect 5396 12804 5400 12836
rect 5360 12756 5400 12804
rect 5360 12724 5364 12756
rect 5396 12724 5400 12756
rect 5360 12676 5400 12724
rect 5360 12644 5364 12676
rect 5396 12644 5400 12676
rect 5360 12596 5400 12644
rect 5360 12564 5364 12596
rect 5396 12564 5400 12596
rect 5360 12516 5400 12564
rect 5360 12484 5364 12516
rect 5396 12484 5400 12516
rect 5360 12436 5400 12484
rect 5360 12404 5364 12436
rect 5396 12404 5400 12436
rect 5360 12356 5400 12404
rect 5360 12324 5364 12356
rect 5396 12324 5400 12356
rect 5360 12276 5400 12324
rect 5360 12244 5364 12276
rect 5396 12244 5400 12276
rect 5360 12196 5400 12244
rect 5360 12164 5364 12196
rect 5396 12164 5400 12196
rect 5360 12116 5400 12164
rect 5360 12084 5364 12116
rect 5396 12084 5400 12116
rect 5360 12036 5400 12084
rect 5360 12004 5364 12036
rect 5396 12004 5400 12036
rect 5360 11956 5400 12004
rect 5360 11924 5364 11956
rect 5396 11924 5400 11956
rect 5360 11876 5400 11924
rect 5360 11844 5364 11876
rect 5396 11844 5400 11876
rect 5360 11796 5400 11844
rect 5360 11764 5364 11796
rect 5396 11764 5400 11796
rect 5360 11716 5400 11764
rect 5360 11684 5364 11716
rect 5396 11684 5400 11716
rect 5360 11636 5400 11684
rect 5360 11604 5364 11636
rect 5396 11604 5400 11636
rect 5360 11556 5400 11604
rect 5360 11524 5364 11556
rect 5396 11524 5400 11556
rect 5360 11476 5400 11524
rect 5360 11444 5364 11476
rect 5396 11444 5400 11476
rect 5360 11396 5400 11444
rect 5360 11364 5364 11396
rect 5396 11364 5400 11396
rect 5360 11316 5400 11364
rect 5360 11284 5364 11316
rect 5396 11284 5400 11316
rect 5360 11236 5400 11284
rect 5360 11204 5364 11236
rect 5396 11204 5400 11236
rect 5360 11156 5400 11204
rect 5360 11124 5364 11156
rect 5396 11124 5400 11156
rect 5360 11076 5400 11124
rect 5360 11044 5364 11076
rect 5396 11044 5400 11076
rect 5360 10996 5400 11044
rect 5360 10964 5364 10996
rect 5396 10964 5400 10996
rect 5360 10916 5400 10964
rect 5360 10884 5364 10916
rect 5396 10884 5400 10916
rect 5360 10836 5400 10884
rect 5360 10804 5364 10836
rect 5396 10804 5400 10836
rect 5360 10756 5400 10804
rect 5360 10724 5364 10756
rect 5396 10724 5400 10756
rect 5360 10676 5400 10724
rect 5360 10644 5364 10676
rect 5396 10644 5400 10676
rect 5360 10596 5400 10644
rect 5360 10564 5364 10596
rect 5396 10564 5400 10596
rect 5360 10516 5400 10564
rect 5360 10484 5364 10516
rect 5396 10484 5400 10516
rect 5360 10436 5400 10484
rect 5360 10404 5364 10436
rect 5396 10404 5400 10436
rect 5360 10356 5400 10404
rect 5360 10324 5364 10356
rect 5396 10324 5400 10356
rect 5360 10276 5400 10324
rect 5360 10244 5364 10276
rect 5396 10244 5400 10276
rect 5360 10196 5400 10244
rect 5360 10164 5364 10196
rect 5396 10164 5400 10196
rect 5360 10116 5400 10164
rect 5360 10084 5364 10116
rect 5396 10084 5400 10116
rect 5360 10036 5400 10084
rect 5360 10004 5364 10036
rect 5396 10004 5400 10036
rect 5360 9956 5400 10004
rect 5360 9924 5364 9956
rect 5396 9924 5400 9956
rect 5360 9876 5400 9924
rect 5360 9844 5364 9876
rect 5396 9844 5400 9876
rect 5360 9796 5400 9844
rect 5360 9764 5364 9796
rect 5396 9764 5400 9796
rect 5360 9716 5400 9764
rect 5360 9684 5364 9716
rect 5396 9684 5400 9716
rect 5360 9636 5400 9684
rect 5360 9604 5364 9636
rect 5396 9604 5400 9636
rect 5360 9556 5400 9604
rect 5360 9524 5364 9556
rect 5396 9524 5400 9556
rect 5360 9476 5400 9524
rect 5360 9444 5364 9476
rect 5396 9444 5400 9476
rect 5360 9396 5400 9444
rect 5360 9364 5364 9396
rect 5396 9364 5400 9396
rect 5360 9316 5400 9364
rect 5360 9284 5364 9316
rect 5396 9284 5400 9316
rect 5360 9236 5400 9284
rect 5360 9204 5364 9236
rect 5396 9204 5400 9236
rect 5360 9156 5400 9204
rect 5360 9124 5364 9156
rect 5396 9124 5400 9156
rect 5360 9076 5400 9124
rect 5360 9044 5364 9076
rect 5396 9044 5400 9076
rect 5360 8996 5400 9044
rect 5360 8964 5364 8996
rect 5396 8964 5400 8996
rect 5360 8916 5400 8964
rect 5360 8884 5364 8916
rect 5396 8884 5400 8916
rect 5360 8836 5400 8884
rect 5360 8804 5364 8836
rect 5396 8804 5400 8836
rect 5360 8756 5400 8804
rect 5360 8724 5364 8756
rect 5396 8724 5400 8756
rect 5360 8676 5400 8724
rect 5360 8644 5364 8676
rect 5396 8644 5400 8676
rect 5360 8596 5400 8644
rect 5360 8564 5364 8596
rect 5396 8564 5400 8596
rect 5360 8516 5400 8564
rect 5360 8484 5364 8516
rect 5396 8484 5400 8516
rect 5360 8436 5400 8484
rect 5360 8404 5364 8436
rect 5396 8404 5400 8436
rect 5360 8356 5400 8404
rect 5360 8324 5364 8356
rect 5396 8324 5400 8356
rect 5360 8276 5400 8324
rect 5360 8244 5364 8276
rect 5396 8244 5400 8276
rect 5360 8196 5400 8244
rect 5360 8164 5364 8196
rect 5396 8164 5400 8196
rect 5360 8116 5400 8164
rect 5360 8084 5364 8116
rect 5396 8084 5400 8116
rect 5360 8036 5400 8084
rect 5360 8004 5364 8036
rect 5396 8004 5400 8036
rect 5360 7956 5400 8004
rect 5360 7924 5364 7956
rect 5396 7924 5400 7956
rect 5360 7876 5400 7924
rect 5360 7844 5364 7876
rect 5396 7844 5400 7876
rect 5360 7796 5400 7844
rect 5360 7764 5364 7796
rect 5396 7764 5400 7796
rect 5360 7716 5400 7764
rect 5360 7684 5364 7716
rect 5396 7684 5400 7716
rect 5360 7636 5400 7684
rect 5360 7604 5364 7636
rect 5396 7604 5400 7636
rect 5360 7556 5400 7604
rect 5360 7524 5364 7556
rect 5396 7524 5400 7556
rect 5360 7476 5400 7524
rect 5360 7444 5364 7476
rect 5396 7444 5400 7476
rect 5360 7396 5400 7444
rect 5360 7364 5364 7396
rect 5396 7364 5400 7396
rect 5360 7316 5400 7364
rect 5360 7284 5364 7316
rect 5396 7284 5400 7316
rect 5360 7236 5400 7284
rect 5360 7204 5364 7236
rect 5396 7204 5400 7236
rect 5360 7156 5400 7204
rect 5360 7124 5364 7156
rect 5396 7124 5400 7156
rect 5360 7076 5400 7124
rect 5360 7044 5364 7076
rect 5396 7044 5400 7076
rect 5360 6996 5400 7044
rect 5360 6964 5364 6996
rect 5396 6964 5400 6996
rect 5360 6916 5400 6964
rect 5360 6884 5364 6916
rect 5396 6884 5400 6916
rect 5360 6836 5400 6884
rect 5360 6804 5364 6836
rect 5396 6804 5400 6836
rect 5360 6756 5400 6804
rect 5360 6724 5364 6756
rect 5396 6724 5400 6756
rect 5360 6676 5400 6724
rect 5360 6644 5364 6676
rect 5396 6644 5400 6676
rect 5360 6596 5400 6644
rect 5360 6564 5364 6596
rect 5396 6564 5400 6596
rect 5360 6516 5400 6564
rect 5360 6484 5364 6516
rect 5396 6484 5400 6516
rect 5360 6436 5400 6484
rect 5360 6404 5364 6436
rect 5396 6404 5400 6436
rect 5360 6356 5400 6404
rect 5360 6324 5364 6356
rect 5396 6324 5400 6356
rect 5360 6276 5400 6324
rect 5360 6244 5364 6276
rect 5396 6244 5400 6276
rect 5360 6196 5400 6244
rect 5360 6164 5364 6196
rect 5396 6164 5400 6196
rect 5360 6116 5400 6164
rect 5360 6084 5364 6116
rect 5396 6084 5400 6116
rect 5360 6036 5400 6084
rect 5360 6004 5364 6036
rect 5396 6004 5400 6036
rect 5360 5956 5400 6004
rect 5360 5924 5364 5956
rect 5396 5924 5400 5956
rect 5360 5876 5400 5924
rect 5360 5844 5364 5876
rect 5396 5844 5400 5876
rect 5360 5796 5400 5844
rect 5360 5764 5364 5796
rect 5396 5764 5400 5796
rect 5360 5716 5400 5764
rect 5360 5684 5364 5716
rect 5396 5684 5400 5716
rect 5360 5636 5400 5684
rect 5360 5604 5364 5636
rect 5396 5604 5400 5636
rect 5360 5556 5400 5604
rect 5360 5524 5364 5556
rect 5396 5524 5400 5556
rect 5360 5476 5400 5524
rect 5360 5444 5364 5476
rect 5396 5444 5400 5476
rect 5360 5396 5400 5444
rect 5360 5364 5364 5396
rect 5396 5364 5400 5396
rect 5360 5316 5400 5364
rect 5360 5284 5364 5316
rect 5396 5284 5400 5316
rect 5360 5236 5400 5284
rect 5360 5204 5364 5236
rect 5396 5204 5400 5236
rect 5360 5156 5400 5204
rect 5360 5124 5364 5156
rect 5396 5124 5400 5156
rect 5360 5076 5400 5124
rect 5360 5044 5364 5076
rect 5396 5044 5400 5076
rect 5360 4996 5400 5044
rect 5360 4964 5364 4996
rect 5396 4964 5400 4996
rect 5360 4916 5400 4964
rect 5360 4884 5364 4916
rect 5396 4884 5400 4916
rect 5360 4836 5400 4884
rect 5360 4804 5364 4836
rect 5396 4804 5400 4836
rect 5360 4756 5400 4804
rect 5360 4724 5364 4756
rect 5396 4724 5400 4756
rect 5360 4676 5400 4724
rect 5360 4644 5364 4676
rect 5396 4644 5400 4676
rect 5360 4596 5400 4644
rect 5360 4564 5364 4596
rect 5396 4564 5400 4596
rect 5360 4516 5400 4564
rect 5360 4484 5364 4516
rect 5396 4484 5400 4516
rect 5360 4436 5400 4484
rect 5360 4404 5364 4436
rect 5396 4404 5400 4436
rect 5360 4356 5400 4404
rect 5360 4324 5364 4356
rect 5396 4324 5400 4356
rect 5360 4276 5400 4324
rect 5360 4244 5364 4276
rect 5396 4244 5400 4276
rect 5360 4196 5400 4244
rect 5360 4164 5364 4196
rect 5396 4164 5400 4196
rect 5360 4116 5400 4164
rect 5360 4084 5364 4116
rect 5396 4084 5400 4116
rect 5360 4036 5400 4084
rect 5360 4004 5364 4036
rect 5396 4004 5400 4036
rect 5360 3956 5400 4004
rect 5360 3924 5364 3956
rect 5396 3924 5400 3956
rect 5360 3876 5400 3924
rect 5360 3844 5364 3876
rect 5396 3844 5400 3876
rect 5360 3796 5400 3844
rect 5360 3764 5364 3796
rect 5396 3764 5400 3796
rect 5360 3716 5400 3764
rect 5360 3684 5364 3716
rect 5396 3684 5400 3716
rect 5360 3636 5400 3684
rect 5360 3604 5364 3636
rect 5396 3604 5400 3636
rect 5360 3556 5400 3604
rect 5360 3524 5364 3556
rect 5396 3524 5400 3556
rect 5360 3476 5400 3524
rect 5360 3444 5364 3476
rect 5396 3444 5400 3476
rect 5360 3396 5400 3444
rect 5360 3364 5364 3396
rect 5396 3364 5400 3396
rect 5360 3316 5400 3364
rect 5360 3284 5364 3316
rect 5396 3284 5400 3316
rect 5360 3236 5400 3284
rect 5360 3204 5364 3236
rect 5396 3204 5400 3236
rect 5360 3156 5400 3204
rect 5360 3124 5364 3156
rect 5396 3124 5400 3156
rect 5360 3076 5400 3124
rect 5360 3044 5364 3076
rect 5396 3044 5400 3076
rect 5360 2996 5400 3044
rect 5360 2964 5364 2996
rect 5396 2964 5400 2996
rect 5360 2916 5400 2964
rect 5360 2884 5364 2916
rect 5396 2884 5400 2916
rect 5360 2836 5400 2884
rect 5360 2804 5364 2836
rect 5396 2804 5400 2836
rect 5360 2756 5400 2804
rect 5360 2724 5364 2756
rect 5396 2724 5400 2756
rect 5360 2676 5400 2724
rect 5360 2644 5364 2676
rect 5396 2644 5400 2676
rect 5360 2596 5400 2644
rect 5360 2564 5364 2596
rect 5396 2564 5400 2596
rect 5360 2516 5400 2564
rect 5360 2484 5364 2516
rect 5396 2484 5400 2516
rect 5360 2436 5400 2484
rect 5360 2404 5364 2436
rect 5396 2404 5400 2436
rect 5360 2356 5400 2404
rect 5360 2324 5364 2356
rect 5396 2324 5400 2356
rect 5360 2276 5400 2324
rect 5360 2244 5364 2276
rect 5396 2244 5400 2276
rect 5360 2196 5400 2244
rect 5360 2164 5364 2196
rect 5396 2164 5400 2196
rect 5360 2116 5400 2164
rect 5360 2084 5364 2116
rect 5396 2084 5400 2116
rect 5360 2036 5400 2084
rect 5360 2004 5364 2036
rect 5396 2004 5400 2036
rect 5360 1956 5400 2004
rect 5360 1924 5364 1956
rect 5396 1924 5400 1956
rect 5360 1876 5400 1924
rect 5360 1844 5364 1876
rect 5396 1844 5400 1876
rect 5360 1796 5400 1844
rect 5360 1764 5364 1796
rect 5396 1764 5400 1796
rect 5360 1716 5400 1764
rect 5360 1684 5364 1716
rect 5396 1684 5400 1716
rect 5360 1636 5400 1684
rect 5360 1604 5364 1636
rect 5396 1604 5400 1636
rect 5360 1556 5400 1604
rect 5360 1524 5364 1556
rect 5396 1524 5400 1556
rect 5360 1476 5400 1524
rect 5360 1444 5364 1476
rect 5396 1444 5400 1476
rect 5360 1396 5400 1444
rect 5360 1364 5364 1396
rect 5396 1364 5400 1396
rect 5360 1316 5400 1364
rect 5360 1284 5364 1316
rect 5396 1284 5400 1316
rect 5360 1236 5400 1284
rect 5360 1204 5364 1236
rect 5396 1204 5400 1236
rect 5360 1156 5400 1204
rect 5360 1124 5364 1156
rect 5396 1124 5400 1156
rect 5360 1076 5400 1124
rect 5360 1044 5364 1076
rect 5396 1044 5400 1076
rect 5360 996 5400 1044
rect 5360 964 5364 996
rect 5396 964 5400 996
rect 5360 916 5400 964
rect 5360 884 5364 916
rect 5396 884 5400 916
rect 5360 836 5400 884
rect 5360 804 5364 836
rect 5396 804 5400 836
rect 5360 756 5400 804
rect 5360 724 5364 756
rect 5396 724 5400 756
rect 5360 676 5400 724
rect 5360 644 5364 676
rect 5396 644 5400 676
rect 5360 596 5400 644
rect 5360 564 5364 596
rect 5396 564 5400 596
rect 5360 516 5400 564
rect 5360 484 5364 516
rect 5396 484 5400 516
rect 5360 436 5400 484
rect 5360 404 5364 436
rect 5396 404 5400 436
rect 5360 356 5400 404
rect 5360 324 5364 356
rect 5396 324 5400 356
rect 5360 276 5400 324
rect 5360 244 5364 276
rect 5396 244 5400 276
rect 5360 196 5400 244
rect 5360 164 5364 196
rect 5396 164 5400 196
rect 5360 116 5400 164
rect 5360 84 5364 116
rect 5396 84 5400 116
rect 5360 36 5400 84
rect 5360 4 5364 36
rect 5396 4 5400 36
rect 5200 -716 5204 -524
rect 5236 -716 5240 -524
rect 5200 -960 5240 -716
rect 5360 -524 5400 4
rect 5440 14155 5480 15760
rect 5440 14125 5445 14155
rect 5475 14125 5480 14155
rect 5440 9115 5480 14125
rect 5440 9085 5445 9115
rect 5475 9085 5480 9115
rect 5440 5995 5480 9085
rect 5440 5965 5445 5995
rect 5475 5965 5480 5995
rect 5440 0 5480 5965
rect 5520 15716 5560 15760
rect 5520 15684 5524 15716
rect 5556 15684 5560 15716
rect 5520 15636 5560 15684
rect 5520 15604 5524 15636
rect 5556 15604 5560 15636
rect 5520 15556 5560 15604
rect 5520 15524 5524 15556
rect 5556 15524 5560 15556
rect 5520 15476 5560 15524
rect 5520 15444 5524 15476
rect 5556 15444 5560 15476
rect 5520 15396 5560 15444
rect 5520 15364 5524 15396
rect 5556 15364 5560 15396
rect 5520 15316 5560 15364
rect 5520 15284 5524 15316
rect 5556 15284 5560 15316
rect 5520 15236 5560 15284
rect 5520 15204 5524 15236
rect 5556 15204 5560 15236
rect 5520 15156 5560 15204
rect 5520 15124 5524 15156
rect 5556 15124 5560 15156
rect 5520 15076 5560 15124
rect 5520 15044 5524 15076
rect 5556 15044 5560 15076
rect 5520 14996 5560 15044
rect 5520 14964 5524 14996
rect 5556 14964 5560 14996
rect 5520 14916 5560 14964
rect 5520 14884 5524 14916
rect 5556 14884 5560 14916
rect 5520 14836 5560 14884
rect 5520 14804 5524 14836
rect 5556 14804 5560 14836
rect 5520 14756 5560 14804
rect 5520 14724 5524 14756
rect 5556 14724 5560 14756
rect 5520 14676 5560 14724
rect 5520 14644 5524 14676
rect 5556 14644 5560 14676
rect 5520 14596 5560 14644
rect 5520 14564 5524 14596
rect 5556 14564 5560 14596
rect 5520 14516 5560 14564
rect 5520 14484 5524 14516
rect 5556 14484 5560 14516
rect 5520 14436 5560 14484
rect 5520 14404 5524 14436
rect 5556 14404 5560 14436
rect 5520 14356 5560 14404
rect 5520 14324 5524 14356
rect 5556 14324 5560 14356
rect 5520 14276 5560 14324
rect 5520 14244 5524 14276
rect 5556 14244 5560 14276
rect 5520 14196 5560 14244
rect 5520 14164 5524 14196
rect 5556 14164 5560 14196
rect 5520 14116 5560 14164
rect 5520 14084 5524 14116
rect 5556 14084 5560 14116
rect 5520 14036 5560 14084
rect 5520 14004 5524 14036
rect 5556 14004 5560 14036
rect 5520 13956 5560 14004
rect 5520 13924 5524 13956
rect 5556 13924 5560 13956
rect 5520 13876 5560 13924
rect 5520 13844 5524 13876
rect 5556 13844 5560 13876
rect 5520 13796 5560 13844
rect 5520 13764 5524 13796
rect 5556 13764 5560 13796
rect 5520 13716 5560 13764
rect 5520 13684 5524 13716
rect 5556 13684 5560 13716
rect 5520 13636 5560 13684
rect 5520 13604 5524 13636
rect 5556 13604 5560 13636
rect 5520 13556 5560 13604
rect 5520 13524 5524 13556
rect 5556 13524 5560 13556
rect 5520 13476 5560 13524
rect 5520 13444 5524 13476
rect 5556 13444 5560 13476
rect 5520 13396 5560 13444
rect 5520 13364 5524 13396
rect 5556 13364 5560 13396
rect 5520 13316 5560 13364
rect 5520 13284 5524 13316
rect 5556 13284 5560 13316
rect 5520 13236 5560 13284
rect 5520 13204 5524 13236
rect 5556 13204 5560 13236
rect 5520 13156 5560 13204
rect 5520 13124 5524 13156
rect 5556 13124 5560 13156
rect 5520 13076 5560 13124
rect 5520 13044 5524 13076
rect 5556 13044 5560 13076
rect 5520 12996 5560 13044
rect 5520 12964 5524 12996
rect 5556 12964 5560 12996
rect 5520 12916 5560 12964
rect 5520 12884 5524 12916
rect 5556 12884 5560 12916
rect 5520 12836 5560 12884
rect 5520 12804 5524 12836
rect 5556 12804 5560 12836
rect 5520 12756 5560 12804
rect 5520 12724 5524 12756
rect 5556 12724 5560 12756
rect 5520 12676 5560 12724
rect 5520 12644 5524 12676
rect 5556 12644 5560 12676
rect 5520 12596 5560 12644
rect 5520 12564 5524 12596
rect 5556 12564 5560 12596
rect 5520 12516 5560 12564
rect 5520 12484 5524 12516
rect 5556 12484 5560 12516
rect 5520 12436 5560 12484
rect 5520 12404 5524 12436
rect 5556 12404 5560 12436
rect 5520 12356 5560 12404
rect 5520 12324 5524 12356
rect 5556 12324 5560 12356
rect 5520 12276 5560 12324
rect 5520 12244 5524 12276
rect 5556 12244 5560 12276
rect 5520 12196 5560 12244
rect 5520 12164 5524 12196
rect 5556 12164 5560 12196
rect 5520 12116 5560 12164
rect 5520 12084 5524 12116
rect 5556 12084 5560 12116
rect 5520 12036 5560 12084
rect 5520 12004 5524 12036
rect 5556 12004 5560 12036
rect 5520 11956 5560 12004
rect 5520 11924 5524 11956
rect 5556 11924 5560 11956
rect 5520 11876 5560 11924
rect 5520 11844 5524 11876
rect 5556 11844 5560 11876
rect 5520 11796 5560 11844
rect 5520 11764 5524 11796
rect 5556 11764 5560 11796
rect 5520 11716 5560 11764
rect 5520 11684 5524 11716
rect 5556 11684 5560 11716
rect 5520 11636 5560 11684
rect 5520 11604 5524 11636
rect 5556 11604 5560 11636
rect 5520 11556 5560 11604
rect 5520 11524 5524 11556
rect 5556 11524 5560 11556
rect 5520 11476 5560 11524
rect 5520 11444 5524 11476
rect 5556 11444 5560 11476
rect 5520 11396 5560 11444
rect 5520 11364 5524 11396
rect 5556 11364 5560 11396
rect 5520 11316 5560 11364
rect 5520 11284 5524 11316
rect 5556 11284 5560 11316
rect 5520 11236 5560 11284
rect 5520 11204 5524 11236
rect 5556 11204 5560 11236
rect 5520 11156 5560 11204
rect 5520 11124 5524 11156
rect 5556 11124 5560 11156
rect 5520 11076 5560 11124
rect 5520 11044 5524 11076
rect 5556 11044 5560 11076
rect 5520 10996 5560 11044
rect 5520 10964 5524 10996
rect 5556 10964 5560 10996
rect 5520 10916 5560 10964
rect 5520 10884 5524 10916
rect 5556 10884 5560 10916
rect 5520 10836 5560 10884
rect 5520 10804 5524 10836
rect 5556 10804 5560 10836
rect 5520 10756 5560 10804
rect 5520 10724 5524 10756
rect 5556 10724 5560 10756
rect 5520 10676 5560 10724
rect 5520 10644 5524 10676
rect 5556 10644 5560 10676
rect 5520 10596 5560 10644
rect 5520 10564 5524 10596
rect 5556 10564 5560 10596
rect 5520 10516 5560 10564
rect 5520 10484 5524 10516
rect 5556 10484 5560 10516
rect 5520 10436 5560 10484
rect 5520 10404 5524 10436
rect 5556 10404 5560 10436
rect 5520 10356 5560 10404
rect 5520 10324 5524 10356
rect 5556 10324 5560 10356
rect 5520 10276 5560 10324
rect 5520 10244 5524 10276
rect 5556 10244 5560 10276
rect 5520 10196 5560 10244
rect 5520 10164 5524 10196
rect 5556 10164 5560 10196
rect 5520 10116 5560 10164
rect 5520 10084 5524 10116
rect 5556 10084 5560 10116
rect 5520 10036 5560 10084
rect 5520 10004 5524 10036
rect 5556 10004 5560 10036
rect 5520 9956 5560 10004
rect 5520 9924 5524 9956
rect 5556 9924 5560 9956
rect 5520 9876 5560 9924
rect 5520 9844 5524 9876
rect 5556 9844 5560 9876
rect 5520 9796 5560 9844
rect 5520 9764 5524 9796
rect 5556 9764 5560 9796
rect 5520 9716 5560 9764
rect 5520 9684 5524 9716
rect 5556 9684 5560 9716
rect 5520 9636 5560 9684
rect 5520 9604 5524 9636
rect 5556 9604 5560 9636
rect 5520 9556 5560 9604
rect 5520 9524 5524 9556
rect 5556 9524 5560 9556
rect 5520 9476 5560 9524
rect 5520 9444 5524 9476
rect 5556 9444 5560 9476
rect 5520 9396 5560 9444
rect 5520 9364 5524 9396
rect 5556 9364 5560 9396
rect 5520 9316 5560 9364
rect 5520 9284 5524 9316
rect 5556 9284 5560 9316
rect 5520 9236 5560 9284
rect 5520 9204 5524 9236
rect 5556 9204 5560 9236
rect 5520 9156 5560 9204
rect 5520 9124 5524 9156
rect 5556 9124 5560 9156
rect 5520 9076 5560 9124
rect 5520 9044 5524 9076
rect 5556 9044 5560 9076
rect 5520 8996 5560 9044
rect 5520 8964 5524 8996
rect 5556 8964 5560 8996
rect 5520 8916 5560 8964
rect 5520 8884 5524 8916
rect 5556 8884 5560 8916
rect 5520 8836 5560 8884
rect 5520 8804 5524 8836
rect 5556 8804 5560 8836
rect 5520 8756 5560 8804
rect 5520 8724 5524 8756
rect 5556 8724 5560 8756
rect 5520 8676 5560 8724
rect 5520 8644 5524 8676
rect 5556 8644 5560 8676
rect 5520 8596 5560 8644
rect 5520 8564 5524 8596
rect 5556 8564 5560 8596
rect 5520 8516 5560 8564
rect 5520 8484 5524 8516
rect 5556 8484 5560 8516
rect 5520 8436 5560 8484
rect 5520 8404 5524 8436
rect 5556 8404 5560 8436
rect 5520 8356 5560 8404
rect 5520 8324 5524 8356
rect 5556 8324 5560 8356
rect 5520 8276 5560 8324
rect 5520 8244 5524 8276
rect 5556 8244 5560 8276
rect 5520 8196 5560 8244
rect 5520 8164 5524 8196
rect 5556 8164 5560 8196
rect 5520 8116 5560 8164
rect 5520 8084 5524 8116
rect 5556 8084 5560 8116
rect 5520 8036 5560 8084
rect 5520 8004 5524 8036
rect 5556 8004 5560 8036
rect 5520 7956 5560 8004
rect 5520 7924 5524 7956
rect 5556 7924 5560 7956
rect 5520 7876 5560 7924
rect 5520 7844 5524 7876
rect 5556 7844 5560 7876
rect 5520 7796 5560 7844
rect 5520 7764 5524 7796
rect 5556 7764 5560 7796
rect 5520 7716 5560 7764
rect 5520 7684 5524 7716
rect 5556 7684 5560 7716
rect 5520 7636 5560 7684
rect 5520 7604 5524 7636
rect 5556 7604 5560 7636
rect 5520 7556 5560 7604
rect 5520 7524 5524 7556
rect 5556 7524 5560 7556
rect 5520 7476 5560 7524
rect 5520 7444 5524 7476
rect 5556 7444 5560 7476
rect 5520 7396 5560 7444
rect 5520 7364 5524 7396
rect 5556 7364 5560 7396
rect 5520 7316 5560 7364
rect 5520 7284 5524 7316
rect 5556 7284 5560 7316
rect 5520 7236 5560 7284
rect 5520 7204 5524 7236
rect 5556 7204 5560 7236
rect 5520 7156 5560 7204
rect 5520 7124 5524 7156
rect 5556 7124 5560 7156
rect 5520 7076 5560 7124
rect 5520 7044 5524 7076
rect 5556 7044 5560 7076
rect 5520 6996 5560 7044
rect 5520 6964 5524 6996
rect 5556 6964 5560 6996
rect 5520 6916 5560 6964
rect 5520 6884 5524 6916
rect 5556 6884 5560 6916
rect 5520 6836 5560 6884
rect 5520 6804 5524 6836
rect 5556 6804 5560 6836
rect 5520 6756 5560 6804
rect 5520 6724 5524 6756
rect 5556 6724 5560 6756
rect 5520 6676 5560 6724
rect 5520 6644 5524 6676
rect 5556 6644 5560 6676
rect 5520 6596 5560 6644
rect 5520 6564 5524 6596
rect 5556 6564 5560 6596
rect 5520 6516 5560 6564
rect 5520 6484 5524 6516
rect 5556 6484 5560 6516
rect 5520 6436 5560 6484
rect 5520 6404 5524 6436
rect 5556 6404 5560 6436
rect 5520 6356 5560 6404
rect 5520 6324 5524 6356
rect 5556 6324 5560 6356
rect 5520 6276 5560 6324
rect 5520 6244 5524 6276
rect 5556 6244 5560 6276
rect 5520 6196 5560 6244
rect 5520 6164 5524 6196
rect 5556 6164 5560 6196
rect 5520 6116 5560 6164
rect 5520 6084 5524 6116
rect 5556 6084 5560 6116
rect 5520 6036 5560 6084
rect 5520 6004 5524 6036
rect 5556 6004 5560 6036
rect 5520 5956 5560 6004
rect 5520 5924 5524 5956
rect 5556 5924 5560 5956
rect 5520 5876 5560 5924
rect 5520 5844 5524 5876
rect 5556 5844 5560 5876
rect 5520 5796 5560 5844
rect 5520 5764 5524 5796
rect 5556 5764 5560 5796
rect 5520 5716 5560 5764
rect 5520 5684 5524 5716
rect 5556 5684 5560 5716
rect 5520 5636 5560 5684
rect 5520 5604 5524 5636
rect 5556 5604 5560 5636
rect 5520 5556 5560 5604
rect 5520 5524 5524 5556
rect 5556 5524 5560 5556
rect 5520 5476 5560 5524
rect 5520 5444 5524 5476
rect 5556 5444 5560 5476
rect 5520 5396 5560 5444
rect 5520 5364 5524 5396
rect 5556 5364 5560 5396
rect 5520 5316 5560 5364
rect 5520 5284 5524 5316
rect 5556 5284 5560 5316
rect 5520 5236 5560 5284
rect 5520 5204 5524 5236
rect 5556 5204 5560 5236
rect 5520 5156 5560 5204
rect 5520 5124 5524 5156
rect 5556 5124 5560 5156
rect 5520 5076 5560 5124
rect 5520 5044 5524 5076
rect 5556 5044 5560 5076
rect 5520 4996 5560 5044
rect 5520 4964 5524 4996
rect 5556 4964 5560 4996
rect 5520 4916 5560 4964
rect 5520 4884 5524 4916
rect 5556 4884 5560 4916
rect 5520 4836 5560 4884
rect 5520 4804 5524 4836
rect 5556 4804 5560 4836
rect 5520 4756 5560 4804
rect 5520 4724 5524 4756
rect 5556 4724 5560 4756
rect 5520 4676 5560 4724
rect 5520 4644 5524 4676
rect 5556 4644 5560 4676
rect 5520 4596 5560 4644
rect 5520 4564 5524 4596
rect 5556 4564 5560 4596
rect 5520 4516 5560 4564
rect 5520 4484 5524 4516
rect 5556 4484 5560 4516
rect 5520 4436 5560 4484
rect 5520 4404 5524 4436
rect 5556 4404 5560 4436
rect 5520 4356 5560 4404
rect 5520 4324 5524 4356
rect 5556 4324 5560 4356
rect 5520 4276 5560 4324
rect 5520 4244 5524 4276
rect 5556 4244 5560 4276
rect 5520 4196 5560 4244
rect 5520 4164 5524 4196
rect 5556 4164 5560 4196
rect 5520 4116 5560 4164
rect 5520 4084 5524 4116
rect 5556 4084 5560 4116
rect 5520 4036 5560 4084
rect 5520 4004 5524 4036
rect 5556 4004 5560 4036
rect 5520 3956 5560 4004
rect 5520 3924 5524 3956
rect 5556 3924 5560 3956
rect 5520 3876 5560 3924
rect 5520 3844 5524 3876
rect 5556 3844 5560 3876
rect 5520 3796 5560 3844
rect 5520 3764 5524 3796
rect 5556 3764 5560 3796
rect 5520 3716 5560 3764
rect 5520 3684 5524 3716
rect 5556 3684 5560 3716
rect 5520 3636 5560 3684
rect 5520 3604 5524 3636
rect 5556 3604 5560 3636
rect 5520 3556 5560 3604
rect 5520 3524 5524 3556
rect 5556 3524 5560 3556
rect 5520 3476 5560 3524
rect 5520 3444 5524 3476
rect 5556 3444 5560 3476
rect 5520 3396 5560 3444
rect 5520 3364 5524 3396
rect 5556 3364 5560 3396
rect 5520 3316 5560 3364
rect 5520 3284 5524 3316
rect 5556 3284 5560 3316
rect 5520 3236 5560 3284
rect 5520 3204 5524 3236
rect 5556 3204 5560 3236
rect 5520 3156 5560 3204
rect 5520 3124 5524 3156
rect 5556 3124 5560 3156
rect 5520 3076 5560 3124
rect 5520 3044 5524 3076
rect 5556 3044 5560 3076
rect 5520 2996 5560 3044
rect 5520 2964 5524 2996
rect 5556 2964 5560 2996
rect 5520 2916 5560 2964
rect 5520 2884 5524 2916
rect 5556 2884 5560 2916
rect 5520 2836 5560 2884
rect 5520 2804 5524 2836
rect 5556 2804 5560 2836
rect 5520 2756 5560 2804
rect 5520 2724 5524 2756
rect 5556 2724 5560 2756
rect 5520 2676 5560 2724
rect 5520 2644 5524 2676
rect 5556 2644 5560 2676
rect 5520 2596 5560 2644
rect 5520 2564 5524 2596
rect 5556 2564 5560 2596
rect 5520 2516 5560 2564
rect 5520 2484 5524 2516
rect 5556 2484 5560 2516
rect 5520 2436 5560 2484
rect 5520 2404 5524 2436
rect 5556 2404 5560 2436
rect 5520 2356 5560 2404
rect 5520 2324 5524 2356
rect 5556 2324 5560 2356
rect 5520 2276 5560 2324
rect 5520 2244 5524 2276
rect 5556 2244 5560 2276
rect 5520 2196 5560 2244
rect 5520 2164 5524 2196
rect 5556 2164 5560 2196
rect 5520 2116 5560 2164
rect 5520 2084 5524 2116
rect 5556 2084 5560 2116
rect 5520 2036 5560 2084
rect 5520 2004 5524 2036
rect 5556 2004 5560 2036
rect 5520 1956 5560 2004
rect 5520 1924 5524 1956
rect 5556 1924 5560 1956
rect 5520 1876 5560 1924
rect 5520 1844 5524 1876
rect 5556 1844 5560 1876
rect 5520 1796 5560 1844
rect 5520 1764 5524 1796
rect 5556 1764 5560 1796
rect 5520 1716 5560 1764
rect 5520 1684 5524 1716
rect 5556 1684 5560 1716
rect 5520 1636 5560 1684
rect 5520 1604 5524 1636
rect 5556 1604 5560 1636
rect 5520 1556 5560 1604
rect 5520 1524 5524 1556
rect 5556 1524 5560 1556
rect 5520 1476 5560 1524
rect 5520 1444 5524 1476
rect 5556 1444 5560 1476
rect 5520 1396 5560 1444
rect 5520 1364 5524 1396
rect 5556 1364 5560 1396
rect 5520 1316 5560 1364
rect 5520 1284 5524 1316
rect 5556 1284 5560 1316
rect 5520 1236 5560 1284
rect 5520 1204 5524 1236
rect 5556 1204 5560 1236
rect 5520 1156 5560 1204
rect 5520 1124 5524 1156
rect 5556 1124 5560 1156
rect 5520 1076 5560 1124
rect 5520 1044 5524 1076
rect 5556 1044 5560 1076
rect 5520 996 5560 1044
rect 5520 964 5524 996
rect 5556 964 5560 996
rect 5520 916 5560 964
rect 5520 884 5524 916
rect 5556 884 5560 916
rect 5520 836 5560 884
rect 5520 804 5524 836
rect 5556 804 5560 836
rect 5520 756 5560 804
rect 5520 724 5524 756
rect 5556 724 5560 756
rect 5520 676 5560 724
rect 5520 644 5524 676
rect 5556 644 5560 676
rect 5520 596 5560 644
rect 5520 564 5524 596
rect 5556 564 5560 596
rect 5520 516 5560 564
rect 5520 484 5524 516
rect 5556 484 5560 516
rect 5520 436 5560 484
rect 5520 404 5524 436
rect 5556 404 5560 436
rect 5520 356 5560 404
rect 5520 324 5524 356
rect 5556 324 5560 356
rect 5520 276 5560 324
rect 5520 244 5524 276
rect 5556 244 5560 276
rect 5520 196 5560 244
rect 5520 164 5524 196
rect 5556 164 5560 196
rect 5520 116 5560 164
rect 5520 84 5524 116
rect 5556 84 5560 116
rect 5520 36 5560 84
rect 5520 4 5524 36
rect 5556 4 5560 36
rect 5360 -716 5364 -524
rect 5396 -716 5400 -524
rect 5360 -960 5400 -716
rect 5520 -524 5560 4
rect 5600 6155 5640 15760
rect 5600 6125 5605 6155
rect 5635 6125 5640 6155
rect 5600 0 5640 6125
rect 5680 15716 5720 15760
rect 5680 15684 5684 15716
rect 5716 15684 5720 15716
rect 5680 15636 5720 15684
rect 5680 15604 5684 15636
rect 5716 15604 5720 15636
rect 5680 15556 5720 15604
rect 5680 15524 5684 15556
rect 5716 15524 5720 15556
rect 5680 15476 5720 15524
rect 5680 15444 5684 15476
rect 5716 15444 5720 15476
rect 5680 15396 5720 15444
rect 5680 15364 5684 15396
rect 5716 15364 5720 15396
rect 5680 15316 5720 15364
rect 5680 15284 5684 15316
rect 5716 15284 5720 15316
rect 5680 15236 5720 15284
rect 5680 15204 5684 15236
rect 5716 15204 5720 15236
rect 5680 15156 5720 15204
rect 5680 15124 5684 15156
rect 5716 15124 5720 15156
rect 5680 15076 5720 15124
rect 5680 15044 5684 15076
rect 5716 15044 5720 15076
rect 5680 14996 5720 15044
rect 5680 14964 5684 14996
rect 5716 14964 5720 14996
rect 5680 14916 5720 14964
rect 5680 14884 5684 14916
rect 5716 14884 5720 14916
rect 5680 14836 5720 14884
rect 5680 14804 5684 14836
rect 5716 14804 5720 14836
rect 5680 14756 5720 14804
rect 5680 14724 5684 14756
rect 5716 14724 5720 14756
rect 5680 14676 5720 14724
rect 5680 14644 5684 14676
rect 5716 14644 5720 14676
rect 5680 14596 5720 14644
rect 5680 14564 5684 14596
rect 5716 14564 5720 14596
rect 5680 14516 5720 14564
rect 5680 14484 5684 14516
rect 5716 14484 5720 14516
rect 5680 14436 5720 14484
rect 5680 14404 5684 14436
rect 5716 14404 5720 14436
rect 5680 14356 5720 14404
rect 5680 14324 5684 14356
rect 5716 14324 5720 14356
rect 5680 14276 5720 14324
rect 5680 14244 5684 14276
rect 5716 14244 5720 14276
rect 5680 14196 5720 14244
rect 5680 14164 5684 14196
rect 5716 14164 5720 14196
rect 5680 14116 5720 14164
rect 5680 14084 5684 14116
rect 5716 14084 5720 14116
rect 5680 14036 5720 14084
rect 5680 14004 5684 14036
rect 5716 14004 5720 14036
rect 5680 13956 5720 14004
rect 5680 13924 5684 13956
rect 5716 13924 5720 13956
rect 5680 13876 5720 13924
rect 5680 13844 5684 13876
rect 5716 13844 5720 13876
rect 5680 13796 5720 13844
rect 5680 13764 5684 13796
rect 5716 13764 5720 13796
rect 5680 13716 5720 13764
rect 5680 13684 5684 13716
rect 5716 13684 5720 13716
rect 5680 13636 5720 13684
rect 5680 13604 5684 13636
rect 5716 13604 5720 13636
rect 5680 13556 5720 13604
rect 5680 13524 5684 13556
rect 5716 13524 5720 13556
rect 5680 13476 5720 13524
rect 5680 13444 5684 13476
rect 5716 13444 5720 13476
rect 5680 13396 5720 13444
rect 5680 13364 5684 13396
rect 5716 13364 5720 13396
rect 5680 13316 5720 13364
rect 5680 13284 5684 13316
rect 5716 13284 5720 13316
rect 5680 13236 5720 13284
rect 5680 13204 5684 13236
rect 5716 13204 5720 13236
rect 5680 13156 5720 13204
rect 5680 13124 5684 13156
rect 5716 13124 5720 13156
rect 5680 13076 5720 13124
rect 5680 13044 5684 13076
rect 5716 13044 5720 13076
rect 5680 12996 5720 13044
rect 5680 12964 5684 12996
rect 5716 12964 5720 12996
rect 5680 12916 5720 12964
rect 5680 12884 5684 12916
rect 5716 12884 5720 12916
rect 5680 12836 5720 12884
rect 5680 12804 5684 12836
rect 5716 12804 5720 12836
rect 5680 12756 5720 12804
rect 5680 12724 5684 12756
rect 5716 12724 5720 12756
rect 5680 12676 5720 12724
rect 5680 12644 5684 12676
rect 5716 12644 5720 12676
rect 5680 12596 5720 12644
rect 5680 12564 5684 12596
rect 5716 12564 5720 12596
rect 5680 12516 5720 12564
rect 5680 12484 5684 12516
rect 5716 12484 5720 12516
rect 5680 12436 5720 12484
rect 5680 12404 5684 12436
rect 5716 12404 5720 12436
rect 5680 12356 5720 12404
rect 5680 12324 5684 12356
rect 5716 12324 5720 12356
rect 5680 12276 5720 12324
rect 5680 12244 5684 12276
rect 5716 12244 5720 12276
rect 5680 12196 5720 12244
rect 5680 12164 5684 12196
rect 5716 12164 5720 12196
rect 5680 12116 5720 12164
rect 5680 12084 5684 12116
rect 5716 12084 5720 12116
rect 5680 12036 5720 12084
rect 5680 12004 5684 12036
rect 5716 12004 5720 12036
rect 5680 11956 5720 12004
rect 5680 11924 5684 11956
rect 5716 11924 5720 11956
rect 5680 11876 5720 11924
rect 5680 11844 5684 11876
rect 5716 11844 5720 11876
rect 5680 11796 5720 11844
rect 5680 11764 5684 11796
rect 5716 11764 5720 11796
rect 5680 11716 5720 11764
rect 5680 11684 5684 11716
rect 5716 11684 5720 11716
rect 5680 11636 5720 11684
rect 5680 11604 5684 11636
rect 5716 11604 5720 11636
rect 5680 11556 5720 11604
rect 5680 11524 5684 11556
rect 5716 11524 5720 11556
rect 5680 11476 5720 11524
rect 5680 11444 5684 11476
rect 5716 11444 5720 11476
rect 5680 11396 5720 11444
rect 5680 11364 5684 11396
rect 5716 11364 5720 11396
rect 5680 11316 5720 11364
rect 5680 11284 5684 11316
rect 5716 11284 5720 11316
rect 5680 11236 5720 11284
rect 5680 11204 5684 11236
rect 5716 11204 5720 11236
rect 5680 11156 5720 11204
rect 5680 11124 5684 11156
rect 5716 11124 5720 11156
rect 5680 11076 5720 11124
rect 5680 11044 5684 11076
rect 5716 11044 5720 11076
rect 5680 10996 5720 11044
rect 5680 10964 5684 10996
rect 5716 10964 5720 10996
rect 5680 10916 5720 10964
rect 5680 10884 5684 10916
rect 5716 10884 5720 10916
rect 5680 10836 5720 10884
rect 5680 10804 5684 10836
rect 5716 10804 5720 10836
rect 5680 10756 5720 10804
rect 5680 10724 5684 10756
rect 5716 10724 5720 10756
rect 5680 10676 5720 10724
rect 5680 10644 5684 10676
rect 5716 10644 5720 10676
rect 5680 10596 5720 10644
rect 5680 10564 5684 10596
rect 5716 10564 5720 10596
rect 5680 10516 5720 10564
rect 5680 10484 5684 10516
rect 5716 10484 5720 10516
rect 5680 10436 5720 10484
rect 5680 10404 5684 10436
rect 5716 10404 5720 10436
rect 5680 10356 5720 10404
rect 5680 10324 5684 10356
rect 5716 10324 5720 10356
rect 5680 10276 5720 10324
rect 5680 10244 5684 10276
rect 5716 10244 5720 10276
rect 5680 10196 5720 10244
rect 5680 10164 5684 10196
rect 5716 10164 5720 10196
rect 5680 10116 5720 10164
rect 5680 10084 5684 10116
rect 5716 10084 5720 10116
rect 5680 10036 5720 10084
rect 5680 10004 5684 10036
rect 5716 10004 5720 10036
rect 5680 9956 5720 10004
rect 5680 9924 5684 9956
rect 5716 9924 5720 9956
rect 5680 9876 5720 9924
rect 5680 9844 5684 9876
rect 5716 9844 5720 9876
rect 5680 9796 5720 9844
rect 5680 9764 5684 9796
rect 5716 9764 5720 9796
rect 5680 9716 5720 9764
rect 5680 9684 5684 9716
rect 5716 9684 5720 9716
rect 5680 9636 5720 9684
rect 5680 9604 5684 9636
rect 5716 9604 5720 9636
rect 5680 9556 5720 9604
rect 5680 9524 5684 9556
rect 5716 9524 5720 9556
rect 5680 9476 5720 9524
rect 5680 9444 5684 9476
rect 5716 9444 5720 9476
rect 5680 9396 5720 9444
rect 5680 9364 5684 9396
rect 5716 9364 5720 9396
rect 5680 9316 5720 9364
rect 5680 9284 5684 9316
rect 5716 9284 5720 9316
rect 5680 9236 5720 9284
rect 5680 9204 5684 9236
rect 5716 9204 5720 9236
rect 5680 9156 5720 9204
rect 5680 9124 5684 9156
rect 5716 9124 5720 9156
rect 5680 9076 5720 9124
rect 5680 9044 5684 9076
rect 5716 9044 5720 9076
rect 5680 8996 5720 9044
rect 5680 8964 5684 8996
rect 5716 8964 5720 8996
rect 5680 8916 5720 8964
rect 5680 8884 5684 8916
rect 5716 8884 5720 8916
rect 5680 8836 5720 8884
rect 5680 8804 5684 8836
rect 5716 8804 5720 8836
rect 5680 8756 5720 8804
rect 5680 8724 5684 8756
rect 5716 8724 5720 8756
rect 5680 8676 5720 8724
rect 5680 8644 5684 8676
rect 5716 8644 5720 8676
rect 5680 8596 5720 8644
rect 5680 8564 5684 8596
rect 5716 8564 5720 8596
rect 5680 8516 5720 8564
rect 5680 8484 5684 8516
rect 5716 8484 5720 8516
rect 5680 8436 5720 8484
rect 5680 8404 5684 8436
rect 5716 8404 5720 8436
rect 5680 8356 5720 8404
rect 5680 8324 5684 8356
rect 5716 8324 5720 8356
rect 5680 8276 5720 8324
rect 5680 8244 5684 8276
rect 5716 8244 5720 8276
rect 5680 8196 5720 8244
rect 5680 8164 5684 8196
rect 5716 8164 5720 8196
rect 5680 8116 5720 8164
rect 5680 8084 5684 8116
rect 5716 8084 5720 8116
rect 5680 8036 5720 8084
rect 5680 8004 5684 8036
rect 5716 8004 5720 8036
rect 5680 7956 5720 8004
rect 5680 7924 5684 7956
rect 5716 7924 5720 7956
rect 5680 7876 5720 7924
rect 5680 7844 5684 7876
rect 5716 7844 5720 7876
rect 5680 7796 5720 7844
rect 5680 7764 5684 7796
rect 5716 7764 5720 7796
rect 5680 7716 5720 7764
rect 5680 7684 5684 7716
rect 5716 7684 5720 7716
rect 5680 7636 5720 7684
rect 5680 7604 5684 7636
rect 5716 7604 5720 7636
rect 5680 7556 5720 7604
rect 5680 7524 5684 7556
rect 5716 7524 5720 7556
rect 5680 7476 5720 7524
rect 5680 7444 5684 7476
rect 5716 7444 5720 7476
rect 5680 7396 5720 7444
rect 5680 7364 5684 7396
rect 5716 7364 5720 7396
rect 5680 7316 5720 7364
rect 5680 7284 5684 7316
rect 5716 7284 5720 7316
rect 5680 7236 5720 7284
rect 5680 7204 5684 7236
rect 5716 7204 5720 7236
rect 5680 7156 5720 7204
rect 5680 7124 5684 7156
rect 5716 7124 5720 7156
rect 5680 7076 5720 7124
rect 5680 7044 5684 7076
rect 5716 7044 5720 7076
rect 5680 6996 5720 7044
rect 5680 6964 5684 6996
rect 5716 6964 5720 6996
rect 5680 6916 5720 6964
rect 5680 6884 5684 6916
rect 5716 6884 5720 6916
rect 5680 6836 5720 6884
rect 5680 6804 5684 6836
rect 5716 6804 5720 6836
rect 5680 6756 5720 6804
rect 5680 6724 5684 6756
rect 5716 6724 5720 6756
rect 5680 6676 5720 6724
rect 5680 6644 5684 6676
rect 5716 6644 5720 6676
rect 5680 6596 5720 6644
rect 5680 6564 5684 6596
rect 5716 6564 5720 6596
rect 5680 6516 5720 6564
rect 5680 6484 5684 6516
rect 5716 6484 5720 6516
rect 5680 6436 5720 6484
rect 5680 6404 5684 6436
rect 5716 6404 5720 6436
rect 5680 6356 5720 6404
rect 5680 6324 5684 6356
rect 5716 6324 5720 6356
rect 5680 6276 5720 6324
rect 5680 6244 5684 6276
rect 5716 6244 5720 6276
rect 5680 6196 5720 6244
rect 5680 6164 5684 6196
rect 5716 6164 5720 6196
rect 5680 6116 5720 6164
rect 5680 6084 5684 6116
rect 5716 6084 5720 6116
rect 5680 6036 5720 6084
rect 5680 6004 5684 6036
rect 5716 6004 5720 6036
rect 5680 5956 5720 6004
rect 5680 5924 5684 5956
rect 5716 5924 5720 5956
rect 5680 5876 5720 5924
rect 5680 5844 5684 5876
rect 5716 5844 5720 5876
rect 5680 5796 5720 5844
rect 5680 5764 5684 5796
rect 5716 5764 5720 5796
rect 5680 5716 5720 5764
rect 5680 5684 5684 5716
rect 5716 5684 5720 5716
rect 5680 5636 5720 5684
rect 5680 5604 5684 5636
rect 5716 5604 5720 5636
rect 5680 5556 5720 5604
rect 5680 5524 5684 5556
rect 5716 5524 5720 5556
rect 5680 5476 5720 5524
rect 5680 5444 5684 5476
rect 5716 5444 5720 5476
rect 5680 5396 5720 5444
rect 5680 5364 5684 5396
rect 5716 5364 5720 5396
rect 5680 5316 5720 5364
rect 5680 5284 5684 5316
rect 5716 5284 5720 5316
rect 5680 5236 5720 5284
rect 5680 5204 5684 5236
rect 5716 5204 5720 5236
rect 5680 5156 5720 5204
rect 5680 5124 5684 5156
rect 5716 5124 5720 5156
rect 5680 5076 5720 5124
rect 5680 5044 5684 5076
rect 5716 5044 5720 5076
rect 5680 4996 5720 5044
rect 5680 4964 5684 4996
rect 5716 4964 5720 4996
rect 5680 4916 5720 4964
rect 5680 4884 5684 4916
rect 5716 4884 5720 4916
rect 5680 4836 5720 4884
rect 5680 4804 5684 4836
rect 5716 4804 5720 4836
rect 5680 4756 5720 4804
rect 5680 4724 5684 4756
rect 5716 4724 5720 4756
rect 5680 4676 5720 4724
rect 5680 4644 5684 4676
rect 5716 4644 5720 4676
rect 5680 4596 5720 4644
rect 5680 4564 5684 4596
rect 5716 4564 5720 4596
rect 5680 4516 5720 4564
rect 5680 4484 5684 4516
rect 5716 4484 5720 4516
rect 5680 4436 5720 4484
rect 5680 4404 5684 4436
rect 5716 4404 5720 4436
rect 5680 4356 5720 4404
rect 5680 4324 5684 4356
rect 5716 4324 5720 4356
rect 5680 4276 5720 4324
rect 5680 4244 5684 4276
rect 5716 4244 5720 4276
rect 5680 4196 5720 4244
rect 5680 4164 5684 4196
rect 5716 4164 5720 4196
rect 5680 4116 5720 4164
rect 5680 4084 5684 4116
rect 5716 4084 5720 4116
rect 5680 4036 5720 4084
rect 5680 4004 5684 4036
rect 5716 4004 5720 4036
rect 5680 3956 5720 4004
rect 5680 3924 5684 3956
rect 5716 3924 5720 3956
rect 5680 3876 5720 3924
rect 5680 3844 5684 3876
rect 5716 3844 5720 3876
rect 5680 3796 5720 3844
rect 5680 3764 5684 3796
rect 5716 3764 5720 3796
rect 5680 3716 5720 3764
rect 5680 3684 5684 3716
rect 5716 3684 5720 3716
rect 5680 3636 5720 3684
rect 5680 3604 5684 3636
rect 5716 3604 5720 3636
rect 5680 3556 5720 3604
rect 5680 3524 5684 3556
rect 5716 3524 5720 3556
rect 5680 3476 5720 3524
rect 5680 3444 5684 3476
rect 5716 3444 5720 3476
rect 5680 3396 5720 3444
rect 5680 3364 5684 3396
rect 5716 3364 5720 3396
rect 5680 3316 5720 3364
rect 5680 3284 5684 3316
rect 5716 3284 5720 3316
rect 5680 3236 5720 3284
rect 5680 3204 5684 3236
rect 5716 3204 5720 3236
rect 5680 3156 5720 3204
rect 5680 3124 5684 3156
rect 5716 3124 5720 3156
rect 5680 3076 5720 3124
rect 5680 3044 5684 3076
rect 5716 3044 5720 3076
rect 5680 2996 5720 3044
rect 5680 2964 5684 2996
rect 5716 2964 5720 2996
rect 5680 2916 5720 2964
rect 5680 2884 5684 2916
rect 5716 2884 5720 2916
rect 5680 2836 5720 2884
rect 5680 2804 5684 2836
rect 5716 2804 5720 2836
rect 5680 2756 5720 2804
rect 5680 2724 5684 2756
rect 5716 2724 5720 2756
rect 5680 2676 5720 2724
rect 5680 2644 5684 2676
rect 5716 2644 5720 2676
rect 5680 2596 5720 2644
rect 5680 2564 5684 2596
rect 5716 2564 5720 2596
rect 5680 2516 5720 2564
rect 5680 2484 5684 2516
rect 5716 2484 5720 2516
rect 5680 2436 5720 2484
rect 5680 2404 5684 2436
rect 5716 2404 5720 2436
rect 5680 2356 5720 2404
rect 5680 2324 5684 2356
rect 5716 2324 5720 2356
rect 5680 2276 5720 2324
rect 5680 2244 5684 2276
rect 5716 2244 5720 2276
rect 5680 2196 5720 2244
rect 5680 2164 5684 2196
rect 5716 2164 5720 2196
rect 5680 2116 5720 2164
rect 5680 2084 5684 2116
rect 5716 2084 5720 2116
rect 5680 2036 5720 2084
rect 5680 2004 5684 2036
rect 5716 2004 5720 2036
rect 5680 1956 5720 2004
rect 5680 1924 5684 1956
rect 5716 1924 5720 1956
rect 5680 1876 5720 1924
rect 5680 1844 5684 1876
rect 5716 1844 5720 1876
rect 5680 1796 5720 1844
rect 5680 1764 5684 1796
rect 5716 1764 5720 1796
rect 5680 1716 5720 1764
rect 5680 1684 5684 1716
rect 5716 1684 5720 1716
rect 5680 1636 5720 1684
rect 5680 1604 5684 1636
rect 5716 1604 5720 1636
rect 5680 1556 5720 1604
rect 5680 1524 5684 1556
rect 5716 1524 5720 1556
rect 5680 1476 5720 1524
rect 5680 1444 5684 1476
rect 5716 1444 5720 1476
rect 5680 1396 5720 1444
rect 5680 1364 5684 1396
rect 5716 1364 5720 1396
rect 5680 1316 5720 1364
rect 5680 1284 5684 1316
rect 5716 1284 5720 1316
rect 5680 1236 5720 1284
rect 5680 1204 5684 1236
rect 5716 1204 5720 1236
rect 5680 1156 5720 1204
rect 5680 1124 5684 1156
rect 5716 1124 5720 1156
rect 5680 1076 5720 1124
rect 5680 1044 5684 1076
rect 5716 1044 5720 1076
rect 5680 996 5720 1044
rect 5680 964 5684 996
rect 5716 964 5720 996
rect 5680 916 5720 964
rect 5680 884 5684 916
rect 5716 884 5720 916
rect 5680 836 5720 884
rect 5680 804 5684 836
rect 5716 804 5720 836
rect 5680 756 5720 804
rect 5680 724 5684 756
rect 5716 724 5720 756
rect 5680 676 5720 724
rect 5680 644 5684 676
rect 5716 644 5720 676
rect 5680 596 5720 644
rect 5680 564 5684 596
rect 5716 564 5720 596
rect 5680 516 5720 564
rect 5680 484 5684 516
rect 5716 484 5720 516
rect 5680 436 5720 484
rect 5680 404 5684 436
rect 5716 404 5720 436
rect 5680 356 5720 404
rect 5680 324 5684 356
rect 5716 324 5720 356
rect 5680 276 5720 324
rect 5680 244 5684 276
rect 5716 244 5720 276
rect 5680 196 5720 244
rect 5680 164 5684 196
rect 5716 164 5720 196
rect 5680 116 5720 164
rect 5680 84 5684 116
rect 5716 84 5720 116
rect 5680 36 5720 84
rect 5680 4 5684 36
rect 5716 4 5720 36
rect 5520 -716 5524 -524
rect 5556 -716 5560 -524
rect 5520 -960 5560 -716
rect 5680 -524 5720 4
rect 5680 -716 5684 -524
rect 5716 -716 5720 -524
rect 5680 -960 5720 -716
rect 5760 15716 5800 15760
rect 5760 15684 5764 15716
rect 5796 15684 5800 15716
rect 5760 15636 5800 15684
rect 5760 15604 5764 15636
rect 5796 15604 5800 15636
rect 5760 15556 5800 15604
rect 5760 15524 5764 15556
rect 5796 15524 5800 15556
rect 5760 15476 5800 15524
rect 5760 15444 5764 15476
rect 5796 15444 5800 15476
rect 5760 15396 5800 15444
rect 5760 15364 5764 15396
rect 5796 15364 5800 15396
rect 5760 15316 5800 15364
rect 5760 15284 5764 15316
rect 5796 15284 5800 15316
rect 5760 15236 5800 15284
rect 5760 15204 5764 15236
rect 5796 15204 5800 15236
rect 5760 15156 5800 15204
rect 5760 15124 5764 15156
rect 5796 15124 5800 15156
rect 5760 15076 5800 15124
rect 5760 15044 5764 15076
rect 5796 15044 5800 15076
rect 5760 14996 5800 15044
rect 5760 14964 5764 14996
rect 5796 14964 5800 14996
rect 5760 14916 5800 14964
rect 5760 14884 5764 14916
rect 5796 14884 5800 14916
rect 5760 14836 5800 14884
rect 5760 14804 5764 14836
rect 5796 14804 5800 14836
rect 5760 14756 5800 14804
rect 5760 14724 5764 14756
rect 5796 14724 5800 14756
rect 5760 14676 5800 14724
rect 5760 14644 5764 14676
rect 5796 14644 5800 14676
rect 5760 14596 5800 14644
rect 5760 14564 5764 14596
rect 5796 14564 5800 14596
rect 5760 14516 5800 14564
rect 5760 14484 5764 14516
rect 5796 14484 5800 14516
rect 5760 14436 5800 14484
rect 5760 14404 5764 14436
rect 5796 14404 5800 14436
rect 5760 14356 5800 14404
rect 5760 14324 5764 14356
rect 5796 14324 5800 14356
rect 5760 14276 5800 14324
rect 5760 14244 5764 14276
rect 5796 14244 5800 14276
rect 5760 14196 5800 14244
rect 5760 14164 5764 14196
rect 5796 14164 5800 14196
rect 5760 14116 5800 14164
rect 5760 14084 5764 14116
rect 5796 14084 5800 14116
rect 5760 14036 5800 14084
rect 5760 14004 5764 14036
rect 5796 14004 5800 14036
rect 5760 13956 5800 14004
rect 5760 13924 5764 13956
rect 5796 13924 5800 13956
rect 5760 13876 5800 13924
rect 5760 13844 5764 13876
rect 5796 13844 5800 13876
rect 5760 13796 5800 13844
rect 5760 13764 5764 13796
rect 5796 13764 5800 13796
rect 5760 13716 5800 13764
rect 5760 13684 5764 13716
rect 5796 13684 5800 13716
rect 5760 13636 5800 13684
rect 5760 13604 5764 13636
rect 5796 13604 5800 13636
rect 5760 13556 5800 13604
rect 5760 13524 5764 13556
rect 5796 13524 5800 13556
rect 5760 13476 5800 13524
rect 5760 13444 5764 13476
rect 5796 13444 5800 13476
rect 5760 13396 5800 13444
rect 5760 13364 5764 13396
rect 5796 13364 5800 13396
rect 5760 13316 5800 13364
rect 5760 13284 5764 13316
rect 5796 13284 5800 13316
rect 5760 13236 5800 13284
rect 5760 13204 5764 13236
rect 5796 13204 5800 13236
rect 5760 13156 5800 13204
rect 5760 13124 5764 13156
rect 5796 13124 5800 13156
rect 5760 13076 5800 13124
rect 5760 13044 5764 13076
rect 5796 13044 5800 13076
rect 5760 12996 5800 13044
rect 5760 12964 5764 12996
rect 5796 12964 5800 12996
rect 5760 12916 5800 12964
rect 5760 12884 5764 12916
rect 5796 12884 5800 12916
rect 5760 12836 5800 12884
rect 5760 12804 5764 12836
rect 5796 12804 5800 12836
rect 5760 12756 5800 12804
rect 5760 12724 5764 12756
rect 5796 12724 5800 12756
rect 5760 12676 5800 12724
rect 5760 12644 5764 12676
rect 5796 12644 5800 12676
rect 5760 12596 5800 12644
rect 5760 12564 5764 12596
rect 5796 12564 5800 12596
rect 5760 12516 5800 12564
rect 5760 12484 5764 12516
rect 5796 12484 5800 12516
rect 5760 12436 5800 12484
rect 5760 12404 5764 12436
rect 5796 12404 5800 12436
rect 5760 12356 5800 12404
rect 5760 12324 5764 12356
rect 5796 12324 5800 12356
rect 5760 12276 5800 12324
rect 5760 12244 5764 12276
rect 5796 12244 5800 12276
rect 5760 12196 5800 12244
rect 5760 12164 5764 12196
rect 5796 12164 5800 12196
rect 5760 12116 5800 12164
rect 5760 12084 5764 12116
rect 5796 12084 5800 12116
rect 5760 12036 5800 12084
rect 5760 12004 5764 12036
rect 5796 12004 5800 12036
rect 5760 11956 5800 12004
rect 5760 11924 5764 11956
rect 5796 11924 5800 11956
rect 5760 11876 5800 11924
rect 5760 11844 5764 11876
rect 5796 11844 5800 11876
rect 5760 11796 5800 11844
rect 5760 11764 5764 11796
rect 5796 11764 5800 11796
rect 5760 11716 5800 11764
rect 5760 11684 5764 11716
rect 5796 11684 5800 11716
rect 5760 11636 5800 11684
rect 5760 11604 5764 11636
rect 5796 11604 5800 11636
rect 5760 11556 5800 11604
rect 5760 11524 5764 11556
rect 5796 11524 5800 11556
rect 5760 11476 5800 11524
rect 5760 11444 5764 11476
rect 5796 11444 5800 11476
rect 5760 11396 5800 11444
rect 5760 11364 5764 11396
rect 5796 11364 5800 11396
rect 5760 11316 5800 11364
rect 5760 11284 5764 11316
rect 5796 11284 5800 11316
rect 5760 11236 5800 11284
rect 5760 11204 5764 11236
rect 5796 11204 5800 11236
rect 5760 11156 5800 11204
rect 5760 11124 5764 11156
rect 5796 11124 5800 11156
rect 5760 11076 5800 11124
rect 5760 11044 5764 11076
rect 5796 11044 5800 11076
rect 5760 10996 5800 11044
rect 5760 10964 5764 10996
rect 5796 10964 5800 10996
rect 5760 10916 5800 10964
rect 5760 10884 5764 10916
rect 5796 10884 5800 10916
rect 5760 10836 5800 10884
rect 5760 10804 5764 10836
rect 5796 10804 5800 10836
rect 5760 10756 5800 10804
rect 5760 10724 5764 10756
rect 5796 10724 5800 10756
rect 5760 10676 5800 10724
rect 5760 10644 5764 10676
rect 5796 10644 5800 10676
rect 5760 10596 5800 10644
rect 5760 10564 5764 10596
rect 5796 10564 5800 10596
rect 5760 10516 5800 10564
rect 5760 10484 5764 10516
rect 5796 10484 5800 10516
rect 5760 10436 5800 10484
rect 5760 10404 5764 10436
rect 5796 10404 5800 10436
rect 5760 10356 5800 10404
rect 5760 10324 5764 10356
rect 5796 10324 5800 10356
rect 5760 10276 5800 10324
rect 5760 10244 5764 10276
rect 5796 10244 5800 10276
rect 5760 10196 5800 10244
rect 5760 10164 5764 10196
rect 5796 10164 5800 10196
rect 5760 10116 5800 10164
rect 5760 10084 5764 10116
rect 5796 10084 5800 10116
rect 5760 10036 5800 10084
rect 5760 10004 5764 10036
rect 5796 10004 5800 10036
rect 5760 9956 5800 10004
rect 5760 9924 5764 9956
rect 5796 9924 5800 9956
rect 5760 9876 5800 9924
rect 5760 9844 5764 9876
rect 5796 9844 5800 9876
rect 5760 9796 5800 9844
rect 5760 9764 5764 9796
rect 5796 9764 5800 9796
rect 5760 9716 5800 9764
rect 5760 9684 5764 9716
rect 5796 9684 5800 9716
rect 5760 9636 5800 9684
rect 5760 9604 5764 9636
rect 5796 9604 5800 9636
rect 5760 9556 5800 9604
rect 5760 9524 5764 9556
rect 5796 9524 5800 9556
rect 5760 9476 5800 9524
rect 5760 9444 5764 9476
rect 5796 9444 5800 9476
rect 5760 9396 5800 9444
rect 5760 9364 5764 9396
rect 5796 9364 5800 9396
rect 5760 9316 5800 9364
rect 5760 9284 5764 9316
rect 5796 9284 5800 9316
rect 5760 9236 5800 9284
rect 5760 9204 5764 9236
rect 5796 9204 5800 9236
rect 5760 9156 5800 9204
rect 5760 9124 5764 9156
rect 5796 9124 5800 9156
rect 5760 9076 5800 9124
rect 5760 9044 5764 9076
rect 5796 9044 5800 9076
rect 5760 8996 5800 9044
rect 5760 8964 5764 8996
rect 5796 8964 5800 8996
rect 5760 8916 5800 8964
rect 5760 8884 5764 8916
rect 5796 8884 5800 8916
rect 5760 8836 5800 8884
rect 5760 8804 5764 8836
rect 5796 8804 5800 8836
rect 5760 8756 5800 8804
rect 5760 8724 5764 8756
rect 5796 8724 5800 8756
rect 5760 8676 5800 8724
rect 5760 8644 5764 8676
rect 5796 8644 5800 8676
rect 5760 8596 5800 8644
rect 5760 8564 5764 8596
rect 5796 8564 5800 8596
rect 5760 8516 5800 8564
rect 5760 8484 5764 8516
rect 5796 8484 5800 8516
rect 5760 8436 5800 8484
rect 5760 8404 5764 8436
rect 5796 8404 5800 8436
rect 5760 8356 5800 8404
rect 5760 8324 5764 8356
rect 5796 8324 5800 8356
rect 5760 8276 5800 8324
rect 5760 8244 5764 8276
rect 5796 8244 5800 8276
rect 5760 8196 5800 8244
rect 5760 8164 5764 8196
rect 5796 8164 5800 8196
rect 5760 8116 5800 8164
rect 5760 8084 5764 8116
rect 5796 8084 5800 8116
rect 5760 8036 5800 8084
rect 5760 8004 5764 8036
rect 5796 8004 5800 8036
rect 5760 7956 5800 8004
rect 5760 7924 5764 7956
rect 5796 7924 5800 7956
rect 5760 7876 5800 7924
rect 5760 7844 5764 7876
rect 5796 7844 5800 7876
rect 5760 7796 5800 7844
rect 5760 7764 5764 7796
rect 5796 7764 5800 7796
rect 5760 7716 5800 7764
rect 5760 7684 5764 7716
rect 5796 7684 5800 7716
rect 5760 7636 5800 7684
rect 5760 7604 5764 7636
rect 5796 7604 5800 7636
rect 5760 7556 5800 7604
rect 5760 7524 5764 7556
rect 5796 7524 5800 7556
rect 5760 7476 5800 7524
rect 5760 7444 5764 7476
rect 5796 7444 5800 7476
rect 5760 7396 5800 7444
rect 5760 7364 5764 7396
rect 5796 7364 5800 7396
rect 5760 7316 5800 7364
rect 5760 7284 5764 7316
rect 5796 7284 5800 7316
rect 5760 7236 5800 7284
rect 5760 7204 5764 7236
rect 5796 7204 5800 7236
rect 5760 7156 5800 7204
rect 5760 7124 5764 7156
rect 5796 7124 5800 7156
rect 5760 7076 5800 7124
rect 5760 7044 5764 7076
rect 5796 7044 5800 7076
rect 5760 6996 5800 7044
rect 5760 6964 5764 6996
rect 5796 6964 5800 6996
rect 5760 6916 5800 6964
rect 5760 6884 5764 6916
rect 5796 6884 5800 6916
rect 5760 6836 5800 6884
rect 5760 6804 5764 6836
rect 5796 6804 5800 6836
rect 5760 6756 5800 6804
rect 5760 6724 5764 6756
rect 5796 6724 5800 6756
rect 5760 6676 5800 6724
rect 5760 6644 5764 6676
rect 5796 6644 5800 6676
rect 5760 6596 5800 6644
rect 5760 6564 5764 6596
rect 5796 6564 5800 6596
rect 5760 6516 5800 6564
rect 5760 6484 5764 6516
rect 5796 6484 5800 6516
rect 5760 6436 5800 6484
rect 5760 6404 5764 6436
rect 5796 6404 5800 6436
rect 5760 6356 5800 6404
rect 5760 6324 5764 6356
rect 5796 6324 5800 6356
rect 5760 6276 5800 6324
rect 5760 6244 5764 6276
rect 5796 6244 5800 6276
rect 5760 6196 5800 6244
rect 5760 6164 5764 6196
rect 5796 6164 5800 6196
rect 5760 6116 5800 6164
rect 5760 6084 5764 6116
rect 5796 6084 5800 6116
rect 5760 6036 5800 6084
rect 5760 6004 5764 6036
rect 5796 6004 5800 6036
rect 5760 5956 5800 6004
rect 5760 5924 5764 5956
rect 5796 5924 5800 5956
rect 5760 5876 5800 5924
rect 5760 5844 5764 5876
rect 5796 5844 5800 5876
rect 5760 5796 5800 5844
rect 5760 5764 5764 5796
rect 5796 5764 5800 5796
rect 5760 5716 5800 5764
rect 5760 5684 5764 5716
rect 5796 5684 5800 5716
rect 5760 5636 5800 5684
rect 5760 5604 5764 5636
rect 5796 5604 5800 5636
rect 5760 5556 5800 5604
rect 5760 5524 5764 5556
rect 5796 5524 5800 5556
rect 5760 5476 5800 5524
rect 5760 5444 5764 5476
rect 5796 5444 5800 5476
rect 5760 5396 5800 5444
rect 5760 5364 5764 5396
rect 5796 5364 5800 5396
rect 5760 5316 5800 5364
rect 5760 5284 5764 5316
rect 5796 5284 5800 5316
rect 5760 5236 5800 5284
rect 5760 5204 5764 5236
rect 5796 5204 5800 5236
rect 5760 5156 5800 5204
rect 5760 5124 5764 5156
rect 5796 5124 5800 5156
rect 5760 5076 5800 5124
rect 5760 5044 5764 5076
rect 5796 5044 5800 5076
rect 5760 4996 5800 5044
rect 5760 4964 5764 4996
rect 5796 4964 5800 4996
rect 5760 4916 5800 4964
rect 5760 4884 5764 4916
rect 5796 4884 5800 4916
rect 5760 4836 5800 4884
rect 5760 4804 5764 4836
rect 5796 4804 5800 4836
rect 5760 4756 5800 4804
rect 5760 4724 5764 4756
rect 5796 4724 5800 4756
rect 5760 4676 5800 4724
rect 5760 4644 5764 4676
rect 5796 4644 5800 4676
rect 5760 4596 5800 4644
rect 5760 4564 5764 4596
rect 5796 4564 5800 4596
rect 5760 4516 5800 4564
rect 5760 4484 5764 4516
rect 5796 4484 5800 4516
rect 5760 4436 5800 4484
rect 5760 4404 5764 4436
rect 5796 4404 5800 4436
rect 5760 4356 5800 4404
rect 5760 4324 5764 4356
rect 5796 4324 5800 4356
rect 5760 4276 5800 4324
rect 5760 4244 5764 4276
rect 5796 4244 5800 4276
rect 5760 4196 5800 4244
rect 5760 4164 5764 4196
rect 5796 4164 5800 4196
rect 5760 4116 5800 4164
rect 5760 4084 5764 4116
rect 5796 4084 5800 4116
rect 5760 4036 5800 4084
rect 5760 4004 5764 4036
rect 5796 4004 5800 4036
rect 5760 3956 5800 4004
rect 5760 3924 5764 3956
rect 5796 3924 5800 3956
rect 5760 3876 5800 3924
rect 5760 3844 5764 3876
rect 5796 3844 5800 3876
rect 5760 3796 5800 3844
rect 5760 3764 5764 3796
rect 5796 3764 5800 3796
rect 5760 3716 5800 3764
rect 5760 3684 5764 3716
rect 5796 3684 5800 3716
rect 5760 3636 5800 3684
rect 5760 3604 5764 3636
rect 5796 3604 5800 3636
rect 5760 3556 5800 3604
rect 5760 3524 5764 3556
rect 5796 3524 5800 3556
rect 5760 3476 5800 3524
rect 5760 3444 5764 3476
rect 5796 3444 5800 3476
rect 5760 3396 5800 3444
rect 5760 3364 5764 3396
rect 5796 3364 5800 3396
rect 5760 3316 5800 3364
rect 5760 3284 5764 3316
rect 5796 3284 5800 3316
rect 5760 3236 5800 3284
rect 5760 3204 5764 3236
rect 5796 3204 5800 3236
rect 5760 3156 5800 3204
rect 5760 3124 5764 3156
rect 5796 3124 5800 3156
rect 5760 3076 5800 3124
rect 5760 3044 5764 3076
rect 5796 3044 5800 3076
rect 5760 2996 5800 3044
rect 5760 2964 5764 2996
rect 5796 2964 5800 2996
rect 5760 2916 5800 2964
rect 5760 2884 5764 2916
rect 5796 2884 5800 2916
rect 5760 2836 5800 2884
rect 5760 2804 5764 2836
rect 5796 2804 5800 2836
rect 5760 2756 5800 2804
rect 5760 2724 5764 2756
rect 5796 2724 5800 2756
rect 5760 2676 5800 2724
rect 5760 2644 5764 2676
rect 5796 2644 5800 2676
rect 5760 2596 5800 2644
rect 5760 2564 5764 2596
rect 5796 2564 5800 2596
rect 5760 2516 5800 2564
rect 5760 2484 5764 2516
rect 5796 2484 5800 2516
rect 5760 2436 5800 2484
rect 5760 2404 5764 2436
rect 5796 2404 5800 2436
rect 5760 2356 5800 2404
rect 5760 2324 5764 2356
rect 5796 2324 5800 2356
rect 5760 2276 5800 2324
rect 5760 2244 5764 2276
rect 5796 2244 5800 2276
rect 5760 2196 5800 2244
rect 5760 2164 5764 2196
rect 5796 2164 5800 2196
rect 5760 2116 5800 2164
rect 5760 2084 5764 2116
rect 5796 2084 5800 2116
rect 5760 2036 5800 2084
rect 5760 2004 5764 2036
rect 5796 2004 5800 2036
rect 5760 1956 5800 2004
rect 5760 1924 5764 1956
rect 5796 1924 5800 1956
rect 5760 1876 5800 1924
rect 5760 1844 5764 1876
rect 5796 1844 5800 1876
rect 5760 1796 5800 1844
rect 5760 1764 5764 1796
rect 5796 1764 5800 1796
rect 5760 1716 5800 1764
rect 5760 1684 5764 1716
rect 5796 1684 5800 1716
rect 5760 1636 5800 1684
rect 5760 1604 5764 1636
rect 5796 1604 5800 1636
rect 5760 1556 5800 1604
rect 5760 1524 5764 1556
rect 5796 1524 5800 1556
rect 5760 1476 5800 1524
rect 5760 1444 5764 1476
rect 5796 1444 5800 1476
rect 5760 1396 5800 1444
rect 5760 1364 5764 1396
rect 5796 1364 5800 1396
rect 5760 1316 5800 1364
rect 5760 1284 5764 1316
rect 5796 1284 5800 1316
rect 5760 1236 5800 1284
rect 5760 1204 5764 1236
rect 5796 1204 5800 1236
rect 5760 1156 5800 1204
rect 5760 1124 5764 1156
rect 5796 1124 5800 1156
rect 5760 1076 5800 1124
rect 5760 1044 5764 1076
rect 5796 1044 5800 1076
rect 5760 996 5800 1044
rect 5760 964 5764 996
rect 5796 964 5800 996
rect 5760 916 5800 964
rect 5760 884 5764 916
rect 5796 884 5800 916
rect 5760 836 5800 884
rect 5760 804 5764 836
rect 5796 804 5800 836
rect 5760 756 5800 804
rect 5760 724 5764 756
rect 5796 724 5800 756
rect 5760 676 5800 724
rect 5760 644 5764 676
rect 5796 644 5800 676
rect 5760 596 5800 644
rect 5760 564 5764 596
rect 5796 564 5800 596
rect 5760 516 5800 564
rect 5760 484 5764 516
rect 5796 484 5800 516
rect 5760 436 5800 484
rect 5760 404 5764 436
rect 5796 404 5800 436
rect 5760 356 5800 404
rect 5760 324 5764 356
rect 5796 324 5800 356
rect 5760 276 5800 324
rect 5760 244 5764 276
rect 5796 244 5800 276
rect 5760 196 5800 244
rect 5760 164 5764 196
rect 5796 164 5800 196
rect 5760 116 5800 164
rect 5760 84 5764 116
rect 5796 84 5800 116
rect 5760 36 5800 84
rect 5760 4 5764 36
rect 5796 4 5800 36
rect 5760 -44 5800 4
rect 5840 4835 5880 15760
rect 5840 4805 5845 4835
rect 5875 4805 5880 4835
rect 5840 3315 5880 4805
rect 5840 3285 5845 3315
rect 5875 3285 5880 3315
rect 5840 0 5880 3285
rect 5920 15716 5960 15760
rect 5920 15684 5924 15716
rect 5956 15684 5960 15716
rect 5920 15636 5960 15684
rect 5920 15604 5924 15636
rect 5956 15604 5960 15636
rect 5920 15556 5960 15604
rect 5920 15524 5924 15556
rect 5956 15524 5960 15556
rect 5920 15476 5960 15524
rect 5920 15444 5924 15476
rect 5956 15444 5960 15476
rect 5920 15396 5960 15444
rect 5920 15364 5924 15396
rect 5956 15364 5960 15396
rect 5920 15316 5960 15364
rect 5920 15284 5924 15316
rect 5956 15284 5960 15316
rect 5920 15236 5960 15284
rect 5920 15204 5924 15236
rect 5956 15204 5960 15236
rect 5920 15156 5960 15204
rect 5920 15124 5924 15156
rect 5956 15124 5960 15156
rect 5920 15076 5960 15124
rect 5920 15044 5924 15076
rect 5956 15044 5960 15076
rect 5920 14996 5960 15044
rect 5920 14964 5924 14996
rect 5956 14964 5960 14996
rect 5920 14916 5960 14964
rect 5920 14884 5924 14916
rect 5956 14884 5960 14916
rect 5920 14836 5960 14884
rect 5920 14804 5924 14836
rect 5956 14804 5960 14836
rect 5920 14756 5960 14804
rect 5920 14724 5924 14756
rect 5956 14724 5960 14756
rect 5920 14676 5960 14724
rect 5920 14644 5924 14676
rect 5956 14644 5960 14676
rect 5920 14596 5960 14644
rect 5920 14564 5924 14596
rect 5956 14564 5960 14596
rect 5920 14516 5960 14564
rect 5920 14484 5924 14516
rect 5956 14484 5960 14516
rect 5920 14436 5960 14484
rect 5920 14404 5924 14436
rect 5956 14404 5960 14436
rect 5920 14356 5960 14404
rect 5920 14324 5924 14356
rect 5956 14324 5960 14356
rect 5920 14276 5960 14324
rect 5920 14244 5924 14276
rect 5956 14244 5960 14276
rect 5920 14196 5960 14244
rect 5920 14164 5924 14196
rect 5956 14164 5960 14196
rect 5920 14116 5960 14164
rect 5920 14084 5924 14116
rect 5956 14084 5960 14116
rect 5920 14036 5960 14084
rect 5920 14004 5924 14036
rect 5956 14004 5960 14036
rect 5920 13956 5960 14004
rect 5920 13924 5924 13956
rect 5956 13924 5960 13956
rect 5920 13876 5960 13924
rect 5920 13844 5924 13876
rect 5956 13844 5960 13876
rect 5920 13796 5960 13844
rect 5920 13764 5924 13796
rect 5956 13764 5960 13796
rect 5920 13716 5960 13764
rect 5920 13684 5924 13716
rect 5956 13684 5960 13716
rect 5920 13636 5960 13684
rect 5920 13604 5924 13636
rect 5956 13604 5960 13636
rect 5920 13556 5960 13604
rect 5920 13524 5924 13556
rect 5956 13524 5960 13556
rect 5920 13476 5960 13524
rect 5920 13444 5924 13476
rect 5956 13444 5960 13476
rect 5920 13396 5960 13444
rect 5920 13364 5924 13396
rect 5956 13364 5960 13396
rect 5920 13316 5960 13364
rect 5920 13284 5924 13316
rect 5956 13284 5960 13316
rect 5920 13236 5960 13284
rect 5920 13204 5924 13236
rect 5956 13204 5960 13236
rect 5920 13156 5960 13204
rect 5920 13124 5924 13156
rect 5956 13124 5960 13156
rect 5920 13076 5960 13124
rect 5920 13044 5924 13076
rect 5956 13044 5960 13076
rect 5920 12996 5960 13044
rect 5920 12964 5924 12996
rect 5956 12964 5960 12996
rect 5920 12916 5960 12964
rect 5920 12884 5924 12916
rect 5956 12884 5960 12916
rect 5920 12836 5960 12884
rect 5920 12804 5924 12836
rect 5956 12804 5960 12836
rect 5920 12756 5960 12804
rect 5920 12724 5924 12756
rect 5956 12724 5960 12756
rect 5920 12676 5960 12724
rect 5920 12644 5924 12676
rect 5956 12644 5960 12676
rect 5920 12596 5960 12644
rect 5920 12564 5924 12596
rect 5956 12564 5960 12596
rect 5920 12516 5960 12564
rect 5920 12484 5924 12516
rect 5956 12484 5960 12516
rect 5920 12436 5960 12484
rect 5920 12404 5924 12436
rect 5956 12404 5960 12436
rect 5920 12356 5960 12404
rect 5920 12324 5924 12356
rect 5956 12324 5960 12356
rect 5920 12276 5960 12324
rect 5920 12244 5924 12276
rect 5956 12244 5960 12276
rect 5920 12196 5960 12244
rect 5920 12164 5924 12196
rect 5956 12164 5960 12196
rect 5920 12116 5960 12164
rect 5920 12084 5924 12116
rect 5956 12084 5960 12116
rect 5920 12036 5960 12084
rect 5920 12004 5924 12036
rect 5956 12004 5960 12036
rect 5920 11956 5960 12004
rect 5920 11924 5924 11956
rect 5956 11924 5960 11956
rect 5920 11876 5960 11924
rect 5920 11844 5924 11876
rect 5956 11844 5960 11876
rect 5920 11796 5960 11844
rect 5920 11764 5924 11796
rect 5956 11764 5960 11796
rect 5920 11716 5960 11764
rect 5920 11684 5924 11716
rect 5956 11684 5960 11716
rect 5920 11636 5960 11684
rect 5920 11604 5924 11636
rect 5956 11604 5960 11636
rect 5920 11556 5960 11604
rect 5920 11524 5924 11556
rect 5956 11524 5960 11556
rect 5920 11476 5960 11524
rect 5920 11444 5924 11476
rect 5956 11444 5960 11476
rect 5920 11396 5960 11444
rect 5920 11364 5924 11396
rect 5956 11364 5960 11396
rect 5920 11316 5960 11364
rect 5920 11284 5924 11316
rect 5956 11284 5960 11316
rect 5920 11236 5960 11284
rect 5920 11204 5924 11236
rect 5956 11204 5960 11236
rect 5920 11156 5960 11204
rect 5920 11124 5924 11156
rect 5956 11124 5960 11156
rect 5920 11076 5960 11124
rect 5920 11044 5924 11076
rect 5956 11044 5960 11076
rect 5920 10996 5960 11044
rect 5920 10964 5924 10996
rect 5956 10964 5960 10996
rect 5920 10916 5960 10964
rect 5920 10884 5924 10916
rect 5956 10884 5960 10916
rect 5920 10836 5960 10884
rect 5920 10804 5924 10836
rect 5956 10804 5960 10836
rect 5920 10756 5960 10804
rect 5920 10724 5924 10756
rect 5956 10724 5960 10756
rect 5920 10676 5960 10724
rect 5920 10644 5924 10676
rect 5956 10644 5960 10676
rect 5920 10596 5960 10644
rect 5920 10564 5924 10596
rect 5956 10564 5960 10596
rect 5920 10516 5960 10564
rect 5920 10484 5924 10516
rect 5956 10484 5960 10516
rect 5920 10436 5960 10484
rect 5920 10404 5924 10436
rect 5956 10404 5960 10436
rect 5920 10356 5960 10404
rect 5920 10324 5924 10356
rect 5956 10324 5960 10356
rect 5920 10276 5960 10324
rect 5920 10244 5924 10276
rect 5956 10244 5960 10276
rect 5920 10196 5960 10244
rect 5920 10164 5924 10196
rect 5956 10164 5960 10196
rect 5920 10116 5960 10164
rect 5920 10084 5924 10116
rect 5956 10084 5960 10116
rect 5920 10036 5960 10084
rect 5920 10004 5924 10036
rect 5956 10004 5960 10036
rect 5920 9956 5960 10004
rect 5920 9924 5924 9956
rect 5956 9924 5960 9956
rect 5920 9876 5960 9924
rect 5920 9844 5924 9876
rect 5956 9844 5960 9876
rect 5920 9796 5960 9844
rect 5920 9764 5924 9796
rect 5956 9764 5960 9796
rect 5920 9716 5960 9764
rect 5920 9684 5924 9716
rect 5956 9684 5960 9716
rect 5920 9636 5960 9684
rect 5920 9604 5924 9636
rect 5956 9604 5960 9636
rect 5920 9556 5960 9604
rect 5920 9524 5924 9556
rect 5956 9524 5960 9556
rect 5920 9476 5960 9524
rect 5920 9444 5924 9476
rect 5956 9444 5960 9476
rect 5920 9396 5960 9444
rect 5920 9364 5924 9396
rect 5956 9364 5960 9396
rect 5920 9316 5960 9364
rect 5920 9284 5924 9316
rect 5956 9284 5960 9316
rect 5920 9236 5960 9284
rect 5920 9204 5924 9236
rect 5956 9204 5960 9236
rect 5920 9156 5960 9204
rect 5920 9124 5924 9156
rect 5956 9124 5960 9156
rect 5920 9076 5960 9124
rect 5920 9044 5924 9076
rect 5956 9044 5960 9076
rect 5920 8996 5960 9044
rect 5920 8964 5924 8996
rect 5956 8964 5960 8996
rect 5920 8916 5960 8964
rect 5920 8884 5924 8916
rect 5956 8884 5960 8916
rect 5920 8836 5960 8884
rect 5920 8804 5924 8836
rect 5956 8804 5960 8836
rect 5920 8756 5960 8804
rect 5920 8724 5924 8756
rect 5956 8724 5960 8756
rect 5920 8676 5960 8724
rect 5920 8644 5924 8676
rect 5956 8644 5960 8676
rect 5920 8596 5960 8644
rect 5920 8564 5924 8596
rect 5956 8564 5960 8596
rect 5920 8516 5960 8564
rect 5920 8484 5924 8516
rect 5956 8484 5960 8516
rect 5920 8436 5960 8484
rect 5920 8404 5924 8436
rect 5956 8404 5960 8436
rect 5920 8356 5960 8404
rect 5920 8324 5924 8356
rect 5956 8324 5960 8356
rect 5920 8276 5960 8324
rect 5920 8244 5924 8276
rect 5956 8244 5960 8276
rect 5920 8196 5960 8244
rect 5920 8164 5924 8196
rect 5956 8164 5960 8196
rect 5920 8116 5960 8164
rect 5920 8084 5924 8116
rect 5956 8084 5960 8116
rect 5920 8036 5960 8084
rect 5920 8004 5924 8036
rect 5956 8004 5960 8036
rect 5920 7956 5960 8004
rect 5920 7924 5924 7956
rect 5956 7924 5960 7956
rect 5920 7876 5960 7924
rect 5920 7844 5924 7876
rect 5956 7844 5960 7876
rect 5920 7796 5960 7844
rect 5920 7764 5924 7796
rect 5956 7764 5960 7796
rect 5920 7716 5960 7764
rect 5920 7684 5924 7716
rect 5956 7684 5960 7716
rect 5920 7636 5960 7684
rect 5920 7604 5924 7636
rect 5956 7604 5960 7636
rect 5920 7556 5960 7604
rect 5920 7524 5924 7556
rect 5956 7524 5960 7556
rect 5920 7476 5960 7524
rect 5920 7444 5924 7476
rect 5956 7444 5960 7476
rect 5920 7396 5960 7444
rect 5920 7364 5924 7396
rect 5956 7364 5960 7396
rect 5920 7316 5960 7364
rect 5920 7284 5924 7316
rect 5956 7284 5960 7316
rect 5920 7236 5960 7284
rect 5920 7204 5924 7236
rect 5956 7204 5960 7236
rect 5920 7156 5960 7204
rect 5920 7124 5924 7156
rect 5956 7124 5960 7156
rect 5920 7076 5960 7124
rect 5920 7044 5924 7076
rect 5956 7044 5960 7076
rect 5920 6996 5960 7044
rect 5920 6964 5924 6996
rect 5956 6964 5960 6996
rect 5920 6916 5960 6964
rect 5920 6884 5924 6916
rect 5956 6884 5960 6916
rect 5920 6836 5960 6884
rect 5920 6804 5924 6836
rect 5956 6804 5960 6836
rect 5920 6756 5960 6804
rect 5920 6724 5924 6756
rect 5956 6724 5960 6756
rect 5920 6676 5960 6724
rect 5920 6644 5924 6676
rect 5956 6644 5960 6676
rect 5920 6596 5960 6644
rect 5920 6564 5924 6596
rect 5956 6564 5960 6596
rect 5920 6516 5960 6564
rect 5920 6484 5924 6516
rect 5956 6484 5960 6516
rect 5920 6436 5960 6484
rect 5920 6404 5924 6436
rect 5956 6404 5960 6436
rect 5920 6356 5960 6404
rect 5920 6324 5924 6356
rect 5956 6324 5960 6356
rect 5920 6276 5960 6324
rect 5920 6244 5924 6276
rect 5956 6244 5960 6276
rect 5920 6196 5960 6244
rect 5920 6164 5924 6196
rect 5956 6164 5960 6196
rect 5920 6116 5960 6164
rect 5920 6084 5924 6116
rect 5956 6084 5960 6116
rect 5920 6036 5960 6084
rect 5920 6004 5924 6036
rect 5956 6004 5960 6036
rect 5920 5956 5960 6004
rect 5920 5924 5924 5956
rect 5956 5924 5960 5956
rect 5920 5876 5960 5924
rect 5920 5844 5924 5876
rect 5956 5844 5960 5876
rect 5920 5796 5960 5844
rect 5920 5764 5924 5796
rect 5956 5764 5960 5796
rect 5920 5716 5960 5764
rect 5920 5684 5924 5716
rect 5956 5684 5960 5716
rect 5920 5636 5960 5684
rect 5920 5604 5924 5636
rect 5956 5604 5960 5636
rect 5920 5556 5960 5604
rect 5920 5524 5924 5556
rect 5956 5524 5960 5556
rect 5920 5476 5960 5524
rect 5920 5444 5924 5476
rect 5956 5444 5960 5476
rect 5920 5396 5960 5444
rect 5920 5364 5924 5396
rect 5956 5364 5960 5396
rect 5920 5316 5960 5364
rect 5920 5284 5924 5316
rect 5956 5284 5960 5316
rect 5920 5236 5960 5284
rect 5920 5204 5924 5236
rect 5956 5204 5960 5236
rect 5920 5156 5960 5204
rect 5920 5124 5924 5156
rect 5956 5124 5960 5156
rect 5920 5076 5960 5124
rect 5920 5044 5924 5076
rect 5956 5044 5960 5076
rect 5920 4996 5960 5044
rect 5920 4964 5924 4996
rect 5956 4964 5960 4996
rect 5920 4916 5960 4964
rect 5920 4884 5924 4916
rect 5956 4884 5960 4916
rect 5920 4836 5960 4884
rect 5920 4804 5924 4836
rect 5956 4804 5960 4836
rect 5920 4756 5960 4804
rect 5920 4724 5924 4756
rect 5956 4724 5960 4756
rect 5920 4676 5960 4724
rect 5920 4644 5924 4676
rect 5956 4644 5960 4676
rect 5920 4596 5960 4644
rect 5920 4564 5924 4596
rect 5956 4564 5960 4596
rect 5920 4516 5960 4564
rect 5920 4484 5924 4516
rect 5956 4484 5960 4516
rect 5920 4436 5960 4484
rect 5920 4404 5924 4436
rect 5956 4404 5960 4436
rect 5920 4356 5960 4404
rect 5920 4324 5924 4356
rect 5956 4324 5960 4356
rect 5920 4276 5960 4324
rect 5920 4244 5924 4276
rect 5956 4244 5960 4276
rect 5920 4196 5960 4244
rect 5920 4164 5924 4196
rect 5956 4164 5960 4196
rect 5920 4116 5960 4164
rect 5920 4084 5924 4116
rect 5956 4084 5960 4116
rect 5920 4036 5960 4084
rect 5920 4004 5924 4036
rect 5956 4004 5960 4036
rect 5920 3956 5960 4004
rect 5920 3924 5924 3956
rect 5956 3924 5960 3956
rect 5920 3876 5960 3924
rect 5920 3844 5924 3876
rect 5956 3844 5960 3876
rect 5920 3796 5960 3844
rect 5920 3764 5924 3796
rect 5956 3764 5960 3796
rect 5920 3716 5960 3764
rect 5920 3684 5924 3716
rect 5956 3684 5960 3716
rect 5920 3636 5960 3684
rect 5920 3604 5924 3636
rect 5956 3604 5960 3636
rect 5920 3556 5960 3604
rect 5920 3524 5924 3556
rect 5956 3524 5960 3556
rect 5920 3476 5960 3524
rect 5920 3444 5924 3476
rect 5956 3444 5960 3476
rect 5920 3396 5960 3444
rect 5920 3364 5924 3396
rect 5956 3364 5960 3396
rect 5920 3316 5960 3364
rect 5920 3284 5924 3316
rect 5956 3284 5960 3316
rect 5920 3236 5960 3284
rect 5920 3204 5924 3236
rect 5956 3204 5960 3236
rect 5920 3156 5960 3204
rect 5920 3124 5924 3156
rect 5956 3124 5960 3156
rect 5920 3076 5960 3124
rect 5920 3044 5924 3076
rect 5956 3044 5960 3076
rect 5920 2996 5960 3044
rect 5920 2964 5924 2996
rect 5956 2964 5960 2996
rect 5920 2916 5960 2964
rect 5920 2884 5924 2916
rect 5956 2884 5960 2916
rect 5920 2836 5960 2884
rect 5920 2804 5924 2836
rect 5956 2804 5960 2836
rect 5920 2756 5960 2804
rect 5920 2724 5924 2756
rect 5956 2724 5960 2756
rect 5920 2676 5960 2724
rect 5920 2644 5924 2676
rect 5956 2644 5960 2676
rect 5920 2596 5960 2644
rect 5920 2564 5924 2596
rect 5956 2564 5960 2596
rect 5920 2516 5960 2564
rect 5920 2484 5924 2516
rect 5956 2484 5960 2516
rect 5920 2436 5960 2484
rect 5920 2404 5924 2436
rect 5956 2404 5960 2436
rect 5920 2356 5960 2404
rect 5920 2324 5924 2356
rect 5956 2324 5960 2356
rect 5920 2276 5960 2324
rect 5920 2244 5924 2276
rect 5956 2244 5960 2276
rect 5920 2196 5960 2244
rect 5920 2164 5924 2196
rect 5956 2164 5960 2196
rect 5920 2116 5960 2164
rect 5920 2084 5924 2116
rect 5956 2084 5960 2116
rect 5920 2036 5960 2084
rect 5920 2004 5924 2036
rect 5956 2004 5960 2036
rect 5920 1956 5960 2004
rect 5920 1924 5924 1956
rect 5956 1924 5960 1956
rect 5920 1876 5960 1924
rect 5920 1844 5924 1876
rect 5956 1844 5960 1876
rect 5920 1796 5960 1844
rect 5920 1764 5924 1796
rect 5956 1764 5960 1796
rect 5920 1716 5960 1764
rect 5920 1684 5924 1716
rect 5956 1684 5960 1716
rect 5920 1636 5960 1684
rect 5920 1604 5924 1636
rect 5956 1604 5960 1636
rect 5920 1556 5960 1604
rect 5920 1524 5924 1556
rect 5956 1524 5960 1556
rect 5920 1476 5960 1524
rect 5920 1444 5924 1476
rect 5956 1444 5960 1476
rect 5920 1396 5960 1444
rect 5920 1364 5924 1396
rect 5956 1364 5960 1396
rect 5920 1316 5960 1364
rect 5920 1284 5924 1316
rect 5956 1284 5960 1316
rect 5920 1236 5960 1284
rect 5920 1204 5924 1236
rect 5956 1204 5960 1236
rect 5920 1156 5960 1204
rect 5920 1124 5924 1156
rect 5956 1124 5960 1156
rect 5920 1076 5960 1124
rect 5920 1044 5924 1076
rect 5956 1044 5960 1076
rect 5920 996 5960 1044
rect 5920 964 5924 996
rect 5956 964 5960 996
rect 5920 916 5960 964
rect 5920 884 5924 916
rect 5956 884 5960 916
rect 5920 836 5960 884
rect 5920 804 5924 836
rect 5956 804 5960 836
rect 5920 756 5960 804
rect 5920 724 5924 756
rect 5956 724 5960 756
rect 5920 676 5960 724
rect 5920 644 5924 676
rect 5956 644 5960 676
rect 5920 596 5960 644
rect 5920 564 5924 596
rect 5956 564 5960 596
rect 5920 516 5960 564
rect 5920 484 5924 516
rect 5956 484 5960 516
rect 5920 436 5960 484
rect 5920 404 5924 436
rect 5956 404 5960 436
rect 5920 356 5960 404
rect 5920 324 5924 356
rect 5956 324 5960 356
rect 5920 276 5960 324
rect 5920 244 5924 276
rect 5956 244 5960 276
rect 5920 196 5960 244
rect 5920 164 5924 196
rect 5956 164 5960 196
rect 5920 116 5960 164
rect 5920 84 5924 116
rect 5956 84 5960 116
rect 5920 36 5960 84
rect 5920 4 5924 36
rect 5956 4 5960 36
rect 5760 -236 5764 -44
rect 5796 -236 5800 -44
rect 5760 -960 5800 -236
rect 5920 -44 5960 4
rect 5920 -236 5924 -44
rect 5956 -236 5960 -44
rect 5920 -960 5960 -236
rect 6000 15716 6040 15760
rect 6000 15684 6004 15716
rect 6036 15684 6040 15716
rect 6000 15636 6040 15684
rect 6000 15604 6004 15636
rect 6036 15604 6040 15636
rect 6000 15556 6040 15604
rect 6000 15524 6004 15556
rect 6036 15524 6040 15556
rect 6000 15476 6040 15524
rect 6000 15444 6004 15476
rect 6036 15444 6040 15476
rect 6000 15396 6040 15444
rect 6000 15364 6004 15396
rect 6036 15364 6040 15396
rect 6000 15316 6040 15364
rect 6000 15284 6004 15316
rect 6036 15284 6040 15316
rect 6000 15236 6040 15284
rect 6000 15204 6004 15236
rect 6036 15204 6040 15236
rect 6000 15156 6040 15204
rect 6000 15124 6004 15156
rect 6036 15124 6040 15156
rect 6000 15076 6040 15124
rect 6000 15044 6004 15076
rect 6036 15044 6040 15076
rect 6000 14996 6040 15044
rect 6000 14964 6004 14996
rect 6036 14964 6040 14996
rect 6000 14916 6040 14964
rect 6000 14884 6004 14916
rect 6036 14884 6040 14916
rect 6000 14836 6040 14884
rect 6000 14804 6004 14836
rect 6036 14804 6040 14836
rect 6000 14756 6040 14804
rect 6000 14724 6004 14756
rect 6036 14724 6040 14756
rect 6000 14676 6040 14724
rect 6000 14644 6004 14676
rect 6036 14644 6040 14676
rect 6000 14596 6040 14644
rect 6000 14564 6004 14596
rect 6036 14564 6040 14596
rect 6000 14516 6040 14564
rect 6000 14484 6004 14516
rect 6036 14484 6040 14516
rect 6000 14436 6040 14484
rect 6000 14404 6004 14436
rect 6036 14404 6040 14436
rect 6000 14356 6040 14404
rect 6000 14324 6004 14356
rect 6036 14324 6040 14356
rect 6000 14276 6040 14324
rect 6000 14244 6004 14276
rect 6036 14244 6040 14276
rect 6000 14196 6040 14244
rect 6000 14164 6004 14196
rect 6036 14164 6040 14196
rect 6000 14116 6040 14164
rect 6000 14084 6004 14116
rect 6036 14084 6040 14116
rect 6000 14036 6040 14084
rect 6000 14004 6004 14036
rect 6036 14004 6040 14036
rect 6000 13956 6040 14004
rect 6000 13924 6004 13956
rect 6036 13924 6040 13956
rect 6000 13876 6040 13924
rect 6000 13844 6004 13876
rect 6036 13844 6040 13876
rect 6000 13796 6040 13844
rect 6000 13764 6004 13796
rect 6036 13764 6040 13796
rect 6000 13716 6040 13764
rect 6000 13684 6004 13716
rect 6036 13684 6040 13716
rect 6000 13636 6040 13684
rect 6000 13604 6004 13636
rect 6036 13604 6040 13636
rect 6000 13556 6040 13604
rect 6000 13524 6004 13556
rect 6036 13524 6040 13556
rect 6000 13476 6040 13524
rect 6000 13444 6004 13476
rect 6036 13444 6040 13476
rect 6000 13396 6040 13444
rect 6000 13364 6004 13396
rect 6036 13364 6040 13396
rect 6000 13316 6040 13364
rect 6000 13284 6004 13316
rect 6036 13284 6040 13316
rect 6000 13236 6040 13284
rect 6000 13204 6004 13236
rect 6036 13204 6040 13236
rect 6000 13156 6040 13204
rect 6000 13124 6004 13156
rect 6036 13124 6040 13156
rect 6000 13076 6040 13124
rect 6000 13044 6004 13076
rect 6036 13044 6040 13076
rect 6000 12996 6040 13044
rect 6000 12964 6004 12996
rect 6036 12964 6040 12996
rect 6000 12916 6040 12964
rect 6000 12884 6004 12916
rect 6036 12884 6040 12916
rect 6000 12836 6040 12884
rect 6000 12804 6004 12836
rect 6036 12804 6040 12836
rect 6000 12756 6040 12804
rect 6000 12724 6004 12756
rect 6036 12724 6040 12756
rect 6000 12676 6040 12724
rect 6000 12644 6004 12676
rect 6036 12644 6040 12676
rect 6000 12596 6040 12644
rect 6000 12564 6004 12596
rect 6036 12564 6040 12596
rect 6000 12516 6040 12564
rect 6000 12484 6004 12516
rect 6036 12484 6040 12516
rect 6000 12436 6040 12484
rect 6000 12404 6004 12436
rect 6036 12404 6040 12436
rect 6000 12356 6040 12404
rect 6000 12324 6004 12356
rect 6036 12324 6040 12356
rect 6000 12276 6040 12324
rect 6000 12244 6004 12276
rect 6036 12244 6040 12276
rect 6000 12196 6040 12244
rect 6000 12164 6004 12196
rect 6036 12164 6040 12196
rect 6000 12116 6040 12164
rect 6000 12084 6004 12116
rect 6036 12084 6040 12116
rect 6000 12036 6040 12084
rect 6000 12004 6004 12036
rect 6036 12004 6040 12036
rect 6000 11956 6040 12004
rect 6000 11924 6004 11956
rect 6036 11924 6040 11956
rect 6000 11876 6040 11924
rect 6000 11844 6004 11876
rect 6036 11844 6040 11876
rect 6000 11796 6040 11844
rect 6000 11764 6004 11796
rect 6036 11764 6040 11796
rect 6000 11716 6040 11764
rect 6000 11684 6004 11716
rect 6036 11684 6040 11716
rect 6000 11636 6040 11684
rect 6000 11604 6004 11636
rect 6036 11604 6040 11636
rect 6000 11556 6040 11604
rect 6000 11524 6004 11556
rect 6036 11524 6040 11556
rect 6000 11476 6040 11524
rect 6000 11444 6004 11476
rect 6036 11444 6040 11476
rect 6000 11396 6040 11444
rect 6000 11364 6004 11396
rect 6036 11364 6040 11396
rect 6000 11316 6040 11364
rect 6000 11284 6004 11316
rect 6036 11284 6040 11316
rect 6000 11236 6040 11284
rect 6000 11204 6004 11236
rect 6036 11204 6040 11236
rect 6000 11156 6040 11204
rect 6000 11124 6004 11156
rect 6036 11124 6040 11156
rect 6000 11076 6040 11124
rect 6000 11044 6004 11076
rect 6036 11044 6040 11076
rect 6000 10996 6040 11044
rect 6000 10964 6004 10996
rect 6036 10964 6040 10996
rect 6000 10916 6040 10964
rect 6000 10884 6004 10916
rect 6036 10884 6040 10916
rect 6000 10836 6040 10884
rect 6000 10804 6004 10836
rect 6036 10804 6040 10836
rect 6000 10756 6040 10804
rect 6000 10724 6004 10756
rect 6036 10724 6040 10756
rect 6000 10676 6040 10724
rect 6000 10644 6004 10676
rect 6036 10644 6040 10676
rect 6000 10596 6040 10644
rect 6000 10564 6004 10596
rect 6036 10564 6040 10596
rect 6000 10516 6040 10564
rect 6000 10484 6004 10516
rect 6036 10484 6040 10516
rect 6000 10436 6040 10484
rect 6000 10404 6004 10436
rect 6036 10404 6040 10436
rect 6000 10356 6040 10404
rect 6000 10324 6004 10356
rect 6036 10324 6040 10356
rect 6000 10276 6040 10324
rect 6000 10244 6004 10276
rect 6036 10244 6040 10276
rect 6000 10196 6040 10244
rect 6000 10164 6004 10196
rect 6036 10164 6040 10196
rect 6000 10116 6040 10164
rect 6000 10084 6004 10116
rect 6036 10084 6040 10116
rect 6000 10036 6040 10084
rect 6000 10004 6004 10036
rect 6036 10004 6040 10036
rect 6000 9956 6040 10004
rect 6000 9924 6004 9956
rect 6036 9924 6040 9956
rect 6000 9876 6040 9924
rect 6000 9844 6004 9876
rect 6036 9844 6040 9876
rect 6000 9796 6040 9844
rect 6000 9764 6004 9796
rect 6036 9764 6040 9796
rect 6000 9716 6040 9764
rect 6000 9684 6004 9716
rect 6036 9684 6040 9716
rect 6000 9636 6040 9684
rect 6000 9604 6004 9636
rect 6036 9604 6040 9636
rect 6000 9556 6040 9604
rect 6000 9524 6004 9556
rect 6036 9524 6040 9556
rect 6000 9476 6040 9524
rect 6000 9444 6004 9476
rect 6036 9444 6040 9476
rect 6000 9396 6040 9444
rect 6000 9364 6004 9396
rect 6036 9364 6040 9396
rect 6000 9316 6040 9364
rect 6000 9284 6004 9316
rect 6036 9284 6040 9316
rect 6000 9236 6040 9284
rect 6000 9204 6004 9236
rect 6036 9204 6040 9236
rect 6000 9156 6040 9204
rect 6000 9124 6004 9156
rect 6036 9124 6040 9156
rect 6000 9076 6040 9124
rect 6000 9044 6004 9076
rect 6036 9044 6040 9076
rect 6000 8996 6040 9044
rect 6000 8964 6004 8996
rect 6036 8964 6040 8996
rect 6000 8916 6040 8964
rect 6000 8884 6004 8916
rect 6036 8884 6040 8916
rect 6000 8836 6040 8884
rect 6000 8804 6004 8836
rect 6036 8804 6040 8836
rect 6000 8756 6040 8804
rect 6000 8724 6004 8756
rect 6036 8724 6040 8756
rect 6000 8676 6040 8724
rect 6000 8644 6004 8676
rect 6036 8644 6040 8676
rect 6000 8596 6040 8644
rect 6000 8564 6004 8596
rect 6036 8564 6040 8596
rect 6000 8516 6040 8564
rect 6000 8484 6004 8516
rect 6036 8484 6040 8516
rect 6000 8436 6040 8484
rect 6000 8404 6004 8436
rect 6036 8404 6040 8436
rect 6000 8356 6040 8404
rect 6000 8324 6004 8356
rect 6036 8324 6040 8356
rect 6000 8276 6040 8324
rect 6000 8244 6004 8276
rect 6036 8244 6040 8276
rect 6000 8196 6040 8244
rect 6000 8164 6004 8196
rect 6036 8164 6040 8196
rect 6000 8116 6040 8164
rect 6000 8084 6004 8116
rect 6036 8084 6040 8116
rect 6000 8036 6040 8084
rect 6000 8004 6004 8036
rect 6036 8004 6040 8036
rect 6000 7956 6040 8004
rect 6000 7924 6004 7956
rect 6036 7924 6040 7956
rect 6000 7876 6040 7924
rect 6000 7844 6004 7876
rect 6036 7844 6040 7876
rect 6000 7796 6040 7844
rect 6000 7764 6004 7796
rect 6036 7764 6040 7796
rect 6000 7716 6040 7764
rect 6000 7684 6004 7716
rect 6036 7684 6040 7716
rect 6000 7636 6040 7684
rect 6000 7604 6004 7636
rect 6036 7604 6040 7636
rect 6000 7556 6040 7604
rect 6000 7524 6004 7556
rect 6036 7524 6040 7556
rect 6000 7476 6040 7524
rect 6000 7444 6004 7476
rect 6036 7444 6040 7476
rect 6000 7396 6040 7444
rect 6000 7364 6004 7396
rect 6036 7364 6040 7396
rect 6000 7316 6040 7364
rect 6000 7284 6004 7316
rect 6036 7284 6040 7316
rect 6000 7236 6040 7284
rect 6000 7204 6004 7236
rect 6036 7204 6040 7236
rect 6000 7156 6040 7204
rect 6000 7124 6004 7156
rect 6036 7124 6040 7156
rect 6000 7076 6040 7124
rect 6000 7044 6004 7076
rect 6036 7044 6040 7076
rect 6000 6996 6040 7044
rect 6000 6964 6004 6996
rect 6036 6964 6040 6996
rect 6000 6916 6040 6964
rect 6000 6884 6004 6916
rect 6036 6884 6040 6916
rect 6000 6836 6040 6884
rect 6000 6804 6004 6836
rect 6036 6804 6040 6836
rect 6000 6756 6040 6804
rect 6000 6724 6004 6756
rect 6036 6724 6040 6756
rect 6000 6676 6040 6724
rect 6000 6644 6004 6676
rect 6036 6644 6040 6676
rect 6000 6596 6040 6644
rect 6000 6564 6004 6596
rect 6036 6564 6040 6596
rect 6000 6516 6040 6564
rect 6000 6484 6004 6516
rect 6036 6484 6040 6516
rect 6000 6436 6040 6484
rect 6000 6404 6004 6436
rect 6036 6404 6040 6436
rect 6000 6356 6040 6404
rect 6000 6324 6004 6356
rect 6036 6324 6040 6356
rect 6000 6276 6040 6324
rect 6000 6244 6004 6276
rect 6036 6244 6040 6276
rect 6000 6196 6040 6244
rect 6000 6164 6004 6196
rect 6036 6164 6040 6196
rect 6000 6116 6040 6164
rect 6000 6084 6004 6116
rect 6036 6084 6040 6116
rect 6000 6036 6040 6084
rect 6000 6004 6004 6036
rect 6036 6004 6040 6036
rect 6000 5956 6040 6004
rect 6000 5924 6004 5956
rect 6036 5924 6040 5956
rect 6000 5876 6040 5924
rect 6000 5844 6004 5876
rect 6036 5844 6040 5876
rect 6000 5796 6040 5844
rect 6000 5764 6004 5796
rect 6036 5764 6040 5796
rect 6000 5716 6040 5764
rect 6000 5684 6004 5716
rect 6036 5684 6040 5716
rect 6000 5636 6040 5684
rect 6000 5604 6004 5636
rect 6036 5604 6040 5636
rect 6000 5556 6040 5604
rect 6000 5524 6004 5556
rect 6036 5524 6040 5556
rect 6000 5476 6040 5524
rect 6000 5444 6004 5476
rect 6036 5444 6040 5476
rect 6000 5396 6040 5444
rect 6000 5364 6004 5396
rect 6036 5364 6040 5396
rect 6000 5316 6040 5364
rect 6000 5284 6004 5316
rect 6036 5284 6040 5316
rect 6000 5236 6040 5284
rect 6000 5204 6004 5236
rect 6036 5204 6040 5236
rect 6000 5156 6040 5204
rect 6000 5124 6004 5156
rect 6036 5124 6040 5156
rect 6000 5076 6040 5124
rect 6000 5044 6004 5076
rect 6036 5044 6040 5076
rect 6000 4996 6040 5044
rect 6000 4964 6004 4996
rect 6036 4964 6040 4996
rect 6000 4916 6040 4964
rect 6000 4884 6004 4916
rect 6036 4884 6040 4916
rect 6000 4836 6040 4884
rect 6000 4804 6004 4836
rect 6036 4804 6040 4836
rect 6000 4756 6040 4804
rect 6000 4724 6004 4756
rect 6036 4724 6040 4756
rect 6000 4676 6040 4724
rect 6000 4644 6004 4676
rect 6036 4644 6040 4676
rect 6000 4596 6040 4644
rect 6000 4564 6004 4596
rect 6036 4564 6040 4596
rect 6000 4516 6040 4564
rect 6000 4484 6004 4516
rect 6036 4484 6040 4516
rect 6000 4436 6040 4484
rect 6000 4404 6004 4436
rect 6036 4404 6040 4436
rect 6000 4356 6040 4404
rect 6000 4324 6004 4356
rect 6036 4324 6040 4356
rect 6000 4276 6040 4324
rect 6000 4244 6004 4276
rect 6036 4244 6040 4276
rect 6000 4196 6040 4244
rect 6000 4164 6004 4196
rect 6036 4164 6040 4196
rect 6000 4116 6040 4164
rect 6000 4084 6004 4116
rect 6036 4084 6040 4116
rect 6000 4036 6040 4084
rect 6000 4004 6004 4036
rect 6036 4004 6040 4036
rect 6000 3956 6040 4004
rect 6000 3924 6004 3956
rect 6036 3924 6040 3956
rect 6000 3876 6040 3924
rect 6000 3844 6004 3876
rect 6036 3844 6040 3876
rect 6000 3796 6040 3844
rect 6000 3764 6004 3796
rect 6036 3764 6040 3796
rect 6000 3716 6040 3764
rect 6000 3684 6004 3716
rect 6036 3684 6040 3716
rect 6000 3636 6040 3684
rect 6000 3604 6004 3636
rect 6036 3604 6040 3636
rect 6000 3556 6040 3604
rect 6000 3524 6004 3556
rect 6036 3524 6040 3556
rect 6000 3476 6040 3524
rect 6000 3444 6004 3476
rect 6036 3444 6040 3476
rect 6000 3396 6040 3444
rect 6000 3364 6004 3396
rect 6036 3364 6040 3396
rect 6000 3316 6040 3364
rect 6000 3284 6004 3316
rect 6036 3284 6040 3316
rect 6000 3236 6040 3284
rect 6000 3204 6004 3236
rect 6036 3204 6040 3236
rect 6000 3156 6040 3204
rect 6000 3124 6004 3156
rect 6036 3124 6040 3156
rect 6000 3076 6040 3124
rect 6000 3044 6004 3076
rect 6036 3044 6040 3076
rect 6000 2996 6040 3044
rect 6000 2964 6004 2996
rect 6036 2964 6040 2996
rect 6000 2916 6040 2964
rect 6000 2884 6004 2916
rect 6036 2884 6040 2916
rect 6000 2836 6040 2884
rect 6000 2804 6004 2836
rect 6036 2804 6040 2836
rect 6000 2756 6040 2804
rect 6000 2724 6004 2756
rect 6036 2724 6040 2756
rect 6000 2676 6040 2724
rect 6000 2644 6004 2676
rect 6036 2644 6040 2676
rect 6000 2596 6040 2644
rect 6000 2564 6004 2596
rect 6036 2564 6040 2596
rect 6000 2516 6040 2564
rect 6000 2484 6004 2516
rect 6036 2484 6040 2516
rect 6000 2436 6040 2484
rect 6000 2404 6004 2436
rect 6036 2404 6040 2436
rect 6000 2356 6040 2404
rect 6000 2324 6004 2356
rect 6036 2324 6040 2356
rect 6000 2276 6040 2324
rect 6000 2244 6004 2276
rect 6036 2244 6040 2276
rect 6000 2196 6040 2244
rect 6000 2164 6004 2196
rect 6036 2164 6040 2196
rect 6000 2116 6040 2164
rect 6000 2084 6004 2116
rect 6036 2084 6040 2116
rect 6000 2036 6040 2084
rect 6000 2004 6004 2036
rect 6036 2004 6040 2036
rect 6000 1956 6040 2004
rect 6000 1924 6004 1956
rect 6036 1924 6040 1956
rect 6000 1876 6040 1924
rect 6000 1844 6004 1876
rect 6036 1844 6040 1876
rect 6000 1796 6040 1844
rect 6000 1764 6004 1796
rect 6036 1764 6040 1796
rect 6000 1716 6040 1764
rect 6000 1684 6004 1716
rect 6036 1684 6040 1716
rect 6000 1636 6040 1684
rect 6000 1604 6004 1636
rect 6036 1604 6040 1636
rect 6000 1556 6040 1604
rect 6000 1524 6004 1556
rect 6036 1524 6040 1556
rect 6000 1476 6040 1524
rect 6000 1444 6004 1476
rect 6036 1444 6040 1476
rect 6000 1396 6040 1444
rect 6000 1364 6004 1396
rect 6036 1364 6040 1396
rect 6000 1316 6040 1364
rect 6000 1284 6004 1316
rect 6036 1284 6040 1316
rect 6000 1236 6040 1284
rect 6000 1204 6004 1236
rect 6036 1204 6040 1236
rect 6000 1156 6040 1204
rect 6000 1124 6004 1156
rect 6036 1124 6040 1156
rect 6000 1076 6040 1124
rect 6000 1044 6004 1076
rect 6036 1044 6040 1076
rect 6000 996 6040 1044
rect 6000 964 6004 996
rect 6036 964 6040 996
rect 6000 916 6040 964
rect 6000 884 6004 916
rect 6036 884 6040 916
rect 6000 836 6040 884
rect 6000 804 6004 836
rect 6036 804 6040 836
rect 6000 756 6040 804
rect 6000 724 6004 756
rect 6036 724 6040 756
rect 6000 676 6040 724
rect 6000 644 6004 676
rect 6036 644 6040 676
rect 6000 596 6040 644
rect 6000 564 6004 596
rect 6036 564 6040 596
rect 6000 516 6040 564
rect 6000 484 6004 516
rect 6036 484 6040 516
rect 6000 436 6040 484
rect 6000 404 6004 436
rect 6036 404 6040 436
rect 6000 356 6040 404
rect 6000 324 6004 356
rect 6036 324 6040 356
rect 6000 276 6040 324
rect 6000 244 6004 276
rect 6036 244 6040 276
rect 6000 196 6040 244
rect 6000 164 6004 196
rect 6036 164 6040 196
rect 6000 116 6040 164
rect 6000 84 6004 116
rect 6036 84 6040 116
rect 6000 36 6040 84
rect 6000 4 6004 36
rect 6036 4 6040 36
rect 6000 -524 6040 4
rect 6080 4595 6120 15760
rect 6080 4565 6085 4595
rect 6115 4565 6120 4595
rect 6080 915 6120 4565
rect 6080 885 6085 915
rect 6115 885 6120 915
rect 6080 0 6120 885
rect 6160 15716 6200 15760
rect 6160 15684 6164 15716
rect 6196 15684 6200 15716
rect 6160 15636 6200 15684
rect 6160 15604 6164 15636
rect 6196 15604 6200 15636
rect 6160 15556 6200 15604
rect 6160 15524 6164 15556
rect 6196 15524 6200 15556
rect 6160 15476 6200 15524
rect 6160 15444 6164 15476
rect 6196 15444 6200 15476
rect 6160 15396 6200 15444
rect 6160 15364 6164 15396
rect 6196 15364 6200 15396
rect 6160 15316 6200 15364
rect 6160 15284 6164 15316
rect 6196 15284 6200 15316
rect 6160 15236 6200 15284
rect 6160 15204 6164 15236
rect 6196 15204 6200 15236
rect 6160 15156 6200 15204
rect 6160 15124 6164 15156
rect 6196 15124 6200 15156
rect 6160 15076 6200 15124
rect 6160 15044 6164 15076
rect 6196 15044 6200 15076
rect 6160 14996 6200 15044
rect 6160 14964 6164 14996
rect 6196 14964 6200 14996
rect 6160 14916 6200 14964
rect 6160 14884 6164 14916
rect 6196 14884 6200 14916
rect 6160 14836 6200 14884
rect 6160 14804 6164 14836
rect 6196 14804 6200 14836
rect 6160 14756 6200 14804
rect 6160 14724 6164 14756
rect 6196 14724 6200 14756
rect 6160 14676 6200 14724
rect 6160 14644 6164 14676
rect 6196 14644 6200 14676
rect 6160 14596 6200 14644
rect 6160 14564 6164 14596
rect 6196 14564 6200 14596
rect 6160 14516 6200 14564
rect 6160 14484 6164 14516
rect 6196 14484 6200 14516
rect 6160 14436 6200 14484
rect 6160 14404 6164 14436
rect 6196 14404 6200 14436
rect 6160 14356 6200 14404
rect 6160 14324 6164 14356
rect 6196 14324 6200 14356
rect 6160 14276 6200 14324
rect 6160 14244 6164 14276
rect 6196 14244 6200 14276
rect 6160 14196 6200 14244
rect 6160 14164 6164 14196
rect 6196 14164 6200 14196
rect 6160 14116 6200 14164
rect 6160 14084 6164 14116
rect 6196 14084 6200 14116
rect 6160 14036 6200 14084
rect 6160 14004 6164 14036
rect 6196 14004 6200 14036
rect 6160 13956 6200 14004
rect 6160 13924 6164 13956
rect 6196 13924 6200 13956
rect 6160 13876 6200 13924
rect 6160 13844 6164 13876
rect 6196 13844 6200 13876
rect 6160 13796 6200 13844
rect 6160 13764 6164 13796
rect 6196 13764 6200 13796
rect 6160 13716 6200 13764
rect 6160 13684 6164 13716
rect 6196 13684 6200 13716
rect 6160 13636 6200 13684
rect 6160 13604 6164 13636
rect 6196 13604 6200 13636
rect 6160 13556 6200 13604
rect 6160 13524 6164 13556
rect 6196 13524 6200 13556
rect 6160 13476 6200 13524
rect 6160 13444 6164 13476
rect 6196 13444 6200 13476
rect 6160 13396 6200 13444
rect 6160 13364 6164 13396
rect 6196 13364 6200 13396
rect 6160 13316 6200 13364
rect 6160 13284 6164 13316
rect 6196 13284 6200 13316
rect 6160 13236 6200 13284
rect 6160 13204 6164 13236
rect 6196 13204 6200 13236
rect 6160 13156 6200 13204
rect 6160 13124 6164 13156
rect 6196 13124 6200 13156
rect 6160 13076 6200 13124
rect 6160 13044 6164 13076
rect 6196 13044 6200 13076
rect 6160 12996 6200 13044
rect 6160 12964 6164 12996
rect 6196 12964 6200 12996
rect 6160 12916 6200 12964
rect 6160 12884 6164 12916
rect 6196 12884 6200 12916
rect 6160 12836 6200 12884
rect 6160 12804 6164 12836
rect 6196 12804 6200 12836
rect 6160 12756 6200 12804
rect 6160 12724 6164 12756
rect 6196 12724 6200 12756
rect 6160 12676 6200 12724
rect 6160 12644 6164 12676
rect 6196 12644 6200 12676
rect 6160 12596 6200 12644
rect 6160 12564 6164 12596
rect 6196 12564 6200 12596
rect 6160 12516 6200 12564
rect 6160 12484 6164 12516
rect 6196 12484 6200 12516
rect 6160 12436 6200 12484
rect 6160 12404 6164 12436
rect 6196 12404 6200 12436
rect 6160 12356 6200 12404
rect 6160 12324 6164 12356
rect 6196 12324 6200 12356
rect 6160 12276 6200 12324
rect 6160 12244 6164 12276
rect 6196 12244 6200 12276
rect 6160 12196 6200 12244
rect 6160 12164 6164 12196
rect 6196 12164 6200 12196
rect 6160 12116 6200 12164
rect 6160 12084 6164 12116
rect 6196 12084 6200 12116
rect 6160 12036 6200 12084
rect 6160 12004 6164 12036
rect 6196 12004 6200 12036
rect 6160 11956 6200 12004
rect 6160 11924 6164 11956
rect 6196 11924 6200 11956
rect 6160 11876 6200 11924
rect 6160 11844 6164 11876
rect 6196 11844 6200 11876
rect 6160 11796 6200 11844
rect 6160 11764 6164 11796
rect 6196 11764 6200 11796
rect 6160 11716 6200 11764
rect 6160 11684 6164 11716
rect 6196 11684 6200 11716
rect 6160 11636 6200 11684
rect 6160 11604 6164 11636
rect 6196 11604 6200 11636
rect 6160 11556 6200 11604
rect 6160 11524 6164 11556
rect 6196 11524 6200 11556
rect 6160 11476 6200 11524
rect 6160 11444 6164 11476
rect 6196 11444 6200 11476
rect 6160 11396 6200 11444
rect 6160 11364 6164 11396
rect 6196 11364 6200 11396
rect 6160 11316 6200 11364
rect 6160 11284 6164 11316
rect 6196 11284 6200 11316
rect 6160 11236 6200 11284
rect 6160 11204 6164 11236
rect 6196 11204 6200 11236
rect 6160 11156 6200 11204
rect 6160 11124 6164 11156
rect 6196 11124 6200 11156
rect 6160 11076 6200 11124
rect 6160 11044 6164 11076
rect 6196 11044 6200 11076
rect 6160 10996 6200 11044
rect 6160 10964 6164 10996
rect 6196 10964 6200 10996
rect 6160 10916 6200 10964
rect 6160 10884 6164 10916
rect 6196 10884 6200 10916
rect 6160 10836 6200 10884
rect 6160 10804 6164 10836
rect 6196 10804 6200 10836
rect 6160 10756 6200 10804
rect 6160 10724 6164 10756
rect 6196 10724 6200 10756
rect 6160 10676 6200 10724
rect 6160 10644 6164 10676
rect 6196 10644 6200 10676
rect 6160 10596 6200 10644
rect 6160 10564 6164 10596
rect 6196 10564 6200 10596
rect 6160 10516 6200 10564
rect 6160 10484 6164 10516
rect 6196 10484 6200 10516
rect 6160 10436 6200 10484
rect 6160 10404 6164 10436
rect 6196 10404 6200 10436
rect 6160 10356 6200 10404
rect 6160 10324 6164 10356
rect 6196 10324 6200 10356
rect 6160 10276 6200 10324
rect 6160 10244 6164 10276
rect 6196 10244 6200 10276
rect 6160 10196 6200 10244
rect 6160 10164 6164 10196
rect 6196 10164 6200 10196
rect 6160 10116 6200 10164
rect 6160 10084 6164 10116
rect 6196 10084 6200 10116
rect 6160 10036 6200 10084
rect 6160 10004 6164 10036
rect 6196 10004 6200 10036
rect 6160 9956 6200 10004
rect 6160 9924 6164 9956
rect 6196 9924 6200 9956
rect 6160 9876 6200 9924
rect 6160 9844 6164 9876
rect 6196 9844 6200 9876
rect 6160 9796 6200 9844
rect 6160 9764 6164 9796
rect 6196 9764 6200 9796
rect 6160 9716 6200 9764
rect 6160 9684 6164 9716
rect 6196 9684 6200 9716
rect 6160 9636 6200 9684
rect 6160 9604 6164 9636
rect 6196 9604 6200 9636
rect 6160 9556 6200 9604
rect 6160 9524 6164 9556
rect 6196 9524 6200 9556
rect 6160 9476 6200 9524
rect 6160 9444 6164 9476
rect 6196 9444 6200 9476
rect 6160 9396 6200 9444
rect 6160 9364 6164 9396
rect 6196 9364 6200 9396
rect 6160 9316 6200 9364
rect 6160 9284 6164 9316
rect 6196 9284 6200 9316
rect 6160 9236 6200 9284
rect 6160 9204 6164 9236
rect 6196 9204 6200 9236
rect 6160 9156 6200 9204
rect 6160 9124 6164 9156
rect 6196 9124 6200 9156
rect 6160 9076 6200 9124
rect 6160 9044 6164 9076
rect 6196 9044 6200 9076
rect 6160 8996 6200 9044
rect 6160 8964 6164 8996
rect 6196 8964 6200 8996
rect 6160 8916 6200 8964
rect 6160 8884 6164 8916
rect 6196 8884 6200 8916
rect 6160 8836 6200 8884
rect 6160 8804 6164 8836
rect 6196 8804 6200 8836
rect 6160 8756 6200 8804
rect 6160 8724 6164 8756
rect 6196 8724 6200 8756
rect 6160 8676 6200 8724
rect 6160 8644 6164 8676
rect 6196 8644 6200 8676
rect 6160 8596 6200 8644
rect 6160 8564 6164 8596
rect 6196 8564 6200 8596
rect 6160 8516 6200 8564
rect 6160 8484 6164 8516
rect 6196 8484 6200 8516
rect 6160 8436 6200 8484
rect 6160 8404 6164 8436
rect 6196 8404 6200 8436
rect 6160 8356 6200 8404
rect 6160 8324 6164 8356
rect 6196 8324 6200 8356
rect 6160 8276 6200 8324
rect 6160 8244 6164 8276
rect 6196 8244 6200 8276
rect 6160 8196 6200 8244
rect 6160 8164 6164 8196
rect 6196 8164 6200 8196
rect 6160 8116 6200 8164
rect 6160 8084 6164 8116
rect 6196 8084 6200 8116
rect 6160 8036 6200 8084
rect 6160 8004 6164 8036
rect 6196 8004 6200 8036
rect 6160 7956 6200 8004
rect 6160 7924 6164 7956
rect 6196 7924 6200 7956
rect 6160 7876 6200 7924
rect 6160 7844 6164 7876
rect 6196 7844 6200 7876
rect 6160 7796 6200 7844
rect 6160 7764 6164 7796
rect 6196 7764 6200 7796
rect 6160 7716 6200 7764
rect 6160 7684 6164 7716
rect 6196 7684 6200 7716
rect 6160 7636 6200 7684
rect 6160 7604 6164 7636
rect 6196 7604 6200 7636
rect 6160 7556 6200 7604
rect 6160 7524 6164 7556
rect 6196 7524 6200 7556
rect 6160 7476 6200 7524
rect 6160 7444 6164 7476
rect 6196 7444 6200 7476
rect 6160 7396 6200 7444
rect 6160 7364 6164 7396
rect 6196 7364 6200 7396
rect 6160 7316 6200 7364
rect 6160 7284 6164 7316
rect 6196 7284 6200 7316
rect 6160 7236 6200 7284
rect 6160 7204 6164 7236
rect 6196 7204 6200 7236
rect 6160 7156 6200 7204
rect 6160 7124 6164 7156
rect 6196 7124 6200 7156
rect 6160 7076 6200 7124
rect 6160 7044 6164 7076
rect 6196 7044 6200 7076
rect 6160 6996 6200 7044
rect 6160 6964 6164 6996
rect 6196 6964 6200 6996
rect 6160 6916 6200 6964
rect 6160 6884 6164 6916
rect 6196 6884 6200 6916
rect 6160 6836 6200 6884
rect 6160 6804 6164 6836
rect 6196 6804 6200 6836
rect 6160 6756 6200 6804
rect 6160 6724 6164 6756
rect 6196 6724 6200 6756
rect 6160 6676 6200 6724
rect 6160 6644 6164 6676
rect 6196 6644 6200 6676
rect 6160 6596 6200 6644
rect 6160 6564 6164 6596
rect 6196 6564 6200 6596
rect 6160 6516 6200 6564
rect 6160 6484 6164 6516
rect 6196 6484 6200 6516
rect 6160 6436 6200 6484
rect 6160 6404 6164 6436
rect 6196 6404 6200 6436
rect 6160 6356 6200 6404
rect 6160 6324 6164 6356
rect 6196 6324 6200 6356
rect 6160 6276 6200 6324
rect 6160 6244 6164 6276
rect 6196 6244 6200 6276
rect 6160 6196 6200 6244
rect 6160 6164 6164 6196
rect 6196 6164 6200 6196
rect 6160 6116 6200 6164
rect 6160 6084 6164 6116
rect 6196 6084 6200 6116
rect 6160 6036 6200 6084
rect 6160 6004 6164 6036
rect 6196 6004 6200 6036
rect 6160 5956 6200 6004
rect 6160 5924 6164 5956
rect 6196 5924 6200 5956
rect 6160 5876 6200 5924
rect 6160 5844 6164 5876
rect 6196 5844 6200 5876
rect 6160 5796 6200 5844
rect 6160 5764 6164 5796
rect 6196 5764 6200 5796
rect 6160 5716 6200 5764
rect 6160 5684 6164 5716
rect 6196 5684 6200 5716
rect 6160 5636 6200 5684
rect 6160 5604 6164 5636
rect 6196 5604 6200 5636
rect 6160 5556 6200 5604
rect 6160 5524 6164 5556
rect 6196 5524 6200 5556
rect 6160 5476 6200 5524
rect 6160 5444 6164 5476
rect 6196 5444 6200 5476
rect 6160 5396 6200 5444
rect 6160 5364 6164 5396
rect 6196 5364 6200 5396
rect 6160 5316 6200 5364
rect 6160 5284 6164 5316
rect 6196 5284 6200 5316
rect 6160 5236 6200 5284
rect 6160 5204 6164 5236
rect 6196 5204 6200 5236
rect 6160 5156 6200 5204
rect 6160 5124 6164 5156
rect 6196 5124 6200 5156
rect 6160 5076 6200 5124
rect 6160 5044 6164 5076
rect 6196 5044 6200 5076
rect 6160 4996 6200 5044
rect 6160 4964 6164 4996
rect 6196 4964 6200 4996
rect 6160 4916 6200 4964
rect 6160 4884 6164 4916
rect 6196 4884 6200 4916
rect 6160 4836 6200 4884
rect 6160 4804 6164 4836
rect 6196 4804 6200 4836
rect 6160 4756 6200 4804
rect 6160 4724 6164 4756
rect 6196 4724 6200 4756
rect 6160 4676 6200 4724
rect 6160 4644 6164 4676
rect 6196 4644 6200 4676
rect 6160 4596 6200 4644
rect 6160 4564 6164 4596
rect 6196 4564 6200 4596
rect 6160 4516 6200 4564
rect 6160 4484 6164 4516
rect 6196 4484 6200 4516
rect 6160 4436 6200 4484
rect 6160 4404 6164 4436
rect 6196 4404 6200 4436
rect 6160 4356 6200 4404
rect 6160 4324 6164 4356
rect 6196 4324 6200 4356
rect 6160 4276 6200 4324
rect 6160 4244 6164 4276
rect 6196 4244 6200 4276
rect 6160 4196 6200 4244
rect 6160 4164 6164 4196
rect 6196 4164 6200 4196
rect 6160 4116 6200 4164
rect 6160 4084 6164 4116
rect 6196 4084 6200 4116
rect 6160 4036 6200 4084
rect 6160 4004 6164 4036
rect 6196 4004 6200 4036
rect 6160 3956 6200 4004
rect 6160 3924 6164 3956
rect 6196 3924 6200 3956
rect 6160 3876 6200 3924
rect 6160 3844 6164 3876
rect 6196 3844 6200 3876
rect 6160 3796 6200 3844
rect 6160 3764 6164 3796
rect 6196 3764 6200 3796
rect 6160 3716 6200 3764
rect 6160 3684 6164 3716
rect 6196 3684 6200 3716
rect 6160 3636 6200 3684
rect 6160 3604 6164 3636
rect 6196 3604 6200 3636
rect 6160 3556 6200 3604
rect 6160 3524 6164 3556
rect 6196 3524 6200 3556
rect 6160 3476 6200 3524
rect 6160 3444 6164 3476
rect 6196 3444 6200 3476
rect 6160 3396 6200 3444
rect 6160 3364 6164 3396
rect 6196 3364 6200 3396
rect 6160 3316 6200 3364
rect 6160 3284 6164 3316
rect 6196 3284 6200 3316
rect 6160 3236 6200 3284
rect 6160 3204 6164 3236
rect 6196 3204 6200 3236
rect 6160 3156 6200 3204
rect 6160 3124 6164 3156
rect 6196 3124 6200 3156
rect 6160 3076 6200 3124
rect 6160 3044 6164 3076
rect 6196 3044 6200 3076
rect 6160 2996 6200 3044
rect 6160 2964 6164 2996
rect 6196 2964 6200 2996
rect 6160 2916 6200 2964
rect 6160 2884 6164 2916
rect 6196 2884 6200 2916
rect 6160 2836 6200 2884
rect 6160 2804 6164 2836
rect 6196 2804 6200 2836
rect 6160 2756 6200 2804
rect 6160 2724 6164 2756
rect 6196 2724 6200 2756
rect 6160 2676 6200 2724
rect 6160 2644 6164 2676
rect 6196 2644 6200 2676
rect 6160 2596 6200 2644
rect 6160 2564 6164 2596
rect 6196 2564 6200 2596
rect 6160 2516 6200 2564
rect 6160 2484 6164 2516
rect 6196 2484 6200 2516
rect 6160 2436 6200 2484
rect 6160 2404 6164 2436
rect 6196 2404 6200 2436
rect 6160 2356 6200 2404
rect 6160 2324 6164 2356
rect 6196 2324 6200 2356
rect 6160 2276 6200 2324
rect 6160 2244 6164 2276
rect 6196 2244 6200 2276
rect 6160 2196 6200 2244
rect 6160 2164 6164 2196
rect 6196 2164 6200 2196
rect 6160 2116 6200 2164
rect 6160 2084 6164 2116
rect 6196 2084 6200 2116
rect 6160 2036 6200 2084
rect 6160 2004 6164 2036
rect 6196 2004 6200 2036
rect 6160 1956 6200 2004
rect 6160 1924 6164 1956
rect 6196 1924 6200 1956
rect 6160 1876 6200 1924
rect 6160 1844 6164 1876
rect 6196 1844 6200 1876
rect 6160 1796 6200 1844
rect 6160 1764 6164 1796
rect 6196 1764 6200 1796
rect 6160 1716 6200 1764
rect 6160 1684 6164 1716
rect 6196 1684 6200 1716
rect 6160 1636 6200 1684
rect 6160 1604 6164 1636
rect 6196 1604 6200 1636
rect 6160 1556 6200 1604
rect 6160 1524 6164 1556
rect 6196 1524 6200 1556
rect 6160 1476 6200 1524
rect 6160 1444 6164 1476
rect 6196 1444 6200 1476
rect 6160 1396 6200 1444
rect 6160 1364 6164 1396
rect 6196 1364 6200 1396
rect 6160 1316 6200 1364
rect 6160 1284 6164 1316
rect 6196 1284 6200 1316
rect 6160 1236 6200 1284
rect 6160 1204 6164 1236
rect 6196 1204 6200 1236
rect 6160 1156 6200 1204
rect 6160 1124 6164 1156
rect 6196 1124 6200 1156
rect 6160 1076 6200 1124
rect 6160 1044 6164 1076
rect 6196 1044 6200 1076
rect 6160 996 6200 1044
rect 6160 964 6164 996
rect 6196 964 6200 996
rect 6160 916 6200 964
rect 6160 884 6164 916
rect 6196 884 6200 916
rect 6160 836 6200 884
rect 6160 804 6164 836
rect 6196 804 6200 836
rect 6160 756 6200 804
rect 6160 724 6164 756
rect 6196 724 6200 756
rect 6160 676 6200 724
rect 6160 644 6164 676
rect 6196 644 6200 676
rect 6160 596 6200 644
rect 6160 564 6164 596
rect 6196 564 6200 596
rect 6160 516 6200 564
rect 6160 484 6164 516
rect 6196 484 6200 516
rect 6160 436 6200 484
rect 6160 404 6164 436
rect 6196 404 6200 436
rect 6160 356 6200 404
rect 6160 324 6164 356
rect 6196 324 6200 356
rect 6160 276 6200 324
rect 6160 244 6164 276
rect 6196 244 6200 276
rect 6160 196 6200 244
rect 6160 164 6164 196
rect 6196 164 6200 196
rect 6160 116 6200 164
rect 6160 84 6164 116
rect 6196 84 6200 116
rect 6160 36 6200 84
rect 6160 4 6164 36
rect 6196 4 6200 36
rect 6000 -716 6004 -524
rect 6036 -716 6040 -524
rect 6000 -960 6040 -716
rect 6160 -524 6200 4
rect 6160 -716 6164 -524
rect 6196 -716 6200 -524
rect 6160 -960 6200 -716
rect 4640 -1036 4644 -1004
rect 4676 -1036 4680 -1004
rect 4640 -1040 4680 -1036
rect 10280 -1004 10320 -1000
rect 10280 -1036 10284 -1004
rect 10316 -1036 10320 -1004
rect 240 -1084 280 -1080
rect 240 -1116 244 -1084
rect 276 -1116 280 -1084
rect 240 -1160 280 -1116
rect 1200 -1084 1240 -1080
rect 1200 -1116 1204 -1084
rect 1236 -1116 1240 -1084
rect 1200 -1160 1240 -1116
rect 240 -2240 1240 -1160
rect 1360 -1084 1400 -1080
rect 1360 -1116 1364 -1084
rect 1396 -1116 1400 -1084
rect 1360 -1160 1400 -1116
rect 2320 -1084 2360 -1080
rect 2320 -1116 2324 -1084
rect 2356 -1116 2360 -1084
rect 2320 -1160 2360 -1116
rect 1360 -2240 2360 -1160
rect 2480 -1084 2520 -1080
rect 2480 -1116 2484 -1084
rect 2516 -1116 2520 -1084
rect 2480 -1160 2520 -1116
rect 3440 -1084 3480 -1080
rect 3440 -1116 3444 -1084
rect 3476 -1116 3480 -1084
rect 3440 -1160 3480 -1116
rect 2480 -2240 3480 -1160
rect 3600 -1084 4600 -1080
rect 3600 -1116 3604 -1084
rect 3636 -1116 4564 -1084
rect 4596 -1116 4600 -1084
rect 3600 -2240 4600 -1116
rect 4720 -1084 4760 -1080
rect 4720 -1116 4724 -1084
rect 4756 -1116 4760 -1084
rect 4720 -1160 4760 -1116
rect 5680 -1084 5720 -1080
rect 5680 -1116 5684 -1084
rect 5716 -1116 5720 -1084
rect 5680 -1160 5720 -1116
rect 4720 -2240 5720 -1160
rect 5840 -1084 6840 -1080
rect 5840 -1116 5844 -1084
rect 5876 -1116 6804 -1084
rect 6836 -1116 6840 -1084
rect 5840 -2240 6840 -1116
rect 6960 -1084 7000 -1080
rect 6960 -1116 6964 -1084
rect 6996 -1116 7000 -1084
rect 6960 -1160 7000 -1116
rect 7920 -1084 7960 -1080
rect 7920 -1116 7924 -1084
rect 7956 -1116 7960 -1084
rect 7920 -1160 7960 -1116
rect 6960 -2240 7960 -1160
rect 8080 -1084 8120 -1080
rect 8080 -1116 8084 -1084
rect 8116 -1116 8120 -1084
rect 8080 -1160 8120 -1116
rect 9040 -1084 9080 -1080
rect 9040 -1116 9044 -1084
rect 9076 -1116 9080 -1084
rect 9040 -1160 9080 -1116
rect 8080 -2240 9080 -1160
rect 9200 -1084 9240 -1080
rect 9200 -1116 9204 -1084
rect 9236 -1116 9240 -1084
rect 9200 -1160 9240 -1116
rect 10160 -1084 10200 -1080
rect 10160 -1116 10164 -1084
rect 10196 -1116 10200 -1084
rect 10160 -1160 10200 -1116
rect 9200 -2240 10200 -1160
rect 120 -2316 124 -2284
rect 156 -2316 160 -2284
rect 120 -2320 160 -2316
rect 10280 -2284 10320 -1036
rect 10280 -2316 10284 -2284
rect 10316 -2316 10320 -2284
rect 10280 -2320 10320 -2316
<< via3 >>
rect 4244 15715 4276 15716
rect 4244 15685 4245 15715
rect 4245 15685 4275 15715
rect 4275 15685 4276 15715
rect 4244 15684 4276 15685
rect 4244 15635 4276 15636
rect 4244 15605 4245 15635
rect 4245 15605 4275 15635
rect 4275 15605 4276 15635
rect 4244 15604 4276 15605
rect 4244 15555 4276 15556
rect 4244 15525 4245 15555
rect 4245 15525 4275 15555
rect 4275 15525 4276 15555
rect 4244 15524 4276 15525
rect 4244 15475 4276 15476
rect 4244 15445 4245 15475
rect 4245 15445 4275 15475
rect 4275 15445 4276 15475
rect 4244 15444 4276 15445
rect 4244 15395 4276 15396
rect 4244 15365 4245 15395
rect 4245 15365 4275 15395
rect 4275 15365 4276 15395
rect 4244 15364 4276 15365
rect 4244 15315 4276 15316
rect 4244 15285 4245 15315
rect 4245 15285 4275 15315
rect 4275 15285 4276 15315
rect 4244 15284 4276 15285
rect 4244 15235 4276 15236
rect 4244 15205 4245 15235
rect 4245 15205 4275 15235
rect 4275 15205 4276 15235
rect 4244 15204 4276 15205
rect 4244 15155 4276 15156
rect 4244 15125 4245 15155
rect 4245 15125 4275 15155
rect 4275 15125 4276 15155
rect 4244 15124 4276 15125
rect 4244 15044 4276 15076
rect 4244 14995 4276 14996
rect 4244 14965 4245 14995
rect 4245 14965 4275 14995
rect 4275 14965 4276 14995
rect 4244 14964 4276 14965
rect 4244 14915 4276 14916
rect 4244 14885 4245 14915
rect 4245 14885 4275 14915
rect 4275 14885 4276 14915
rect 4244 14884 4276 14885
rect 4244 14835 4276 14836
rect 4244 14805 4245 14835
rect 4245 14805 4275 14835
rect 4275 14805 4276 14835
rect 4244 14804 4276 14805
rect 4244 14755 4276 14756
rect 4244 14725 4245 14755
rect 4245 14725 4275 14755
rect 4275 14725 4276 14755
rect 4244 14724 4276 14725
rect 4244 14675 4276 14676
rect 4244 14645 4245 14675
rect 4245 14645 4275 14675
rect 4275 14645 4276 14675
rect 4244 14644 4276 14645
rect 4244 14595 4276 14596
rect 4244 14565 4245 14595
rect 4245 14565 4275 14595
rect 4275 14565 4276 14595
rect 4244 14564 4276 14565
rect 4244 14515 4276 14516
rect 4244 14485 4245 14515
rect 4245 14485 4275 14515
rect 4275 14485 4276 14515
rect 4244 14484 4276 14485
rect 4244 14435 4276 14436
rect 4244 14405 4245 14435
rect 4245 14405 4275 14435
rect 4275 14405 4276 14435
rect 4244 14404 4276 14405
rect 4244 14324 4276 14356
rect 4244 14244 4276 14276
rect 4244 14164 4276 14196
rect 4244 14084 4276 14116
rect 4244 14035 4276 14036
rect 4244 14005 4245 14035
rect 4245 14005 4275 14035
rect 4275 14005 4276 14035
rect 4244 14004 4276 14005
rect 4244 13955 4276 13956
rect 4244 13925 4245 13955
rect 4245 13925 4275 13955
rect 4275 13925 4276 13955
rect 4244 13924 4276 13925
rect 4244 13875 4276 13876
rect 4244 13845 4245 13875
rect 4245 13845 4275 13875
rect 4275 13845 4276 13875
rect 4244 13844 4276 13845
rect 4244 13795 4276 13796
rect 4244 13765 4245 13795
rect 4245 13765 4275 13795
rect 4275 13765 4276 13795
rect 4244 13764 4276 13765
rect 4244 13715 4276 13716
rect 4244 13685 4245 13715
rect 4245 13685 4275 13715
rect 4275 13685 4276 13715
rect 4244 13684 4276 13685
rect 4244 13635 4276 13636
rect 4244 13605 4245 13635
rect 4245 13605 4275 13635
rect 4275 13605 4276 13635
rect 4244 13604 4276 13605
rect 4244 13555 4276 13556
rect 4244 13525 4245 13555
rect 4245 13525 4275 13555
rect 4275 13525 4276 13555
rect 4244 13524 4276 13525
rect 4244 13475 4276 13476
rect 4244 13445 4245 13475
rect 4245 13445 4275 13475
rect 4275 13445 4276 13475
rect 4244 13444 4276 13445
rect 4244 13364 4276 13396
rect 4244 13284 4276 13316
rect 4244 13204 4276 13236
rect 4244 13124 4276 13156
rect 4244 13075 4276 13076
rect 4244 13045 4245 13075
rect 4245 13045 4275 13075
rect 4275 13045 4276 13075
rect 4244 13044 4276 13045
rect 4244 12995 4276 12996
rect 4244 12965 4245 12995
rect 4245 12965 4275 12995
rect 4275 12965 4276 12995
rect 4244 12964 4276 12965
rect 4244 12915 4276 12916
rect 4244 12885 4245 12915
rect 4245 12885 4275 12915
rect 4275 12885 4276 12915
rect 4244 12884 4276 12885
rect 4244 12835 4276 12836
rect 4244 12805 4245 12835
rect 4245 12805 4275 12835
rect 4275 12805 4276 12835
rect 4244 12804 4276 12805
rect 4244 12755 4276 12756
rect 4244 12725 4245 12755
rect 4245 12725 4275 12755
rect 4275 12725 4276 12755
rect 4244 12724 4276 12725
rect 4244 12675 4276 12676
rect 4244 12645 4245 12675
rect 4245 12645 4275 12675
rect 4275 12645 4276 12675
rect 4244 12644 4276 12645
rect 4244 12595 4276 12596
rect 4244 12565 4245 12595
rect 4245 12565 4275 12595
rect 4275 12565 4276 12595
rect 4244 12564 4276 12565
rect 4244 12515 4276 12516
rect 4244 12485 4245 12515
rect 4245 12485 4275 12515
rect 4275 12485 4276 12515
rect 4244 12484 4276 12485
rect 4244 12404 4276 12436
rect 4244 12355 4276 12356
rect 4244 12325 4245 12355
rect 4245 12325 4275 12355
rect 4275 12325 4276 12355
rect 4244 12324 4276 12325
rect 4244 12275 4276 12276
rect 4244 12245 4245 12275
rect 4245 12245 4275 12275
rect 4275 12245 4276 12275
rect 4244 12244 4276 12245
rect 4244 12195 4276 12196
rect 4244 12165 4245 12195
rect 4245 12165 4275 12195
rect 4275 12165 4276 12195
rect 4244 12164 4276 12165
rect 4244 12115 4276 12116
rect 4244 12085 4245 12115
rect 4245 12085 4275 12115
rect 4275 12085 4276 12115
rect 4244 12084 4276 12085
rect 4244 12035 4276 12036
rect 4244 12005 4245 12035
rect 4245 12005 4275 12035
rect 4275 12005 4276 12035
rect 4244 12004 4276 12005
rect 4244 11955 4276 11956
rect 4244 11925 4245 11955
rect 4245 11925 4275 11955
rect 4275 11925 4276 11955
rect 4244 11924 4276 11925
rect 4244 11875 4276 11876
rect 4244 11845 4245 11875
rect 4245 11845 4275 11875
rect 4275 11845 4276 11875
rect 4244 11844 4276 11845
rect 4244 11795 4276 11796
rect 4244 11765 4245 11795
rect 4245 11765 4275 11795
rect 4275 11765 4276 11795
rect 4244 11764 4276 11765
rect 4244 11715 4276 11716
rect 4244 11685 4245 11715
rect 4245 11685 4275 11715
rect 4275 11685 4276 11715
rect 4244 11684 4276 11685
rect 4244 11635 4276 11636
rect 4244 11605 4245 11635
rect 4245 11605 4275 11635
rect 4275 11605 4276 11635
rect 4244 11604 4276 11605
rect 4244 11555 4276 11556
rect 4244 11525 4245 11555
rect 4245 11525 4275 11555
rect 4275 11525 4276 11555
rect 4244 11524 4276 11525
rect 4244 11475 4276 11476
rect 4244 11445 4245 11475
rect 4245 11445 4275 11475
rect 4275 11445 4276 11475
rect 4244 11444 4276 11445
rect 4244 11395 4276 11396
rect 4244 11365 4245 11395
rect 4245 11365 4275 11395
rect 4275 11365 4276 11395
rect 4244 11364 4276 11365
rect 4244 11315 4276 11316
rect 4244 11285 4245 11315
rect 4245 11285 4275 11315
rect 4275 11285 4276 11315
rect 4244 11284 4276 11285
rect 4244 11235 4276 11236
rect 4244 11205 4245 11235
rect 4245 11205 4275 11235
rect 4275 11205 4276 11235
rect 4244 11204 4276 11205
rect 4244 11155 4276 11156
rect 4244 11125 4245 11155
rect 4245 11125 4275 11155
rect 4275 11125 4276 11155
rect 4244 11124 4276 11125
rect 4244 11075 4276 11076
rect 4244 11045 4245 11075
rect 4245 11045 4275 11075
rect 4275 11045 4276 11075
rect 4244 11044 4276 11045
rect 4244 10964 4276 10996
rect 4244 10915 4276 10916
rect 4244 10885 4245 10915
rect 4245 10885 4275 10915
rect 4275 10885 4276 10915
rect 4244 10884 4276 10885
rect 4244 10835 4276 10836
rect 4244 10805 4245 10835
rect 4245 10805 4275 10835
rect 4275 10805 4276 10835
rect 4244 10804 4276 10805
rect 4244 10755 4276 10756
rect 4244 10725 4245 10755
rect 4245 10725 4275 10755
rect 4275 10725 4276 10755
rect 4244 10724 4276 10725
rect 4244 10675 4276 10676
rect 4244 10645 4245 10675
rect 4245 10645 4275 10675
rect 4275 10645 4276 10675
rect 4244 10644 4276 10645
rect 4244 10595 4276 10596
rect 4244 10565 4245 10595
rect 4245 10565 4275 10595
rect 4275 10565 4276 10595
rect 4244 10564 4276 10565
rect 4244 10515 4276 10516
rect 4244 10485 4245 10515
rect 4245 10485 4275 10515
rect 4275 10485 4276 10515
rect 4244 10484 4276 10485
rect 4244 10435 4276 10436
rect 4244 10405 4245 10435
rect 4245 10405 4275 10435
rect 4275 10405 4276 10435
rect 4244 10404 4276 10405
rect 4244 10355 4276 10356
rect 4244 10325 4245 10355
rect 4245 10325 4275 10355
rect 4275 10325 4276 10355
rect 4244 10324 4276 10325
rect 4244 10244 4276 10276
rect 4244 10164 4276 10196
rect 4244 10084 4276 10116
rect 4244 10004 4276 10036
rect 4244 9955 4276 9956
rect 4244 9925 4245 9955
rect 4245 9925 4275 9955
rect 4275 9925 4276 9955
rect 4244 9924 4276 9925
rect 4244 9875 4276 9876
rect 4244 9845 4245 9875
rect 4245 9845 4275 9875
rect 4275 9845 4276 9875
rect 4244 9844 4276 9845
rect 4244 9795 4276 9796
rect 4244 9765 4245 9795
rect 4245 9765 4275 9795
rect 4275 9765 4276 9795
rect 4244 9764 4276 9765
rect 4244 9715 4276 9716
rect 4244 9685 4245 9715
rect 4245 9685 4275 9715
rect 4275 9685 4276 9715
rect 4244 9684 4276 9685
rect 4244 9635 4276 9636
rect 4244 9605 4245 9635
rect 4245 9605 4275 9635
rect 4275 9605 4276 9635
rect 4244 9604 4276 9605
rect 4244 9555 4276 9556
rect 4244 9525 4245 9555
rect 4245 9525 4275 9555
rect 4275 9525 4276 9555
rect 4244 9524 4276 9525
rect 4244 9475 4276 9476
rect 4244 9445 4245 9475
rect 4245 9445 4275 9475
rect 4275 9445 4276 9475
rect 4244 9444 4276 9445
rect 4244 9395 4276 9396
rect 4244 9365 4245 9395
rect 4245 9365 4275 9395
rect 4275 9365 4276 9395
rect 4244 9364 4276 9365
rect 4244 9284 4276 9316
rect 4244 9204 4276 9236
rect 4244 9124 4276 9156
rect 4244 9044 4276 9076
rect 4244 8995 4276 8996
rect 4244 8965 4245 8995
rect 4245 8965 4275 8995
rect 4275 8965 4276 8995
rect 4244 8964 4276 8965
rect 4244 8915 4276 8916
rect 4244 8885 4245 8915
rect 4245 8885 4275 8915
rect 4275 8885 4276 8915
rect 4244 8884 4276 8885
rect 4244 8835 4276 8836
rect 4244 8805 4245 8835
rect 4245 8805 4275 8835
rect 4275 8805 4276 8835
rect 4244 8804 4276 8805
rect 4244 8755 4276 8756
rect 4244 8725 4245 8755
rect 4245 8725 4275 8755
rect 4275 8725 4276 8755
rect 4244 8724 4276 8725
rect 4244 8675 4276 8676
rect 4244 8645 4245 8675
rect 4245 8645 4275 8675
rect 4275 8645 4276 8675
rect 4244 8644 4276 8645
rect 4244 8595 4276 8596
rect 4244 8565 4245 8595
rect 4245 8565 4275 8595
rect 4275 8565 4276 8595
rect 4244 8564 4276 8565
rect 4244 8515 4276 8516
rect 4244 8485 4245 8515
rect 4245 8485 4275 8515
rect 4275 8485 4276 8515
rect 4244 8484 4276 8485
rect 4244 8435 4276 8436
rect 4244 8405 4245 8435
rect 4245 8405 4275 8435
rect 4275 8405 4276 8435
rect 4244 8404 4276 8405
rect 4244 8324 4276 8356
rect 4244 8275 4276 8276
rect 4244 8245 4245 8275
rect 4245 8245 4275 8275
rect 4275 8245 4276 8275
rect 4244 8244 4276 8245
rect 4244 8195 4276 8196
rect 4244 8165 4245 8195
rect 4245 8165 4275 8195
rect 4275 8165 4276 8195
rect 4244 8164 4276 8165
rect 4244 8115 4276 8116
rect 4244 8085 4245 8115
rect 4245 8085 4275 8115
rect 4275 8085 4276 8115
rect 4244 8084 4276 8085
rect 4244 8035 4276 8036
rect 4244 8005 4245 8035
rect 4245 8005 4275 8035
rect 4275 8005 4276 8035
rect 4244 8004 4276 8005
rect 4244 7955 4276 7956
rect 4244 7925 4245 7955
rect 4245 7925 4275 7955
rect 4275 7925 4276 7955
rect 4244 7924 4276 7925
rect 4244 7875 4276 7876
rect 4244 7845 4245 7875
rect 4245 7845 4275 7875
rect 4275 7845 4276 7875
rect 4244 7844 4276 7845
rect 4244 7795 4276 7796
rect 4244 7765 4245 7795
rect 4245 7765 4275 7795
rect 4275 7765 4276 7795
rect 4244 7764 4276 7765
rect 4244 7715 4276 7716
rect 4244 7685 4245 7715
rect 4245 7685 4275 7715
rect 4275 7685 4276 7715
rect 4244 7684 4276 7685
rect 4244 7635 4276 7636
rect 4244 7605 4245 7635
rect 4245 7605 4275 7635
rect 4275 7605 4276 7635
rect 4244 7604 4276 7605
rect 4244 7555 4276 7556
rect 4244 7525 4245 7555
rect 4245 7525 4275 7555
rect 4275 7525 4276 7555
rect 4244 7524 4276 7525
rect 4244 7475 4276 7476
rect 4244 7445 4245 7475
rect 4245 7445 4275 7475
rect 4275 7445 4276 7475
rect 4244 7444 4276 7445
rect 4244 7395 4276 7396
rect 4244 7365 4245 7395
rect 4245 7365 4275 7395
rect 4275 7365 4276 7395
rect 4244 7364 4276 7365
rect 4244 7315 4276 7316
rect 4244 7285 4245 7315
rect 4245 7285 4275 7315
rect 4275 7285 4276 7315
rect 4244 7284 4276 7285
rect 4244 7235 4276 7236
rect 4244 7205 4245 7235
rect 4245 7205 4275 7235
rect 4275 7205 4276 7235
rect 4244 7204 4276 7205
rect 4244 7155 4276 7156
rect 4244 7125 4245 7155
rect 4245 7125 4275 7155
rect 4275 7125 4276 7155
rect 4244 7124 4276 7125
rect 4244 7075 4276 7076
rect 4244 7045 4245 7075
rect 4245 7045 4275 7075
rect 4275 7045 4276 7075
rect 4244 7044 4276 7045
rect 4244 6995 4276 6996
rect 4244 6965 4245 6995
rect 4245 6965 4275 6995
rect 4275 6965 4276 6995
rect 4244 6964 4276 6965
rect 4244 6884 4276 6916
rect 4244 6835 4276 6836
rect 4244 6805 4245 6835
rect 4245 6805 4275 6835
rect 4275 6805 4276 6835
rect 4244 6804 4276 6805
rect 4244 6755 4276 6756
rect 4244 6725 4245 6755
rect 4245 6725 4275 6755
rect 4275 6725 4276 6755
rect 4244 6724 4276 6725
rect 4244 6675 4276 6676
rect 4244 6645 4245 6675
rect 4245 6645 4275 6675
rect 4275 6645 4276 6675
rect 4244 6644 4276 6645
rect 4244 6595 4276 6596
rect 4244 6565 4245 6595
rect 4245 6565 4275 6595
rect 4275 6565 4276 6595
rect 4244 6564 4276 6565
rect 4244 6515 4276 6516
rect 4244 6485 4245 6515
rect 4245 6485 4275 6515
rect 4275 6485 4276 6515
rect 4244 6484 4276 6485
rect 4244 6435 4276 6436
rect 4244 6405 4245 6435
rect 4245 6405 4275 6435
rect 4275 6405 4276 6435
rect 4244 6404 4276 6405
rect 4244 6355 4276 6356
rect 4244 6325 4245 6355
rect 4245 6325 4275 6355
rect 4275 6325 4276 6355
rect 4244 6324 4276 6325
rect 4244 6275 4276 6276
rect 4244 6245 4245 6275
rect 4245 6245 4275 6275
rect 4275 6245 4276 6275
rect 4244 6244 4276 6245
rect 4244 6164 4276 6196
rect 4244 6084 4276 6116
rect 4244 6004 4276 6036
rect 4244 5924 4276 5956
rect 4244 5875 4276 5876
rect 4244 5845 4245 5875
rect 4245 5845 4275 5875
rect 4275 5845 4276 5875
rect 4244 5844 4276 5845
rect 4244 5795 4276 5796
rect 4244 5765 4245 5795
rect 4245 5765 4275 5795
rect 4275 5765 4276 5795
rect 4244 5764 4276 5765
rect 4244 5715 4276 5716
rect 4244 5685 4245 5715
rect 4245 5685 4275 5715
rect 4275 5685 4276 5715
rect 4244 5684 4276 5685
rect 4244 5635 4276 5636
rect 4244 5605 4245 5635
rect 4245 5605 4275 5635
rect 4275 5605 4276 5635
rect 4244 5604 4276 5605
rect 4244 5555 4276 5556
rect 4244 5525 4245 5555
rect 4245 5525 4275 5555
rect 4275 5525 4276 5555
rect 4244 5524 4276 5525
rect 4244 5475 4276 5476
rect 4244 5445 4245 5475
rect 4245 5445 4275 5475
rect 4275 5445 4276 5475
rect 4244 5444 4276 5445
rect 4244 5395 4276 5396
rect 4244 5365 4245 5395
rect 4245 5365 4275 5395
rect 4275 5365 4276 5395
rect 4244 5364 4276 5365
rect 4244 5315 4276 5316
rect 4244 5285 4245 5315
rect 4245 5285 4275 5315
rect 4275 5285 4276 5315
rect 4244 5284 4276 5285
rect 4244 5235 4276 5236
rect 4244 5205 4245 5235
rect 4245 5205 4275 5235
rect 4275 5205 4276 5235
rect 4244 5204 4276 5205
rect 4244 5155 4276 5156
rect 4244 5125 4245 5155
rect 4245 5125 4275 5155
rect 4275 5125 4276 5155
rect 4244 5124 4276 5125
rect 4244 5075 4276 5076
rect 4244 5045 4245 5075
rect 4245 5045 4275 5075
rect 4275 5045 4276 5075
rect 4244 5044 4276 5045
rect 4244 4995 4276 4996
rect 4244 4965 4245 4995
rect 4245 4965 4275 4995
rect 4275 4965 4276 4995
rect 4244 4964 4276 4965
rect 4244 4915 4276 4916
rect 4244 4885 4245 4915
rect 4245 4885 4275 4915
rect 4275 4885 4276 4915
rect 4244 4884 4276 4885
rect 4244 4804 4276 4836
rect 4244 4755 4276 4756
rect 4244 4725 4245 4755
rect 4245 4725 4275 4755
rect 4275 4725 4276 4755
rect 4244 4724 4276 4725
rect 4244 4675 4276 4676
rect 4244 4645 4245 4675
rect 4245 4645 4275 4675
rect 4275 4645 4276 4675
rect 4244 4644 4276 4645
rect 4244 4564 4276 4596
rect 4244 4515 4276 4516
rect 4244 4485 4245 4515
rect 4245 4485 4275 4515
rect 4275 4485 4276 4515
rect 4244 4484 4276 4485
rect 4244 4435 4276 4436
rect 4244 4405 4245 4435
rect 4245 4405 4275 4435
rect 4275 4405 4276 4435
rect 4244 4404 4276 4405
rect 4244 4355 4276 4356
rect 4244 4325 4245 4355
rect 4245 4325 4275 4355
rect 4275 4325 4276 4355
rect 4244 4324 4276 4325
rect 4244 4275 4276 4276
rect 4244 4245 4245 4275
rect 4245 4245 4275 4275
rect 4275 4245 4276 4275
rect 4244 4244 4276 4245
rect 4244 4195 4276 4196
rect 4244 4165 4245 4195
rect 4245 4165 4275 4195
rect 4275 4165 4276 4195
rect 4244 4164 4276 4165
rect 4244 4115 4276 4116
rect 4244 4085 4245 4115
rect 4245 4085 4275 4115
rect 4275 4085 4276 4115
rect 4244 4084 4276 4085
rect 4244 4035 4276 4036
rect 4244 4005 4245 4035
rect 4245 4005 4275 4035
rect 4275 4005 4276 4035
rect 4244 4004 4276 4005
rect 4244 3955 4276 3956
rect 4244 3925 4245 3955
rect 4245 3925 4275 3955
rect 4275 3925 4276 3955
rect 4244 3924 4276 3925
rect 4244 3875 4276 3876
rect 4244 3845 4245 3875
rect 4245 3845 4275 3875
rect 4275 3845 4276 3875
rect 4244 3844 4276 3845
rect 4244 3764 4276 3796
rect 4244 3715 4276 3716
rect 4244 3685 4245 3715
rect 4245 3685 4275 3715
rect 4275 3685 4276 3715
rect 4244 3684 4276 3685
rect 4244 3635 4276 3636
rect 4244 3605 4245 3635
rect 4245 3605 4275 3635
rect 4275 3605 4276 3635
rect 4244 3604 4276 3605
rect 4244 3524 4276 3556
rect 4244 3475 4276 3476
rect 4244 3445 4245 3475
rect 4245 3445 4275 3475
rect 4275 3445 4276 3475
rect 4244 3444 4276 3445
rect 4244 3395 4276 3396
rect 4244 3365 4245 3395
rect 4245 3365 4275 3395
rect 4275 3365 4276 3395
rect 4244 3364 4276 3365
rect 4244 3284 4276 3316
rect 4244 3235 4276 3236
rect 4244 3205 4245 3235
rect 4245 3205 4275 3235
rect 4275 3205 4276 3235
rect 4244 3204 4276 3205
rect 4244 3155 4276 3156
rect 4244 3125 4245 3155
rect 4245 3125 4275 3155
rect 4275 3125 4276 3155
rect 4244 3124 4276 3125
rect 4244 3075 4276 3076
rect 4244 3045 4245 3075
rect 4245 3045 4275 3075
rect 4275 3045 4276 3075
rect 4244 3044 4276 3045
rect 4244 2995 4276 2996
rect 4244 2965 4245 2995
rect 4245 2965 4275 2995
rect 4275 2965 4276 2995
rect 4244 2964 4276 2965
rect 4244 2915 4276 2916
rect 4244 2885 4245 2915
rect 4245 2885 4275 2915
rect 4275 2885 4276 2915
rect 4244 2884 4276 2885
rect 4244 2835 4276 2836
rect 4244 2805 4245 2835
rect 4245 2805 4275 2835
rect 4275 2805 4276 2835
rect 4244 2804 4276 2805
rect 4244 2755 4276 2756
rect 4244 2725 4245 2755
rect 4245 2725 4275 2755
rect 4275 2725 4276 2755
rect 4244 2724 4276 2725
rect 4244 2675 4276 2676
rect 4244 2645 4245 2675
rect 4245 2645 4275 2675
rect 4275 2645 4276 2675
rect 4244 2644 4276 2645
rect 4244 2595 4276 2596
rect 4244 2565 4245 2595
rect 4245 2565 4275 2595
rect 4275 2565 4276 2595
rect 4244 2564 4276 2565
rect 4244 2515 4276 2516
rect 4244 2485 4245 2515
rect 4245 2485 4275 2515
rect 4275 2485 4276 2515
rect 4244 2484 4276 2485
rect 4244 2435 4276 2436
rect 4244 2405 4245 2435
rect 4245 2405 4275 2435
rect 4275 2405 4276 2435
rect 4244 2404 4276 2405
rect 4244 2355 4276 2356
rect 4244 2325 4245 2355
rect 4245 2325 4275 2355
rect 4275 2325 4276 2355
rect 4244 2324 4276 2325
rect 4244 2275 4276 2276
rect 4244 2245 4245 2275
rect 4245 2245 4275 2275
rect 4275 2245 4276 2275
rect 4244 2244 4276 2245
rect 4244 2195 4276 2196
rect 4244 2165 4245 2195
rect 4245 2165 4275 2195
rect 4275 2165 4276 2195
rect 4244 2164 4276 2165
rect 4244 2115 4276 2116
rect 4244 2085 4245 2115
rect 4245 2085 4275 2115
rect 4275 2085 4276 2115
rect 4244 2084 4276 2085
rect 4244 2035 4276 2036
rect 4244 2005 4245 2035
rect 4245 2005 4275 2035
rect 4275 2005 4276 2035
rect 4244 2004 4276 2005
rect 4244 1955 4276 1956
rect 4244 1925 4245 1955
rect 4245 1925 4275 1955
rect 4275 1925 4276 1955
rect 4244 1924 4276 1925
rect 4244 1844 4276 1876
rect 4244 1764 4276 1796
rect 4244 1715 4276 1716
rect 4244 1685 4245 1715
rect 4245 1685 4275 1715
rect 4275 1685 4276 1715
rect 4244 1684 4276 1685
rect 4244 1635 4276 1636
rect 4244 1605 4245 1635
rect 4245 1605 4275 1635
rect 4275 1605 4276 1635
rect 4244 1604 4276 1605
rect 4244 1555 4276 1556
rect 4244 1525 4245 1555
rect 4245 1525 4275 1555
rect 4275 1525 4276 1555
rect 4244 1524 4276 1525
rect 4244 1475 4276 1476
rect 4244 1445 4245 1475
rect 4245 1445 4275 1475
rect 4275 1445 4276 1475
rect 4244 1444 4276 1445
rect 4244 1395 4276 1396
rect 4244 1365 4245 1395
rect 4245 1365 4275 1395
rect 4275 1365 4276 1395
rect 4244 1364 4276 1365
rect 4244 1315 4276 1316
rect 4244 1285 4245 1315
rect 4245 1285 4275 1315
rect 4275 1285 4276 1315
rect 4244 1284 4276 1285
rect 4244 1235 4276 1236
rect 4244 1205 4245 1235
rect 4245 1205 4275 1235
rect 4275 1205 4276 1235
rect 4244 1204 4276 1205
rect 4244 1155 4276 1156
rect 4244 1125 4245 1155
rect 4245 1125 4275 1155
rect 4275 1125 4276 1155
rect 4244 1124 4276 1125
rect 4244 1075 4276 1076
rect 4244 1045 4245 1075
rect 4245 1045 4275 1075
rect 4275 1045 4276 1075
rect 4244 1044 4276 1045
rect 4244 995 4276 996
rect 4244 965 4245 995
rect 4245 965 4275 995
rect 4275 965 4276 995
rect 4244 964 4276 965
rect 4244 884 4276 916
rect 4244 835 4276 836
rect 4244 805 4245 835
rect 4245 805 4275 835
rect 4275 805 4276 835
rect 4244 804 4276 805
rect 4244 755 4276 756
rect 4244 725 4245 755
rect 4245 725 4275 755
rect 4275 725 4276 755
rect 4244 724 4276 725
rect 4244 675 4276 676
rect 4244 645 4245 675
rect 4245 645 4275 675
rect 4275 645 4276 675
rect 4244 644 4276 645
rect 4244 595 4276 596
rect 4244 565 4245 595
rect 4245 565 4275 595
rect 4275 565 4276 595
rect 4244 564 4276 565
rect 4244 515 4276 516
rect 4244 485 4245 515
rect 4245 485 4275 515
rect 4275 485 4276 515
rect 4244 484 4276 485
rect 4244 404 4276 436
rect 4244 324 4276 356
rect 4244 275 4276 276
rect 4244 245 4245 275
rect 4245 245 4275 275
rect 4275 245 4276 275
rect 4244 244 4276 245
rect 4244 195 4276 196
rect 4244 165 4245 195
rect 4245 165 4275 195
rect 4275 165 4276 195
rect 4244 164 4276 165
rect 4244 115 4276 116
rect 4244 85 4245 115
rect 4245 85 4275 115
rect 4275 85 4276 115
rect 4244 84 4276 85
rect 4244 35 4276 36
rect 4244 5 4245 35
rect 4245 5 4275 35
rect 4275 5 4276 35
rect 4244 4 4276 5
rect 4404 15715 4436 15716
rect 4404 15685 4405 15715
rect 4405 15685 4435 15715
rect 4435 15685 4436 15715
rect 4404 15684 4436 15685
rect 4404 15635 4436 15636
rect 4404 15605 4405 15635
rect 4405 15605 4435 15635
rect 4435 15605 4436 15635
rect 4404 15604 4436 15605
rect 4404 15555 4436 15556
rect 4404 15525 4405 15555
rect 4405 15525 4435 15555
rect 4435 15525 4436 15555
rect 4404 15524 4436 15525
rect 4404 15475 4436 15476
rect 4404 15445 4405 15475
rect 4405 15445 4435 15475
rect 4435 15445 4436 15475
rect 4404 15444 4436 15445
rect 4404 15395 4436 15396
rect 4404 15365 4405 15395
rect 4405 15365 4435 15395
rect 4435 15365 4436 15395
rect 4404 15364 4436 15365
rect 4404 15315 4436 15316
rect 4404 15285 4405 15315
rect 4405 15285 4435 15315
rect 4435 15285 4436 15315
rect 4404 15284 4436 15285
rect 4404 15235 4436 15236
rect 4404 15205 4405 15235
rect 4405 15205 4435 15235
rect 4435 15205 4436 15235
rect 4404 15204 4436 15205
rect 4404 15155 4436 15156
rect 4404 15125 4405 15155
rect 4405 15125 4435 15155
rect 4435 15125 4436 15155
rect 4404 15124 4436 15125
rect 4404 15044 4436 15076
rect 4404 14995 4436 14996
rect 4404 14965 4405 14995
rect 4405 14965 4435 14995
rect 4435 14965 4436 14995
rect 4404 14964 4436 14965
rect 4404 14915 4436 14916
rect 4404 14885 4405 14915
rect 4405 14885 4435 14915
rect 4435 14885 4436 14915
rect 4404 14884 4436 14885
rect 4404 14835 4436 14836
rect 4404 14805 4405 14835
rect 4405 14805 4435 14835
rect 4435 14805 4436 14835
rect 4404 14804 4436 14805
rect 4404 14755 4436 14756
rect 4404 14725 4405 14755
rect 4405 14725 4435 14755
rect 4435 14725 4436 14755
rect 4404 14724 4436 14725
rect 4404 14675 4436 14676
rect 4404 14645 4405 14675
rect 4405 14645 4435 14675
rect 4435 14645 4436 14675
rect 4404 14644 4436 14645
rect 4404 14595 4436 14596
rect 4404 14565 4405 14595
rect 4405 14565 4435 14595
rect 4435 14565 4436 14595
rect 4404 14564 4436 14565
rect 4404 14515 4436 14516
rect 4404 14485 4405 14515
rect 4405 14485 4435 14515
rect 4435 14485 4436 14515
rect 4404 14484 4436 14485
rect 4404 14435 4436 14436
rect 4404 14405 4405 14435
rect 4405 14405 4435 14435
rect 4435 14405 4436 14435
rect 4404 14404 4436 14405
rect 4404 14324 4436 14356
rect 4404 14244 4436 14276
rect 4404 14164 4436 14196
rect 4404 14084 4436 14116
rect 4404 14035 4436 14036
rect 4404 14005 4405 14035
rect 4405 14005 4435 14035
rect 4435 14005 4436 14035
rect 4404 14004 4436 14005
rect 4404 13955 4436 13956
rect 4404 13925 4405 13955
rect 4405 13925 4435 13955
rect 4435 13925 4436 13955
rect 4404 13924 4436 13925
rect 4404 13875 4436 13876
rect 4404 13845 4405 13875
rect 4405 13845 4435 13875
rect 4435 13845 4436 13875
rect 4404 13844 4436 13845
rect 4404 13795 4436 13796
rect 4404 13765 4405 13795
rect 4405 13765 4435 13795
rect 4435 13765 4436 13795
rect 4404 13764 4436 13765
rect 4404 13715 4436 13716
rect 4404 13685 4405 13715
rect 4405 13685 4435 13715
rect 4435 13685 4436 13715
rect 4404 13684 4436 13685
rect 4404 13635 4436 13636
rect 4404 13605 4405 13635
rect 4405 13605 4435 13635
rect 4435 13605 4436 13635
rect 4404 13604 4436 13605
rect 4404 13555 4436 13556
rect 4404 13525 4405 13555
rect 4405 13525 4435 13555
rect 4435 13525 4436 13555
rect 4404 13524 4436 13525
rect 4404 13475 4436 13476
rect 4404 13445 4405 13475
rect 4405 13445 4435 13475
rect 4435 13445 4436 13475
rect 4404 13444 4436 13445
rect 4404 13364 4436 13396
rect 4404 13284 4436 13316
rect 4404 13204 4436 13236
rect 4404 13124 4436 13156
rect 4404 13075 4436 13076
rect 4404 13045 4405 13075
rect 4405 13045 4435 13075
rect 4435 13045 4436 13075
rect 4404 13044 4436 13045
rect 4404 12995 4436 12996
rect 4404 12965 4405 12995
rect 4405 12965 4435 12995
rect 4435 12965 4436 12995
rect 4404 12964 4436 12965
rect 4404 12915 4436 12916
rect 4404 12885 4405 12915
rect 4405 12885 4435 12915
rect 4435 12885 4436 12915
rect 4404 12884 4436 12885
rect 4404 12835 4436 12836
rect 4404 12805 4405 12835
rect 4405 12805 4435 12835
rect 4435 12805 4436 12835
rect 4404 12804 4436 12805
rect 4404 12755 4436 12756
rect 4404 12725 4405 12755
rect 4405 12725 4435 12755
rect 4435 12725 4436 12755
rect 4404 12724 4436 12725
rect 4404 12675 4436 12676
rect 4404 12645 4405 12675
rect 4405 12645 4435 12675
rect 4435 12645 4436 12675
rect 4404 12644 4436 12645
rect 4404 12595 4436 12596
rect 4404 12565 4405 12595
rect 4405 12565 4435 12595
rect 4435 12565 4436 12595
rect 4404 12564 4436 12565
rect 4404 12515 4436 12516
rect 4404 12485 4405 12515
rect 4405 12485 4435 12515
rect 4435 12485 4436 12515
rect 4404 12484 4436 12485
rect 4404 12404 4436 12436
rect 4404 12355 4436 12356
rect 4404 12325 4405 12355
rect 4405 12325 4435 12355
rect 4435 12325 4436 12355
rect 4404 12324 4436 12325
rect 4404 12275 4436 12276
rect 4404 12245 4405 12275
rect 4405 12245 4435 12275
rect 4435 12245 4436 12275
rect 4404 12244 4436 12245
rect 4404 12195 4436 12196
rect 4404 12165 4405 12195
rect 4405 12165 4435 12195
rect 4435 12165 4436 12195
rect 4404 12164 4436 12165
rect 4404 12115 4436 12116
rect 4404 12085 4405 12115
rect 4405 12085 4435 12115
rect 4435 12085 4436 12115
rect 4404 12084 4436 12085
rect 4404 12035 4436 12036
rect 4404 12005 4405 12035
rect 4405 12005 4435 12035
rect 4435 12005 4436 12035
rect 4404 12004 4436 12005
rect 4404 11955 4436 11956
rect 4404 11925 4405 11955
rect 4405 11925 4435 11955
rect 4435 11925 4436 11955
rect 4404 11924 4436 11925
rect 4404 11875 4436 11876
rect 4404 11845 4405 11875
rect 4405 11845 4435 11875
rect 4435 11845 4436 11875
rect 4404 11844 4436 11845
rect 4404 11795 4436 11796
rect 4404 11765 4405 11795
rect 4405 11765 4435 11795
rect 4435 11765 4436 11795
rect 4404 11764 4436 11765
rect 4404 11715 4436 11716
rect 4404 11685 4405 11715
rect 4405 11685 4435 11715
rect 4435 11685 4436 11715
rect 4404 11684 4436 11685
rect 4404 11635 4436 11636
rect 4404 11605 4405 11635
rect 4405 11605 4435 11635
rect 4435 11605 4436 11635
rect 4404 11604 4436 11605
rect 4404 11555 4436 11556
rect 4404 11525 4405 11555
rect 4405 11525 4435 11555
rect 4435 11525 4436 11555
rect 4404 11524 4436 11525
rect 4404 11475 4436 11476
rect 4404 11445 4405 11475
rect 4405 11445 4435 11475
rect 4435 11445 4436 11475
rect 4404 11444 4436 11445
rect 4404 11395 4436 11396
rect 4404 11365 4405 11395
rect 4405 11365 4435 11395
rect 4435 11365 4436 11395
rect 4404 11364 4436 11365
rect 4404 11315 4436 11316
rect 4404 11285 4405 11315
rect 4405 11285 4435 11315
rect 4435 11285 4436 11315
rect 4404 11284 4436 11285
rect 4404 11235 4436 11236
rect 4404 11205 4405 11235
rect 4405 11205 4435 11235
rect 4435 11205 4436 11235
rect 4404 11204 4436 11205
rect 4404 11155 4436 11156
rect 4404 11125 4405 11155
rect 4405 11125 4435 11155
rect 4435 11125 4436 11155
rect 4404 11124 4436 11125
rect 4404 11075 4436 11076
rect 4404 11045 4405 11075
rect 4405 11045 4435 11075
rect 4435 11045 4436 11075
rect 4404 11044 4436 11045
rect 4404 10964 4436 10996
rect 4404 10915 4436 10916
rect 4404 10885 4405 10915
rect 4405 10885 4435 10915
rect 4435 10885 4436 10915
rect 4404 10884 4436 10885
rect 4404 10835 4436 10836
rect 4404 10805 4405 10835
rect 4405 10805 4435 10835
rect 4435 10805 4436 10835
rect 4404 10804 4436 10805
rect 4404 10755 4436 10756
rect 4404 10725 4405 10755
rect 4405 10725 4435 10755
rect 4435 10725 4436 10755
rect 4404 10724 4436 10725
rect 4404 10675 4436 10676
rect 4404 10645 4405 10675
rect 4405 10645 4435 10675
rect 4435 10645 4436 10675
rect 4404 10644 4436 10645
rect 4404 10595 4436 10596
rect 4404 10565 4405 10595
rect 4405 10565 4435 10595
rect 4435 10565 4436 10595
rect 4404 10564 4436 10565
rect 4404 10515 4436 10516
rect 4404 10485 4405 10515
rect 4405 10485 4435 10515
rect 4435 10485 4436 10515
rect 4404 10484 4436 10485
rect 4404 10435 4436 10436
rect 4404 10405 4405 10435
rect 4405 10405 4435 10435
rect 4435 10405 4436 10435
rect 4404 10404 4436 10405
rect 4404 10355 4436 10356
rect 4404 10325 4405 10355
rect 4405 10325 4435 10355
rect 4435 10325 4436 10355
rect 4404 10324 4436 10325
rect 4404 10244 4436 10276
rect 4404 10164 4436 10196
rect 4404 10084 4436 10116
rect 4404 10004 4436 10036
rect 4404 9955 4436 9956
rect 4404 9925 4405 9955
rect 4405 9925 4435 9955
rect 4435 9925 4436 9955
rect 4404 9924 4436 9925
rect 4404 9875 4436 9876
rect 4404 9845 4405 9875
rect 4405 9845 4435 9875
rect 4435 9845 4436 9875
rect 4404 9844 4436 9845
rect 4404 9795 4436 9796
rect 4404 9765 4405 9795
rect 4405 9765 4435 9795
rect 4435 9765 4436 9795
rect 4404 9764 4436 9765
rect 4404 9715 4436 9716
rect 4404 9685 4405 9715
rect 4405 9685 4435 9715
rect 4435 9685 4436 9715
rect 4404 9684 4436 9685
rect 4404 9635 4436 9636
rect 4404 9605 4405 9635
rect 4405 9605 4435 9635
rect 4435 9605 4436 9635
rect 4404 9604 4436 9605
rect 4404 9555 4436 9556
rect 4404 9525 4405 9555
rect 4405 9525 4435 9555
rect 4435 9525 4436 9555
rect 4404 9524 4436 9525
rect 4404 9475 4436 9476
rect 4404 9445 4405 9475
rect 4405 9445 4435 9475
rect 4435 9445 4436 9475
rect 4404 9444 4436 9445
rect 4404 9395 4436 9396
rect 4404 9365 4405 9395
rect 4405 9365 4435 9395
rect 4435 9365 4436 9395
rect 4404 9364 4436 9365
rect 4404 9284 4436 9316
rect 4404 9204 4436 9236
rect 4404 9124 4436 9156
rect 4404 9044 4436 9076
rect 4404 8995 4436 8996
rect 4404 8965 4405 8995
rect 4405 8965 4435 8995
rect 4435 8965 4436 8995
rect 4404 8964 4436 8965
rect 4404 8915 4436 8916
rect 4404 8885 4405 8915
rect 4405 8885 4435 8915
rect 4435 8885 4436 8915
rect 4404 8884 4436 8885
rect 4404 8835 4436 8836
rect 4404 8805 4405 8835
rect 4405 8805 4435 8835
rect 4435 8805 4436 8835
rect 4404 8804 4436 8805
rect 4404 8755 4436 8756
rect 4404 8725 4405 8755
rect 4405 8725 4435 8755
rect 4435 8725 4436 8755
rect 4404 8724 4436 8725
rect 4404 8675 4436 8676
rect 4404 8645 4405 8675
rect 4405 8645 4435 8675
rect 4435 8645 4436 8675
rect 4404 8644 4436 8645
rect 4404 8595 4436 8596
rect 4404 8565 4405 8595
rect 4405 8565 4435 8595
rect 4435 8565 4436 8595
rect 4404 8564 4436 8565
rect 4404 8515 4436 8516
rect 4404 8485 4405 8515
rect 4405 8485 4435 8515
rect 4435 8485 4436 8515
rect 4404 8484 4436 8485
rect 4404 8435 4436 8436
rect 4404 8405 4405 8435
rect 4405 8405 4435 8435
rect 4435 8405 4436 8435
rect 4404 8404 4436 8405
rect 4404 8324 4436 8356
rect 4404 8275 4436 8276
rect 4404 8245 4405 8275
rect 4405 8245 4435 8275
rect 4435 8245 4436 8275
rect 4404 8244 4436 8245
rect 4404 8195 4436 8196
rect 4404 8165 4405 8195
rect 4405 8165 4435 8195
rect 4435 8165 4436 8195
rect 4404 8164 4436 8165
rect 4404 8115 4436 8116
rect 4404 8085 4405 8115
rect 4405 8085 4435 8115
rect 4435 8085 4436 8115
rect 4404 8084 4436 8085
rect 4404 8035 4436 8036
rect 4404 8005 4405 8035
rect 4405 8005 4435 8035
rect 4435 8005 4436 8035
rect 4404 8004 4436 8005
rect 4404 7955 4436 7956
rect 4404 7925 4405 7955
rect 4405 7925 4435 7955
rect 4435 7925 4436 7955
rect 4404 7924 4436 7925
rect 4404 7875 4436 7876
rect 4404 7845 4405 7875
rect 4405 7845 4435 7875
rect 4435 7845 4436 7875
rect 4404 7844 4436 7845
rect 4404 7795 4436 7796
rect 4404 7765 4405 7795
rect 4405 7765 4435 7795
rect 4435 7765 4436 7795
rect 4404 7764 4436 7765
rect 4404 7715 4436 7716
rect 4404 7685 4405 7715
rect 4405 7685 4435 7715
rect 4435 7685 4436 7715
rect 4404 7684 4436 7685
rect 4404 7635 4436 7636
rect 4404 7605 4405 7635
rect 4405 7605 4435 7635
rect 4435 7605 4436 7635
rect 4404 7604 4436 7605
rect 4404 7555 4436 7556
rect 4404 7525 4405 7555
rect 4405 7525 4435 7555
rect 4435 7525 4436 7555
rect 4404 7524 4436 7525
rect 4404 7475 4436 7476
rect 4404 7445 4405 7475
rect 4405 7445 4435 7475
rect 4435 7445 4436 7475
rect 4404 7444 4436 7445
rect 4404 7395 4436 7396
rect 4404 7365 4405 7395
rect 4405 7365 4435 7395
rect 4435 7365 4436 7395
rect 4404 7364 4436 7365
rect 4404 7315 4436 7316
rect 4404 7285 4405 7315
rect 4405 7285 4435 7315
rect 4435 7285 4436 7315
rect 4404 7284 4436 7285
rect 4404 7235 4436 7236
rect 4404 7205 4405 7235
rect 4405 7205 4435 7235
rect 4435 7205 4436 7235
rect 4404 7204 4436 7205
rect 4404 7155 4436 7156
rect 4404 7125 4405 7155
rect 4405 7125 4435 7155
rect 4435 7125 4436 7155
rect 4404 7124 4436 7125
rect 4404 7075 4436 7076
rect 4404 7045 4405 7075
rect 4405 7045 4435 7075
rect 4435 7045 4436 7075
rect 4404 7044 4436 7045
rect 4404 6995 4436 6996
rect 4404 6965 4405 6995
rect 4405 6965 4435 6995
rect 4435 6965 4436 6995
rect 4404 6964 4436 6965
rect 4404 6884 4436 6916
rect 4404 6835 4436 6836
rect 4404 6805 4405 6835
rect 4405 6805 4435 6835
rect 4435 6805 4436 6835
rect 4404 6804 4436 6805
rect 4404 6755 4436 6756
rect 4404 6725 4405 6755
rect 4405 6725 4435 6755
rect 4435 6725 4436 6755
rect 4404 6724 4436 6725
rect 4404 6675 4436 6676
rect 4404 6645 4405 6675
rect 4405 6645 4435 6675
rect 4435 6645 4436 6675
rect 4404 6644 4436 6645
rect 4404 6595 4436 6596
rect 4404 6565 4405 6595
rect 4405 6565 4435 6595
rect 4435 6565 4436 6595
rect 4404 6564 4436 6565
rect 4404 6515 4436 6516
rect 4404 6485 4405 6515
rect 4405 6485 4435 6515
rect 4435 6485 4436 6515
rect 4404 6484 4436 6485
rect 4404 6435 4436 6436
rect 4404 6405 4405 6435
rect 4405 6405 4435 6435
rect 4435 6405 4436 6435
rect 4404 6404 4436 6405
rect 4404 6355 4436 6356
rect 4404 6325 4405 6355
rect 4405 6325 4435 6355
rect 4435 6325 4436 6355
rect 4404 6324 4436 6325
rect 4404 6275 4436 6276
rect 4404 6245 4405 6275
rect 4405 6245 4435 6275
rect 4435 6245 4436 6275
rect 4404 6244 4436 6245
rect 4404 6164 4436 6196
rect 4404 6084 4436 6116
rect 4404 6004 4436 6036
rect 4404 5924 4436 5956
rect 4404 5875 4436 5876
rect 4404 5845 4405 5875
rect 4405 5845 4435 5875
rect 4435 5845 4436 5875
rect 4404 5844 4436 5845
rect 4404 5795 4436 5796
rect 4404 5765 4405 5795
rect 4405 5765 4435 5795
rect 4435 5765 4436 5795
rect 4404 5764 4436 5765
rect 4404 5715 4436 5716
rect 4404 5685 4405 5715
rect 4405 5685 4435 5715
rect 4435 5685 4436 5715
rect 4404 5684 4436 5685
rect 4404 5635 4436 5636
rect 4404 5605 4405 5635
rect 4405 5605 4435 5635
rect 4435 5605 4436 5635
rect 4404 5604 4436 5605
rect 4404 5555 4436 5556
rect 4404 5525 4405 5555
rect 4405 5525 4435 5555
rect 4435 5525 4436 5555
rect 4404 5524 4436 5525
rect 4404 5475 4436 5476
rect 4404 5445 4405 5475
rect 4405 5445 4435 5475
rect 4435 5445 4436 5475
rect 4404 5444 4436 5445
rect 4404 5395 4436 5396
rect 4404 5365 4405 5395
rect 4405 5365 4435 5395
rect 4435 5365 4436 5395
rect 4404 5364 4436 5365
rect 4404 5315 4436 5316
rect 4404 5285 4405 5315
rect 4405 5285 4435 5315
rect 4435 5285 4436 5315
rect 4404 5284 4436 5285
rect 4404 5235 4436 5236
rect 4404 5205 4405 5235
rect 4405 5205 4435 5235
rect 4435 5205 4436 5235
rect 4404 5204 4436 5205
rect 4404 5155 4436 5156
rect 4404 5125 4405 5155
rect 4405 5125 4435 5155
rect 4435 5125 4436 5155
rect 4404 5124 4436 5125
rect 4404 5075 4436 5076
rect 4404 5045 4405 5075
rect 4405 5045 4435 5075
rect 4435 5045 4436 5075
rect 4404 5044 4436 5045
rect 4404 4995 4436 4996
rect 4404 4965 4405 4995
rect 4405 4965 4435 4995
rect 4435 4965 4436 4995
rect 4404 4964 4436 4965
rect 4404 4915 4436 4916
rect 4404 4885 4405 4915
rect 4405 4885 4435 4915
rect 4435 4885 4436 4915
rect 4404 4884 4436 4885
rect 4404 4804 4436 4836
rect 4404 4755 4436 4756
rect 4404 4725 4405 4755
rect 4405 4725 4435 4755
rect 4435 4725 4436 4755
rect 4404 4724 4436 4725
rect 4404 4675 4436 4676
rect 4404 4645 4405 4675
rect 4405 4645 4435 4675
rect 4435 4645 4436 4675
rect 4404 4644 4436 4645
rect 4404 4564 4436 4596
rect 4404 4515 4436 4516
rect 4404 4485 4405 4515
rect 4405 4485 4435 4515
rect 4435 4485 4436 4515
rect 4404 4484 4436 4485
rect 4404 4435 4436 4436
rect 4404 4405 4405 4435
rect 4405 4405 4435 4435
rect 4435 4405 4436 4435
rect 4404 4404 4436 4405
rect 4404 4355 4436 4356
rect 4404 4325 4405 4355
rect 4405 4325 4435 4355
rect 4435 4325 4436 4355
rect 4404 4324 4436 4325
rect 4404 4275 4436 4276
rect 4404 4245 4405 4275
rect 4405 4245 4435 4275
rect 4435 4245 4436 4275
rect 4404 4244 4436 4245
rect 4404 4195 4436 4196
rect 4404 4165 4405 4195
rect 4405 4165 4435 4195
rect 4435 4165 4436 4195
rect 4404 4164 4436 4165
rect 4404 4115 4436 4116
rect 4404 4085 4405 4115
rect 4405 4085 4435 4115
rect 4435 4085 4436 4115
rect 4404 4084 4436 4085
rect 4404 4035 4436 4036
rect 4404 4005 4405 4035
rect 4405 4005 4435 4035
rect 4435 4005 4436 4035
rect 4404 4004 4436 4005
rect 4404 3955 4436 3956
rect 4404 3925 4405 3955
rect 4405 3925 4435 3955
rect 4435 3925 4436 3955
rect 4404 3924 4436 3925
rect 4404 3875 4436 3876
rect 4404 3845 4405 3875
rect 4405 3845 4435 3875
rect 4435 3845 4436 3875
rect 4404 3844 4436 3845
rect 4404 3764 4436 3796
rect 4404 3715 4436 3716
rect 4404 3685 4405 3715
rect 4405 3685 4435 3715
rect 4435 3685 4436 3715
rect 4404 3684 4436 3685
rect 4404 3635 4436 3636
rect 4404 3605 4405 3635
rect 4405 3605 4435 3635
rect 4435 3605 4436 3635
rect 4404 3604 4436 3605
rect 4404 3524 4436 3556
rect 4404 3475 4436 3476
rect 4404 3445 4405 3475
rect 4405 3445 4435 3475
rect 4435 3445 4436 3475
rect 4404 3444 4436 3445
rect 4404 3395 4436 3396
rect 4404 3365 4405 3395
rect 4405 3365 4435 3395
rect 4435 3365 4436 3395
rect 4404 3364 4436 3365
rect 4404 3284 4436 3316
rect 4404 3235 4436 3236
rect 4404 3205 4405 3235
rect 4405 3205 4435 3235
rect 4435 3205 4436 3235
rect 4404 3204 4436 3205
rect 4404 3155 4436 3156
rect 4404 3125 4405 3155
rect 4405 3125 4435 3155
rect 4435 3125 4436 3155
rect 4404 3124 4436 3125
rect 4404 3075 4436 3076
rect 4404 3045 4405 3075
rect 4405 3045 4435 3075
rect 4435 3045 4436 3075
rect 4404 3044 4436 3045
rect 4404 2995 4436 2996
rect 4404 2965 4405 2995
rect 4405 2965 4435 2995
rect 4435 2965 4436 2995
rect 4404 2964 4436 2965
rect 4404 2915 4436 2916
rect 4404 2885 4405 2915
rect 4405 2885 4435 2915
rect 4435 2885 4436 2915
rect 4404 2884 4436 2885
rect 4404 2835 4436 2836
rect 4404 2805 4405 2835
rect 4405 2805 4435 2835
rect 4435 2805 4436 2835
rect 4404 2804 4436 2805
rect 4404 2755 4436 2756
rect 4404 2725 4405 2755
rect 4405 2725 4435 2755
rect 4435 2725 4436 2755
rect 4404 2724 4436 2725
rect 4404 2675 4436 2676
rect 4404 2645 4405 2675
rect 4405 2645 4435 2675
rect 4435 2645 4436 2675
rect 4404 2644 4436 2645
rect 4404 2595 4436 2596
rect 4404 2565 4405 2595
rect 4405 2565 4435 2595
rect 4435 2565 4436 2595
rect 4404 2564 4436 2565
rect 4404 2515 4436 2516
rect 4404 2485 4405 2515
rect 4405 2485 4435 2515
rect 4435 2485 4436 2515
rect 4404 2484 4436 2485
rect 4404 2435 4436 2436
rect 4404 2405 4405 2435
rect 4405 2405 4435 2435
rect 4435 2405 4436 2435
rect 4404 2404 4436 2405
rect 4404 2355 4436 2356
rect 4404 2325 4405 2355
rect 4405 2325 4435 2355
rect 4435 2325 4436 2355
rect 4404 2324 4436 2325
rect 4404 2275 4436 2276
rect 4404 2245 4405 2275
rect 4405 2245 4435 2275
rect 4435 2245 4436 2275
rect 4404 2244 4436 2245
rect 4404 2195 4436 2196
rect 4404 2165 4405 2195
rect 4405 2165 4435 2195
rect 4435 2165 4436 2195
rect 4404 2164 4436 2165
rect 4404 2115 4436 2116
rect 4404 2085 4405 2115
rect 4405 2085 4435 2115
rect 4435 2085 4436 2115
rect 4404 2084 4436 2085
rect 4404 2035 4436 2036
rect 4404 2005 4405 2035
rect 4405 2005 4435 2035
rect 4435 2005 4436 2035
rect 4404 2004 4436 2005
rect 4404 1955 4436 1956
rect 4404 1925 4405 1955
rect 4405 1925 4435 1955
rect 4435 1925 4436 1955
rect 4404 1924 4436 1925
rect 4404 1844 4436 1876
rect 4404 1764 4436 1796
rect 4404 1715 4436 1716
rect 4404 1685 4405 1715
rect 4405 1685 4435 1715
rect 4435 1685 4436 1715
rect 4404 1684 4436 1685
rect 4404 1635 4436 1636
rect 4404 1605 4405 1635
rect 4405 1605 4435 1635
rect 4435 1605 4436 1635
rect 4404 1604 4436 1605
rect 4404 1555 4436 1556
rect 4404 1525 4405 1555
rect 4405 1525 4435 1555
rect 4435 1525 4436 1555
rect 4404 1524 4436 1525
rect 4404 1475 4436 1476
rect 4404 1445 4405 1475
rect 4405 1445 4435 1475
rect 4435 1445 4436 1475
rect 4404 1444 4436 1445
rect 4404 1395 4436 1396
rect 4404 1365 4405 1395
rect 4405 1365 4435 1395
rect 4435 1365 4436 1395
rect 4404 1364 4436 1365
rect 4404 1315 4436 1316
rect 4404 1285 4405 1315
rect 4405 1285 4435 1315
rect 4435 1285 4436 1315
rect 4404 1284 4436 1285
rect 4404 1235 4436 1236
rect 4404 1205 4405 1235
rect 4405 1205 4435 1235
rect 4435 1205 4436 1235
rect 4404 1204 4436 1205
rect 4404 1155 4436 1156
rect 4404 1125 4405 1155
rect 4405 1125 4435 1155
rect 4435 1125 4436 1155
rect 4404 1124 4436 1125
rect 4404 1075 4436 1076
rect 4404 1045 4405 1075
rect 4405 1045 4435 1075
rect 4435 1045 4436 1075
rect 4404 1044 4436 1045
rect 4404 995 4436 996
rect 4404 965 4405 995
rect 4405 965 4435 995
rect 4435 965 4436 995
rect 4404 964 4436 965
rect 4404 884 4436 916
rect 4404 835 4436 836
rect 4404 805 4405 835
rect 4405 805 4435 835
rect 4435 805 4436 835
rect 4404 804 4436 805
rect 4404 755 4436 756
rect 4404 725 4405 755
rect 4405 725 4435 755
rect 4435 725 4436 755
rect 4404 724 4436 725
rect 4404 675 4436 676
rect 4404 645 4405 675
rect 4405 645 4435 675
rect 4435 645 4436 675
rect 4404 644 4436 645
rect 4404 595 4436 596
rect 4404 565 4405 595
rect 4405 565 4435 595
rect 4435 565 4436 595
rect 4404 564 4436 565
rect 4404 515 4436 516
rect 4404 485 4405 515
rect 4405 485 4435 515
rect 4435 485 4436 515
rect 4404 484 4436 485
rect 4404 404 4436 436
rect 4404 324 4436 356
rect 4404 275 4436 276
rect 4404 245 4405 275
rect 4405 245 4435 275
rect 4435 245 4436 275
rect 4404 244 4436 245
rect 4404 195 4436 196
rect 4404 165 4405 195
rect 4405 165 4435 195
rect 4435 165 4436 195
rect 4404 164 4436 165
rect 4404 115 4436 116
rect 4404 85 4405 115
rect 4405 85 4435 115
rect 4435 85 4436 115
rect 4404 84 4436 85
rect 4404 35 4436 36
rect 4404 5 4405 35
rect 4405 5 4435 35
rect 4435 5 4436 35
rect 4404 4 4436 5
rect 4244 -956 4276 -764
rect 4404 -956 4436 -764
rect 4484 15715 4516 15716
rect 4484 15685 4485 15715
rect 4485 15685 4515 15715
rect 4515 15685 4516 15715
rect 4484 15684 4516 15685
rect 4484 15635 4516 15636
rect 4484 15605 4485 15635
rect 4485 15605 4515 15635
rect 4515 15605 4516 15635
rect 4484 15604 4516 15605
rect 4484 15555 4516 15556
rect 4484 15525 4485 15555
rect 4485 15525 4515 15555
rect 4515 15525 4516 15555
rect 4484 15524 4516 15525
rect 4484 15475 4516 15476
rect 4484 15445 4485 15475
rect 4485 15445 4515 15475
rect 4515 15445 4516 15475
rect 4484 15444 4516 15445
rect 4484 15395 4516 15396
rect 4484 15365 4485 15395
rect 4485 15365 4515 15395
rect 4515 15365 4516 15395
rect 4484 15364 4516 15365
rect 4484 15315 4516 15316
rect 4484 15285 4485 15315
rect 4485 15285 4515 15315
rect 4515 15285 4516 15315
rect 4484 15284 4516 15285
rect 4484 15235 4516 15236
rect 4484 15205 4485 15235
rect 4485 15205 4515 15235
rect 4515 15205 4516 15235
rect 4484 15204 4516 15205
rect 4484 15155 4516 15156
rect 4484 15125 4485 15155
rect 4485 15125 4515 15155
rect 4515 15125 4516 15155
rect 4484 15124 4516 15125
rect 4484 15044 4516 15076
rect 4484 14995 4516 14996
rect 4484 14965 4485 14995
rect 4485 14965 4515 14995
rect 4515 14965 4516 14995
rect 4484 14964 4516 14965
rect 4484 14915 4516 14916
rect 4484 14885 4485 14915
rect 4485 14885 4515 14915
rect 4515 14885 4516 14915
rect 4484 14884 4516 14885
rect 4484 14835 4516 14836
rect 4484 14805 4485 14835
rect 4485 14805 4515 14835
rect 4515 14805 4516 14835
rect 4484 14804 4516 14805
rect 4484 14755 4516 14756
rect 4484 14725 4485 14755
rect 4485 14725 4515 14755
rect 4515 14725 4516 14755
rect 4484 14724 4516 14725
rect 4484 14675 4516 14676
rect 4484 14645 4485 14675
rect 4485 14645 4515 14675
rect 4515 14645 4516 14675
rect 4484 14644 4516 14645
rect 4484 14595 4516 14596
rect 4484 14565 4485 14595
rect 4485 14565 4515 14595
rect 4515 14565 4516 14595
rect 4484 14564 4516 14565
rect 4484 14515 4516 14516
rect 4484 14485 4485 14515
rect 4485 14485 4515 14515
rect 4515 14485 4516 14515
rect 4484 14484 4516 14485
rect 4484 14435 4516 14436
rect 4484 14405 4485 14435
rect 4485 14405 4515 14435
rect 4515 14405 4516 14435
rect 4484 14404 4516 14405
rect 4484 14324 4516 14356
rect 4484 14244 4516 14276
rect 4484 14164 4516 14196
rect 4484 14084 4516 14116
rect 4484 14035 4516 14036
rect 4484 14005 4485 14035
rect 4485 14005 4515 14035
rect 4515 14005 4516 14035
rect 4484 14004 4516 14005
rect 4484 13955 4516 13956
rect 4484 13925 4485 13955
rect 4485 13925 4515 13955
rect 4515 13925 4516 13955
rect 4484 13924 4516 13925
rect 4484 13875 4516 13876
rect 4484 13845 4485 13875
rect 4485 13845 4515 13875
rect 4515 13845 4516 13875
rect 4484 13844 4516 13845
rect 4484 13795 4516 13796
rect 4484 13765 4485 13795
rect 4485 13765 4515 13795
rect 4515 13765 4516 13795
rect 4484 13764 4516 13765
rect 4484 13715 4516 13716
rect 4484 13685 4485 13715
rect 4485 13685 4515 13715
rect 4515 13685 4516 13715
rect 4484 13684 4516 13685
rect 4484 13635 4516 13636
rect 4484 13605 4485 13635
rect 4485 13605 4515 13635
rect 4515 13605 4516 13635
rect 4484 13604 4516 13605
rect 4484 13555 4516 13556
rect 4484 13525 4485 13555
rect 4485 13525 4515 13555
rect 4515 13525 4516 13555
rect 4484 13524 4516 13525
rect 4484 13475 4516 13476
rect 4484 13445 4485 13475
rect 4485 13445 4515 13475
rect 4515 13445 4516 13475
rect 4484 13444 4516 13445
rect 4484 13364 4516 13396
rect 4484 13284 4516 13316
rect 4484 13204 4516 13236
rect 4484 13124 4516 13156
rect 4484 13075 4516 13076
rect 4484 13045 4485 13075
rect 4485 13045 4515 13075
rect 4515 13045 4516 13075
rect 4484 13044 4516 13045
rect 4484 12995 4516 12996
rect 4484 12965 4485 12995
rect 4485 12965 4515 12995
rect 4515 12965 4516 12995
rect 4484 12964 4516 12965
rect 4484 12915 4516 12916
rect 4484 12885 4485 12915
rect 4485 12885 4515 12915
rect 4515 12885 4516 12915
rect 4484 12884 4516 12885
rect 4484 12835 4516 12836
rect 4484 12805 4485 12835
rect 4485 12805 4515 12835
rect 4515 12805 4516 12835
rect 4484 12804 4516 12805
rect 4484 12755 4516 12756
rect 4484 12725 4485 12755
rect 4485 12725 4515 12755
rect 4515 12725 4516 12755
rect 4484 12724 4516 12725
rect 4484 12675 4516 12676
rect 4484 12645 4485 12675
rect 4485 12645 4515 12675
rect 4515 12645 4516 12675
rect 4484 12644 4516 12645
rect 4484 12595 4516 12596
rect 4484 12565 4485 12595
rect 4485 12565 4515 12595
rect 4515 12565 4516 12595
rect 4484 12564 4516 12565
rect 4484 12515 4516 12516
rect 4484 12485 4485 12515
rect 4485 12485 4515 12515
rect 4515 12485 4516 12515
rect 4484 12484 4516 12485
rect 4484 12404 4516 12436
rect 4484 12355 4516 12356
rect 4484 12325 4485 12355
rect 4485 12325 4515 12355
rect 4515 12325 4516 12355
rect 4484 12324 4516 12325
rect 4484 12275 4516 12276
rect 4484 12245 4485 12275
rect 4485 12245 4515 12275
rect 4515 12245 4516 12275
rect 4484 12244 4516 12245
rect 4484 12195 4516 12196
rect 4484 12165 4485 12195
rect 4485 12165 4515 12195
rect 4515 12165 4516 12195
rect 4484 12164 4516 12165
rect 4484 12115 4516 12116
rect 4484 12085 4485 12115
rect 4485 12085 4515 12115
rect 4515 12085 4516 12115
rect 4484 12084 4516 12085
rect 4484 12035 4516 12036
rect 4484 12005 4485 12035
rect 4485 12005 4515 12035
rect 4515 12005 4516 12035
rect 4484 12004 4516 12005
rect 4484 11955 4516 11956
rect 4484 11925 4485 11955
rect 4485 11925 4515 11955
rect 4515 11925 4516 11955
rect 4484 11924 4516 11925
rect 4484 11875 4516 11876
rect 4484 11845 4485 11875
rect 4485 11845 4515 11875
rect 4515 11845 4516 11875
rect 4484 11844 4516 11845
rect 4484 11795 4516 11796
rect 4484 11765 4485 11795
rect 4485 11765 4515 11795
rect 4515 11765 4516 11795
rect 4484 11764 4516 11765
rect 4484 11715 4516 11716
rect 4484 11685 4485 11715
rect 4485 11685 4515 11715
rect 4515 11685 4516 11715
rect 4484 11684 4516 11685
rect 4484 11635 4516 11636
rect 4484 11605 4485 11635
rect 4485 11605 4515 11635
rect 4515 11605 4516 11635
rect 4484 11604 4516 11605
rect 4484 11555 4516 11556
rect 4484 11525 4485 11555
rect 4485 11525 4515 11555
rect 4515 11525 4516 11555
rect 4484 11524 4516 11525
rect 4484 11475 4516 11476
rect 4484 11445 4485 11475
rect 4485 11445 4515 11475
rect 4515 11445 4516 11475
rect 4484 11444 4516 11445
rect 4484 11395 4516 11396
rect 4484 11365 4485 11395
rect 4485 11365 4515 11395
rect 4515 11365 4516 11395
rect 4484 11364 4516 11365
rect 4484 11315 4516 11316
rect 4484 11285 4485 11315
rect 4485 11285 4515 11315
rect 4515 11285 4516 11315
rect 4484 11284 4516 11285
rect 4484 11235 4516 11236
rect 4484 11205 4485 11235
rect 4485 11205 4515 11235
rect 4515 11205 4516 11235
rect 4484 11204 4516 11205
rect 4484 11155 4516 11156
rect 4484 11125 4485 11155
rect 4485 11125 4515 11155
rect 4515 11125 4516 11155
rect 4484 11124 4516 11125
rect 4484 11075 4516 11076
rect 4484 11045 4485 11075
rect 4485 11045 4515 11075
rect 4515 11045 4516 11075
rect 4484 11044 4516 11045
rect 4484 10964 4516 10996
rect 4484 10915 4516 10916
rect 4484 10885 4485 10915
rect 4485 10885 4515 10915
rect 4515 10885 4516 10915
rect 4484 10884 4516 10885
rect 4484 10835 4516 10836
rect 4484 10805 4485 10835
rect 4485 10805 4515 10835
rect 4515 10805 4516 10835
rect 4484 10804 4516 10805
rect 4484 10755 4516 10756
rect 4484 10725 4485 10755
rect 4485 10725 4515 10755
rect 4515 10725 4516 10755
rect 4484 10724 4516 10725
rect 4484 10675 4516 10676
rect 4484 10645 4485 10675
rect 4485 10645 4515 10675
rect 4515 10645 4516 10675
rect 4484 10644 4516 10645
rect 4484 10595 4516 10596
rect 4484 10565 4485 10595
rect 4485 10565 4515 10595
rect 4515 10565 4516 10595
rect 4484 10564 4516 10565
rect 4484 10515 4516 10516
rect 4484 10485 4485 10515
rect 4485 10485 4515 10515
rect 4515 10485 4516 10515
rect 4484 10484 4516 10485
rect 4484 10435 4516 10436
rect 4484 10405 4485 10435
rect 4485 10405 4515 10435
rect 4515 10405 4516 10435
rect 4484 10404 4516 10405
rect 4484 10355 4516 10356
rect 4484 10325 4485 10355
rect 4485 10325 4515 10355
rect 4515 10325 4516 10355
rect 4484 10324 4516 10325
rect 4484 10244 4516 10276
rect 4484 10164 4516 10196
rect 4484 10084 4516 10116
rect 4484 10004 4516 10036
rect 4484 9955 4516 9956
rect 4484 9925 4485 9955
rect 4485 9925 4515 9955
rect 4515 9925 4516 9955
rect 4484 9924 4516 9925
rect 4484 9875 4516 9876
rect 4484 9845 4485 9875
rect 4485 9845 4515 9875
rect 4515 9845 4516 9875
rect 4484 9844 4516 9845
rect 4484 9795 4516 9796
rect 4484 9765 4485 9795
rect 4485 9765 4515 9795
rect 4515 9765 4516 9795
rect 4484 9764 4516 9765
rect 4484 9715 4516 9716
rect 4484 9685 4485 9715
rect 4485 9685 4515 9715
rect 4515 9685 4516 9715
rect 4484 9684 4516 9685
rect 4484 9635 4516 9636
rect 4484 9605 4485 9635
rect 4485 9605 4515 9635
rect 4515 9605 4516 9635
rect 4484 9604 4516 9605
rect 4484 9555 4516 9556
rect 4484 9525 4485 9555
rect 4485 9525 4515 9555
rect 4515 9525 4516 9555
rect 4484 9524 4516 9525
rect 4484 9475 4516 9476
rect 4484 9445 4485 9475
rect 4485 9445 4515 9475
rect 4515 9445 4516 9475
rect 4484 9444 4516 9445
rect 4484 9395 4516 9396
rect 4484 9365 4485 9395
rect 4485 9365 4515 9395
rect 4515 9365 4516 9395
rect 4484 9364 4516 9365
rect 4484 9284 4516 9316
rect 4484 9204 4516 9236
rect 4484 9124 4516 9156
rect 4484 9044 4516 9076
rect 4484 8995 4516 8996
rect 4484 8965 4485 8995
rect 4485 8965 4515 8995
rect 4515 8965 4516 8995
rect 4484 8964 4516 8965
rect 4484 8915 4516 8916
rect 4484 8885 4485 8915
rect 4485 8885 4515 8915
rect 4515 8885 4516 8915
rect 4484 8884 4516 8885
rect 4484 8835 4516 8836
rect 4484 8805 4485 8835
rect 4485 8805 4515 8835
rect 4515 8805 4516 8835
rect 4484 8804 4516 8805
rect 4484 8755 4516 8756
rect 4484 8725 4485 8755
rect 4485 8725 4515 8755
rect 4515 8725 4516 8755
rect 4484 8724 4516 8725
rect 4484 8675 4516 8676
rect 4484 8645 4485 8675
rect 4485 8645 4515 8675
rect 4515 8645 4516 8675
rect 4484 8644 4516 8645
rect 4484 8595 4516 8596
rect 4484 8565 4485 8595
rect 4485 8565 4515 8595
rect 4515 8565 4516 8595
rect 4484 8564 4516 8565
rect 4484 8515 4516 8516
rect 4484 8485 4485 8515
rect 4485 8485 4515 8515
rect 4515 8485 4516 8515
rect 4484 8484 4516 8485
rect 4484 8435 4516 8436
rect 4484 8405 4485 8435
rect 4485 8405 4515 8435
rect 4515 8405 4516 8435
rect 4484 8404 4516 8405
rect 4484 8324 4516 8356
rect 4484 8275 4516 8276
rect 4484 8245 4485 8275
rect 4485 8245 4515 8275
rect 4515 8245 4516 8275
rect 4484 8244 4516 8245
rect 4484 8195 4516 8196
rect 4484 8165 4485 8195
rect 4485 8165 4515 8195
rect 4515 8165 4516 8195
rect 4484 8164 4516 8165
rect 4484 8115 4516 8116
rect 4484 8085 4485 8115
rect 4485 8085 4515 8115
rect 4515 8085 4516 8115
rect 4484 8084 4516 8085
rect 4484 8035 4516 8036
rect 4484 8005 4485 8035
rect 4485 8005 4515 8035
rect 4515 8005 4516 8035
rect 4484 8004 4516 8005
rect 4484 7955 4516 7956
rect 4484 7925 4485 7955
rect 4485 7925 4515 7955
rect 4515 7925 4516 7955
rect 4484 7924 4516 7925
rect 4484 7875 4516 7876
rect 4484 7845 4485 7875
rect 4485 7845 4515 7875
rect 4515 7845 4516 7875
rect 4484 7844 4516 7845
rect 4484 7795 4516 7796
rect 4484 7765 4485 7795
rect 4485 7765 4515 7795
rect 4515 7765 4516 7795
rect 4484 7764 4516 7765
rect 4484 7715 4516 7716
rect 4484 7685 4485 7715
rect 4485 7685 4515 7715
rect 4515 7685 4516 7715
rect 4484 7684 4516 7685
rect 4484 7635 4516 7636
rect 4484 7605 4485 7635
rect 4485 7605 4515 7635
rect 4515 7605 4516 7635
rect 4484 7604 4516 7605
rect 4484 7555 4516 7556
rect 4484 7525 4485 7555
rect 4485 7525 4515 7555
rect 4515 7525 4516 7555
rect 4484 7524 4516 7525
rect 4484 7475 4516 7476
rect 4484 7445 4485 7475
rect 4485 7445 4515 7475
rect 4515 7445 4516 7475
rect 4484 7444 4516 7445
rect 4484 7395 4516 7396
rect 4484 7365 4485 7395
rect 4485 7365 4515 7395
rect 4515 7365 4516 7395
rect 4484 7364 4516 7365
rect 4484 7315 4516 7316
rect 4484 7285 4485 7315
rect 4485 7285 4515 7315
rect 4515 7285 4516 7315
rect 4484 7284 4516 7285
rect 4484 7235 4516 7236
rect 4484 7205 4485 7235
rect 4485 7205 4515 7235
rect 4515 7205 4516 7235
rect 4484 7204 4516 7205
rect 4484 7155 4516 7156
rect 4484 7125 4485 7155
rect 4485 7125 4515 7155
rect 4515 7125 4516 7155
rect 4484 7124 4516 7125
rect 4484 7075 4516 7076
rect 4484 7045 4485 7075
rect 4485 7045 4515 7075
rect 4515 7045 4516 7075
rect 4484 7044 4516 7045
rect 4484 6995 4516 6996
rect 4484 6965 4485 6995
rect 4485 6965 4515 6995
rect 4515 6965 4516 6995
rect 4484 6964 4516 6965
rect 4484 6884 4516 6916
rect 4484 6835 4516 6836
rect 4484 6805 4485 6835
rect 4485 6805 4515 6835
rect 4515 6805 4516 6835
rect 4484 6804 4516 6805
rect 4484 6755 4516 6756
rect 4484 6725 4485 6755
rect 4485 6725 4515 6755
rect 4515 6725 4516 6755
rect 4484 6724 4516 6725
rect 4484 6675 4516 6676
rect 4484 6645 4485 6675
rect 4485 6645 4515 6675
rect 4515 6645 4516 6675
rect 4484 6644 4516 6645
rect 4484 6595 4516 6596
rect 4484 6565 4485 6595
rect 4485 6565 4515 6595
rect 4515 6565 4516 6595
rect 4484 6564 4516 6565
rect 4484 6515 4516 6516
rect 4484 6485 4485 6515
rect 4485 6485 4515 6515
rect 4515 6485 4516 6515
rect 4484 6484 4516 6485
rect 4484 6435 4516 6436
rect 4484 6405 4485 6435
rect 4485 6405 4515 6435
rect 4515 6405 4516 6435
rect 4484 6404 4516 6405
rect 4484 6355 4516 6356
rect 4484 6325 4485 6355
rect 4485 6325 4515 6355
rect 4515 6325 4516 6355
rect 4484 6324 4516 6325
rect 4484 6275 4516 6276
rect 4484 6245 4485 6275
rect 4485 6245 4515 6275
rect 4515 6245 4516 6275
rect 4484 6244 4516 6245
rect 4484 6164 4516 6196
rect 4484 6084 4516 6116
rect 4484 6004 4516 6036
rect 4484 5924 4516 5956
rect 4484 5875 4516 5876
rect 4484 5845 4485 5875
rect 4485 5845 4515 5875
rect 4515 5845 4516 5875
rect 4484 5844 4516 5845
rect 4484 5795 4516 5796
rect 4484 5765 4485 5795
rect 4485 5765 4515 5795
rect 4515 5765 4516 5795
rect 4484 5764 4516 5765
rect 4484 5715 4516 5716
rect 4484 5685 4485 5715
rect 4485 5685 4515 5715
rect 4515 5685 4516 5715
rect 4484 5684 4516 5685
rect 4484 5635 4516 5636
rect 4484 5605 4485 5635
rect 4485 5605 4515 5635
rect 4515 5605 4516 5635
rect 4484 5604 4516 5605
rect 4484 5555 4516 5556
rect 4484 5525 4485 5555
rect 4485 5525 4515 5555
rect 4515 5525 4516 5555
rect 4484 5524 4516 5525
rect 4484 5475 4516 5476
rect 4484 5445 4485 5475
rect 4485 5445 4515 5475
rect 4515 5445 4516 5475
rect 4484 5444 4516 5445
rect 4484 5395 4516 5396
rect 4484 5365 4485 5395
rect 4485 5365 4515 5395
rect 4515 5365 4516 5395
rect 4484 5364 4516 5365
rect 4484 5315 4516 5316
rect 4484 5285 4485 5315
rect 4485 5285 4515 5315
rect 4515 5285 4516 5315
rect 4484 5284 4516 5285
rect 4484 5235 4516 5236
rect 4484 5205 4485 5235
rect 4485 5205 4515 5235
rect 4515 5205 4516 5235
rect 4484 5204 4516 5205
rect 4484 5155 4516 5156
rect 4484 5125 4485 5155
rect 4485 5125 4515 5155
rect 4515 5125 4516 5155
rect 4484 5124 4516 5125
rect 4484 5075 4516 5076
rect 4484 5045 4485 5075
rect 4485 5045 4515 5075
rect 4515 5045 4516 5075
rect 4484 5044 4516 5045
rect 4484 4995 4516 4996
rect 4484 4965 4485 4995
rect 4485 4965 4515 4995
rect 4515 4965 4516 4995
rect 4484 4964 4516 4965
rect 4484 4915 4516 4916
rect 4484 4885 4485 4915
rect 4485 4885 4515 4915
rect 4515 4885 4516 4915
rect 4484 4884 4516 4885
rect 4484 4804 4516 4836
rect 4484 4755 4516 4756
rect 4484 4725 4485 4755
rect 4485 4725 4515 4755
rect 4515 4725 4516 4755
rect 4484 4724 4516 4725
rect 4484 4675 4516 4676
rect 4484 4645 4485 4675
rect 4485 4645 4515 4675
rect 4515 4645 4516 4675
rect 4484 4644 4516 4645
rect 4484 4564 4516 4596
rect 4484 4515 4516 4516
rect 4484 4485 4485 4515
rect 4485 4485 4515 4515
rect 4515 4485 4516 4515
rect 4484 4484 4516 4485
rect 4484 4435 4516 4436
rect 4484 4405 4485 4435
rect 4485 4405 4515 4435
rect 4515 4405 4516 4435
rect 4484 4404 4516 4405
rect 4484 4355 4516 4356
rect 4484 4325 4485 4355
rect 4485 4325 4515 4355
rect 4515 4325 4516 4355
rect 4484 4324 4516 4325
rect 4484 4275 4516 4276
rect 4484 4245 4485 4275
rect 4485 4245 4515 4275
rect 4515 4245 4516 4275
rect 4484 4244 4516 4245
rect 4484 4195 4516 4196
rect 4484 4165 4485 4195
rect 4485 4165 4515 4195
rect 4515 4165 4516 4195
rect 4484 4164 4516 4165
rect 4484 4115 4516 4116
rect 4484 4085 4485 4115
rect 4485 4085 4515 4115
rect 4515 4085 4516 4115
rect 4484 4084 4516 4085
rect 4484 4035 4516 4036
rect 4484 4005 4485 4035
rect 4485 4005 4515 4035
rect 4515 4005 4516 4035
rect 4484 4004 4516 4005
rect 4484 3955 4516 3956
rect 4484 3925 4485 3955
rect 4485 3925 4515 3955
rect 4515 3925 4516 3955
rect 4484 3924 4516 3925
rect 4484 3875 4516 3876
rect 4484 3845 4485 3875
rect 4485 3845 4515 3875
rect 4515 3845 4516 3875
rect 4484 3844 4516 3845
rect 4484 3764 4516 3796
rect 4484 3715 4516 3716
rect 4484 3685 4485 3715
rect 4485 3685 4515 3715
rect 4515 3685 4516 3715
rect 4484 3684 4516 3685
rect 4484 3635 4516 3636
rect 4484 3605 4485 3635
rect 4485 3605 4515 3635
rect 4515 3605 4516 3635
rect 4484 3604 4516 3605
rect 4484 3524 4516 3556
rect 4484 3475 4516 3476
rect 4484 3445 4485 3475
rect 4485 3445 4515 3475
rect 4515 3445 4516 3475
rect 4484 3444 4516 3445
rect 4484 3395 4516 3396
rect 4484 3365 4485 3395
rect 4485 3365 4515 3395
rect 4515 3365 4516 3395
rect 4484 3364 4516 3365
rect 4484 3284 4516 3316
rect 4484 3235 4516 3236
rect 4484 3205 4485 3235
rect 4485 3205 4515 3235
rect 4515 3205 4516 3235
rect 4484 3204 4516 3205
rect 4484 3155 4516 3156
rect 4484 3125 4485 3155
rect 4485 3125 4515 3155
rect 4515 3125 4516 3155
rect 4484 3124 4516 3125
rect 4484 3075 4516 3076
rect 4484 3045 4485 3075
rect 4485 3045 4515 3075
rect 4515 3045 4516 3075
rect 4484 3044 4516 3045
rect 4484 2995 4516 2996
rect 4484 2965 4485 2995
rect 4485 2965 4515 2995
rect 4515 2965 4516 2995
rect 4484 2964 4516 2965
rect 4484 2915 4516 2916
rect 4484 2885 4485 2915
rect 4485 2885 4515 2915
rect 4515 2885 4516 2915
rect 4484 2884 4516 2885
rect 4484 2835 4516 2836
rect 4484 2805 4485 2835
rect 4485 2805 4515 2835
rect 4515 2805 4516 2835
rect 4484 2804 4516 2805
rect 4484 2755 4516 2756
rect 4484 2725 4485 2755
rect 4485 2725 4515 2755
rect 4515 2725 4516 2755
rect 4484 2724 4516 2725
rect 4484 2675 4516 2676
rect 4484 2645 4485 2675
rect 4485 2645 4515 2675
rect 4515 2645 4516 2675
rect 4484 2644 4516 2645
rect 4484 2595 4516 2596
rect 4484 2565 4485 2595
rect 4485 2565 4515 2595
rect 4515 2565 4516 2595
rect 4484 2564 4516 2565
rect 4484 2515 4516 2516
rect 4484 2485 4485 2515
rect 4485 2485 4515 2515
rect 4515 2485 4516 2515
rect 4484 2484 4516 2485
rect 4484 2435 4516 2436
rect 4484 2405 4485 2435
rect 4485 2405 4515 2435
rect 4515 2405 4516 2435
rect 4484 2404 4516 2405
rect 4484 2355 4516 2356
rect 4484 2325 4485 2355
rect 4485 2325 4515 2355
rect 4515 2325 4516 2355
rect 4484 2324 4516 2325
rect 4484 2275 4516 2276
rect 4484 2245 4485 2275
rect 4485 2245 4515 2275
rect 4515 2245 4516 2275
rect 4484 2244 4516 2245
rect 4484 2195 4516 2196
rect 4484 2165 4485 2195
rect 4485 2165 4515 2195
rect 4515 2165 4516 2195
rect 4484 2164 4516 2165
rect 4484 2115 4516 2116
rect 4484 2085 4485 2115
rect 4485 2085 4515 2115
rect 4515 2085 4516 2115
rect 4484 2084 4516 2085
rect 4484 2035 4516 2036
rect 4484 2005 4485 2035
rect 4485 2005 4515 2035
rect 4515 2005 4516 2035
rect 4484 2004 4516 2005
rect 4484 1955 4516 1956
rect 4484 1925 4485 1955
rect 4485 1925 4515 1955
rect 4515 1925 4516 1955
rect 4484 1924 4516 1925
rect 4484 1844 4516 1876
rect 4484 1764 4516 1796
rect 4484 1715 4516 1716
rect 4484 1685 4485 1715
rect 4485 1685 4515 1715
rect 4515 1685 4516 1715
rect 4484 1684 4516 1685
rect 4484 1635 4516 1636
rect 4484 1605 4485 1635
rect 4485 1605 4515 1635
rect 4515 1605 4516 1635
rect 4484 1604 4516 1605
rect 4484 1555 4516 1556
rect 4484 1525 4485 1555
rect 4485 1525 4515 1555
rect 4515 1525 4516 1555
rect 4484 1524 4516 1525
rect 4484 1475 4516 1476
rect 4484 1445 4485 1475
rect 4485 1445 4515 1475
rect 4515 1445 4516 1475
rect 4484 1444 4516 1445
rect 4484 1395 4516 1396
rect 4484 1365 4485 1395
rect 4485 1365 4515 1395
rect 4515 1365 4516 1395
rect 4484 1364 4516 1365
rect 4484 1315 4516 1316
rect 4484 1285 4485 1315
rect 4485 1285 4515 1315
rect 4515 1285 4516 1315
rect 4484 1284 4516 1285
rect 4484 1235 4516 1236
rect 4484 1205 4485 1235
rect 4485 1205 4515 1235
rect 4515 1205 4516 1235
rect 4484 1204 4516 1205
rect 4484 1155 4516 1156
rect 4484 1125 4485 1155
rect 4485 1125 4515 1155
rect 4515 1125 4516 1155
rect 4484 1124 4516 1125
rect 4484 1075 4516 1076
rect 4484 1045 4485 1075
rect 4485 1045 4515 1075
rect 4515 1045 4516 1075
rect 4484 1044 4516 1045
rect 4484 995 4516 996
rect 4484 965 4485 995
rect 4485 965 4515 995
rect 4515 965 4516 995
rect 4484 964 4516 965
rect 4484 884 4516 916
rect 4484 835 4516 836
rect 4484 805 4485 835
rect 4485 805 4515 835
rect 4515 805 4516 835
rect 4484 804 4516 805
rect 4484 755 4516 756
rect 4484 725 4485 755
rect 4485 725 4515 755
rect 4515 725 4516 755
rect 4484 724 4516 725
rect 4484 675 4516 676
rect 4484 645 4485 675
rect 4485 645 4515 675
rect 4515 645 4516 675
rect 4484 644 4516 645
rect 4484 595 4516 596
rect 4484 565 4485 595
rect 4485 565 4515 595
rect 4515 565 4516 595
rect 4484 564 4516 565
rect 4484 515 4516 516
rect 4484 485 4485 515
rect 4485 485 4515 515
rect 4515 485 4516 515
rect 4484 484 4516 485
rect 4484 404 4516 436
rect 4484 324 4516 356
rect 4484 275 4516 276
rect 4484 245 4485 275
rect 4485 245 4515 275
rect 4515 245 4516 275
rect 4484 244 4516 245
rect 4484 195 4516 196
rect 4484 165 4485 195
rect 4485 165 4515 195
rect 4515 165 4516 195
rect 4484 164 4516 165
rect 4484 115 4516 116
rect 4484 85 4485 115
rect 4485 85 4515 115
rect 4515 85 4516 115
rect 4484 84 4516 85
rect 4484 35 4516 36
rect 4484 5 4485 35
rect 4485 5 4515 35
rect 4515 5 4516 35
rect 4484 4 4516 5
rect 4484 -476 4516 -284
rect 124 -1036 156 -1004
rect 4484 -1036 4516 -1004
rect 4644 15715 4676 15716
rect 4644 15685 4645 15715
rect 4645 15685 4675 15715
rect 4675 15685 4676 15715
rect 4644 15684 4676 15685
rect 4644 15635 4676 15636
rect 4644 15605 4645 15635
rect 4645 15605 4675 15635
rect 4675 15605 4676 15635
rect 4644 15604 4676 15605
rect 4644 15555 4676 15556
rect 4644 15525 4645 15555
rect 4645 15525 4675 15555
rect 4675 15525 4676 15555
rect 4644 15524 4676 15525
rect 4644 15475 4676 15476
rect 4644 15445 4645 15475
rect 4645 15445 4675 15475
rect 4675 15445 4676 15475
rect 4644 15444 4676 15445
rect 4644 15395 4676 15396
rect 4644 15365 4645 15395
rect 4645 15365 4675 15395
rect 4675 15365 4676 15395
rect 4644 15364 4676 15365
rect 4644 15315 4676 15316
rect 4644 15285 4645 15315
rect 4645 15285 4675 15315
rect 4675 15285 4676 15315
rect 4644 15284 4676 15285
rect 4644 15235 4676 15236
rect 4644 15205 4645 15235
rect 4645 15205 4675 15235
rect 4675 15205 4676 15235
rect 4644 15204 4676 15205
rect 4644 15155 4676 15156
rect 4644 15125 4645 15155
rect 4645 15125 4675 15155
rect 4675 15125 4676 15155
rect 4644 15124 4676 15125
rect 4644 15044 4676 15076
rect 4644 14995 4676 14996
rect 4644 14965 4645 14995
rect 4645 14965 4675 14995
rect 4675 14965 4676 14995
rect 4644 14964 4676 14965
rect 4644 14915 4676 14916
rect 4644 14885 4645 14915
rect 4645 14885 4675 14915
rect 4675 14885 4676 14915
rect 4644 14884 4676 14885
rect 4644 14835 4676 14836
rect 4644 14805 4645 14835
rect 4645 14805 4675 14835
rect 4675 14805 4676 14835
rect 4644 14804 4676 14805
rect 4644 14755 4676 14756
rect 4644 14725 4645 14755
rect 4645 14725 4675 14755
rect 4675 14725 4676 14755
rect 4644 14724 4676 14725
rect 4644 14675 4676 14676
rect 4644 14645 4645 14675
rect 4645 14645 4675 14675
rect 4675 14645 4676 14675
rect 4644 14644 4676 14645
rect 4644 14595 4676 14596
rect 4644 14565 4645 14595
rect 4645 14565 4675 14595
rect 4675 14565 4676 14595
rect 4644 14564 4676 14565
rect 4644 14515 4676 14516
rect 4644 14485 4645 14515
rect 4645 14485 4675 14515
rect 4675 14485 4676 14515
rect 4644 14484 4676 14485
rect 4644 14435 4676 14436
rect 4644 14405 4645 14435
rect 4645 14405 4675 14435
rect 4675 14405 4676 14435
rect 4644 14404 4676 14405
rect 4644 14324 4676 14356
rect 4644 14244 4676 14276
rect 4644 14164 4676 14196
rect 4644 14084 4676 14116
rect 4644 14035 4676 14036
rect 4644 14005 4645 14035
rect 4645 14005 4675 14035
rect 4675 14005 4676 14035
rect 4644 14004 4676 14005
rect 4644 13955 4676 13956
rect 4644 13925 4645 13955
rect 4645 13925 4675 13955
rect 4675 13925 4676 13955
rect 4644 13924 4676 13925
rect 4644 13875 4676 13876
rect 4644 13845 4645 13875
rect 4645 13845 4675 13875
rect 4675 13845 4676 13875
rect 4644 13844 4676 13845
rect 4644 13795 4676 13796
rect 4644 13765 4645 13795
rect 4645 13765 4675 13795
rect 4675 13765 4676 13795
rect 4644 13764 4676 13765
rect 4644 13715 4676 13716
rect 4644 13685 4645 13715
rect 4645 13685 4675 13715
rect 4675 13685 4676 13715
rect 4644 13684 4676 13685
rect 4644 13635 4676 13636
rect 4644 13605 4645 13635
rect 4645 13605 4675 13635
rect 4675 13605 4676 13635
rect 4644 13604 4676 13605
rect 4644 13555 4676 13556
rect 4644 13525 4645 13555
rect 4645 13525 4675 13555
rect 4675 13525 4676 13555
rect 4644 13524 4676 13525
rect 4644 13475 4676 13476
rect 4644 13445 4645 13475
rect 4645 13445 4675 13475
rect 4675 13445 4676 13475
rect 4644 13444 4676 13445
rect 4644 13364 4676 13396
rect 4644 13284 4676 13316
rect 4644 13204 4676 13236
rect 4644 13124 4676 13156
rect 4644 13075 4676 13076
rect 4644 13045 4645 13075
rect 4645 13045 4675 13075
rect 4675 13045 4676 13075
rect 4644 13044 4676 13045
rect 4644 12995 4676 12996
rect 4644 12965 4645 12995
rect 4645 12965 4675 12995
rect 4675 12965 4676 12995
rect 4644 12964 4676 12965
rect 4644 12915 4676 12916
rect 4644 12885 4645 12915
rect 4645 12885 4675 12915
rect 4675 12885 4676 12915
rect 4644 12884 4676 12885
rect 4644 12835 4676 12836
rect 4644 12805 4645 12835
rect 4645 12805 4675 12835
rect 4675 12805 4676 12835
rect 4644 12804 4676 12805
rect 4644 12755 4676 12756
rect 4644 12725 4645 12755
rect 4645 12725 4675 12755
rect 4675 12725 4676 12755
rect 4644 12724 4676 12725
rect 4644 12675 4676 12676
rect 4644 12645 4645 12675
rect 4645 12645 4675 12675
rect 4675 12645 4676 12675
rect 4644 12644 4676 12645
rect 4644 12595 4676 12596
rect 4644 12565 4645 12595
rect 4645 12565 4675 12595
rect 4675 12565 4676 12595
rect 4644 12564 4676 12565
rect 4644 12515 4676 12516
rect 4644 12485 4645 12515
rect 4645 12485 4675 12515
rect 4675 12485 4676 12515
rect 4644 12484 4676 12485
rect 4644 12404 4676 12436
rect 4644 12355 4676 12356
rect 4644 12325 4645 12355
rect 4645 12325 4675 12355
rect 4675 12325 4676 12355
rect 4644 12324 4676 12325
rect 4644 12275 4676 12276
rect 4644 12245 4645 12275
rect 4645 12245 4675 12275
rect 4675 12245 4676 12275
rect 4644 12244 4676 12245
rect 4644 12195 4676 12196
rect 4644 12165 4645 12195
rect 4645 12165 4675 12195
rect 4675 12165 4676 12195
rect 4644 12164 4676 12165
rect 4644 12115 4676 12116
rect 4644 12085 4645 12115
rect 4645 12085 4675 12115
rect 4675 12085 4676 12115
rect 4644 12084 4676 12085
rect 4644 12035 4676 12036
rect 4644 12005 4645 12035
rect 4645 12005 4675 12035
rect 4675 12005 4676 12035
rect 4644 12004 4676 12005
rect 4644 11955 4676 11956
rect 4644 11925 4645 11955
rect 4645 11925 4675 11955
rect 4675 11925 4676 11955
rect 4644 11924 4676 11925
rect 4644 11875 4676 11876
rect 4644 11845 4645 11875
rect 4645 11845 4675 11875
rect 4675 11845 4676 11875
rect 4644 11844 4676 11845
rect 4644 11795 4676 11796
rect 4644 11765 4645 11795
rect 4645 11765 4675 11795
rect 4675 11765 4676 11795
rect 4644 11764 4676 11765
rect 4644 11715 4676 11716
rect 4644 11685 4645 11715
rect 4645 11685 4675 11715
rect 4675 11685 4676 11715
rect 4644 11684 4676 11685
rect 4644 11635 4676 11636
rect 4644 11605 4645 11635
rect 4645 11605 4675 11635
rect 4675 11605 4676 11635
rect 4644 11604 4676 11605
rect 4644 11555 4676 11556
rect 4644 11525 4645 11555
rect 4645 11525 4675 11555
rect 4675 11525 4676 11555
rect 4644 11524 4676 11525
rect 4644 11475 4676 11476
rect 4644 11445 4645 11475
rect 4645 11445 4675 11475
rect 4675 11445 4676 11475
rect 4644 11444 4676 11445
rect 4644 11395 4676 11396
rect 4644 11365 4645 11395
rect 4645 11365 4675 11395
rect 4675 11365 4676 11395
rect 4644 11364 4676 11365
rect 4644 11315 4676 11316
rect 4644 11285 4645 11315
rect 4645 11285 4675 11315
rect 4675 11285 4676 11315
rect 4644 11284 4676 11285
rect 4644 11235 4676 11236
rect 4644 11205 4645 11235
rect 4645 11205 4675 11235
rect 4675 11205 4676 11235
rect 4644 11204 4676 11205
rect 4644 11155 4676 11156
rect 4644 11125 4645 11155
rect 4645 11125 4675 11155
rect 4675 11125 4676 11155
rect 4644 11124 4676 11125
rect 4644 11075 4676 11076
rect 4644 11045 4645 11075
rect 4645 11045 4675 11075
rect 4675 11045 4676 11075
rect 4644 11044 4676 11045
rect 4644 10964 4676 10996
rect 4644 10915 4676 10916
rect 4644 10885 4645 10915
rect 4645 10885 4675 10915
rect 4675 10885 4676 10915
rect 4644 10884 4676 10885
rect 4644 10835 4676 10836
rect 4644 10805 4645 10835
rect 4645 10805 4675 10835
rect 4675 10805 4676 10835
rect 4644 10804 4676 10805
rect 4644 10755 4676 10756
rect 4644 10725 4645 10755
rect 4645 10725 4675 10755
rect 4675 10725 4676 10755
rect 4644 10724 4676 10725
rect 4644 10675 4676 10676
rect 4644 10645 4645 10675
rect 4645 10645 4675 10675
rect 4675 10645 4676 10675
rect 4644 10644 4676 10645
rect 4644 10595 4676 10596
rect 4644 10565 4645 10595
rect 4645 10565 4675 10595
rect 4675 10565 4676 10595
rect 4644 10564 4676 10565
rect 4644 10515 4676 10516
rect 4644 10485 4645 10515
rect 4645 10485 4675 10515
rect 4675 10485 4676 10515
rect 4644 10484 4676 10485
rect 4644 10435 4676 10436
rect 4644 10405 4645 10435
rect 4645 10405 4675 10435
rect 4675 10405 4676 10435
rect 4644 10404 4676 10405
rect 4644 10355 4676 10356
rect 4644 10325 4645 10355
rect 4645 10325 4675 10355
rect 4675 10325 4676 10355
rect 4644 10324 4676 10325
rect 4644 10244 4676 10276
rect 4644 10164 4676 10196
rect 4644 10084 4676 10116
rect 4644 10004 4676 10036
rect 4644 9955 4676 9956
rect 4644 9925 4645 9955
rect 4645 9925 4675 9955
rect 4675 9925 4676 9955
rect 4644 9924 4676 9925
rect 4644 9875 4676 9876
rect 4644 9845 4645 9875
rect 4645 9845 4675 9875
rect 4675 9845 4676 9875
rect 4644 9844 4676 9845
rect 4644 9795 4676 9796
rect 4644 9765 4645 9795
rect 4645 9765 4675 9795
rect 4675 9765 4676 9795
rect 4644 9764 4676 9765
rect 4644 9715 4676 9716
rect 4644 9685 4645 9715
rect 4645 9685 4675 9715
rect 4675 9685 4676 9715
rect 4644 9684 4676 9685
rect 4644 9635 4676 9636
rect 4644 9605 4645 9635
rect 4645 9605 4675 9635
rect 4675 9605 4676 9635
rect 4644 9604 4676 9605
rect 4644 9555 4676 9556
rect 4644 9525 4645 9555
rect 4645 9525 4675 9555
rect 4675 9525 4676 9555
rect 4644 9524 4676 9525
rect 4644 9475 4676 9476
rect 4644 9445 4645 9475
rect 4645 9445 4675 9475
rect 4675 9445 4676 9475
rect 4644 9444 4676 9445
rect 4644 9395 4676 9396
rect 4644 9365 4645 9395
rect 4645 9365 4675 9395
rect 4675 9365 4676 9395
rect 4644 9364 4676 9365
rect 4644 9284 4676 9316
rect 4644 9204 4676 9236
rect 4644 9124 4676 9156
rect 4644 9044 4676 9076
rect 4644 8995 4676 8996
rect 4644 8965 4645 8995
rect 4645 8965 4675 8995
rect 4675 8965 4676 8995
rect 4644 8964 4676 8965
rect 4644 8915 4676 8916
rect 4644 8885 4645 8915
rect 4645 8885 4675 8915
rect 4675 8885 4676 8915
rect 4644 8884 4676 8885
rect 4644 8835 4676 8836
rect 4644 8805 4645 8835
rect 4645 8805 4675 8835
rect 4675 8805 4676 8835
rect 4644 8804 4676 8805
rect 4644 8755 4676 8756
rect 4644 8725 4645 8755
rect 4645 8725 4675 8755
rect 4675 8725 4676 8755
rect 4644 8724 4676 8725
rect 4644 8675 4676 8676
rect 4644 8645 4645 8675
rect 4645 8645 4675 8675
rect 4675 8645 4676 8675
rect 4644 8644 4676 8645
rect 4644 8595 4676 8596
rect 4644 8565 4645 8595
rect 4645 8565 4675 8595
rect 4675 8565 4676 8595
rect 4644 8564 4676 8565
rect 4644 8515 4676 8516
rect 4644 8485 4645 8515
rect 4645 8485 4675 8515
rect 4675 8485 4676 8515
rect 4644 8484 4676 8485
rect 4644 8435 4676 8436
rect 4644 8405 4645 8435
rect 4645 8405 4675 8435
rect 4675 8405 4676 8435
rect 4644 8404 4676 8405
rect 4644 8324 4676 8356
rect 4644 8275 4676 8276
rect 4644 8245 4645 8275
rect 4645 8245 4675 8275
rect 4675 8245 4676 8275
rect 4644 8244 4676 8245
rect 4644 8195 4676 8196
rect 4644 8165 4645 8195
rect 4645 8165 4675 8195
rect 4675 8165 4676 8195
rect 4644 8164 4676 8165
rect 4644 8115 4676 8116
rect 4644 8085 4645 8115
rect 4645 8085 4675 8115
rect 4675 8085 4676 8115
rect 4644 8084 4676 8085
rect 4644 8035 4676 8036
rect 4644 8005 4645 8035
rect 4645 8005 4675 8035
rect 4675 8005 4676 8035
rect 4644 8004 4676 8005
rect 4644 7955 4676 7956
rect 4644 7925 4645 7955
rect 4645 7925 4675 7955
rect 4675 7925 4676 7955
rect 4644 7924 4676 7925
rect 4644 7875 4676 7876
rect 4644 7845 4645 7875
rect 4645 7845 4675 7875
rect 4675 7845 4676 7875
rect 4644 7844 4676 7845
rect 4644 7795 4676 7796
rect 4644 7765 4645 7795
rect 4645 7765 4675 7795
rect 4675 7765 4676 7795
rect 4644 7764 4676 7765
rect 4644 7715 4676 7716
rect 4644 7685 4645 7715
rect 4645 7685 4675 7715
rect 4675 7685 4676 7715
rect 4644 7684 4676 7685
rect 4644 7635 4676 7636
rect 4644 7605 4645 7635
rect 4645 7605 4675 7635
rect 4675 7605 4676 7635
rect 4644 7604 4676 7605
rect 4644 7555 4676 7556
rect 4644 7525 4645 7555
rect 4645 7525 4675 7555
rect 4675 7525 4676 7555
rect 4644 7524 4676 7525
rect 4644 7475 4676 7476
rect 4644 7445 4645 7475
rect 4645 7445 4675 7475
rect 4675 7445 4676 7475
rect 4644 7444 4676 7445
rect 4644 7395 4676 7396
rect 4644 7365 4645 7395
rect 4645 7365 4675 7395
rect 4675 7365 4676 7395
rect 4644 7364 4676 7365
rect 4644 7315 4676 7316
rect 4644 7285 4645 7315
rect 4645 7285 4675 7315
rect 4675 7285 4676 7315
rect 4644 7284 4676 7285
rect 4644 7235 4676 7236
rect 4644 7205 4645 7235
rect 4645 7205 4675 7235
rect 4675 7205 4676 7235
rect 4644 7204 4676 7205
rect 4644 7155 4676 7156
rect 4644 7125 4645 7155
rect 4645 7125 4675 7155
rect 4675 7125 4676 7155
rect 4644 7124 4676 7125
rect 4644 7075 4676 7076
rect 4644 7045 4645 7075
rect 4645 7045 4675 7075
rect 4675 7045 4676 7075
rect 4644 7044 4676 7045
rect 4644 6995 4676 6996
rect 4644 6965 4645 6995
rect 4645 6965 4675 6995
rect 4675 6965 4676 6995
rect 4644 6964 4676 6965
rect 4644 6884 4676 6916
rect 4644 6835 4676 6836
rect 4644 6805 4645 6835
rect 4645 6805 4675 6835
rect 4675 6805 4676 6835
rect 4644 6804 4676 6805
rect 4644 6755 4676 6756
rect 4644 6725 4645 6755
rect 4645 6725 4675 6755
rect 4675 6725 4676 6755
rect 4644 6724 4676 6725
rect 4644 6675 4676 6676
rect 4644 6645 4645 6675
rect 4645 6645 4675 6675
rect 4675 6645 4676 6675
rect 4644 6644 4676 6645
rect 4644 6595 4676 6596
rect 4644 6565 4645 6595
rect 4645 6565 4675 6595
rect 4675 6565 4676 6595
rect 4644 6564 4676 6565
rect 4644 6515 4676 6516
rect 4644 6485 4645 6515
rect 4645 6485 4675 6515
rect 4675 6485 4676 6515
rect 4644 6484 4676 6485
rect 4644 6435 4676 6436
rect 4644 6405 4645 6435
rect 4645 6405 4675 6435
rect 4675 6405 4676 6435
rect 4644 6404 4676 6405
rect 4644 6355 4676 6356
rect 4644 6325 4645 6355
rect 4645 6325 4675 6355
rect 4675 6325 4676 6355
rect 4644 6324 4676 6325
rect 4644 6275 4676 6276
rect 4644 6245 4645 6275
rect 4645 6245 4675 6275
rect 4675 6245 4676 6275
rect 4644 6244 4676 6245
rect 4644 6164 4676 6196
rect 4644 6084 4676 6116
rect 4644 6004 4676 6036
rect 4644 5924 4676 5956
rect 4644 5875 4676 5876
rect 4644 5845 4645 5875
rect 4645 5845 4675 5875
rect 4675 5845 4676 5875
rect 4644 5844 4676 5845
rect 4644 5795 4676 5796
rect 4644 5765 4645 5795
rect 4645 5765 4675 5795
rect 4675 5765 4676 5795
rect 4644 5764 4676 5765
rect 4644 5715 4676 5716
rect 4644 5685 4645 5715
rect 4645 5685 4675 5715
rect 4675 5685 4676 5715
rect 4644 5684 4676 5685
rect 4644 5635 4676 5636
rect 4644 5605 4645 5635
rect 4645 5605 4675 5635
rect 4675 5605 4676 5635
rect 4644 5604 4676 5605
rect 4644 5555 4676 5556
rect 4644 5525 4645 5555
rect 4645 5525 4675 5555
rect 4675 5525 4676 5555
rect 4644 5524 4676 5525
rect 4644 5475 4676 5476
rect 4644 5445 4645 5475
rect 4645 5445 4675 5475
rect 4675 5445 4676 5475
rect 4644 5444 4676 5445
rect 4644 5395 4676 5396
rect 4644 5365 4645 5395
rect 4645 5365 4675 5395
rect 4675 5365 4676 5395
rect 4644 5364 4676 5365
rect 4644 5315 4676 5316
rect 4644 5285 4645 5315
rect 4645 5285 4675 5315
rect 4675 5285 4676 5315
rect 4644 5284 4676 5285
rect 4644 5235 4676 5236
rect 4644 5205 4645 5235
rect 4645 5205 4675 5235
rect 4675 5205 4676 5235
rect 4644 5204 4676 5205
rect 4644 5155 4676 5156
rect 4644 5125 4645 5155
rect 4645 5125 4675 5155
rect 4675 5125 4676 5155
rect 4644 5124 4676 5125
rect 4644 5075 4676 5076
rect 4644 5045 4645 5075
rect 4645 5045 4675 5075
rect 4675 5045 4676 5075
rect 4644 5044 4676 5045
rect 4644 4995 4676 4996
rect 4644 4965 4645 4995
rect 4645 4965 4675 4995
rect 4675 4965 4676 4995
rect 4644 4964 4676 4965
rect 4644 4915 4676 4916
rect 4644 4885 4645 4915
rect 4645 4885 4675 4915
rect 4675 4885 4676 4915
rect 4644 4884 4676 4885
rect 4644 4804 4676 4836
rect 4644 4755 4676 4756
rect 4644 4725 4645 4755
rect 4645 4725 4675 4755
rect 4675 4725 4676 4755
rect 4644 4724 4676 4725
rect 4644 4675 4676 4676
rect 4644 4645 4645 4675
rect 4645 4645 4675 4675
rect 4675 4645 4676 4675
rect 4644 4644 4676 4645
rect 4644 4564 4676 4596
rect 4644 4515 4676 4516
rect 4644 4485 4645 4515
rect 4645 4485 4675 4515
rect 4675 4485 4676 4515
rect 4644 4484 4676 4485
rect 4644 4435 4676 4436
rect 4644 4405 4645 4435
rect 4645 4405 4675 4435
rect 4675 4405 4676 4435
rect 4644 4404 4676 4405
rect 4644 4355 4676 4356
rect 4644 4325 4645 4355
rect 4645 4325 4675 4355
rect 4675 4325 4676 4355
rect 4644 4324 4676 4325
rect 4644 4275 4676 4276
rect 4644 4245 4645 4275
rect 4645 4245 4675 4275
rect 4675 4245 4676 4275
rect 4644 4244 4676 4245
rect 4644 4195 4676 4196
rect 4644 4165 4645 4195
rect 4645 4165 4675 4195
rect 4675 4165 4676 4195
rect 4644 4164 4676 4165
rect 4644 4115 4676 4116
rect 4644 4085 4645 4115
rect 4645 4085 4675 4115
rect 4675 4085 4676 4115
rect 4644 4084 4676 4085
rect 4644 4035 4676 4036
rect 4644 4005 4645 4035
rect 4645 4005 4675 4035
rect 4675 4005 4676 4035
rect 4644 4004 4676 4005
rect 4644 3955 4676 3956
rect 4644 3925 4645 3955
rect 4645 3925 4675 3955
rect 4675 3925 4676 3955
rect 4644 3924 4676 3925
rect 4644 3875 4676 3876
rect 4644 3845 4645 3875
rect 4645 3845 4675 3875
rect 4675 3845 4676 3875
rect 4644 3844 4676 3845
rect 4644 3764 4676 3796
rect 4644 3715 4676 3716
rect 4644 3685 4645 3715
rect 4645 3685 4675 3715
rect 4675 3685 4676 3715
rect 4644 3684 4676 3685
rect 4644 3635 4676 3636
rect 4644 3605 4645 3635
rect 4645 3605 4675 3635
rect 4675 3605 4676 3635
rect 4644 3604 4676 3605
rect 4644 3524 4676 3556
rect 4644 3475 4676 3476
rect 4644 3445 4645 3475
rect 4645 3445 4675 3475
rect 4675 3445 4676 3475
rect 4644 3444 4676 3445
rect 4644 3395 4676 3396
rect 4644 3365 4645 3395
rect 4645 3365 4675 3395
rect 4675 3365 4676 3395
rect 4644 3364 4676 3365
rect 4644 3284 4676 3316
rect 4644 3235 4676 3236
rect 4644 3205 4645 3235
rect 4645 3205 4675 3235
rect 4675 3205 4676 3235
rect 4644 3204 4676 3205
rect 4644 3155 4676 3156
rect 4644 3125 4645 3155
rect 4645 3125 4675 3155
rect 4675 3125 4676 3155
rect 4644 3124 4676 3125
rect 4644 3075 4676 3076
rect 4644 3045 4645 3075
rect 4645 3045 4675 3075
rect 4675 3045 4676 3075
rect 4644 3044 4676 3045
rect 4644 2995 4676 2996
rect 4644 2965 4645 2995
rect 4645 2965 4675 2995
rect 4675 2965 4676 2995
rect 4644 2964 4676 2965
rect 4644 2915 4676 2916
rect 4644 2885 4645 2915
rect 4645 2885 4675 2915
rect 4675 2885 4676 2915
rect 4644 2884 4676 2885
rect 4644 2835 4676 2836
rect 4644 2805 4645 2835
rect 4645 2805 4675 2835
rect 4675 2805 4676 2835
rect 4644 2804 4676 2805
rect 4644 2755 4676 2756
rect 4644 2725 4645 2755
rect 4645 2725 4675 2755
rect 4675 2725 4676 2755
rect 4644 2724 4676 2725
rect 4644 2675 4676 2676
rect 4644 2645 4645 2675
rect 4645 2645 4675 2675
rect 4675 2645 4676 2675
rect 4644 2644 4676 2645
rect 4644 2595 4676 2596
rect 4644 2565 4645 2595
rect 4645 2565 4675 2595
rect 4675 2565 4676 2595
rect 4644 2564 4676 2565
rect 4644 2515 4676 2516
rect 4644 2485 4645 2515
rect 4645 2485 4675 2515
rect 4675 2485 4676 2515
rect 4644 2484 4676 2485
rect 4644 2435 4676 2436
rect 4644 2405 4645 2435
rect 4645 2405 4675 2435
rect 4675 2405 4676 2435
rect 4644 2404 4676 2405
rect 4644 2355 4676 2356
rect 4644 2325 4645 2355
rect 4645 2325 4675 2355
rect 4675 2325 4676 2355
rect 4644 2324 4676 2325
rect 4644 2275 4676 2276
rect 4644 2245 4645 2275
rect 4645 2245 4675 2275
rect 4675 2245 4676 2275
rect 4644 2244 4676 2245
rect 4644 2195 4676 2196
rect 4644 2165 4645 2195
rect 4645 2165 4675 2195
rect 4675 2165 4676 2195
rect 4644 2164 4676 2165
rect 4644 2115 4676 2116
rect 4644 2085 4645 2115
rect 4645 2085 4675 2115
rect 4675 2085 4676 2115
rect 4644 2084 4676 2085
rect 4644 2035 4676 2036
rect 4644 2005 4645 2035
rect 4645 2005 4675 2035
rect 4675 2005 4676 2035
rect 4644 2004 4676 2005
rect 4644 1955 4676 1956
rect 4644 1925 4645 1955
rect 4645 1925 4675 1955
rect 4675 1925 4676 1955
rect 4644 1924 4676 1925
rect 4644 1844 4676 1876
rect 4644 1764 4676 1796
rect 4644 1715 4676 1716
rect 4644 1685 4645 1715
rect 4645 1685 4675 1715
rect 4675 1685 4676 1715
rect 4644 1684 4676 1685
rect 4644 1635 4676 1636
rect 4644 1605 4645 1635
rect 4645 1605 4675 1635
rect 4675 1605 4676 1635
rect 4644 1604 4676 1605
rect 4644 1555 4676 1556
rect 4644 1525 4645 1555
rect 4645 1525 4675 1555
rect 4675 1525 4676 1555
rect 4644 1524 4676 1525
rect 4644 1475 4676 1476
rect 4644 1445 4645 1475
rect 4645 1445 4675 1475
rect 4675 1445 4676 1475
rect 4644 1444 4676 1445
rect 4644 1395 4676 1396
rect 4644 1365 4645 1395
rect 4645 1365 4675 1395
rect 4675 1365 4676 1395
rect 4644 1364 4676 1365
rect 4644 1315 4676 1316
rect 4644 1285 4645 1315
rect 4645 1285 4675 1315
rect 4675 1285 4676 1315
rect 4644 1284 4676 1285
rect 4644 1235 4676 1236
rect 4644 1205 4645 1235
rect 4645 1205 4675 1235
rect 4675 1205 4676 1235
rect 4644 1204 4676 1205
rect 4644 1155 4676 1156
rect 4644 1125 4645 1155
rect 4645 1125 4675 1155
rect 4675 1125 4676 1155
rect 4644 1124 4676 1125
rect 4644 1075 4676 1076
rect 4644 1045 4645 1075
rect 4645 1045 4675 1075
rect 4675 1045 4676 1075
rect 4644 1044 4676 1045
rect 4644 995 4676 996
rect 4644 965 4645 995
rect 4645 965 4675 995
rect 4675 965 4676 995
rect 4644 964 4676 965
rect 4644 884 4676 916
rect 4644 835 4676 836
rect 4644 805 4645 835
rect 4645 805 4675 835
rect 4675 805 4676 835
rect 4644 804 4676 805
rect 4644 755 4676 756
rect 4644 725 4645 755
rect 4645 725 4675 755
rect 4675 725 4676 755
rect 4644 724 4676 725
rect 4644 675 4676 676
rect 4644 645 4645 675
rect 4645 645 4675 675
rect 4675 645 4676 675
rect 4644 644 4676 645
rect 4644 595 4676 596
rect 4644 565 4645 595
rect 4645 565 4675 595
rect 4675 565 4676 595
rect 4644 564 4676 565
rect 4644 515 4676 516
rect 4644 485 4645 515
rect 4645 485 4675 515
rect 4675 485 4676 515
rect 4644 484 4676 485
rect 4644 404 4676 436
rect 4644 324 4676 356
rect 4644 275 4676 276
rect 4644 245 4645 275
rect 4645 245 4675 275
rect 4675 245 4676 275
rect 4644 244 4676 245
rect 4644 195 4676 196
rect 4644 165 4645 195
rect 4645 165 4675 195
rect 4675 165 4676 195
rect 4644 164 4676 165
rect 4644 115 4676 116
rect 4644 85 4645 115
rect 4645 85 4675 115
rect 4675 85 4676 115
rect 4644 84 4676 85
rect 4644 35 4676 36
rect 4644 5 4645 35
rect 4645 5 4675 35
rect 4675 5 4676 35
rect 4644 4 4676 5
rect 4644 -476 4676 -284
rect 4724 15715 4756 15716
rect 4724 15685 4725 15715
rect 4725 15685 4755 15715
rect 4755 15685 4756 15715
rect 4724 15684 4756 15685
rect 4724 15635 4756 15636
rect 4724 15605 4725 15635
rect 4725 15605 4755 15635
rect 4755 15605 4756 15635
rect 4724 15604 4756 15605
rect 4724 15555 4756 15556
rect 4724 15525 4725 15555
rect 4725 15525 4755 15555
rect 4755 15525 4756 15555
rect 4724 15524 4756 15525
rect 4724 15475 4756 15476
rect 4724 15445 4725 15475
rect 4725 15445 4755 15475
rect 4755 15445 4756 15475
rect 4724 15444 4756 15445
rect 4724 15395 4756 15396
rect 4724 15365 4725 15395
rect 4725 15365 4755 15395
rect 4755 15365 4756 15395
rect 4724 15364 4756 15365
rect 4724 15315 4756 15316
rect 4724 15285 4725 15315
rect 4725 15285 4755 15315
rect 4755 15285 4756 15315
rect 4724 15284 4756 15285
rect 4724 15235 4756 15236
rect 4724 15205 4725 15235
rect 4725 15205 4755 15235
rect 4755 15205 4756 15235
rect 4724 15204 4756 15205
rect 4724 15155 4756 15156
rect 4724 15125 4725 15155
rect 4725 15125 4755 15155
rect 4755 15125 4756 15155
rect 4724 15124 4756 15125
rect 4724 15044 4756 15076
rect 4724 14995 4756 14996
rect 4724 14965 4725 14995
rect 4725 14965 4755 14995
rect 4755 14965 4756 14995
rect 4724 14964 4756 14965
rect 4724 14915 4756 14916
rect 4724 14885 4725 14915
rect 4725 14885 4755 14915
rect 4755 14885 4756 14915
rect 4724 14884 4756 14885
rect 4724 14835 4756 14836
rect 4724 14805 4725 14835
rect 4725 14805 4755 14835
rect 4755 14805 4756 14835
rect 4724 14804 4756 14805
rect 4724 14755 4756 14756
rect 4724 14725 4725 14755
rect 4725 14725 4755 14755
rect 4755 14725 4756 14755
rect 4724 14724 4756 14725
rect 4724 14675 4756 14676
rect 4724 14645 4725 14675
rect 4725 14645 4755 14675
rect 4755 14645 4756 14675
rect 4724 14644 4756 14645
rect 4724 14595 4756 14596
rect 4724 14565 4725 14595
rect 4725 14565 4755 14595
rect 4755 14565 4756 14595
rect 4724 14564 4756 14565
rect 4724 14515 4756 14516
rect 4724 14485 4725 14515
rect 4725 14485 4755 14515
rect 4755 14485 4756 14515
rect 4724 14484 4756 14485
rect 4724 14435 4756 14436
rect 4724 14405 4725 14435
rect 4725 14405 4755 14435
rect 4755 14405 4756 14435
rect 4724 14404 4756 14405
rect 4724 14324 4756 14356
rect 4724 14244 4756 14276
rect 4724 14164 4756 14196
rect 4724 14084 4756 14116
rect 4724 14035 4756 14036
rect 4724 14005 4725 14035
rect 4725 14005 4755 14035
rect 4755 14005 4756 14035
rect 4724 14004 4756 14005
rect 4724 13955 4756 13956
rect 4724 13925 4725 13955
rect 4725 13925 4755 13955
rect 4755 13925 4756 13955
rect 4724 13924 4756 13925
rect 4724 13875 4756 13876
rect 4724 13845 4725 13875
rect 4725 13845 4755 13875
rect 4755 13845 4756 13875
rect 4724 13844 4756 13845
rect 4724 13795 4756 13796
rect 4724 13765 4725 13795
rect 4725 13765 4755 13795
rect 4755 13765 4756 13795
rect 4724 13764 4756 13765
rect 4724 13715 4756 13716
rect 4724 13685 4725 13715
rect 4725 13685 4755 13715
rect 4755 13685 4756 13715
rect 4724 13684 4756 13685
rect 4724 13635 4756 13636
rect 4724 13605 4725 13635
rect 4725 13605 4755 13635
rect 4755 13605 4756 13635
rect 4724 13604 4756 13605
rect 4724 13555 4756 13556
rect 4724 13525 4725 13555
rect 4725 13525 4755 13555
rect 4755 13525 4756 13555
rect 4724 13524 4756 13525
rect 4724 13475 4756 13476
rect 4724 13445 4725 13475
rect 4725 13445 4755 13475
rect 4755 13445 4756 13475
rect 4724 13444 4756 13445
rect 4724 13364 4756 13396
rect 4724 13284 4756 13316
rect 4724 13204 4756 13236
rect 4724 13124 4756 13156
rect 4724 13075 4756 13076
rect 4724 13045 4725 13075
rect 4725 13045 4755 13075
rect 4755 13045 4756 13075
rect 4724 13044 4756 13045
rect 4724 12995 4756 12996
rect 4724 12965 4725 12995
rect 4725 12965 4755 12995
rect 4755 12965 4756 12995
rect 4724 12964 4756 12965
rect 4724 12915 4756 12916
rect 4724 12885 4725 12915
rect 4725 12885 4755 12915
rect 4755 12885 4756 12915
rect 4724 12884 4756 12885
rect 4724 12835 4756 12836
rect 4724 12805 4725 12835
rect 4725 12805 4755 12835
rect 4755 12805 4756 12835
rect 4724 12804 4756 12805
rect 4724 12755 4756 12756
rect 4724 12725 4725 12755
rect 4725 12725 4755 12755
rect 4755 12725 4756 12755
rect 4724 12724 4756 12725
rect 4724 12675 4756 12676
rect 4724 12645 4725 12675
rect 4725 12645 4755 12675
rect 4755 12645 4756 12675
rect 4724 12644 4756 12645
rect 4724 12595 4756 12596
rect 4724 12565 4725 12595
rect 4725 12565 4755 12595
rect 4755 12565 4756 12595
rect 4724 12564 4756 12565
rect 4724 12515 4756 12516
rect 4724 12485 4725 12515
rect 4725 12485 4755 12515
rect 4755 12485 4756 12515
rect 4724 12484 4756 12485
rect 4724 12404 4756 12436
rect 4724 12355 4756 12356
rect 4724 12325 4725 12355
rect 4725 12325 4755 12355
rect 4755 12325 4756 12355
rect 4724 12324 4756 12325
rect 4724 12275 4756 12276
rect 4724 12245 4725 12275
rect 4725 12245 4755 12275
rect 4755 12245 4756 12275
rect 4724 12244 4756 12245
rect 4724 12195 4756 12196
rect 4724 12165 4725 12195
rect 4725 12165 4755 12195
rect 4755 12165 4756 12195
rect 4724 12164 4756 12165
rect 4724 12115 4756 12116
rect 4724 12085 4725 12115
rect 4725 12085 4755 12115
rect 4755 12085 4756 12115
rect 4724 12084 4756 12085
rect 4724 12035 4756 12036
rect 4724 12005 4725 12035
rect 4725 12005 4755 12035
rect 4755 12005 4756 12035
rect 4724 12004 4756 12005
rect 4724 11955 4756 11956
rect 4724 11925 4725 11955
rect 4725 11925 4755 11955
rect 4755 11925 4756 11955
rect 4724 11924 4756 11925
rect 4724 11875 4756 11876
rect 4724 11845 4725 11875
rect 4725 11845 4755 11875
rect 4755 11845 4756 11875
rect 4724 11844 4756 11845
rect 4724 11795 4756 11796
rect 4724 11765 4725 11795
rect 4725 11765 4755 11795
rect 4755 11765 4756 11795
rect 4724 11764 4756 11765
rect 4724 11715 4756 11716
rect 4724 11685 4725 11715
rect 4725 11685 4755 11715
rect 4755 11685 4756 11715
rect 4724 11684 4756 11685
rect 4724 11635 4756 11636
rect 4724 11605 4725 11635
rect 4725 11605 4755 11635
rect 4755 11605 4756 11635
rect 4724 11604 4756 11605
rect 4724 11555 4756 11556
rect 4724 11525 4725 11555
rect 4725 11525 4755 11555
rect 4755 11525 4756 11555
rect 4724 11524 4756 11525
rect 4724 11475 4756 11476
rect 4724 11445 4725 11475
rect 4725 11445 4755 11475
rect 4755 11445 4756 11475
rect 4724 11444 4756 11445
rect 4724 11395 4756 11396
rect 4724 11365 4725 11395
rect 4725 11365 4755 11395
rect 4755 11365 4756 11395
rect 4724 11364 4756 11365
rect 4724 11315 4756 11316
rect 4724 11285 4725 11315
rect 4725 11285 4755 11315
rect 4755 11285 4756 11315
rect 4724 11284 4756 11285
rect 4724 11235 4756 11236
rect 4724 11205 4725 11235
rect 4725 11205 4755 11235
rect 4755 11205 4756 11235
rect 4724 11204 4756 11205
rect 4724 11155 4756 11156
rect 4724 11125 4725 11155
rect 4725 11125 4755 11155
rect 4755 11125 4756 11155
rect 4724 11124 4756 11125
rect 4724 11075 4756 11076
rect 4724 11045 4725 11075
rect 4725 11045 4755 11075
rect 4755 11045 4756 11075
rect 4724 11044 4756 11045
rect 4724 10964 4756 10996
rect 4724 10915 4756 10916
rect 4724 10885 4725 10915
rect 4725 10885 4755 10915
rect 4755 10885 4756 10915
rect 4724 10884 4756 10885
rect 4724 10835 4756 10836
rect 4724 10805 4725 10835
rect 4725 10805 4755 10835
rect 4755 10805 4756 10835
rect 4724 10804 4756 10805
rect 4724 10755 4756 10756
rect 4724 10725 4725 10755
rect 4725 10725 4755 10755
rect 4755 10725 4756 10755
rect 4724 10724 4756 10725
rect 4724 10675 4756 10676
rect 4724 10645 4725 10675
rect 4725 10645 4755 10675
rect 4755 10645 4756 10675
rect 4724 10644 4756 10645
rect 4724 10595 4756 10596
rect 4724 10565 4725 10595
rect 4725 10565 4755 10595
rect 4755 10565 4756 10595
rect 4724 10564 4756 10565
rect 4724 10515 4756 10516
rect 4724 10485 4725 10515
rect 4725 10485 4755 10515
rect 4755 10485 4756 10515
rect 4724 10484 4756 10485
rect 4724 10435 4756 10436
rect 4724 10405 4725 10435
rect 4725 10405 4755 10435
rect 4755 10405 4756 10435
rect 4724 10404 4756 10405
rect 4724 10355 4756 10356
rect 4724 10325 4725 10355
rect 4725 10325 4755 10355
rect 4755 10325 4756 10355
rect 4724 10324 4756 10325
rect 4724 10244 4756 10276
rect 4724 10164 4756 10196
rect 4724 10084 4756 10116
rect 4724 10004 4756 10036
rect 4724 9955 4756 9956
rect 4724 9925 4725 9955
rect 4725 9925 4755 9955
rect 4755 9925 4756 9955
rect 4724 9924 4756 9925
rect 4724 9875 4756 9876
rect 4724 9845 4725 9875
rect 4725 9845 4755 9875
rect 4755 9845 4756 9875
rect 4724 9844 4756 9845
rect 4724 9795 4756 9796
rect 4724 9765 4725 9795
rect 4725 9765 4755 9795
rect 4755 9765 4756 9795
rect 4724 9764 4756 9765
rect 4724 9715 4756 9716
rect 4724 9685 4725 9715
rect 4725 9685 4755 9715
rect 4755 9685 4756 9715
rect 4724 9684 4756 9685
rect 4724 9635 4756 9636
rect 4724 9605 4725 9635
rect 4725 9605 4755 9635
rect 4755 9605 4756 9635
rect 4724 9604 4756 9605
rect 4724 9555 4756 9556
rect 4724 9525 4725 9555
rect 4725 9525 4755 9555
rect 4755 9525 4756 9555
rect 4724 9524 4756 9525
rect 4724 9475 4756 9476
rect 4724 9445 4725 9475
rect 4725 9445 4755 9475
rect 4755 9445 4756 9475
rect 4724 9444 4756 9445
rect 4724 9395 4756 9396
rect 4724 9365 4725 9395
rect 4725 9365 4755 9395
rect 4755 9365 4756 9395
rect 4724 9364 4756 9365
rect 4724 9284 4756 9316
rect 4724 9204 4756 9236
rect 4724 9124 4756 9156
rect 4724 9044 4756 9076
rect 4724 8995 4756 8996
rect 4724 8965 4725 8995
rect 4725 8965 4755 8995
rect 4755 8965 4756 8995
rect 4724 8964 4756 8965
rect 4724 8915 4756 8916
rect 4724 8885 4725 8915
rect 4725 8885 4755 8915
rect 4755 8885 4756 8915
rect 4724 8884 4756 8885
rect 4724 8835 4756 8836
rect 4724 8805 4725 8835
rect 4725 8805 4755 8835
rect 4755 8805 4756 8835
rect 4724 8804 4756 8805
rect 4724 8755 4756 8756
rect 4724 8725 4725 8755
rect 4725 8725 4755 8755
rect 4755 8725 4756 8755
rect 4724 8724 4756 8725
rect 4724 8675 4756 8676
rect 4724 8645 4725 8675
rect 4725 8645 4755 8675
rect 4755 8645 4756 8675
rect 4724 8644 4756 8645
rect 4724 8595 4756 8596
rect 4724 8565 4725 8595
rect 4725 8565 4755 8595
rect 4755 8565 4756 8595
rect 4724 8564 4756 8565
rect 4724 8515 4756 8516
rect 4724 8485 4725 8515
rect 4725 8485 4755 8515
rect 4755 8485 4756 8515
rect 4724 8484 4756 8485
rect 4724 8435 4756 8436
rect 4724 8405 4725 8435
rect 4725 8405 4755 8435
rect 4755 8405 4756 8435
rect 4724 8404 4756 8405
rect 4724 8324 4756 8356
rect 4724 8275 4756 8276
rect 4724 8245 4725 8275
rect 4725 8245 4755 8275
rect 4755 8245 4756 8275
rect 4724 8244 4756 8245
rect 4724 8195 4756 8196
rect 4724 8165 4725 8195
rect 4725 8165 4755 8195
rect 4755 8165 4756 8195
rect 4724 8164 4756 8165
rect 4724 8115 4756 8116
rect 4724 8085 4725 8115
rect 4725 8085 4755 8115
rect 4755 8085 4756 8115
rect 4724 8084 4756 8085
rect 4724 8035 4756 8036
rect 4724 8005 4725 8035
rect 4725 8005 4755 8035
rect 4755 8005 4756 8035
rect 4724 8004 4756 8005
rect 4724 7955 4756 7956
rect 4724 7925 4725 7955
rect 4725 7925 4755 7955
rect 4755 7925 4756 7955
rect 4724 7924 4756 7925
rect 4724 7875 4756 7876
rect 4724 7845 4725 7875
rect 4725 7845 4755 7875
rect 4755 7845 4756 7875
rect 4724 7844 4756 7845
rect 4724 7795 4756 7796
rect 4724 7765 4725 7795
rect 4725 7765 4755 7795
rect 4755 7765 4756 7795
rect 4724 7764 4756 7765
rect 4724 7715 4756 7716
rect 4724 7685 4725 7715
rect 4725 7685 4755 7715
rect 4755 7685 4756 7715
rect 4724 7684 4756 7685
rect 4724 7635 4756 7636
rect 4724 7605 4725 7635
rect 4725 7605 4755 7635
rect 4755 7605 4756 7635
rect 4724 7604 4756 7605
rect 4724 7555 4756 7556
rect 4724 7525 4725 7555
rect 4725 7525 4755 7555
rect 4755 7525 4756 7555
rect 4724 7524 4756 7525
rect 4724 7475 4756 7476
rect 4724 7445 4725 7475
rect 4725 7445 4755 7475
rect 4755 7445 4756 7475
rect 4724 7444 4756 7445
rect 4724 7395 4756 7396
rect 4724 7365 4725 7395
rect 4725 7365 4755 7395
rect 4755 7365 4756 7395
rect 4724 7364 4756 7365
rect 4724 7315 4756 7316
rect 4724 7285 4725 7315
rect 4725 7285 4755 7315
rect 4755 7285 4756 7315
rect 4724 7284 4756 7285
rect 4724 7235 4756 7236
rect 4724 7205 4725 7235
rect 4725 7205 4755 7235
rect 4755 7205 4756 7235
rect 4724 7204 4756 7205
rect 4724 7155 4756 7156
rect 4724 7125 4725 7155
rect 4725 7125 4755 7155
rect 4755 7125 4756 7155
rect 4724 7124 4756 7125
rect 4724 7075 4756 7076
rect 4724 7045 4725 7075
rect 4725 7045 4755 7075
rect 4755 7045 4756 7075
rect 4724 7044 4756 7045
rect 4724 6995 4756 6996
rect 4724 6965 4725 6995
rect 4725 6965 4755 6995
rect 4755 6965 4756 6995
rect 4724 6964 4756 6965
rect 4724 6884 4756 6916
rect 4724 6835 4756 6836
rect 4724 6805 4725 6835
rect 4725 6805 4755 6835
rect 4755 6805 4756 6835
rect 4724 6804 4756 6805
rect 4724 6755 4756 6756
rect 4724 6725 4725 6755
rect 4725 6725 4755 6755
rect 4755 6725 4756 6755
rect 4724 6724 4756 6725
rect 4724 6675 4756 6676
rect 4724 6645 4725 6675
rect 4725 6645 4755 6675
rect 4755 6645 4756 6675
rect 4724 6644 4756 6645
rect 4724 6595 4756 6596
rect 4724 6565 4725 6595
rect 4725 6565 4755 6595
rect 4755 6565 4756 6595
rect 4724 6564 4756 6565
rect 4724 6515 4756 6516
rect 4724 6485 4725 6515
rect 4725 6485 4755 6515
rect 4755 6485 4756 6515
rect 4724 6484 4756 6485
rect 4724 6435 4756 6436
rect 4724 6405 4725 6435
rect 4725 6405 4755 6435
rect 4755 6405 4756 6435
rect 4724 6404 4756 6405
rect 4724 6355 4756 6356
rect 4724 6325 4725 6355
rect 4725 6325 4755 6355
rect 4755 6325 4756 6355
rect 4724 6324 4756 6325
rect 4724 6275 4756 6276
rect 4724 6245 4725 6275
rect 4725 6245 4755 6275
rect 4755 6245 4756 6275
rect 4724 6244 4756 6245
rect 4724 6164 4756 6196
rect 4724 6084 4756 6116
rect 4724 6004 4756 6036
rect 4724 5924 4756 5956
rect 4724 5875 4756 5876
rect 4724 5845 4725 5875
rect 4725 5845 4755 5875
rect 4755 5845 4756 5875
rect 4724 5844 4756 5845
rect 4724 5795 4756 5796
rect 4724 5765 4725 5795
rect 4725 5765 4755 5795
rect 4755 5765 4756 5795
rect 4724 5764 4756 5765
rect 4724 5715 4756 5716
rect 4724 5685 4725 5715
rect 4725 5685 4755 5715
rect 4755 5685 4756 5715
rect 4724 5684 4756 5685
rect 4724 5635 4756 5636
rect 4724 5605 4725 5635
rect 4725 5605 4755 5635
rect 4755 5605 4756 5635
rect 4724 5604 4756 5605
rect 4724 5555 4756 5556
rect 4724 5525 4725 5555
rect 4725 5525 4755 5555
rect 4755 5525 4756 5555
rect 4724 5524 4756 5525
rect 4724 5475 4756 5476
rect 4724 5445 4725 5475
rect 4725 5445 4755 5475
rect 4755 5445 4756 5475
rect 4724 5444 4756 5445
rect 4724 5395 4756 5396
rect 4724 5365 4725 5395
rect 4725 5365 4755 5395
rect 4755 5365 4756 5395
rect 4724 5364 4756 5365
rect 4724 5315 4756 5316
rect 4724 5285 4725 5315
rect 4725 5285 4755 5315
rect 4755 5285 4756 5315
rect 4724 5284 4756 5285
rect 4724 5235 4756 5236
rect 4724 5205 4725 5235
rect 4725 5205 4755 5235
rect 4755 5205 4756 5235
rect 4724 5204 4756 5205
rect 4724 5155 4756 5156
rect 4724 5125 4725 5155
rect 4725 5125 4755 5155
rect 4755 5125 4756 5155
rect 4724 5124 4756 5125
rect 4724 5075 4756 5076
rect 4724 5045 4725 5075
rect 4725 5045 4755 5075
rect 4755 5045 4756 5075
rect 4724 5044 4756 5045
rect 4724 4995 4756 4996
rect 4724 4965 4725 4995
rect 4725 4965 4755 4995
rect 4755 4965 4756 4995
rect 4724 4964 4756 4965
rect 4724 4915 4756 4916
rect 4724 4885 4725 4915
rect 4725 4885 4755 4915
rect 4755 4885 4756 4915
rect 4724 4884 4756 4885
rect 4724 4804 4756 4836
rect 4724 4755 4756 4756
rect 4724 4725 4725 4755
rect 4725 4725 4755 4755
rect 4755 4725 4756 4755
rect 4724 4724 4756 4725
rect 4724 4675 4756 4676
rect 4724 4645 4725 4675
rect 4725 4645 4755 4675
rect 4755 4645 4756 4675
rect 4724 4644 4756 4645
rect 4724 4564 4756 4596
rect 4724 4515 4756 4516
rect 4724 4485 4725 4515
rect 4725 4485 4755 4515
rect 4755 4485 4756 4515
rect 4724 4484 4756 4485
rect 4724 4435 4756 4436
rect 4724 4405 4725 4435
rect 4725 4405 4755 4435
rect 4755 4405 4756 4435
rect 4724 4404 4756 4405
rect 4724 4355 4756 4356
rect 4724 4325 4725 4355
rect 4725 4325 4755 4355
rect 4755 4325 4756 4355
rect 4724 4324 4756 4325
rect 4724 4275 4756 4276
rect 4724 4245 4725 4275
rect 4725 4245 4755 4275
rect 4755 4245 4756 4275
rect 4724 4244 4756 4245
rect 4724 4195 4756 4196
rect 4724 4165 4725 4195
rect 4725 4165 4755 4195
rect 4755 4165 4756 4195
rect 4724 4164 4756 4165
rect 4724 4115 4756 4116
rect 4724 4085 4725 4115
rect 4725 4085 4755 4115
rect 4755 4085 4756 4115
rect 4724 4084 4756 4085
rect 4724 4035 4756 4036
rect 4724 4005 4725 4035
rect 4725 4005 4755 4035
rect 4755 4005 4756 4035
rect 4724 4004 4756 4005
rect 4724 3955 4756 3956
rect 4724 3925 4725 3955
rect 4725 3925 4755 3955
rect 4755 3925 4756 3955
rect 4724 3924 4756 3925
rect 4724 3875 4756 3876
rect 4724 3845 4725 3875
rect 4725 3845 4755 3875
rect 4755 3845 4756 3875
rect 4724 3844 4756 3845
rect 4724 3764 4756 3796
rect 4724 3715 4756 3716
rect 4724 3685 4725 3715
rect 4725 3685 4755 3715
rect 4755 3685 4756 3715
rect 4724 3684 4756 3685
rect 4724 3635 4756 3636
rect 4724 3605 4725 3635
rect 4725 3605 4755 3635
rect 4755 3605 4756 3635
rect 4724 3604 4756 3605
rect 4724 3524 4756 3556
rect 4724 3475 4756 3476
rect 4724 3445 4725 3475
rect 4725 3445 4755 3475
rect 4755 3445 4756 3475
rect 4724 3444 4756 3445
rect 4724 3395 4756 3396
rect 4724 3365 4725 3395
rect 4725 3365 4755 3395
rect 4755 3365 4756 3395
rect 4724 3364 4756 3365
rect 4724 3284 4756 3316
rect 4724 3235 4756 3236
rect 4724 3205 4725 3235
rect 4725 3205 4755 3235
rect 4755 3205 4756 3235
rect 4724 3204 4756 3205
rect 4724 3155 4756 3156
rect 4724 3125 4725 3155
rect 4725 3125 4755 3155
rect 4755 3125 4756 3155
rect 4724 3124 4756 3125
rect 4724 3075 4756 3076
rect 4724 3045 4725 3075
rect 4725 3045 4755 3075
rect 4755 3045 4756 3075
rect 4724 3044 4756 3045
rect 4724 2995 4756 2996
rect 4724 2965 4725 2995
rect 4725 2965 4755 2995
rect 4755 2965 4756 2995
rect 4724 2964 4756 2965
rect 4724 2915 4756 2916
rect 4724 2885 4725 2915
rect 4725 2885 4755 2915
rect 4755 2885 4756 2915
rect 4724 2884 4756 2885
rect 4724 2835 4756 2836
rect 4724 2805 4725 2835
rect 4725 2805 4755 2835
rect 4755 2805 4756 2835
rect 4724 2804 4756 2805
rect 4724 2755 4756 2756
rect 4724 2725 4725 2755
rect 4725 2725 4755 2755
rect 4755 2725 4756 2755
rect 4724 2724 4756 2725
rect 4724 2675 4756 2676
rect 4724 2645 4725 2675
rect 4725 2645 4755 2675
rect 4755 2645 4756 2675
rect 4724 2644 4756 2645
rect 4724 2595 4756 2596
rect 4724 2565 4725 2595
rect 4725 2565 4755 2595
rect 4755 2565 4756 2595
rect 4724 2564 4756 2565
rect 4724 2515 4756 2516
rect 4724 2485 4725 2515
rect 4725 2485 4755 2515
rect 4755 2485 4756 2515
rect 4724 2484 4756 2485
rect 4724 2435 4756 2436
rect 4724 2405 4725 2435
rect 4725 2405 4755 2435
rect 4755 2405 4756 2435
rect 4724 2404 4756 2405
rect 4724 2355 4756 2356
rect 4724 2325 4725 2355
rect 4725 2325 4755 2355
rect 4755 2325 4756 2355
rect 4724 2324 4756 2325
rect 4724 2275 4756 2276
rect 4724 2245 4725 2275
rect 4725 2245 4755 2275
rect 4755 2245 4756 2275
rect 4724 2244 4756 2245
rect 4724 2195 4756 2196
rect 4724 2165 4725 2195
rect 4725 2165 4755 2195
rect 4755 2165 4756 2195
rect 4724 2164 4756 2165
rect 4724 2115 4756 2116
rect 4724 2085 4725 2115
rect 4725 2085 4755 2115
rect 4755 2085 4756 2115
rect 4724 2084 4756 2085
rect 4724 2035 4756 2036
rect 4724 2005 4725 2035
rect 4725 2005 4755 2035
rect 4755 2005 4756 2035
rect 4724 2004 4756 2005
rect 4724 1955 4756 1956
rect 4724 1925 4725 1955
rect 4725 1925 4755 1955
rect 4755 1925 4756 1955
rect 4724 1924 4756 1925
rect 4724 1844 4756 1876
rect 4724 1764 4756 1796
rect 4724 1715 4756 1716
rect 4724 1685 4725 1715
rect 4725 1685 4755 1715
rect 4755 1685 4756 1715
rect 4724 1684 4756 1685
rect 4724 1635 4756 1636
rect 4724 1605 4725 1635
rect 4725 1605 4755 1635
rect 4755 1605 4756 1635
rect 4724 1604 4756 1605
rect 4724 1555 4756 1556
rect 4724 1525 4725 1555
rect 4725 1525 4755 1555
rect 4755 1525 4756 1555
rect 4724 1524 4756 1525
rect 4724 1475 4756 1476
rect 4724 1445 4725 1475
rect 4725 1445 4755 1475
rect 4755 1445 4756 1475
rect 4724 1444 4756 1445
rect 4724 1395 4756 1396
rect 4724 1365 4725 1395
rect 4725 1365 4755 1395
rect 4755 1365 4756 1395
rect 4724 1364 4756 1365
rect 4724 1315 4756 1316
rect 4724 1285 4725 1315
rect 4725 1285 4755 1315
rect 4755 1285 4756 1315
rect 4724 1284 4756 1285
rect 4724 1235 4756 1236
rect 4724 1205 4725 1235
rect 4725 1205 4755 1235
rect 4755 1205 4756 1235
rect 4724 1204 4756 1205
rect 4724 1155 4756 1156
rect 4724 1125 4725 1155
rect 4725 1125 4755 1155
rect 4755 1125 4756 1155
rect 4724 1124 4756 1125
rect 4724 1075 4756 1076
rect 4724 1045 4725 1075
rect 4725 1045 4755 1075
rect 4755 1045 4756 1075
rect 4724 1044 4756 1045
rect 4724 995 4756 996
rect 4724 965 4725 995
rect 4725 965 4755 995
rect 4755 965 4756 995
rect 4724 964 4756 965
rect 4724 884 4756 916
rect 4724 835 4756 836
rect 4724 805 4725 835
rect 4725 805 4755 835
rect 4755 805 4756 835
rect 4724 804 4756 805
rect 4724 755 4756 756
rect 4724 725 4725 755
rect 4725 725 4755 755
rect 4755 725 4756 755
rect 4724 724 4756 725
rect 4724 675 4756 676
rect 4724 645 4725 675
rect 4725 645 4755 675
rect 4755 645 4756 675
rect 4724 644 4756 645
rect 4724 595 4756 596
rect 4724 565 4725 595
rect 4725 565 4755 595
rect 4755 565 4756 595
rect 4724 564 4756 565
rect 4724 515 4756 516
rect 4724 485 4725 515
rect 4725 485 4755 515
rect 4755 485 4756 515
rect 4724 484 4756 485
rect 4724 404 4756 436
rect 4724 324 4756 356
rect 4724 275 4756 276
rect 4724 245 4725 275
rect 4725 245 4755 275
rect 4755 245 4756 275
rect 4724 244 4756 245
rect 4724 195 4756 196
rect 4724 165 4725 195
rect 4725 165 4755 195
rect 4755 165 4756 195
rect 4724 164 4756 165
rect 4724 115 4756 116
rect 4724 85 4725 115
rect 4725 85 4755 115
rect 4755 85 4756 115
rect 4724 84 4756 85
rect 4724 35 4756 36
rect 4724 5 4725 35
rect 4725 5 4755 35
rect 4755 5 4756 35
rect 4724 4 4756 5
rect 4884 15715 4916 15716
rect 4884 15685 4885 15715
rect 4885 15685 4915 15715
rect 4915 15685 4916 15715
rect 4884 15684 4916 15685
rect 4884 15635 4916 15636
rect 4884 15605 4885 15635
rect 4885 15605 4915 15635
rect 4915 15605 4916 15635
rect 4884 15604 4916 15605
rect 4884 15555 4916 15556
rect 4884 15525 4885 15555
rect 4885 15525 4915 15555
rect 4915 15525 4916 15555
rect 4884 15524 4916 15525
rect 4884 15475 4916 15476
rect 4884 15445 4885 15475
rect 4885 15445 4915 15475
rect 4915 15445 4916 15475
rect 4884 15444 4916 15445
rect 4884 15395 4916 15396
rect 4884 15365 4885 15395
rect 4885 15365 4915 15395
rect 4915 15365 4916 15395
rect 4884 15364 4916 15365
rect 4884 15315 4916 15316
rect 4884 15285 4885 15315
rect 4885 15285 4915 15315
rect 4915 15285 4916 15315
rect 4884 15284 4916 15285
rect 4884 15235 4916 15236
rect 4884 15205 4885 15235
rect 4885 15205 4915 15235
rect 4915 15205 4916 15235
rect 4884 15204 4916 15205
rect 4884 15155 4916 15156
rect 4884 15125 4885 15155
rect 4885 15125 4915 15155
rect 4915 15125 4916 15155
rect 4884 15124 4916 15125
rect 4884 15044 4916 15076
rect 4884 14995 4916 14996
rect 4884 14965 4885 14995
rect 4885 14965 4915 14995
rect 4915 14965 4916 14995
rect 4884 14964 4916 14965
rect 4884 14915 4916 14916
rect 4884 14885 4885 14915
rect 4885 14885 4915 14915
rect 4915 14885 4916 14915
rect 4884 14884 4916 14885
rect 4884 14835 4916 14836
rect 4884 14805 4885 14835
rect 4885 14805 4915 14835
rect 4915 14805 4916 14835
rect 4884 14804 4916 14805
rect 4884 14755 4916 14756
rect 4884 14725 4885 14755
rect 4885 14725 4915 14755
rect 4915 14725 4916 14755
rect 4884 14724 4916 14725
rect 4884 14675 4916 14676
rect 4884 14645 4885 14675
rect 4885 14645 4915 14675
rect 4915 14645 4916 14675
rect 4884 14644 4916 14645
rect 4884 14595 4916 14596
rect 4884 14565 4885 14595
rect 4885 14565 4915 14595
rect 4915 14565 4916 14595
rect 4884 14564 4916 14565
rect 4884 14515 4916 14516
rect 4884 14485 4885 14515
rect 4885 14485 4915 14515
rect 4915 14485 4916 14515
rect 4884 14484 4916 14485
rect 4884 14435 4916 14436
rect 4884 14405 4885 14435
rect 4885 14405 4915 14435
rect 4915 14405 4916 14435
rect 4884 14404 4916 14405
rect 4884 14324 4916 14356
rect 4884 14244 4916 14276
rect 4884 14164 4916 14196
rect 4884 14084 4916 14116
rect 4884 14035 4916 14036
rect 4884 14005 4885 14035
rect 4885 14005 4915 14035
rect 4915 14005 4916 14035
rect 4884 14004 4916 14005
rect 4884 13955 4916 13956
rect 4884 13925 4885 13955
rect 4885 13925 4915 13955
rect 4915 13925 4916 13955
rect 4884 13924 4916 13925
rect 4884 13875 4916 13876
rect 4884 13845 4885 13875
rect 4885 13845 4915 13875
rect 4915 13845 4916 13875
rect 4884 13844 4916 13845
rect 4884 13795 4916 13796
rect 4884 13765 4885 13795
rect 4885 13765 4915 13795
rect 4915 13765 4916 13795
rect 4884 13764 4916 13765
rect 4884 13715 4916 13716
rect 4884 13685 4885 13715
rect 4885 13685 4915 13715
rect 4915 13685 4916 13715
rect 4884 13684 4916 13685
rect 4884 13635 4916 13636
rect 4884 13605 4885 13635
rect 4885 13605 4915 13635
rect 4915 13605 4916 13635
rect 4884 13604 4916 13605
rect 4884 13555 4916 13556
rect 4884 13525 4885 13555
rect 4885 13525 4915 13555
rect 4915 13525 4916 13555
rect 4884 13524 4916 13525
rect 4884 13475 4916 13476
rect 4884 13445 4885 13475
rect 4885 13445 4915 13475
rect 4915 13445 4916 13475
rect 4884 13444 4916 13445
rect 4884 13364 4916 13396
rect 4884 13284 4916 13316
rect 4884 13204 4916 13236
rect 4884 13124 4916 13156
rect 4884 13075 4916 13076
rect 4884 13045 4885 13075
rect 4885 13045 4915 13075
rect 4915 13045 4916 13075
rect 4884 13044 4916 13045
rect 4884 12995 4916 12996
rect 4884 12965 4885 12995
rect 4885 12965 4915 12995
rect 4915 12965 4916 12995
rect 4884 12964 4916 12965
rect 4884 12915 4916 12916
rect 4884 12885 4885 12915
rect 4885 12885 4915 12915
rect 4915 12885 4916 12915
rect 4884 12884 4916 12885
rect 4884 12835 4916 12836
rect 4884 12805 4885 12835
rect 4885 12805 4915 12835
rect 4915 12805 4916 12835
rect 4884 12804 4916 12805
rect 4884 12755 4916 12756
rect 4884 12725 4885 12755
rect 4885 12725 4915 12755
rect 4915 12725 4916 12755
rect 4884 12724 4916 12725
rect 4884 12675 4916 12676
rect 4884 12645 4885 12675
rect 4885 12645 4915 12675
rect 4915 12645 4916 12675
rect 4884 12644 4916 12645
rect 4884 12595 4916 12596
rect 4884 12565 4885 12595
rect 4885 12565 4915 12595
rect 4915 12565 4916 12595
rect 4884 12564 4916 12565
rect 4884 12515 4916 12516
rect 4884 12485 4885 12515
rect 4885 12485 4915 12515
rect 4915 12485 4916 12515
rect 4884 12484 4916 12485
rect 4884 12404 4916 12436
rect 4884 12355 4916 12356
rect 4884 12325 4885 12355
rect 4885 12325 4915 12355
rect 4915 12325 4916 12355
rect 4884 12324 4916 12325
rect 4884 12275 4916 12276
rect 4884 12245 4885 12275
rect 4885 12245 4915 12275
rect 4915 12245 4916 12275
rect 4884 12244 4916 12245
rect 4884 12195 4916 12196
rect 4884 12165 4885 12195
rect 4885 12165 4915 12195
rect 4915 12165 4916 12195
rect 4884 12164 4916 12165
rect 4884 12115 4916 12116
rect 4884 12085 4885 12115
rect 4885 12085 4915 12115
rect 4915 12085 4916 12115
rect 4884 12084 4916 12085
rect 4884 12035 4916 12036
rect 4884 12005 4885 12035
rect 4885 12005 4915 12035
rect 4915 12005 4916 12035
rect 4884 12004 4916 12005
rect 4884 11955 4916 11956
rect 4884 11925 4885 11955
rect 4885 11925 4915 11955
rect 4915 11925 4916 11955
rect 4884 11924 4916 11925
rect 4884 11875 4916 11876
rect 4884 11845 4885 11875
rect 4885 11845 4915 11875
rect 4915 11845 4916 11875
rect 4884 11844 4916 11845
rect 4884 11795 4916 11796
rect 4884 11765 4885 11795
rect 4885 11765 4915 11795
rect 4915 11765 4916 11795
rect 4884 11764 4916 11765
rect 4884 11715 4916 11716
rect 4884 11685 4885 11715
rect 4885 11685 4915 11715
rect 4915 11685 4916 11715
rect 4884 11684 4916 11685
rect 4884 11635 4916 11636
rect 4884 11605 4885 11635
rect 4885 11605 4915 11635
rect 4915 11605 4916 11635
rect 4884 11604 4916 11605
rect 4884 11555 4916 11556
rect 4884 11525 4885 11555
rect 4885 11525 4915 11555
rect 4915 11525 4916 11555
rect 4884 11524 4916 11525
rect 4884 11475 4916 11476
rect 4884 11445 4885 11475
rect 4885 11445 4915 11475
rect 4915 11445 4916 11475
rect 4884 11444 4916 11445
rect 4884 11395 4916 11396
rect 4884 11365 4885 11395
rect 4885 11365 4915 11395
rect 4915 11365 4916 11395
rect 4884 11364 4916 11365
rect 4884 11315 4916 11316
rect 4884 11285 4885 11315
rect 4885 11285 4915 11315
rect 4915 11285 4916 11315
rect 4884 11284 4916 11285
rect 4884 11235 4916 11236
rect 4884 11205 4885 11235
rect 4885 11205 4915 11235
rect 4915 11205 4916 11235
rect 4884 11204 4916 11205
rect 4884 11155 4916 11156
rect 4884 11125 4885 11155
rect 4885 11125 4915 11155
rect 4915 11125 4916 11155
rect 4884 11124 4916 11125
rect 4884 11075 4916 11076
rect 4884 11045 4885 11075
rect 4885 11045 4915 11075
rect 4915 11045 4916 11075
rect 4884 11044 4916 11045
rect 4884 10964 4916 10996
rect 4884 10915 4916 10916
rect 4884 10885 4885 10915
rect 4885 10885 4915 10915
rect 4915 10885 4916 10915
rect 4884 10884 4916 10885
rect 4884 10835 4916 10836
rect 4884 10805 4885 10835
rect 4885 10805 4915 10835
rect 4915 10805 4916 10835
rect 4884 10804 4916 10805
rect 4884 10755 4916 10756
rect 4884 10725 4885 10755
rect 4885 10725 4915 10755
rect 4915 10725 4916 10755
rect 4884 10724 4916 10725
rect 4884 10675 4916 10676
rect 4884 10645 4885 10675
rect 4885 10645 4915 10675
rect 4915 10645 4916 10675
rect 4884 10644 4916 10645
rect 4884 10595 4916 10596
rect 4884 10565 4885 10595
rect 4885 10565 4915 10595
rect 4915 10565 4916 10595
rect 4884 10564 4916 10565
rect 4884 10515 4916 10516
rect 4884 10485 4885 10515
rect 4885 10485 4915 10515
rect 4915 10485 4916 10515
rect 4884 10484 4916 10485
rect 4884 10435 4916 10436
rect 4884 10405 4885 10435
rect 4885 10405 4915 10435
rect 4915 10405 4916 10435
rect 4884 10404 4916 10405
rect 4884 10355 4916 10356
rect 4884 10325 4885 10355
rect 4885 10325 4915 10355
rect 4915 10325 4916 10355
rect 4884 10324 4916 10325
rect 4884 10244 4916 10276
rect 4884 10164 4916 10196
rect 4884 10084 4916 10116
rect 4884 10004 4916 10036
rect 4884 9955 4916 9956
rect 4884 9925 4885 9955
rect 4885 9925 4915 9955
rect 4915 9925 4916 9955
rect 4884 9924 4916 9925
rect 4884 9875 4916 9876
rect 4884 9845 4885 9875
rect 4885 9845 4915 9875
rect 4915 9845 4916 9875
rect 4884 9844 4916 9845
rect 4884 9795 4916 9796
rect 4884 9765 4885 9795
rect 4885 9765 4915 9795
rect 4915 9765 4916 9795
rect 4884 9764 4916 9765
rect 4884 9715 4916 9716
rect 4884 9685 4885 9715
rect 4885 9685 4915 9715
rect 4915 9685 4916 9715
rect 4884 9684 4916 9685
rect 4884 9635 4916 9636
rect 4884 9605 4885 9635
rect 4885 9605 4915 9635
rect 4915 9605 4916 9635
rect 4884 9604 4916 9605
rect 4884 9555 4916 9556
rect 4884 9525 4885 9555
rect 4885 9525 4915 9555
rect 4915 9525 4916 9555
rect 4884 9524 4916 9525
rect 4884 9475 4916 9476
rect 4884 9445 4885 9475
rect 4885 9445 4915 9475
rect 4915 9445 4916 9475
rect 4884 9444 4916 9445
rect 4884 9395 4916 9396
rect 4884 9365 4885 9395
rect 4885 9365 4915 9395
rect 4915 9365 4916 9395
rect 4884 9364 4916 9365
rect 4884 9284 4916 9316
rect 4884 9204 4916 9236
rect 4884 9124 4916 9156
rect 4884 9044 4916 9076
rect 4884 8995 4916 8996
rect 4884 8965 4885 8995
rect 4885 8965 4915 8995
rect 4915 8965 4916 8995
rect 4884 8964 4916 8965
rect 4884 8915 4916 8916
rect 4884 8885 4885 8915
rect 4885 8885 4915 8915
rect 4915 8885 4916 8915
rect 4884 8884 4916 8885
rect 4884 8835 4916 8836
rect 4884 8805 4885 8835
rect 4885 8805 4915 8835
rect 4915 8805 4916 8835
rect 4884 8804 4916 8805
rect 4884 8755 4916 8756
rect 4884 8725 4885 8755
rect 4885 8725 4915 8755
rect 4915 8725 4916 8755
rect 4884 8724 4916 8725
rect 4884 8675 4916 8676
rect 4884 8645 4885 8675
rect 4885 8645 4915 8675
rect 4915 8645 4916 8675
rect 4884 8644 4916 8645
rect 4884 8595 4916 8596
rect 4884 8565 4885 8595
rect 4885 8565 4915 8595
rect 4915 8565 4916 8595
rect 4884 8564 4916 8565
rect 4884 8515 4916 8516
rect 4884 8485 4885 8515
rect 4885 8485 4915 8515
rect 4915 8485 4916 8515
rect 4884 8484 4916 8485
rect 4884 8435 4916 8436
rect 4884 8405 4885 8435
rect 4885 8405 4915 8435
rect 4915 8405 4916 8435
rect 4884 8404 4916 8405
rect 4884 8324 4916 8356
rect 4884 8275 4916 8276
rect 4884 8245 4885 8275
rect 4885 8245 4915 8275
rect 4915 8245 4916 8275
rect 4884 8244 4916 8245
rect 4884 8195 4916 8196
rect 4884 8165 4885 8195
rect 4885 8165 4915 8195
rect 4915 8165 4916 8195
rect 4884 8164 4916 8165
rect 4884 8115 4916 8116
rect 4884 8085 4885 8115
rect 4885 8085 4915 8115
rect 4915 8085 4916 8115
rect 4884 8084 4916 8085
rect 4884 8035 4916 8036
rect 4884 8005 4885 8035
rect 4885 8005 4915 8035
rect 4915 8005 4916 8035
rect 4884 8004 4916 8005
rect 4884 7955 4916 7956
rect 4884 7925 4885 7955
rect 4885 7925 4915 7955
rect 4915 7925 4916 7955
rect 4884 7924 4916 7925
rect 4884 7875 4916 7876
rect 4884 7845 4885 7875
rect 4885 7845 4915 7875
rect 4915 7845 4916 7875
rect 4884 7844 4916 7845
rect 4884 7795 4916 7796
rect 4884 7765 4885 7795
rect 4885 7765 4915 7795
rect 4915 7765 4916 7795
rect 4884 7764 4916 7765
rect 4884 7715 4916 7716
rect 4884 7685 4885 7715
rect 4885 7685 4915 7715
rect 4915 7685 4916 7715
rect 4884 7684 4916 7685
rect 4884 7635 4916 7636
rect 4884 7605 4885 7635
rect 4885 7605 4915 7635
rect 4915 7605 4916 7635
rect 4884 7604 4916 7605
rect 4884 7555 4916 7556
rect 4884 7525 4885 7555
rect 4885 7525 4915 7555
rect 4915 7525 4916 7555
rect 4884 7524 4916 7525
rect 4884 7475 4916 7476
rect 4884 7445 4885 7475
rect 4885 7445 4915 7475
rect 4915 7445 4916 7475
rect 4884 7444 4916 7445
rect 4884 7395 4916 7396
rect 4884 7365 4885 7395
rect 4885 7365 4915 7395
rect 4915 7365 4916 7395
rect 4884 7364 4916 7365
rect 4884 7315 4916 7316
rect 4884 7285 4885 7315
rect 4885 7285 4915 7315
rect 4915 7285 4916 7315
rect 4884 7284 4916 7285
rect 4884 7235 4916 7236
rect 4884 7205 4885 7235
rect 4885 7205 4915 7235
rect 4915 7205 4916 7235
rect 4884 7204 4916 7205
rect 4884 7155 4916 7156
rect 4884 7125 4885 7155
rect 4885 7125 4915 7155
rect 4915 7125 4916 7155
rect 4884 7124 4916 7125
rect 4884 7075 4916 7076
rect 4884 7045 4885 7075
rect 4885 7045 4915 7075
rect 4915 7045 4916 7075
rect 4884 7044 4916 7045
rect 4884 6995 4916 6996
rect 4884 6965 4885 6995
rect 4885 6965 4915 6995
rect 4915 6965 4916 6995
rect 4884 6964 4916 6965
rect 4884 6884 4916 6916
rect 4884 6835 4916 6836
rect 4884 6805 4885 6835
rect 4885 6805 4915 6835
rect 4915 6805 4916 6835
rect 4884 6804 4916 6805
rect 4884 6755 4916 6756
rect 4884 6725 4885 6755
rect 4885 6725 4915 6755
rect 4915 6725 4916 6755
rect 4884 6724 4916 6725
rect 4884 6675 4916 6676
rect 4884 6645 4885 6675
rect 4885 6645 4915 6675
rect 4915 6645 4916 6675
rect 4884 6644 4916 6645
rect 4884 6595 4916 6596
rect 4884 6565 4885 6595
rect 4885 6565 4915 6595
rect 4915 6565 4916 6595
rect 4884 6564 4916 6565
rect 4884 6515 4916 6516
rect 4884 6485 4885 6515
rect 4885 6485 4915 6515
rect 4915 6485 4916 6515
rect 4884 6484 4916 6485
rect 4884 6435 4916 6436
rect 4884 6405 4885 6435
rect 4885 6405 4915 6435
rect 4915 6405 4916 6435
rect 4884 6404 4916 6405
rect 4884 6355 4916 6356
rect 4884 6325 4885 6355
rect 4885 6325 4915 6355
rect 4915 6325 4916 6355
rect 4884 6324 4916 6325
rect 4884 6275 4916 6276
rect 4884 6245 4885 6275
rect 4885 6245 4915 6275
rect 4915 6245 4916 6275
rect 4884 6244 4916 6245
rect 4884 6164 4916 6196
rect 4884 6084 4916 6116
rect 4884 6004 4916 6036
rect 4884 5924 4916 5956
rect 4884 5875 4916 5876
rect 4884 5845 4885 5875
rect 4885 5845 4915 5875
rect 4915 5845 4916 5875
rect 4884 5844 4916 5845
rect 4884 5795 4916 5796
rect 4884 5765 4885 5795
rect 4885 5765 4915 5795
rect 4915 5765 4916 5795
rect 4884 5764 4916 5765
rect 4884 5715 4916 5716
rect 4884 5685 4885 5715
rect 4885 5685 4915 5715
rect 4915 5685 4916 5715
rect 4884 5684 4916 5685
rect 4884 5635 4916 5636
rect 4884 5605 4885 5635
rect 4885 5605 4915 5635
rect 4915 5605 4916 5635
rect 4884 5604 4916 5605
rect 4884 5555 4916 5556
rect 4884 5525 4885 5555
rect 4885 5525 4915 5555
rect 4915 5525 4916 5555
rect 4884 5524 4916 5525
rect 4884 5475 4916 5476
rect 4884 5445 4885 5475
rect 4885 5445 4915 5475
rect 4915 5445 4916 5475
rect 4884 5444 4916 5445
rect 4884 5395 4916 5396
rect 4884 5365 4885 5395
rect 4885 5365 4915 5395
rect 4915 5365 4916 5395
rect 4884 5364 4916 5365
rect 4884 5315 4916 5316
rect 4884 5285 4885 5315
rect 4885 5285 4915 5315
rect 4915 5285 4916 5315
rect 4884 5284 4916 5285
rect 4884 5235 4916 5236
rect 4884 5205 4885 5235
rect 4885 5205 4915 5235
rect 4915 5205 4916 5235
rect 4884 5204 4916 5205
rect 4884 5155 4916 5156
rect 4884 5125 4885 5155
rect 4885 5125 4915 5155
rect 4915 5125 4916 5155
rect 4884 5124 4916 5125
rect 4884 5075 4916 5076
rect 4884 5045 4885 5075
rect 4885 5045 4915 5075
rect 4915 5045 4916 5075
rect 4884 5044 4916 5045
rect 4884 4995 4916 4996
rect 4884 4965 4885 4995
rect 4885 4965 4915 4995
rect 4915 4965 4916 4995
rect 4884 4964 4916 4965
rect 4884 4915 4916 4916
rect 4884 4885 4885 4915
rect 4885 4885 4915 4915
rect 4915 4885 4916 4915
rect 4884 4884 4916 4885
rect 4884 4804 4916 4836
rect 4884 4755 4916 4756
rect 4884 4725 4885 4755
rect 4885 4725 4915 4755
rect 4915 4725 4916 4755
rect 4884 4724 4916 4725
rect 4884 4675 4916 4676
rect 4884 4645 4885 4675
rect 4885 4645 4915 4675
rect 4915 4645 4916 4675
rect 4884 4644 4916 4645
rect 4884 4564 4916 4596
rect 4884 4515 4916 4516
rect 4884 4485 4885 4515
rect 4885 4485 4915 4515
rect 4915 4485 4916 4515
rect 4884 4484 4916 4485
rect 4884 4435 4916 4436
rect 4884 4405 4885 4435
rect 4885 4405 4915 4435
rect 4915 4405 4916 4435
rect 4884 4404 4916 4405
rect 4884 4355 4916 4356
rect 4884 4325 4885 4355
rect 4885 4325 4915 4355
rect 4915 4325 4916 4355
rect 4884 4324 4916 4325
rect 4884 4275 4916 4276
rect 4884 4245 4885 4275
rect 4885 4245 4915 4275
rect 4915 4245 4916 4275
rect 4884 4244 4916 4245
rect 4884 4195 4916 4196
rect 4884 4165 4885 4195
rect 4885 4165 4915 4195
rect 4915 4165 4916 4195
rect 4884 4164 4916 4165
rect 4884 4115 4916 4116
rect 4884 4085 4885 4115
rect 4885 4085 4915 4115
rect 4915 4085 4916 4115
rect 4884 4084 4916 4085
rect 4884 4035 4916 4036
rect 4884 4005 4885 4035
rect 4885 4005 4915 4035
rect 4915 4005 4916 4035
rect 4884 4004 4916 4005
rect 4884 3955 4916 3956
rect 4884 3925 4885 3955
rect 4885 3925 4915 3955
rect 4915 3925 4916 3955
rect 4884 3924 4916 3925
rect 4884 3875 4916 3876
rect 4884 3845 4885 3875
rect 4885 3845 4915 3875
rect 4915 3845 4916 3875
rect 4884 3844 4916 3845
rect 4884 3764 4916 3796
rect 4884 3715 4916 3716
rect 4884 3685 4885 3715
rect 4885 3685 4915 3715
rect 4915 3685 4916 3715
rect 4884 3684 4916 3685
rect 4884 3635 4916 3636
rect 4884 3605 4885 3635
rect 4885 3605 4915 3635
rect 4915 3605 4916 3635
rect 4884 3604 4916 3605
rect 4884 3524 4916 3556
rect 4884 3475 4916 3476
rect 4884 3445 4885 3475
rect 4885 3445 4915 3475
rect 4915 3445 4916 3475
rect 4884 3444 4916 3445
rect 4884 3395 4916 3396
rect 4884 3365 4885 3395
rect 4885 3365 4915 3395
rect 4915 3365 4916 3395
rect 4884 3364 4916 3365
rect 4884 3284 4916 3316
rect 4884 3235 4916 3236
rect 4884 3205 4885 3235
rect 4885 3205 4915 3235
rect 4915 3205 4916 3235
rect 4884 3204 4916 3205
rect 4884 3155 4916 3156
rect 4884 3125 4885 3155
rect 4885 3125 4915 3155
rect 4915 3125 4916 3155
rect 4884 3124 4916 3125
rect 4884 3075 4916 3076
rect 4884 3045 4885 3075
rect 4885 3045 4915 3075
rect 4915 3045 4916 3075
rect 4884 3044 4916 3045
rect 4884 2995 4916 2996
rect 4884 2965 4885 2995
rect 4885 2965 4915 2995
rect 4915 2965 4916 2995
rect 4884 2964 4916 2965
rect 4884 2915 4916 2916
rect 4884 2885 4885 2915
rect 4885 2885 4915 2915
rect 4915 2885 4916 2915
rect 4884 2884 4916 2885
rect 4884 2835 4916 2836
rect 4884 2805 4885 2835
rect 4885 2805 4915 2835
rect 4915 2805 4916 2835
rect 4884 2804 4916 2805
rect 4884 2755 4916 2756
rect 4884 2725 4885 2755
rect 4885 2725 4915 2755
rect 4915 2725 4916 2755
rect 4884 2724 4916 2725
rect 4884 2675 4916 2676
rect 4884 2645 4885 2675
rect 4885 2645 4915 2675
rect 4915 2645 4916 2675
rect 4884 2644 4916 2645
rect 4884 2595 4916 2596
rect 4884 2565 4885 2595
rect 4885 2565 4915 2595
rect 4915 2565 4916 2595
rect 4884 2564 4916 2565
rect 4884 2515 4916 2516
rect 4884 2485 4885 2515
rect 4885 2485 4915 2515
rect 4915 2485 4916 2515
rect 4884 2484 4916 2485
rect 4884 2435 4916 2436
rect 4884 2405 4885 2435
rect 4885 2405 4915 2435
rect 4915 2405 4916 2435
rect 4884 2404 4916 2405
rect 4884 2355 4916 2356
rect 4884 2325 4885 2355
rect 4885 2325 4915 2355
rect 4915 2325 4916 2355
rect 4884 2324 4916 2325
rect 4884 2275 4916 2276
rect 4884 2245 4885 2275
rect 4885 2245 4915 2275
rect 4915 2245 4916 2275
rect 4884 2244 4916 2245
rect 4884 2195 4916 2196
rect 4884 2165 4885 2195
rect 4885 2165 4915 2195
rect 4915 2165 4916 2195
rect 4884 2164 4916 2165
rect 4884 2115 4916 2116
rect 4884 2085 4885 2115
rect 4885 2085 4915 2115
rect 4915 2085 4916 2115
rect 4884 2084 4916 2085
rect 4884 2035 4916 2036
rect 4884 2005 4885 2035
rect 4885 2005 4915 2035
rect 4915 2005 4916 2035
rect 4884 2004 4916 2005
rect 4884 1955 4916 1956
rect 4884 1925 4885 1955
rect 4885 1925 4915 1955
rect 4915 1925 4916 1955
rect 4884 1924 4916 1925
rect 4884 1844 4916 1876
rect 4884 1764 4916 1796
rect 4884 1715 4916 1716
rect 4884 1685 4885 1715
rect 4885 1685 4915 1715
rect 4915 1685 4916 1715
rect 4884 1684 4916 1685
rect 4884 1635 4916 1636
rect 4884 1605 4885 1635
rect 4885 1605 4915 1635
rect 4915 1605 4916 1635
rect 4884 1604 4916 1605
rect 4884 1555 4916 1556
rect 4884 1525 4885 1555
rect 4885 1525 4915 1555
rect 4915 1525 4916 1555
rect 4884 1524 4916 1525
rect 4884 1475 4916 1476
rect 4884 1445 4885 1475
rect 4885 1445 4915 1475
rect 4915 1445 4916 1475
rect 4884 1444 4916 1445
rect 4884 1395 4916 1396
rect 4884 1365 4885 1395
rect 4885 1365 4915 1395
rect 4915 1365 4916 1395
rect 4884 1364 4916 1365
rect 4884 1315 4916 1316
rect 4884 1285 4885 1315
rect 4885 1285 4915 1315
rect 4915 1285 4916 1315
rect 4884 1284 4916 1285
rect 4884 1235 4916 1236
rect 4884 1205 4885 1235
rect 4885 1205 4915 1235
rect 4915 1205 4916 1235
rect 4884 1204 4916 1205
rect 4884 1155 4916 1156
rect 4884 1125 4885 1155
rect 4885 1125 4915 1155
rect 4915 1125 4916 1155
rect 4884 1124 4916 1125
rect 4884 1075 4916 1076
rect 4884 1045 4885 1075
rect 4885 1045 4915 1075
rect 4915 1045 4916 1075
rect 4884 1044 4916 1045
rect 4884 995 4916 996
rect 4884 965 4885 995
rect 4885 965 4915 995
rect 4915 965 4916 995
rect 4884 964 4916 965
rect 4884 884 4916 916
rect 4884 835 4916 836
rect 4884 805 4885 835
rect 4885 805 4915 835
rect 4915 805 4916 835
rect 4884 804 4916 805
rect 4884 755 4916 756
rect 4884 725 4885 755
rect 4885 725 4915 755
rect 4915 725 4916 755
rect 4884 724 4916 725
rect 4884 675 4916 676
rect 4884 645 4885 675
rect 4885 645 4915 675
rect 4915 645 4916 675
rect 4884 644 4916 645
rect 4884 595 4916 596
rect 4884 565 4885 595
rect 4885 565 4915 595
rect 4915 565 4916 595
rect 4884 564 4916 565
rect 4884 515 4916 516
rect 4884 485 4885 515
rect 4885 485 4915 515
rect 4915 485 4916 515
rect 4884 484 4916 485
rect 4884 404 4916 436
rect 4884 324 4916 356
rect 4884 275 4916 276
rect 4884 245 4885 275
rect 4885 245 4915 275
rect 4915 245 4916 275
rect 4884 244 4916 245
rect 4884 195 4916 196
rect 4884 165 4885 195
rect 4885 165 4915 195
rect 4915 165 4916 195
rect 4884 164 4916 165
rect 4884 115 4916 116
rect 4884 85 4885 115
rect 4885 85 4915 115
rect 4915 85 4916 115
rect 4884 84 4916 85
rect 4884 35 4916 36
rect 4884 5 4885 35
rect 4885 5 4915 35
rect 4915 5 4916 35
rect 4884 4 4916 5
rect 4724 -716 4756 -524
rect 5044 15715 5076 15716
rect 5044 15685 5045 15715
rect 5045 15685 5075 15715
rect 5075 15685 5076 15715
rect 5044 15684 5076 15685
rect 5044 15635 5076 15636
rect 5044 15605 5045 15635
rect 5045 15605 5075 15635
rect 5075 15605 5076 15635
rect 5044 15604 5076 15605
rect 5044 15555 5076 15556
rect 5044 15525 5045 15555
rect 5045 15525 5075 15555
rect 5075 15525 5076 15555
rect 5044 15524 5076 15525
rect 5044 15475 5076 15476
rect 5044 15445 5045 15475
rect 5045 15445 5075 15475
rect 5075 15445 5076 15475
rect 5044 15444 5076 15445
rect 5044 15395 5076 15396
rect 5044 15365 5045 15395
rect 5045 15365 5075 15395
rect 5075 15365 5076 15395
rect 5044 15364 5076 15365
rect 5044 15315 5076 15316
rect 5044 15285 5045 15315
rect 5045 15285 5075 15315
rect 5075 15285 5076 15315
rect 5044 15284 5076 15285
rect 5044 15235 5076 15236
rect 5044 15205 5045 15235
rect 5045 15205 5075 15235
rect 5075 15205 5076 15235
rect 5044 15204 5076 15205
rect 5044 15155 5076 15156
rect 5044 15125 5045 15155
rect 5045 15125 5075 15155
rect 5075 15125 5076 15155
rect 5044 15124 5076 15125
rect 5044 15044 5076 15076
rect 5044 14995 5076 14996
rect 5044 14965 5045 14995
rect 5045 14965 5075 14995
rect 5075 14965 5076 14995
rect 5044 14964 5076 14965
rect 5044 14915 5076 14916
rect 5044 14885 5045 14915
rect 5045 14885 5075 14915
rect 5075 14885 5076 14915
rect 5044 14884 5076 14885
rect 5044 14835 5076 14836
rect 5044 14805 5045 14835
rect 5045 14805 5075 14835
rect 5075 14805 5076 14835
rect 5044 14804 5076 14805
rect 5044 14755 5076 14756
rect 5044 14725 5045 14755
rect 5045 14725 5075 14755
rect 5075 14725 5076 14755
rect 5044 14724 5076 14725
rect 5044 14675 5076 14676
rect 5044 14645 5045 14675
rect 5045 14645 5075 14675
rect 5075 14645 5076 14675
rect 5044 14644 5076 14645
rect 5044 14595 5076 14596
rect 5044 14565 5045 14595
rect 5045 14565 5075 14595
rect 5075 14565 5076 14595
rect 5044 14564 5076 14565
rect 5044 14515 5076 14516
rect 5044 14485 5045 14515
rect 5045 14485 5075 14515
rect 5075 14485 5076 14515
rect 5044 14484 5076 14485
rect 5044 14435 5076 14436
rect 5044 14405 5045 14435
rect 5045 14405 5075 14435
rect 5075 14405 5076 14435
rect 5044 14404 5076 14405
rect 5044 14324 5076 14356
rect 5044 14244 5076 14276
rect 5044 14164 5076 14196
rect 5044 14084 5076 14116
rect 5044 14035 5076 14036
rect 5044 14005 5045 14035
rect 5045 14005 5075 14035
rect 5075 14005 5076 14035
rect 5044 14004 5076 14005
rect 5044 13955 5076 13956
rect 5044 13925 5045 13955
rect 5045 13925 5075 13955
rect 5075 13925 5076 13955
rect 5044 13924 5076 13925
rect 5044 13875 5076 13876
rect 5044 13845 5045 13875
rect 5045 13845 5075 13875
rect 5075 13845 5076 13875
rect 5044 13844 5076 13845
rect 5044 13795 5076 13796
rect 5044 13765 5045 13795
rect 5045 13765 5075 13795
rect 5075 13765 5076 13795
rect 5044 13764 5076 13765
rect 5044 13715 5076 13716
rect 5044 13685 5045 13715
rect 5045 13685 5075 13715
rect 5075 13685 5076 13715
rect 5044 13684 5076 13685
rect 5044 13635 5076 13636
rect 5044 13605 5045 13635
rect 5045 13605 5075 13635
rect 5075 13605 5076 13635
rect 5044 13604 5076 13605
rect 5044 13555 5076 13556
rect 5044 13525 5045 13555
rect 5045 13525 5075 13555
rect 5075 13525 5076 13555
rect 5044 13524 5076 13525
rect 5044 13475 5076 13476
rect 5044 13445 5045 13475
rect 5045 13445 5075 13475
rect 5075 13445 5076 13475
rect 5044 13444 5076 13445
rect 5044 13364 5076 13396
rect 5044 13284 5076 13316
rect 5044 13204 5076 13236
rect 5044 13124 5076 13156
rect 5044 13075 5076 13076
rect 5044 13045 5045 13075
rect 5045 13045 5075 13075
rect 5075 13045 5076 13075
rect 5044 13044 5076 13045
rect 5044 12995 5076 12996
rect 5044 12965 5045 12995
rect 5045 12965 5075 12995
rect 5075 12965 5076 12995
rect 5044 12964 5076 12965
rect 5044 12915 5076 12916
rect 5044 12885 5045 12915
rect 5045 12885 5075 12915
rect 5075 12885 5076 12915
rect 5044 12884 5076 12885
rect 5044 12835 5076 12836
rect 5044 12805 5045 12835
rect 5045 12805 5075 12835
rect 5075 12805 5076 12835
rect 5044 12804 5076 12805
rect 5044 12755 5076 12756
rect 5044 12725 5045 12755
rect 5045 12725 5075 12755
rect 5075 12725 5076 12755
rect 5044 12724 5076 12725
rect 5044 12675 5076 12676
rect 5044 12645 5045 12675
rect 5045 12645 5075 12675
rect 5075 12645 5076 12675
rect 5044 12644 5076 12645
rect 5044 12595 5076 12596
rect 5044 12565 5045 12595
rect 5045 12565 5075 12595
rect 5075 12565 5076 12595
rect 5044 12564 5076 12565
rect 5044 12515 5076 12516
rect 5044 12485 5045 12515
rect 5045 12485 5075 12515
rect 5075 12485 5076 12515
rect 5044 12484 5076 12485
rect 5044 12404 5076 12436
rect 5044 12355 5076 12356
rect 5044 12325 5045 12355
rect 5045 12325 5075 12355
rect 5075 12325 5076 12355
rect 5044 12324 5076 12325
rect 5044 12275 5076 12276
rect 5044 12245 5045 12275
rect 5045 12245 5075 12275
rect 5075 12245 5076 12275
rect 5044 12244 5076 12245
rect 5044 12195 5076 12196
rect 5044 12165 5045 12195
rect 5045 12165 5075 12195
rect 5075 12165 5076 12195
rect 5044 12164 5076 12165
rect 5044 12115 5076 12116
rect 5044 12085 5045 12115
rect 5045 12085 5075 12115
rect 5075 12085 5076 12115
rect 5044 12084 5076 12085
rect 5044 12035 5076 12036
rect 5044 12005 5045 12035
rect 5045 12005 5075 12035
rect 5075 12005 5076 12035
rect 5044 12004 5076 12005
rect 5044 11955 5076 11956
rect 5044 11925 5045 11955
rect 5045 11925 5075 11955
rect 5075 11925 5076 11955
rect 5044 11924 5076 11925
rect 5044 11875 5076 11876
rect 5044 11845 5045 11875
rect 5045 11845 5075 11875
rect 5075 11845 5076 11875
rect 5044 11844 5076 11845
rect 5044 11795 5076 11796
rect 5044 11765 5045 11795
rect 5045 11765 5075 11795
rect 5075 11765 5076 11795
rect 5044 11764 5076 11765
rect 5044 11715 5076 11716
rect 5044 11685 5045 11715
rect 5045 11685 5075 11715
rect 5075 11685 5076 11715
rect 5044 11684 5076 11685
rect 5044 11635 5076 11636
rect 5044 11605 5045 11635
rect 5045 11605 5075 11635
rect 5075 11605 5076 11635
rect 5044 11604 5076 11605
rect 5044 11555 5076 11556
rect 5044 11525 5045 11555
rect 5045 11525 5075 11555
rect 5075 11525 5076 11555
rect 5044 11524 5076 11525
rect 5044 11475 5076 11476
rect 5044 11445 5045 11475
rect 5045 11445 5075 11475
rect 5075 11445 5076 11475
rect 5044 11444 5076 11445
rect 5044 11395 5076 11396
rect 5044 11365 5045 11395
rect 5045 11365 5075 11395
rect 5075 11365 5076 11395
rect 5044 11364 5076 11365
rect 5044 11315 5076 11316
rect 5044 11285 5045 11315
rect 5045 11285 5075 11315
rect 5075 11285 5076 11315
rect 5044 11284 5076 11285
rect 5044 11235 5076 11236
rect 5044 11205 5045 11235
rect 5045 11205 5075 11235
rect 5075 11205 5076 11235
rect 5044 11204 5076 11205
rect 5044 11155 5076 11156
rect 5044 11125 5045 11155
rect 5045 11125 5075 11155
rect 5075 11125 5076 11155
rect 5044 11124 5076 11125
rect 5044 11075 5076 11076
rect 5044 11045 5045 11075
rect 5045 11045 5075 11075
rect 5075 11045 5076 11075
rect 5044 11044 5076 11045
rect 5044 10964 5076 10996
rect 5044 10915 5076 10916
rect 5044 10885 5045 10915
rect 5045 10885 5075 10915
rect 5075 10885 5076 10915
rect 5044 10884 5076 10885
rect 5044 10835 5076 10836
rect 5044 10805 5045 10835
rect 5045 10805 5075 10835
rect 5075 10805 5076 10835
rect 5044 10804 5076 10805
rect 5044 10755 5076 10756
rect 5044 10725 5045 10755
rect 5045 10725 5075 10755
rect 5075 10725 5076 10755
rect 5044 10724 5076 10725
rect 5044 10675 5076 10676
rect 5044 10645 5045 10675
rect 5045 10645 5075 10675
rect 5075 10645 5076 10675
rect 5044 10644 5076 10645
rect 5044 10595 5076 10596
rect 5044 10565 5045 10595
rect 5045 10565 5075 10595
rect 5075 10565 5076 10595
rect 5044 10564 5076 10565
rect 5044 10515 5076 10516
rect 5044 10485 5045 10515
rect 5045 10485 5075 10515
rect 5075 10485 5076 10515
rect 5044 10484 5076 10485
rect 5044 10435 5076 10436
rect 5044 10405 5045 10435
rect 5045 10405 5075 10435
rect 5075 10405 5076 10435
rect 5044 10404 5076 10405
rect 5044 10355 5076 10356
rect 5044 10325 5045 10355
rect 5045 10325 5075 10355
rect 5075 10325 5076 10355
rect 5044 10324 5076 10325
rect 5044 10244 5076 10276
rect 5044 10164 5076 10196
rect 5044 10084 5076 10116
rect 5044 10004 5076 10036
rect 5044 9955 5076 9956
rect 5044 9925 5045 9955
rect 5045 9925 5075 9955
rect 5075 9925 5076 9955
rect 5044 9924 5076 9925
rect 5044 9875 5076 9876
rect 5044 9845 5045 9875
rect 5045 9845 5075 9875
rect 5075 9845 5076 9875
rect 5044 9844 5076 9845
rect 5044 9795 5076 9796
rect 5044 9765 5045 9795
rect 5045 9765 5075 9795
rect 5075 9765 5076 9795
rect 5044 9764 5076 9765
rect 5044 9715 5076 9716
rect 5044 9685 5045 9715
rect 5045 9685 5075 9715
rect 5075 9685 5076 9715
rect 5044 9684 5076 9685
rect 5044 9635 5076 9636
rect 5044 9605 5045 9635
rect 5045 9605 5075 9635
rect 5075 9605 5076 9635
rect 5044 9604 5076 9605
rect 5044 9555 5076 9556
rect 5044 9525 5045 9555
rect 5045 9525 5075 9555
rect 5075 9525 5076 9555
rect 5044 9524 5076 9525
rect 5044 9475 5076 9476
rect 5044 9445 5045 9475
rect 5045 9445 5075 9475
rect 5075 9445 5076 9475
rect 5044 9444 5076 9445
rect 5044 9395 5076 9396
rect 5044 9365 5045 9395
rect 5045 9365 5075 9395
rect 5075 9365 5076 9395
rect 5044 9364 5076 9365
rect 5044 9284 5076 9316
rect 5044 9204 5076 9236
rect 5044 9124 5076 9156
rect 5044 9044 5076 9076
rect 5044 8995 5076 8996
rect 5044 8965 5045 8995
rect 5045 8965 5075 8995
rect 5075 8965 5076 8995
rect 5044 8964 5076 8965
rect 5044 8915 5076 8916
rect 5044 8885 5045 8915
rect 5045 8885 5075 8915
rect 5075 8885 5076 8915
rect 5044 8884 5076 8885
rect 5044 8835 5076 8836
rect 5044 8805 5045 8835
rect 5045 8805 5075 8835
rect 5075 8805 5076 8835
rect 5044 8804 5076 8805
rect 5044 8755 5076 8756
rect 5044 8725 5045 8755
rect 5045 8725 5075 8755
rect 5075 8725 5076 8755
rect 5044 8724 5076 8725
rect 5044 8675 5076 8676
rect 5044 8645 5045 8675
rect 5045 8645 5075 8675
rect 5075 8645 5076 8675
rect 5044 8644 5076 8645
rect 5044 8595 5076 8596
rect 5044 8565 5045 8595
rect 5045 8565 5075 8595
rect 5075 8565 5076 8595
rect 5044 8564 5076 8565
rect 5044 8515 5076 8516
rect 5044 8485 5045 8515
rect 5045 8485 5075 8515
rect 5075 8485 5076 8515
rect 5044 8484 5076 8485
rect 5044 8435 5076 8436
rect 5044 8405 5045 8435
rect 5045 8405 5075 8435
rect 5075 8405 5076 8435
rect 5044 8404 5076 8405
rect 5044 8324 5076 8356
rect 5044 8275 5076 8276
rect 5044 8245 5045 8275
rect 5045 8245 5075 8275
rect 5075 8245 5076 8275
rect 5044 8244 5076 8245
rect 5044 8195 5076 8196
rect 5044 8165 5045 8195
rect 5045 8165 5075 8195
rect 5075 8165 5076 8195
rect 5044 8164 5076 8165
rect 5044 8115 5076 8116
rect 5044 8085 5045 8115
rect 5045 8085 5075 8115
rect 5075 8085 5076 8115
rect 5044 8084 5076 8085
rect 5044 8035 5076 8036
rect 5044 8005 5045 8035
rect 5045 8005 5075 8035
rect 5075 8005 5076 8035
rect 5044 8004 5076 8005
rect 5044 7955 5076 7956
rect 5044 7925 5045 7955
rect 5045 7925 5075 7955
rect 5075 7925 5076 7955
rect 5044 7924 5076 7925
rect 5044 7875 5076 7876
rect 5044 7845 5045 7875
rect 5045 7845 5075 7875
rect 5075 7845 5076 7875
rect 5044 7844 5076 7845
rect 5044 7795 5076 7796
rect 5044 7765 5045 7795
rect 5045 7765 5075 7795
rect 5075 7765 5076 7795
rect 5044 7764 5076 7765
rect 5044 7715 5076 7716
rect 5044 7685 5045 7715
rect 5045 7685 5075 7715
rect 5075 7685 5076 7715
rect 5044 7684 5076 7685
rect 5044 7635 5076 7636
rect 5044 7605 5045 7635
rect 5045 7605 5075 7635
rect 5075 7605 5076 7635
rect 5044 7604 5076 7605
rect 5044 7555 5076 7556
rect 5044 7525 5045 7555
rect 5045 7525 5075 7555
rect 5075 7525 5076 7555
rect 5044 7524 5076 7525
rect 5044 7475 5076 7476
rect 5044 7445 5045 7475
rect 5045 7445 5075 7475
rect 5075 7445 5076 7475
rect 5044 7444 5076 7445
rect 5044 7395 5076 7396
rect 5044 7365 5045 7395
rect 5045 7365 5075 7395
rect 5075 7365 5076 7395
rect 5044 7364 5076 7365
rect 5044 7315 5076 7316
rect 5044 7285 5045 7315
rect 5045 7285 5075 7315
rect 5075 7285 5076 7315
rect 5044 7284 5076 7285
rect 5044 7235 5076 7236
rect 5044 7205 5045 7235
rect 5045 7205 5075 7235
rect 5075 7205 5076 7235
rect 5044 7204 5076 7205
rect 5044 7155 5076 7156
rect 5044 7125 5045 7155
rect 5045 7125 5075 7155
rect 5075 7125 5076 7155
rect 5044 7124 5076 7125
rect 5044 7075 5076 7076
rect 5044 7045 5045 7075
rect 5045 7045 5075 7075
rect 5075 7045 5076 7075
rect 5044 7044 5076 7045
rect 5044 6995 5076 6996
rect 5044 6965 5045 6995
rect 5045 6965 5075 6995
rect 5075 6965 5076 6995
rect 5044 6964 5076 6965
rect 5044 6884 5076 6916
rect 5044 6835 5076 6836
rect 5044 6805 5045 6835
rect 5045 6805 5075 6835
rect 5075 6805 5076 6835
rect 5044 6804 5076 6805
rect 5044 6755 5076 6756
rect 5044 6725 5045 6755
rect 5045 6725 5075 6755
rect 5075 6725 5076 6755
rect 5044 6724 5076 6725
rect 5044 6675 5076 6676
rect 5044 6645 5045 6675
rect 5045 6645 5075 6675
rect 5075 6645 5076 6675
rect 5044 6644 5076 6645
rect 5044 6595 5076 6596
rect 5044 6565 5045 6595
rect 5045 6565 5075 6595
rect 5075 6565 5076 6595
rect 5044 6564 5076 6565
rect 5044 6515 5076 6516
rect 5044 6485 5045 6515
rect 5045 6485 5075 6515
rect 5075 6485 5076 6515
rect 5044 6484 5076 6485
rect 5044 6435 5076 6436
rect 5044 6405 5045 6435
rect 5045 6405 5075 6435
rect 5075 6405 5076 6435
rect 5044 6404 5076 6405
rect 5044 6355 5076 6356
rect 5044 6325 5045 6355
rect 5045 6325 5075 6355
rect 5075 6325 5076 6355
rect 5044 6324 5076 6325
rect 5044 6275 5076 6276
rect 5044 6245 5045 6275
rect 5045 6245 5075 6275
rect 5075 6245 5076 6275
rect 5044 6244 5076 6245
rect 5044 6164 5076 6196
rect 5044 6084 5076 6116
rect 5044 6004 5076 6036
rect 5044 5924 5076 5956
rect 5044 5875 5076 5876
rect 5044 5845 5045 5875
rect 5045 5845 5075 5875
rect 5075 5845 5076 5875
rect 5044 5844 5076 5845
rect 5044 5795 5076 5796
rect 5044 5765 5045 5795
rect 5045 5765 5075 5795
rect 5075 5765 5076 5795
rect 5044 5764 5076 5765
rect 5044 5715 5076 5716
rect 5044 5685 5045 5715
rect 5045 5685 5075 5715
rect 5075 5685 5076 5715
rect 5044 5684 5076 5685
rect 5044 5635 5076 5636
rect 5044 5605 5045 5635
rect 5045 5605 5075 5635
rect 5075 5605 5076 5635
rect 5044 5604 5076 5605
rect 5044 5555 5076 5556
rect 5044 5525 5045 5555
rect 5045 5525 5075 5555
rect 5075 5525 5076 5555
rect 5044 5524 5076 5525
rect 5044 5475 5076 5476
rect 5044 5445 5045 5475
rect 5045 5445 5075 5475
rect 5075 5445 5076 5475
rect 5044 5444 5076 5445
rect 5044 5395 5076 5396
rect 5044 5365 5045 5395
rect 5045 5365 5075 5395
rect 5075 5365 5076 5395
rect 5044 5364 5076 5365
rect 5044 5315 5076 5316
rect 5044 5285 5045 5315
rect 5045 5285 5075 5315
rect 5075 5285 5076 5315
rect 5044 5284 5076 5285
rect 5044 5235 5076 5236
rect 5044 5205 5045 5235
rect 5045 5205 5075 5235
rect 5075 5205 5076 5235
rect 5044 5204 5076 5205
rect 5044 5155 5076 5156
rect 5044 5125 5045 5155
rect 5045 5125 5075 5155
rect 5075 5125 5076 5155
rect 5044 5124 5076 5125
rect 5044 5075 5076 5076
rect 5044 5045 5045 5075
rect 5045 5045 5075 5075
rect 5075 5045 5076 5075
rect 5044 5044 5076 5045
rect 5044 4995 5076 4996
rect 5044 4965 5045 4995
rect 5045 4965 5075 4995
rect 5075 4965 5076 4995
rect 5044 4964 5076 4965
rect 5044 4915 5076 4916
rect 5044 4885 5045 4915
rect 5045 4885 5075 4915
rect 5075 4885 5076 4915
rect 5044 4884 5076 4885
rect 5044 4804 5076 4836
rect 5044 4755 5076 4756
rect 5044 4725 5045 4755
rect 5045 4725 5075 4755
rect 5075 4725 5076 4755
rect 5044 4724 5076 4725
rect 5044 4675 5076 4676
rect 5044 4645 5045 4675
rect 5045 4645 5075 4675
rect 5075 4645 5076 4675
rect 5044 4644 5076 4645
rect 5044 4564 5076 4596
rect 5044 4515 5076 4516
rect 5044 4485 5045 4515
rect 5045 4485 5075 4515
rect 5075 4485 5076 4515
rect 5044 4484 5076 4485
rect 5044 4435 5076 4436
rect 5044 4405 5045 4435
rect 5045 4405 5075 4435
rect 5075 4405 5076 4435
rect 5044 4404 5076 4405
rect 5044 4355 5076 4356
rect 5044 4325 5045 4355
rect 5045 4325 5075 4355
rect 5075 4325 5076 4355
rect 5044 4324 5076 4325
rect 5044 4275 5076 4276
rect 5044 4245 5045 4275
rect 5045 4245 5075 4275
rect 5075 4245 5076 4275
rect 5044 4244 5076 4245
rect 5044 4195 5076 4196
rect 5044 4165 5045 4195
rect 5045 4165 5075 4195
rect 5075 4165 5076 4195
rect 5044 4164 5076 4165
rect 5044 4115 5076 4116
rect 5044 4085 5045 4115
rect 5045 4085 5075 4115
rect 5075 4085 5076 4115
rect 5044 4084 5076 4085
rect 5044 4035 5076 4036
rect 5044 4005 5045 4035
rect 5045 4005 5075 4035
rect 5075 4005 5076 4035
rect 5044 4004 5076 4005
rect 5044 3955 5076 3956
rect 5044 3925 5045 3955
rect 5045 3925 5075 3955
rect 5075 3925 5076 3955
rect 5044 3924 5076 3925
rect 5044 3875 5076 3876
rect 5044 3845 5045 3875
rect 5045 3845 5075 3875
rect 5075 3845 5076 3875
rect 5044 3844 5076 3845
rect 5044 3764 5076 3796
rect 5044 3715 5076 3716
rect 5044 3685 5045 3715
rect 5045 3685 5075 3715
rect 5075 3685 5076 3715
rect 5044 3684 5076 3685
rect 5044 3635 5076 3636
rect 5044 3605 5045 3635
rect 5045 3605 5075 3635
rect 5075 3605 5076 3635
rect 5044 3604 5076 3605
rect 5044 3524 5076 3556
rect 5044 3475 5076 3476
rect 5044 3445 5045 3475
rect 5045 3445 5075 3475
rect 5075 3445 5076 3475
rect 5044 3444 5076 3445
rect 5044 3395 5076 3396
rect 5044 3365 5045 3395
rect 5045 3365 5075 3395
rect 5075 3365 5076 3395
rect 5044 3364 5076 3365
rect 5044 3284 5076 3316
rect 5044 3235 5076 3236
rect 5044 3205 5045 3235
rect 5045 3205 5075 3235
rect 5075 3205 5076 3235
rect 5044 3204 5076 3205
rect 5044 3155 5076 3156
rect 5044 3125 5045 3155
rect 5045 3125 5075 3155
rect 5075 3125 5076 3155
rect 5044 3124 5076 3125
rect 5044 3075 5076 3076
rect 5044 3045 5045 3075
rect 5045 3045 5075 3075
rect 5075 3045 5076 3075
rect 5044 3044 5076 3045
rect 5044 2995 5076 2996
rect 5044 2965 5045 2995
rect 5045 2965 5075 2995
rect 5075 2965 5076 2995
rect 5044 2964 5076 2965
rect 5044 2915 5076 2916
rect 5044 2885 5045 2915
rect 5045 2885 5075 2915
rect 5075 2885 5076 2915
rect 5044 2884 5076 2885
rect 5044 2835 5076 2836
rect 5044 2805 5045 2835
rect 5045 2805 5075 2835
rect 5075 2805 5076 2835
rect 5044 2804 5076 2805
rect 5044 2755 5076 2756
rect 5044 2725 5045 2755
rect 5045 2725 5075 2755
rect 5075 2725 5076 2755
rect 5044 2724 5076 2725
rect 5044 2675 5076 2676
rect 5044 2645 5045 2675
rect 5045 2645 5075 2675
rect 5075 2645 5076 2675
rect 5044 2644 5076 2645
rect 5044 2595 5076 2596
rect 5044 2565 5045 2595
rect 5045 2565 5075 2595
rect 5075 2565 5076 2595
rect 5044 2564 5076 2565
rect 5044 2515 5076 2516
rect 5044 2485 5045 2515
rect 5045 2485 5075 2515
rect 5075 2485 5076 2515
rect 5044 2484 5076 2485
rect 5044 2435 5076 2436
rect 5044 2405 5045 2435
rect 5045 2405 5075 2435
rect 5075 2405 5076 2435
rect 5044 2404 5076 2405
rect 5044 2355 5076 2356
rect 5044 2325 5045 2355
rect 5045 2325 5075 2355
rect 5075 2325 5076 2355
rect 5044 2324 5076 2325
rect 5044 2275 5076 2276
rect 5044 2245 5045 2275
rect 5045 2245 5075 2275
rect 5075 2245 5076 2275
rect 5044 2244 5076 2245
rect 5044 2195 5076 2196
rect 5044 2165 5045 2195
rect 5045 2165 5075 2195
rect 5075 2165 5076 2195
rect 5044 2164 5076 2165
rect 5044 2115 5076 2116
rect 5044 2085 5045 2115
rect 5045 2085 5075 2115
rect 5075 2085 5076 2115
rect 5044 2084 5076 2085
rect 5044 2035 5076 2036
rect 5044 2005 5045 2035
rect 5045 2005 5075 2035
rect 5075 2005 5076 2035
rect 5044 2004 5076 2005
rect 5044 1955 5076 1956
rect 5044 1925 5045 1955
rect 5045 1925 5075 1955
rect 5075 1925 5076 1955
rect 5044 1924 5076 1925
rect 5044 1844 5076 1876
rect 5044 1764 5076 1796
rect 5044 1715 5076 1716
rect 5044 1685 5045 1715
rect 5045 1685 5075 1715
rect 5075 1685 5076 1715
rect 5044 1684 5076 1685
rect 5044 1635 5076 1636
rect 5044 1605 5045 1635
rect 5045 1605 5075 1635
rect 5075 1605 5076 1635
rect 5044 1604 5076 1605
rect 5044 1555 5076 1556
rect 5044 1525 5045 1555
rect 5045 1525 5075 1555
rect 5075 1525 5076 1555
rect 5044 1524 5076 1525
rect 5044 1475 5076 1476
rect 5044 1445 5045 1475
rect 5045 1445 5075 1475
rect 5075 1445 5076 1475
rect 5044 1444 5076 1445
rect 5044 1395 5076 1396
rect 5044 1365 5045 1395
rect 5045 1365 5075 1395
rect 5075 1365 5076 1395
rect 5044 1364 5076 1365
rect 5044 1315 5076 1316
rect 5044 1285 5045 1315
rect 5045 1285 5075 1315
rect 5075 1285 5076 1315
rect 5044 1284 5076 1285
rect 5044 1235 5076 1236
rect 5044 1205 5045 1235
rect 5045 1205 5075 1235
rect 5075 1205 5076 1235
rect 5044 1204 5076 1205
rect 5044 1155 5076 1156
rect 5044 1125 5045 1155
rect 5045 1125 5075 1155
rect 5075 1125 5076 1155
rect 5044 1124 5076 1125
rect 5044 1075 5076 1076
rect 5044 1045 5045 1075
rect 5045 1045 5075 1075
rect 5075 1045 5076 1075
rect 5044 1044 5076 1045
rect 5044 995 5076 996
rect 5044 965 5045 995
rect 5045 965 5075 995
rect 5075 965 5076 995
rect 5044 964 5076 965
rect 5044 884 5076 916
rect 5044 835 5076 836
rect 5044 805 5045 835
rect 5045 805 5075 835
rect 5075 805 5076 835
rect 5044 804 5076 805
rect 5044 755 5076 756
rect 5044 725 5045 755
rect 5045 725 5075 755
rect 5075 725 5076 755
rect 5044 724 5076 725
rect 5044 675 5076 676
rect 5044 645 5045 675
rect 5045 645 5075 675
rect 5075 645 5076 675
rect 5044 644 5076 645
rect 5044 595 5076 596
rect 5044 565 5045 595
rect 5045 565 5075 595
rect 5075 565 5076 595
rect 5044 564 5076 565
rect 5044 515 5076 516
rect 5044 485 5045 515
rect 5045 485 5075 515
rect 5075 485 5076 515
rect 5044 484 5076 485
rect 5044 404 5076 436
rect 5044 324 5076 356
rect 5044 275 5076 276
rect 5044 245 5045 275
rect 5045 245 5075 275
rect 5075 245 5076 275
rect 5044 244 5076 245
rect 5044 195 5076 196
rect 5044 165 5045 195
rect 5045 165 5075 195
rect 5075 165 5076 195
rect 5044 164 5076 165
rect 5044 115 5076 116
rect 5044 85 5045 115
rect 5045 85 5075 115
rect 5075 85 5076 115
rect 5044 84 5076 85
rect 5044 35 5076 36
rect 5044 5 5045 35
rect 5045 5 5075 35
rect 5075 5 5076 35
rect 5044 4 5076 5
rect 4884 -716 4916 -524
rect 5204 15715 5236 15716
rect 5204 15685 5205 15715
rect 5205 15685 5235 15715
rect 5235 15685 5236 15715
rect 5204 15684 5236 15685
rect 5204 15635 5236 15636
rect 5204 15605 5205 15635
rect 5205 15605 5235 15635
rect 5235 15605 5236 15635
rect 5204 15604 5236 15605
rect 5204 15555 5236 15556
rect 5204 15525 5205 15555
rect 5205 15525 5235 15555
rect 5235 15525 5236 15555
rect 5204 15524 5236 15525
rect 5204 15475 5236 15476
rect 5204 15445 5205 15475
rect 5205 15445 5235 15475
rect 5235 15445 5236 15475
rect 5204 15444 5236 15445
rect 5204 15395 5236 15396
rect 5204 15365 5205 15395
rect 5205 15365 5235 15395
rect 5235 15365 5236 15395
rect 5204 15364 5236 15365
rect 5204 15315 5236 15316
rect 5204 15285 5205 15315
rect 5205 15285 5235 15315
rect 5235 15285 5236 15315
rect 5204 15284 5236 15285
rect 5204 15235 5236 15236
rect 5204 15205 5205 15235
rect 5205 15205 5235 15235
rect 5235 15205 5236 15235
rect 5204 15204 5236 15205
rect 5204 15155 5236 15156
rect 5204 15125 5205 15155
rect 5205 15125 5235 15155
rect 5235 15125 5236 15155
rect 5204 15124 5236 15125
rect 5204 15044 5236 15076
rect 5204 14995 5236 14996
rect 5204 14965 5205 14995
rect 5205 14965 5235 14995
rect 5235 14965 5236 14995
rect 5204 14964 5236 14965
rect 5204 14915 5236 14916
rect 5204 14885 5205 14915
rect 5205 14885 5235 14915
rect 5235 14885 5236 14915
rect 5204 14884 5236 14885
rect 5204 14835 5236 14836
rect 5204 14805 5205 14835
rect 5205 14805 5235 14835
rect 5235 14805 5236 14835
rect 5204 14804 5236 14805
rect 5204 14755 5236 14756
rect 5204 14725 5205 14755
rect 5205 14725 5235 14755
rect 5235 14725 5236 14755
rect 5204 14724 5236 14725
rect 5204 14675 5236 14676
rect 5204 14645 5205 14675
rect 5205 14645 5235 14675
rect 5235 14645 5236 14675
rect 5204 14644 5236 14645
rect 5204 14595 5236 14596
rect 5204 14565 5205 14595
rect 5205 14565 5235 14595
rect 5235 14565 5236 14595
rect 5204 14564 5236 14565
rect 5204 14515 5236 14516
rect 5204 14485 5205 14515
rect 5205 14485 5235 14515
rect 5235 14485 5236 14515
rect 5204 14484 5236 14485
rect 5204 14435 5236 14436
rect 5204 14405 5205 14435
rect 5205 14405 5235 14435
rect 5235 14405 5236 14435
rect 5204 14404 5236 14405
rect 5204 14324 5236 14356
rect 5204 14244 5236 14276
rect 5204 14164 5236 14196
rect 5204 14084 5236 14116
rect 5204 14035 5236 14036
rect 5204 14005 5205 14035
rect 5205 14005 5235 14035
rect 5235 14005 5236 14035
rect 5204 14004 5236 14005
rect 5204 13955 5236 13956
rect 5204 13925 5205 13955
rect 5205 13925 5235 13955
rect 5235 13925 5236 13955
rect 5204 13924 5236 13925
rect 5204 13875 5236 13876
rect 5204 13845 5205 13875
rect 5205 13845 5235 13875
rect 5235 13845 5236 13875
rect 5204 13844 5236 13845
rect 5204 13795 5236 13796
rect 5204 13765 5205 13795
rect 5205 13765 5235 13795
rect 5235 13765 5236 13795
rect 5204 13764 5236 13765
rect 5204 13715 5236 13716
rect 5204 13685 5205 13715
rect 5205 13685 5235 13715
rect 5235 13685 5236 13715
rect 5204 13684 5236 13685
rect 5204 13635 5236 13636
rect 5204 13605 5205 13635
rect 5205 13605 5235 13635
rect 5235 13605 5236 13635
rect 5204 13604 5236 13605
rect 5204 13555 5236 13556
rect 5204 13525 5205 13555
rect 5205 13525 5235 13555
rect 5235 13525 5236 13555
rect 5204 13524 5236 13525
rect 5204 13475 5236 13476
rect 5204 13445 5205 13475
rect 5205 13445 5235 13475
rect 5235 13445 5236 13475
rect 5204 13444 5236 13445
rect 5204 13364 5236 13396
rect 5204 13284 5236 13316
rect 5204 13204 5236 13236
rect 5204 13124 5236 13156
rect 5204 13075 5236 13076
rect 5204 13045 5205 13075
rect 5205 13045 5235 13075
rect 5235 13045 5236 13075
rect 5204 13044 5236 13045
rect 5204 12995 5236 12996
rect 5204 12965 5205 12995
rect 5205 12965 5235 12995
rect 5235 12965 5236 12995
rect 5204 12964 5236 12965
rect 5204 12915 5236 12916
rect 5204 12885 5205 12915
rect 5205 12885 5235 12915
rect 5235 12885 5236 12915
rect 5204 12884 5236 12885
rect 5204 12835 5236 12836
rect 5204 12805 5205 12835
rect 5205 12805 5235 12835
rect 5235 12805 5236 12835
rect 5204 12804 5236 12805
rect 5204 12755 5236 12756
rect 5204 12725 5205 12755
rect 5205 12725 5235 12755
rect 5235 12725 5236 12755
rect 5204 12724 5236 12725
rect 5204 12675 5236 12676
rect 5204 12645 5205 12675
rect 5205 12645 5235 12675
rect 5235 12645 5236 12675
rect 5204 12644 5236 12645
rect 5204 12595 5236 12596
rect 5204 12565 5205 12595
rect 5205 12565 5235 12595
rect 5235 12565 5236 12595
rect 5204 12564 5236 12565
rect 5204 12515 5236 12516
rect 5204 12485 5205 12515
rect 5205 12485 5235 12515
rect 5235 12485 5236 12515
rect 5204 12484 5236 12485
rect 5204 12404 5236 12436
rect 5204 12355 5236 12356
rect 5204 12325 5205 12355
rect 5205 12325 5235 12355
rect 5235 12325 5236 12355
rect 5204 12324 5236 12325
rect 5204 12275 5236 12276
rect 5204 12245 5205 12275
rect 5205 12245 5235 12275
rect 5235 12245 5236 12275
rect 5204 12244 5236 12245
rect 5204 12195 5236 12196
rect 5204 12165 5205 12195
rect 5205 12165 5235 12195
rect 5235 12165 5236 12195
rect 5204 12164 5236 12165
rect 5204 12115 5236 12116
rect 5204 12085 5205 12115
rect 5205 12085 5235 12115
rect 5235 12085 5236 12115
rect 5204 12084 5236 12085
rect 5204 12035 5236 12036
rect 5204 12005 5205 12035
rect 5205 12005 5235 12035
rect 5235 12005 5236 12035
rect 5204 12004 5236 12005
rect 5204 11955 5236 11956
rect 5204 11925 5205 11955
rect 5205 11925 5235 11955
rect 5235 11925 5236 11955
rect 5204 11924 5236 11925
rect 5204 11875 5236 11876
rect 5204 11845 5205 11875
rect 5205 11845 5235 11875
rect 5235 11845 5236 11875
rect 5204 11844 5236 11845
rect 5204 11795 5236 11796
rect 5204 11765 5205 11795
rect 5205 11765 5235 11795
rect 5235 11765 5236 11795
rect 5204 11764 5236 11765
rect 5204 11715 5236 11716
rect 5204 11685 5205 11715
rect 5205 11685 5235 11715
rect 5235 11685 5236 11715
rect 5204 11684 5236 11685
rect 5204 11635 5236 11636
rect 5204 11605 5205 11635
rect 5205 11605 5235 11635
rect 5235 11605 5236 11635
rect 5204 11604 5236 11605
rect 5204 11555 5236 11556
rect 5204 11525 5205 11555
rect 5205 11525 5235 11555
rect 5235 11525 5236 11555
rect 5204 11524 5236 11525
rect 5204 11475 5236 11476
rect 5204 11445 5205 11475
rect 5205 11445 5235 11475
rect 5235 11445 5236 11475
rect 5204 11444 5236 11445
rect 5204 11395 5236 11396
rect 5204 11365 5205 11395
rect 5205 11365 5235 11395
rect 5235 11365 5236 11395
rect 5204 11364 5236 11365
rect 5204 11315 5236 11316
rect 5204 11285 5205 11315
rect 5205 11285 5235 11315
rect 5235 11285 5236 11315
rect 5204 11284 5236 11285
rect 5204 11235 5236 11236
rect 5204 11205 5205 11235
rect 5205 11205 5235 11235
rect 5235 11205 5236 11235
rect 5204 11204 5236 11205
rect 5204 11155 5236 11156
rect 5204 11125 5205 11155
rect 5205 11125 5235 11155
rect 5235 11125 5236 11155
rect 5204 11124 5236 11125
rect 5204 11075 5236 11076
rect 5204 11045 5205 11075
rect 5205 11045 5235 11075
rect 5235 11045 5236 11075
rect 5204 11044 5236 11045
rect 5204 10964 5236 10996
rect 5204 10915 5236 10916
rect 5204 10885 5205 10915
rect 5205 10885 5235 10915
rect 5235 10885 5236 10915
rect 5204 10884 5236 10885
rect 5204 10835 5236 10836
rect 5204 10805 5205 10835
rect 5205 10805 5235 10835
rect 5235 10805 5236 10835
rect 5204 10804 5236 10805
rect 5204 10755 5236 10756
rect 5204 10725 5205 10755
rect 5205 10725 5235 10755
rect 5235 10725 5236 10755
rect 5204 10724 5236 10725
rect 5204 10675 5236 10676
rect 5204 10645 5205 10675
rect 5205 10645 5235 10675
rect 5235 10645 5236 10675
rect 5204 10644 5236 10645
rect 5204 10595 5236 10596
rect 5204 10565 5205 10595
rect 5205 10565 5235 10595
rect 5235 10565 5236 10595
rect 5204 10564 5236 10565
rect 5204 10515 5236 10516
rect 5204 10485 5205 10515
rect 5205 10485 5235 10515
rect 5235 10485 5236 10515
rect 5204 10484 5236 10485
rect 5204 10435 5236 10436
rect 5204 10405 5205 10435
rect 5205 10405 5235 10435
rect 5235 10405 5236 10435
rect 5204 10404 5236 10405
rect 5204 10355 5236 10356
rect 5204 10325 5205 10355
rect 5205 10325 5235 10355
rect 5235 10325 5236 10355
rect 5204 10324 5236 10325
rect 5204 10244 5236 10276
rect 5204 10164 5236 10196
rect 5204 10084 5236 10116
rect 5204 10004 5236 10036
rect 5204 9955 5236 9956
rect 5204 9925 5205 9955
rect 5205 9925 5235 9955
rect 5235 9925 5236 9955
rect 5204 9924 5236 9925
rect 5204 9875 5236 9876
rect 5204 9845 5205 9875
rect 5205 9845 5235 9875
rect 5235 9845 5236 9875
rect 5204 9844 5236 9845
rect 5204 9795 5236 9796
rect 5204 9765 5205 9795
rect 5205 9765 5235 9795
rect 5235 9765 5236 9795
rect 5204 9764 5236 9765
rect 5204 9715 5236 9716
rect 5204 9685 5205 9715
rect 5205 9685 5235 9715
rect 5235 9685 5236 9715
rect 5204 9684 5236 9685
rect 5204 9635 5236 9636
rect 5204 9605 5205 9635
rect 5205 9605 5235 9635
rect 5235 9605 5236 9635
rect 5204 9604 5236 9605
rect 5204 9555 5236 9556
rect 5204 9525 5205 9555
rect 5205 9525 5235 9555
rect 5235 9525 5236 9555
rect 5204 9524 5236 9525
rect 5204 9475 5236 9476
rect 5204 9445 5205 9475
rect 5205 9445 5235 9475
rect 5235 9445 5236 9475
rect 5204 9444 5236 9445
rect 5204 9395 5236 9396
rect 5204 9365 5205 9395
rect 5205 9365 5235 9395
rect 5235 9365 5236 9395
rect 5204 9364 5236 9365
rect 5204 9284 5236 9316
rect 5204 9204 5236 9236
rect 5204 9124 5236 9156
rect 5204 9044 5236 9076
rect 5204 8995 5236 8996
rect 5204 8965 5205 8995
rect 5205 8965 5235 8995
rect 5235 8965 5236 8995
rect 5204 8964 5236 8965
rect 5204 8915 5236 8916
rect 5204 8885 5205 8915
rect 5205 8885 5235 8915
rect 5235 8885 5236 8915
rect 5204 8884 5236 8885
rect 5204 8835 5236 8836
rect 5204 8805 5205 8835
rect 5205 8805 5235 8835
rect 5235 8805 5236 8835
rect 5204 8804 5236 8805
rect 5204 8755 5236 8756
rect 5204 8725 5205 8755
rect 5205 8725 5235 8755
rect 5235 8725 5236 8755
rect 5204 8724 5236 8725
rect 5204 8675 5236 8676
rect 5204 8645 5205 8675
rect 5205 8645 5235 8675
rect 5235 8645 5236 8675
rect 5204 8644 5236 8645
rect 5204 8595 5236 8596
rect 5204 8565 5205 8595
rect 5205 8565 5235 8595
rect 5235 8565 5236 8595
rect 5204 8564 5236 8565
rect 5204 8515 5236 8516
rect 5204 8485 5205 8515
rect 5205 8485 5235 8515
rect 5235 8485 5236 8515
rect 5204 8484 5236 8485
rect 5204 8435 5236 8436
rect 5204 8405 5205 8435
rect 5205 8405 5235 8435
rect 5235 8405 5236 8435
rect 5204 8404 5236 8405
rect 5204 8324 5236 8356
rect 5204 8275 5236 8276
rect 5204 8245 5205 8275
rect 5205 8245 5235 8275
rect 5235 8245 5236 8275
rect 5204 8244 5236 8245
rect 5204 8195 5236 8196
rect 5204 8165 5205 8195
rect 5205 8165 5235 8195
rect 5235 8165 5236 8195
rect 5204 8164 5236 8165
rect 5204 8115 5236 8116
rect 5204 8085 5205 8115
rect 5205 8085 5235 8115
rect 5235 8085 5236 8115
rect 5204 8084 5236 8085
rect 5204 8035 5236 8036
rect 5204 8005 5205 8035
rect 5205 8005 5235 8035
rect 5235 8005 5236 8035
rect 5204 8004 5236 8005
rect 5204 7955 5236 7956
rect 5204 7925 5205 7955
rect 5205 7925 5235 7955
rect 5235 7925 5236 7955
rect 5204 7924 5236 7925
rect 5204 7875 5236 7876
rect 5204 7845 5205 7875
rect 5205 7845 5235 7875
rect 5235 7845 5236 7875
rect 5204 7844 5236 7845
rect 5204 7795 5236 7796
rect 5204 7765 5205 7795
rect 5205 7765 5235 7795
rect 5235 7765 5236 7795
rect 5204 7764 5236 7765
rect 5204 7715 5236 7716
rect 5204 7685 5205 7715
rect 5205 7685 5235 7715
rect 5235 7685 5236 7715
rect 5204 7684 5236 7685
rect 5204 7635 5236 7636
rect 5204 7605 5205 7635
rect 5205 7605 5235 7635
rect 5235 7605 5236 7635
rect 5204 7604 5236 7605
rect 5204 7555 5236 7556
rect 5204 7525 5205 7555
rect 5205 7525 5235 7555
rect 5235 7525 5236 7555
rect 5204 7524 5236 7525
rect 5204 7475 5236 7476
rect 5204 7445 5205 7475
rect 5205 7445 5235 7475
rect 5235 7445 5236 7475
rect 5204 7444 5236 7445
rect 5204 7395 5236 7396
rect 5204 7365 5205 7395
rect 5205 7365 5235 7395
rect 5235 7365 5236 7395
rect 5204 7364 5236 7365
rect 5204 7315 5236 7316
rect 5204 7285 5205 7315
rect 5205 7285 5235 7315
rect 5235 7285 5236 7315
rect 5204 7284 5236 7285
rect 5204 7235 5236 7236
rect 5204 7205 5205 7235
rect 5205 7205 5235 7235
rect 5235 7205 5236 7235
rect 5204 7204 5236 7205
rect 5204 7155 5236 7156
rect 5204 7125 5205 7155
rect 5205 7125 5235 7155
rect 5235 7125 5236 7155
rect 5204 7124 5236 7125
rect 5204 7075 5236 7076
rect 5204 7045 5205 7075
rect 5205 7045 5235 7075
rect 5235 7045 5236 7075
rect 5204 7044 5236 7045
rect 5204 6995 5236 6996
rect 5204 6965 5205 6995
rect 5205 6965 5235 6995
rect 5235 6965 5236 6995
rect 5204 6964 5236 6965
rect 5204 6884 5236 6916
rect 5204 6835 5236 6836
rect 5204 6805 5205 6835
rect 5205 6805 5235 6835
rect 5235 6805 5236 6835
rect 5204 6804 5236 6805
rect 5204 6755 5236 6756
rect 5204 6725 5205 6755
rect 5205 6725 5235 6755
rect 5235 6725 5236 6755
rect 5204 6724 5236 6725
rect 5204 6675 5236 6676
rect 5204 6645 5205 6675
rect 5205 6645 5235 6675
rect 5235 6645 5236 6675
rect 5204 6644 5236 6645
rect 5204 6595 5236 6596
rect 5204 6565 5205 6595
rect 5205 6565 5235 6595
rect 5235 6565 5236 6595
rect 5204 6564 5236 6565
rect 5204 6515 5236 6516
rect 5204 6485 5205 6515
rect 5205 6485 5235 6515
rect 5235 6485 5236 6515
rect 5204 6484 5236 6485
rect 5204 6435 5236 6436
rect 5204 6405 5205 6435
rect 5205 6405 5235 6435
rect 5235 6405 5236 6435
rect 5204 6404 5236 6405
rect 5204 6355 5236 6356
rect 5204 6325 5205 6355
rect 5205 6325 5235 6355
rect 5235 6325 5236 6355
rect 5204 6324 5236 6325
rect 5204 6275 5236 6276
rect 5204 6245 5205 6275
rect 5205 6245 5235 6275
rect 5235 6245 5236 6275
rect 5204 6244 5236 6245
rect 5204 6164 5236 6196
rect 5204 6084 5236 6116
rect 5204 6004 5236 6036
rect 5204 5924 5236 5956
rect 5204 5875 5236 5876
rect 5204 5845 5205 5875
rect 5205 5845 5235 5875
rect 5235 5845 5236 5875
rect 5204 5844 5236 5845
rect 5204 5795 5236 5796
rect 5204 5765 5205 5795
rect 5205 5765 5235 5795
rect 5235 5765 5236 5795
rect 5204 5764 5236 5765
rect 5204 5715 5236 5716
rect 5204 5685 5205 5715
rect 5205 5685 5235 5715
rect 5235 5685 5236 5715
rect 5204 5684 5236 5685
rect 5204 5635 5236 5636
rect 5204 5605 5205 5635
rect 5205 5605 5235 5635
rect 5235 5605 5236 5635
rect 5204 5604 5236 5605
rect 5204 5555 5236 5556
rect 5204 5525 5205 5555
rect 5205 5525 5235 5555
rect 5235 5525 5236 5555
rect 5204 5524 5236 5525
rect 5204 5475 5236 5476
rect 5204 5445 5205 5475
rect 5205 5445 5235 5475
rect 5235 5445 5236 5475
rect 5204 5444 5236 5445
rect 5204 5395 5236 5396
rect 5204 5365 5205 5395
rect 5205 5365 5235 5395
rect 5235 5365 5236 5395
rect 5204 5364 5236 5365
rect 5204 5315 5236 5316
rect 5204 5285 5205 5315
rect 5205 5285 5235 5315
rect 5235 5285 5236 5315
rect 5204 5284 5236 5285
rect 5204 5235 5236 5236
rect 5204 5205 5205 5235
rect 5205 5205 5235 5235
rect 5235 5205 5236 5235
rect 5204 5204 5236 5205
rect 5204 5155 5236 5156
rect 5204 5125 5205 5155
rect 5205 5125 5235 5155
rect 5235 5125 5236 5155
rect 5204 5124 5236 5125
rect 5204 5075 5236 5076
rect 5204 5045 5205 5075
rect 5205 5045 5235 5075
rect 5235 5045 5236 5075
rect 5204 5044 5236 5045
rect 5204 4995 5236 4996
rect 5204 4965 5205 4995
rect 5205 4965 5235 4995
rect 5235 4965 5236 4995
rect 5204 4964 5236 4965
rect 5204 4915 5236 4916
rect 5204 4885 5205 4915
rect 5205 4885 5235 4915
rect 5235 4885 5236 4915
rect 5204 4884 5236 4885
rect 5204 4804 5236 4836
rect 5204 4755 5236 4756
rect 5204 4725 5205 4755
rect 5205 4725 5235 4755
rect 5235 4725 5236 4755
rect 5204 4724 5236 4725
rect 5204 4675 5236 4676
rect 5204 4645 5205 4675
rect 5205 4645 5235 4675
rect 5235 4645 5236 4675
rect 5204 4644 5236 4645
rect 5204 4564 5236 4596
rect 5204 4515 5236 4516
rect 5204 4485 5205 4515
rect 5205 4485 5235 4515
rect 5235 4485 5236 4515
rect 5204 4484 5236 4485
rect 5204 4435 5236 4436
rect 5204 4405 5205 4435
rect 5205 4405 5235 4435
rect 5235 4405 5236 4435
rect 5204 4404 5236 4405
rect 5204 4355 5236 4356
rect 5204 4325 5205 4355
rect 5205 4325 5235 4355
rect 5235 4325 5236 4355
rect 5204 4324 5236 4325
rect 5204 4275 5236 4276
rect 5204 4245 5205 4275
rect 5205 4245 5235 4275
rect 5235 4245 5236 4275
rect 5204 4244 5236 4245
rect 5204 4195 5236 4196
rect 5204 4165 5205 4195
rect 5205 4165 5235 4195
rect 5235 4165 5236 4195
rect 5204 4164 5236 4165
rect 5204 4115 5236 4116
rect 5204 4085 5205 4115
rect 5205 4085 5235 4115
rect 5235 4085 5236 4115
rect 5204 4084 5236 4085
rect 5204 4035 5236 4036
rect 5204 4005 5205 4035
rect 5205 4005 5235 4035
rect 5235 4005 5236 4035
rect 5204 4004 5236 4005
rect 5204 3955 5236 3956
rect 5204 3925 5205 3955
rect 5205 3925 5235 3955
rect 5235 3925 5236 3955
rect 5204 3924 5236 3925
rect 5204 3875 5236 3876
rect 5204 3845 5205 3875
rect 5205 3845 5235 3875
rect 5235 3845 5236 3875
rect 5204 3844 5236 3845
rect 5204 3764 5236 3796
rect 5204 3715 5236 3716
rect 5204 3685 5205 3715
rect 5205 3685 5235 3715
rect 5235 3685 5236 3715
rect 5204 3684 5236 3685
rect 5204 3635 5236 3636
rect 5204 3605 5205 3635
rect 5205 3605 5235 3635
rect 5235 3605 5236 3635
rect 5204 3604 5236 3605
rect 5204 3524 5236 3556
rect 5204 3475 5236 3476
rect 5204 3445 5205 3475
rect 5205 3445 5235 3475
rect 5235 3445 5236 3475
rect 5204 3444 5236 3445
rect 5204 3395 5236 3396
rect 5204 3365 5205 3395
rect 5205 3365 5235 3395
rect 5235 3365 5236 3395
rect 5204 3364 5236 3365
rect 5204 3284 5236 3316
rect 5204 3235 5236 3236
rect 5204 3205 5205 3235
rect 5205 3205 5235 3235
rect 5235 3205 5236 3235
rect 5204 3204 5236 3205
rect 5204 3155 5236 3156
rect 5204 3125 5205 3155
rect 5205 3125 5235 3155
rect 5235 3125 5236 3155
rect 5204 3124 5236 3125
rect 5204 3075 5236 3076
rect 5204 3045 5205 3075
rect 5205 3045 5235 3075
rect 5235 3045 5236 3075
rect 5204 3044 5236 3045
rect 5204 2995 5236 2996
rect 5204 2965 5205 2995
rect 5205 2965 5235 2995
rect 5235 2965 5236 2995
rect 5204 2964 5236 2965
rect 5204 2915 5236 2916
rect 5204 2885 5205 2915
rect 5205 2885 5235 2915
rect 5235 2885 5236 2915
rect 5204 2884 5236 2885
rect 5204 2835 5236 2836
rect 5204 2805 5205 2835
rect 5205 2805 5235 2835
rect 5235 2805 5236 2835
rect 5204 2804 5236 2805
rect 5204 2755 5236 2756
rect 5204 2725 5205 2755
rect 5205 2725 5235 2755
rect 5235 2725 5236 2755
rect 5204 2724 5236 2725
rect 5204 2675 5236 2676
rect 5204 2645 5205 2675
rect 5205 2645 5235 2675
rect 5235 2645 5236 2675
rect 5204 2644 5236 2645
rect 5204 2595 5236 2596
rect 5204 2565 5205 2595
rect 5205 2565 5235 2595
rect 5235 2565 5236 2595
rect 5204 2564 5236 2565
rect 5204 2515 5236 2516
rect 5204 2485 5205 2515
rect 5205 2485 5235 2515
rect 5235 2485 5236 2515
rect 5204 2484 5236 2485
rect 5204 2435 5236 2436
rect 5204 2405 5205 2435
rect 5205 2405 5235 2435
rect 5235 2405 5236 2435
rect 5204 2404 5236 2405
rect 5204 2355 5236 2356
rect 5204 2325 5205 2355
rect 5205 2325 5235 2355
rect 5235 2325 5236 2355
rect 5204 2324 5236 2325
rect 5204 2275 5236 2276
rect 5204 2245 5205 2275
rect 5205 2245 5235 2275
rect 5235 2245 5236 2275
rect 5204 2244 5236 2245
rect 5204 2195 5236 2196
rect 5204 2165 5205 2195
rect 5205 2165 5235 2195
rect 5235 2165 5236 2195
rect 5204 2164 5236 2165
rect 5204 2115 5236 2116
rect 5204 2085 5205 2115
rect 5205 2085 5235 2115
rect 5235 2085 5236 2115
rect 5204 2084 5236 2085
rect 5204 2035 5236 2036
rect 5204 2005 5205 2035
rect 5205 2005 5235 2035
rect 5235 2005 5236 2035
rect 5204 2004 5236 2005
rect 5204 1955 5236 1956
rect 5204 1925 5205 1955
rect 5205 1925 5235 1955
rect 5235 1925 5236 1955
rect 5204 1924 5236 1925
rect 5204 1844 5236 1876
rect 5204 1764 5236 1796
rect 5204 1715 5236 1716
rect 5204 1685 5205 1715
rect 5205 1685 5235 1715
rect 5235 1685 5236 1715
rect 5204 1684 5236 1685
rect 5204 1635 5236 1636
rect 5204 1605 5205 1635
rect 5205 1605 5235 1635
rect 5235 1605 5236 1635
rect 5204 1604 5236 1605
rect 5204 1555 5236 1556
rect 5204 1525 5205 1555
rect 5205 1525 5235 1555
rect 5235 1525 5236 1555
rect 5204 1524 5236 1525
rect 5204 1475 5236 1476
rect 5204 1445 5205 1475
rect 5205 1445 5235 1475
rect 5235 1445 5236 1475
rect 5204 1444 5236 1445
rect 5204 1395 5236 1396
rect 5204 1365 5205 1395
rect 5205 1365 5235 1395
rect 5235 1365 5236 1395
rect 5204 1364 5236 1365
rect 5204 1315 5236 1316
rect 5204 1285 5205 1315
rect 5205 1285 5235 1315
rect 5235 1285 5236 1315
rect 5204 1284 5236 1285
rect 5204 1235 5236 1236
rect 5204 1205 5205 1235
rect 5205 1205 5235 1235
rect 5235 1205 5236 1235
rect 5204 1204 5236 1205
rect 5204 1155 5236 1156
rect 5204 1125 5205 1155
rect 5205 1125 5235 1155
rect 5235 1125 5236 1155
rect 5204 1124 5236 1125
rect 5204 1075 5236 1076
rect 5204 1045 5205 1075
rect 5205 1045 5235 1075
rect 5235 1045 5236 1075
rect 5204 1044 5236 1045
rect 5204 995 5236 996
rect 5204 965 5205 995
rect 5205 965 5235 995
rect 5235 965 5236 995
rect 5204 964 5236 965
rect 5204 884 5236 916
rect 5204 835 5236 836
rect 5204 805 5205 835
rect 5205 805 5235 835
rect 5235 805 5236 835
rect 5204 804 5236 805
rect 5204 755 5236 756
rect 5204 725 5205 755
rect 5205 725 5235 755
rect 5235 725 5236 755
rect 5204 724 5236 725
rect 5204 675 5236 676
rect 5204 645 5205 675
rect 5205 645 5235 675
rect 5235 645 5236 675
rect 5204 644 5236 645
rect 5204 595 5236 596
rect 5204 565 5205 595
rect 5205 565 5235 595
rect 5235 565 5236 595
rect 5204 564 5236 565
rect 5204 515 5236 516
rect 5204 485 5205 515
rect 5205 485 5235 515
rect 5235 485 5236 515
rect 5204 484 5236 485
rect 5204 404 5236 436
rect 5204 324 5236 356
rect 5204 275 5236 276
rect 5204 245 5205 275
rect 5205 245 5235 275
rect 5235 245 5236 275
rect 5204 244 5236 245
rect 5204 195 5236 196
rect 5204 165 5205 195
rect 5205 165 5235 195
rect 5235 165 5236 195
rect 5204 164 5236 165
rect 5204 115 5236 116
rect 5204 85 5205 115
rect 5205 85 5235 115
rect 5235 85 5236 115
rect 5204 84 5236 85
rect 5204 35 5236 36
rect 5204 5 5205 35
rect 5205 5 5235 35
rect 5235 5 5236 35
rect 5204 4 5236 5
rect 5044 -716 5076 -524
rect 5364 15715 5396 15716
rect 5364 15685 5365 15715
rect 5365 15685 5395 15715
rect 5395 15685 5396 15715
rect 5364 15684 5396 15685
rect 5364 15635 5396 15636
rect 5364 15605 5365 15635
rect 5365 15605 5395 15635
rect 5395 15605 5396 15635
rect 5364 15604 5396 15605
rect 5364 15555 5396 15556
rect 5364 15525 5365 15555
rect 5365 15525 5395 15555
rect 5395 15525 5396 15555
rect 5364 15524 5396 15525
rect 5364 15475 5396 15476
rect 5364 15445 5365 15475
rect 5365 15445 5395 15475
rect 5395 15445 5396 15475
rect 5364 15444 5396 15445
rect 5364 15395 5396 15396
rect 5364 15365 5365 15395
rect 5365 15365 5395 15395
rect 5395 15365 5396 15395
rect 5364 15364 5396 15365
rect 5364 15315 5396 15316
rect 5364 15285 5365 15315
rect 5365 15285 5395 15315
rect 5395 15285 5396 15315
rect 5364 15284 5396 15285
rect 5364 15235 5396 15236
rect 5364 15205 5365 15235
rect 5365 15205 5395 15235
rect 5395 15205 5396 15235
rect 5364 15204 5396 15205
rect 5364 15155 5396 15156
rect 5364 15125 5365 15155
rect 5365 15125 5395 15155
rect 5395 15125 5396 15155
rect 5364 15124 5396 15125
rect 5364 15044 5396 15076
rect 5364 14995 5396 14996
rect 5364 14965 5365 14995
rect 5365 14965 5395 14995
rect 5395 14965 5396 14995
rect 5364 14964 5396 14965
rect 5364 14915 5396 14916
rect 5364 14885 5365 14915
rect 5365 14885 5395 14915
rect 5395 14885 5396 14915
rect 5364 14884 5396 14885
rect 5364 14835 5396 14836
rect 5364 14805 5365 14835
rect 5365 14805 5395 14835
rect 5395 14805 5396 14835
rect 5364 14804 5396 14805
rect 5364 14755 5396 14756
rect 5364 14725 5365 14755
rect 5365 14725 5395 14755
rect 5395 14725 5396 14755
rect 5364 14724 5396 14725
rect 5364 14675 5396 14676
rect 5364 14645 5365 14675
rect 5365 14645 5395 14675
rect 5395 14645 5396 14675
rect 5364 14644 5396 14645
rect 5364 14595 5396 14596
rect 5364 14565 5365 14595
rect 5365 14565 5395 14595
rect 5395 14565 5396 14595
rect 5364 14564 5396 14565
rect 5364 14515 5396 14516
rect 5364 14485 5365 14515
rect 5365 14485 5395 14515
rect 5395 14485 5396 14515
rect 5364 14484 5396 14485
rect 5364 14435 5396 14436
rect 5364 14405 5365 14435
rect 5365 14405 5395 14435
rect 5395 14405 5396 14435
rect 5364 14404 5396 14405
rect 5364 14324 5396 14356
rect 5364 14244 5396 14276
rect 5364 14164 5396 14196
rect 5364 14084 5396 14116
rect 5364 14035 5396 14036
rect 5364 14005 5365 14035
rect 5365 14005 5395 14035
rect 5395 14005 5396 14035
rect 5364 14004 5396 14005
rect 5364 13955 5396 13956
rect 5364 13925 5365 13955
rect 5365 13925 5395 13955
rect 5395 13925 5396 13955
rect 5364 13924 5396 13925
rect 5364 13875 5396 13876
rect 5364 13845 5365 13875
rect 5365 13845 5395 13875
rect 5395 13845 5396 13875
rect 5364 13844 5396 13845
rect 5364 13795 5396 13796
rect 5364 13765 5365 13795
rect 5365 13765 5395 13795
rect 5395 13765 5396 13795
rect 5364 13764 5396 13765
rect 5364 13715 5396 13716
rect 5364 13685 5365 13715
rect 5365 13685 5395 13715
rect 5395 13685 5396 13715
rect 5364 13684 5396 13685
rect 5364 13635 5396 13636
rect 5364 13605 5365 13635
rect 5365 13605 5395 13635
rect 5395 13605 5396 13635
rect 5364 13604 5396 13605
rect 5364 13555 5396 13556
rect 5364 13525 5365 13555
rect 5365 13525 5395 13555
rect 5395 13525 5396 13555
rect 5364 13524 5396 13525
rect 5364 13475 5396 13476
rect 5364 13445 5365 13475
rect 5365 13445 5395 13475
rect 5395 13445 5396 13475
rect 5364 13444 5396 13445
rect 5364 13364 5396 13396
rect 5364 13284 5396 13316
rect 5364 13204 5396 13236
rect 5364 13124 5396 13156
rect 5364 13075 5396 13076
rect 5364 13045 5365 13075
rect 5365 13045 5395 13075
rect 5395 13045 5396 13075
rect 5364 13044 5396 13045
rect 5364 12995 5396 12996
rect 5364 12965 5365 12995
rect 5365 12965 5395 12995
rect 5395 12965 5396 12995
rect 5364 12964 5396 12965
rect 5364 12915 5396 12916
rect 5364 12885 5365 12915
rect 5365 12885 5395 12915
rect 5395 12885 5396 12915
rect 5364 12884 5396 12885
rect 5364 12835 5396 12836
rect 5364 12805 5365 12835
rect 5365 12805 5395 12835
rect 5395 12805 5396 12835
rect 5364 12804 5396 12805
rect 5364 12755 5396 12756
rect 5364 12725 5365 12755
rect 5365 12725 5395 12755
rect 5395 12725 5396 12755
rect 5364 12724 5396 12725
rect 5364 12675 5396 12676
rect 5364 12645 5365 12675
rect 5365 12645 5395 12675
rect 5395 12645 5396 12675
rect 5364 12644 5396 12645
rect 5364 12595 5396 12596
rect 5364 12565 5365 12595
rect 5365 12565 5395 12595
rect 5395 12565 5396 12595
rect 5364 12564 5396 12565
rect 5364 12515 5396 12516
rect 5364 12485 5365 12515
rect 5365 12485 5395 12515
rect 5395 12485 5396 12515
rect 5364 12484 5396 12485
rect 5364 12404 5396 12436
rect 5364 12355 5396 12356
rect 5364 12325 5365 12355
rect 5365 12325 5395 12355
rect 5395 12325 5396 12355
rect 5364 12324 5396 12325
rect 5364 12275 5396 12276
rect 5364 12245 5365 12275
rect 5365 12245 5395 12275
rect 5395 12245 5396 12275
rect 5364 12244 5396 12245
rect 5364 12195 5396 12196
rect 5364 12165 5365 12195
rect 5365 12165 5395 12195
rect 5395 12165 5396 12195
rect 5364 12164 5396 12165
rect 5364 12115 5396 12116
rect 5364 12085 5365 12115
rect 5365 12085 5395 12115
rect 5395 12085 5396 12115
rect 5364 12084 5396 12085
rect 5364 12035 5396 12036
rect 5364 12005 5365 12035
rect 5365 12005 5395 12035
rect 5395 12005 5396 12035
rect 5364 12004 5396 12005
rect 5364 11955 5396 11956
rect 5364 11925 5365 11955
rect 5365 11925 5395 11955
rect 5395 11925 5396 11955
rect 5364 11924 5396 11925
rect 5364 11875 5396 11876
rect 5364 11845 5365 11875
rect 5365 11845 5395 11875
rect 5395 11845 5396 11875
rect 5364 11844 5396 11845
rect 5364 11795 5396 11796
rect 5364 11765 5365 11795
rect 5365 11765 5395 11795
rect 5395 11765 5396 11795
rect 5364 11764 5396 11765
rect 5364 11715 5396 11716
rect 5364 11685 5365 11715
rect 5365 11685 5395 11715
rect 5395 11685 5396 11715
rect 5364 11684 5396 11685
rect 5364 11635 5396 11636
rect 5364 11605 5365 11635
rect 5365 11605 5395 11635
rect 5395 11605 5396 11635
rect 5364 11604 5396 11605
rect 5364 11555 5396 11556
rect 5364 11525 5365 11555
rect 5365 11525 5395 11555
rect 5395 11525 5396 11555
rect 5364 11524 5396 11525
rect 5364 11475 5396 11476
rect 5364 11445 5365 11475
rect 5365 11445 5395 11475
rect 5395 11445 5396 11475
rect 5364 11444 5396 11445
rect 5364 11395 5396 11396
rect 5364 11365 5365 11395
rect 5365 11365 5395 11395
rect 5395 11365 5396 11395
rect 5364 11364 5396 11365
rect 5364 11315 5396 11316
rect 5364 11285 5365 11315
rect 5365 11285 5395 11315
rect 5395 11285 5396 11315
rect 5364 11284 5396 11285
rect 5364 11235 5396 11236
rect 5364 11205 5365 11235
rect 5365 11205 5395 11235
rect 5395 11205 5396 11235
rect 5364 11204 5396 11205
rect 5364 11155 5396 11156
rect 5364 11125 5365 11155
rect 5365 11125 5395 11155
rect 5395 11125 5396 11155
rect 5364 11124 5396 11125
rect 5364 11075 5396 11076
rect 5364 11045 5365 11075
rect 5365 11045 5395 11075
rect 5395 11045 5396 11075
rect 5364 11044 5396 11045
rect 5364 10964 5396 10996
rect 5364 10915 5396 10916
rect 5364 10885 5365 10915
rect 5365 10885 5395 10915
rect 5395 10885 5396 10915
rect 5364 10884 5396 10885
rect 5364 10835 5396 10836
rect 5364 10805 5365 10835
rect 5365 10805 5395 10835
rect 5395 10805 5396 10835
rect 5364 10804 5396 10805
rect 5364 10755 5396 10756
rect 5364 10725 5365 10755
rect 5365 10725 5395 10755
rect 5395 10725 5396 10755
rect 5364 10724 5396 10725
rect 5364 10675 5396 10676
rect 5364 10645 5365 10675
rect 5365 10645 5395 10675
rect 5395 10645 5396 10675
rect 5364 10644 5396 10645
rect 5364 10595 5396 10596
rect 5364 10565 5365 10595
rect 5365 10565 5395 10595
rect 5395 10565 5396 10595
rect 5364 10564 5396 10565
rect 5364 10515 5396 10516
rect 5364 10485 5365 10515
rect 5365 10485 5395 10515
rect 5395 10485 5396 10515
rect 5364 10484 5396 10485
rect 5364 10435 5396 10436
rect 5364 10405 5365 10435
rect 5365 10405 5395 10435
rect 5395 10405 5396 10435
rect 5364 10404 5396 10405
rect 5364 10355 5396 10356
rect 5364 10325 5365 10355
rect 5365 10325 5395 10355
rect 5395 10325 5396 10355
rect 5364 10324 5396 10325
rect 5364 10244 5396 10276
rect 5364 10164 5396 10196
rect 5364 10084 5396 10116
rect 5364 10004 5396 10036
rect 5364 9955 5396 9956
rect 5364 9925 5365 9955
rect 5365 9925 5395 9955
rect 5395 9925 5396 9955
rect 5364 9924 5396 9925
rect 5364 9875 5396 9876
rect 5364 9845 5365 9875
rect 5365 9845 5395 9875
rect 5395 9845 5396 9875
rect 5364 9844 5396 9845
rect 5364 9795 5396 9796
rect 5364 9765 5365 9795
rect 5365 9765 5395 9795
rect 5395 9765 5396 9795
rect 5364 9764 5396 9765
rect 5364 9715 5396 9716
rect 5364 9685 5365 9715
rect 5365 9685 5395 9715
rect 5395 9685 5396 9715
rect 5364 9684 5396 9685
rect 5364 9635 5396 9636
rect 5364 9605 5365 9635
rect 5365 9605 5395 9635
rect 5395 9605 5396 9635
rect 5364 9604 5396 9605
rect 5364 9555 5396 9556
rect 5364 9525 5365 9555
rect 5365 9525 5395 9555
rect 5395 9525 5396 9555
rect 5364 9524 5396 9525
rect 5364 9475 5396 9476
rect 5364 9445 5365 9475
rect 5365 9445 5395 9475
rect 5395 9445 5396 9475
rect 5364 9444 5396 9445
rect 5364 9395 5396 9396
rect 5364 9365 5365 9395
rect 5365 9365 5395 9395
rect 5395 9365 5396 9395
rect 5364 9364 5396 9365
rect 5364 9284 5396 9316
rect 5364 9204 5396 9236
rect 5364 9124 5396 9156
rect 5364 9044 5396 9076
rect 5364 8995 5396 8996
rect 5364 8965 5365 8995
rect 5365 8965 5395 8995
rect 5395 8965 5396 8995
rect 5364 8964 5396 8965
rect 5364 8915 5396 8916
rect 5364 8885 5365 8915
rect 5365 8885 5395 8915
rect 5395 8885 5396 8915
rect 5364 8884 5396 8885
rect 5364 8835 5396 8836
rect 5364 8805 5365 8835
rect 5365 8805 5395 8835
rect 5395 8805 5396 8835
rect 5364 8804 5396 8805
rect 5364 8755 5396 8756
rect 5364 8725 5365 8755
rect 5365 8725 5395 8755
rect 5395 8725 5396 8755
rect 5364 8724 5396 8725
rect 5364 8675 5396 8676
rect 5364 8645 5365 8675
rect 5365 8645 5395 8675
rect 5395 8645 5396 8675
rect 5364 8644 5396 8645
rect 5364 8595 5396 8596
rect 5364 8565 5365 8595
rect 5365 8565 5395 8595
rect 5395 8565 5396 8595
rect 5364 8564 5396 8565
rect 5364 8515 5396 8516
rect 5364 8485 5365 8515
rect 5365 8485 5395 8515
rect 5395 8485 5396 8515
rect 5364 8484 5396 8485
rect 5364 8435 5396 8436
rect 5364 8405 5365 8435
rect 5365 8405 5395 8435
rect 5395 8405 5396 8435
rect 5364 8404 5396 8405
rect 5364 8324 5396 8356
rect 5364 8275 5396 8276
rect 5364 8245 5365 8275
rect 5365 8245 5395 8275
rect 5395 8245 5396 8275
rect 5364 8244 5396 8245
rect 5364 8195 5396 8196
rect 5364 8165 5365 8195
rect 5365 8165 5395 8195
rect 5395 8165 5396 8195
rect 5364 8164 5396 8165
rect 5364 8115 5396 8116
rect 5364 8085 5365 8115
rect 5365 8085 5395 8115
rect 5395 8085 5396 8115
rect 5364 8084 5396 8085
rect 5364 8035 5396 8036
rect 5364 8005 5365 8035
rect 5365 8005 5395 8035
rect 5395 8005 5396 8035
rect 5364 8004 5396 8005
rect 5364 7955 5396 7956
rect 5364 7925 5365 7955
rect 5365 7925 5395 7955
rect 5395 7925 5396 7955
rect 5364 7924 5396 7925
rect 5364 7875 5396 7876
rect 5364 7845 5365 7875
rect 5365 7845 5395 7875
rect 5395 7845 5396 7875
rect 5364 7844 5396 7845
rect 5364 7795 5396 7796
rect 5364 7765 5365 7795
rect 5365 7765 5395 7795
rect 5395 7765 5396 7795
rect 5364 7764 5396 7765
rect 5364 7715 5396 7716
rect 5364 7685 5365 7715
rect 5365 7685 5395 7715
rect 5395 7685 5396 7715
rect 5364 7684 5396 7685
rect 5364 7635 5396 7636
rect 5364 7605 5365 7635
rect 5365 7605 5395 7635
rect 5395 7605 5396 7635
rect 5364 7604 5396 7605
rect 5364 7555 5396 7556
rect 5364 7525 5365 7555
rect 5365 7525 5395 7555
rect 5395 7525 5396 7555
rect 5364 7524 5396 7525
rect 5364 7475 5396 7476
rect 5364 7445 5365 7475
rect 5365 7445 5395 7475
rect 5395 7445 5396 7475
rect 5364 7444 5396 7445
rect 5364 7395 5396 7396
rect 5364 7365 5365 7395
rect 5365 7365 5395 7395
rect 5395 7365 5396 7395
rect 5364 7364 5396 7365
rect 5364 7315 5396 7316
rect 5364 7285 5365 7315
rect 5365 7285 5395 7315
rect 5395 7285 5396 7315
rect 5364 7284 5396 7285
rect 5364 7235 5396 7236
rect 5364 7205 5365 7235
rect 5365 7205 5395 7235
rect 5395 7205 5396 7235
rect 5364 7204 5396 7205
rect 5364 7155 5396 7156
rect 5364 7125 5365 7155
rect 5365 7125 5395 7155
rect 5395 7125 5396 7155
rect 5364 7124 5396 7125
rect 5364 7075 5396 7076
rect 5364 7045 5365 7075
rect 5365 7045 5395 7075
rect 5395 7045 5396 7075
rect 5364 7044 5396 7045
rect 5364 6995 5396 6996
rect 5364 6965 5365 6995
rect 5365 6965 5395 6995
rect 5395 6965 5396 6995
rect 5364 6964 5396 6965
rect 5364 6884 5396 6916
rect 5364 6835 5396 6836
rect 5364 6805 5365 6835
rect 5365 6805 5395 6835
rect 5395 6805 5396 6835
rect 5364 6804 5396 6805
rect 5364 6755 5396 6756
rect 5364 6725 5365 6755
rect 5365 6725 5395 6755
rect 5395 6725 5396 6755
rect 5364 6724 5396 6725
rect 5364 6675 5396 6676
rect 5364 6645 5365 6675
rect 5365 6645 5395 6675
rect 5395 6645 5396 6675
rect 5364 6644 5396 6645
rect 5364 6595 5396 6596
rect 5364 6565 5365 6595
rect 5365 6565 5395 6595
rect 5395 6565 5396 6595
rect 5364 6564 5396 6565
rect 5364 6515 5396 6516
rect 5364 6485 5365 6515
rect 5365 6485 5395 6515
rect 5395 6485 5396 6515
rect 5364 6484 5396 6485
rect 5364 6435 5396 6436
rect 5364 6405 5365 6435
rect 5365 6405 5395 6435
rect 5395 6405 5396 6435
rect 5364 6404 5396 6405
rect 5364 6355 5396 6356
rect 5364 6325 5365 6355
rect 5365 6325 5395 6355
rect 5395 6325 5396 6355
rect 5364 6324 5396 6325
rect 5364 6275 5396 6276
rect 5364 6245 5365 6275
rect 5365 6245 5395 6275
rect 5395 6245 5396 6275
rect 5364 6244 5396 6245
rect 5364 6164 5396 6196
rect 5364 6084 5396 6116
rect 5364 6004 5396 6036
rect 5364 5924 5396 5956
rect 5364 5875 5396 5876
rect 5364 5845 5365 5875
rect 5365 5845 5395 5875
rect 5395 5845 5396 5875
rect 5364 5844 5396 5845
rect 5364 5795 5396 5796
rect 5364 5765 5365 5795
rect 5365 5765 5395 5795
rect 5395 5765 5396 5795
rect 5364 5764 5396 5765
rect 5364 5715 5396 5716
rect 5364 5685 5365 5715
rect 5365 5685 5395 5715
rect 5395 5685 5396 5715
rect 5364 5684 5396 5685
rect 5364 5635 5396 5636
rect 5364 5605 5365 5635
rect 5365 5605 5395 5635
rect 5395 5605 5396 5635
rect 5364 5604 5396 5605
rect 5364 5555 5396 5556
rect 5364 5525 5365 5555
rect 5365 5525 5395 5555
rect 5395 5525 5396 5555
rect 5364 5524 5396 5525
rect 5364 5475 5396 5476
rect 5364 5445 5365 5475
rect 5365 5445 5395 5475
rect 5395 5445 5396 5475
rect 5364 5444 5396 5445
rect 5364 5395 5396 5396
rect 5364 5365 5365 5395
rect 5365 5365 5395 5395
rect 5395 5365 5396 5395
rect 5364 5364 5396 5365
rect 5364 5315 5396 5316
rect 5364 5285 5365 5315
rect 5365 5285 5395 5315
rect 5395 5285 5396 5315
rect 5364 5284 5396 5285
rect 5364 5235 5396 5236
rect 5364 5205 5365 5235
rect 5365 5205 5395 5235
rect 5395 5205 5396 5235
rect 5364 5204 5396 5205
rect 5364 5155 5396 5156
rect 5364 5125 5365 5155
rect 5365 5125 5395 5155
rect 5395 5125 5396 5155
rect 5364 5124 5396 5125
rect 5364 5075 5396 5076
rect 5364 5045 5365 5075
rect 5365 5045 5395 5075
rect 5395 5045 5396 5075
rect 5364 5044 5396 5045
rect 5364 4995 5396 4996
rect 5364 4965 5365 4995
rect 5365 4965 5395 4995
rect 5395 4965 5396 4995
rect 5364 4964 5396 4965
rect 5364 4915 5396 4916
rect 5364 4885 5365 4915
rect 5365 4885 5395 4915
rect 5395 4885 5396 4915
rect 5364 4884 5396 4885
rect 5364 4804 5396 4836
rect 5364 4755 5396 4756
rect 5364 4725 5365 4755
rect 5365 4725 5395 4755
rect 5395 4725 5396 4755
rect 5364 4724 5396 4725
rect 5364 4675 5396 4676
rect 5364 4645 5365 4675
rect 5365 4645 5395 4675
rect 5395 4645 5396 4675
rect 5364 4644 5396 4645
rect 5364 4564 5396 4596
rect 5364 4515 5396 4516
rect 5364 4485 5365 4515
rect 5365 4485 5395 4515
rect 5395 4485 5396 4515
rect 5364 4484 5396 4485
rect 5364 4435 5396 4436
rect 5364 4405 5365 4435
rect 5365 4405 5395 4435
rect 5395 4405 5396 4435
rect 5364 4404 5396 4405
rect 5364 4355 5396 4356
rect 5364 4325 5365 4355
rect 5365 4325 5395 4355
rect 5395 4325 5396 4355
rect 5364 4324 5396 4325
rect 5364 4275 5396 4276
rect 5364 4245 5365 4275
rect 5365 4245 5395 4275
rect 5395 4245 5396 4275
rect 5364 4244 5396 4245
rect 5364 4195 5396 4196
rect 5364 4165 5365 4195
rect 5365 4165 5395 4195
rect 5395 4165 5396 4195
rect 5364 4164 5396 4165
rect 5364 4115 5396 4116
rect 5364 4085 5365 4115
rect 5365 4085 5395 4115
rect 5395 4085 5396 4115
rect 5364 4084 5396 4085
rect 5364 4035 5396 4036
rect 5364 4005 5365 4035
rect 5365 4005 5395 4035
rect 5395 4005 5396 4035
rect 5364 4004 5396 4005
rect 5364 3955 5396 3956
rect 5364 3925 5365 3955
rect 5365 3925 5395 3955
rect 5395 3925 5396 3955
rect 5364 3924 5396 3925
rect 5364 3875 5396 3876
rect 5364 3845 5365 3875
rect 5365 3845 5395 3875
rect 5395 3845 5396 3875
rect 5364 3844 5396 3845
rect 5364 3764 5396 3796
rect 5364 3715 5396 3716
rect 5364 3685 5365 3715
rect 5365 3685 5395 3715
rect 5395 3685 5396 3715
rect 5364 3684 5396 3685
rect 5364 3635 5396 3636
rect 5364 3605 5365 3635
rect 5365 3605 5395 3635
rect 5395 3605 5396 3635
rect 5364 3604 5396 3605
rect 5364 3524 5396 3556
rect 5364 3475 5396 3476
rect 5364 3445 5365 3475
rect 5365 3445 5395 3475
rect 5395 3445 5396 3475
rect 5364 3444 5396 3445
rect 5364 3395 5396 3396
rect 5364 3365 5365 3395
rect 5365 3365 5395 3395
rect 5395 3365 5396 3395
rect 5364 3364 5396 3365
rect 5364 3284 5396 3316
rect 5364 3235 5396 3236
rect 5364 3205 5365 3235
rect 5365 3205 5395 3235
rect 5395 3205 5396 3235
rect 5364 3204 5396 3205
rect 5364 3155 5396 3156
rect 5364 3125 5365 3155
rect 5365 3125 5395 3155
rect 5395 3125 5396 3155
rect 5364 3124 5396 3125
rect 5364 3075 5396 3076
rect 5364 3045 5365 3075
rect 5365 3045 5395 3075
rect 5395 3045 5396 3075
rect 5364 3044 5396 3045
rect 5364 2995 5396 2996
rect 5364 2965 5365 2995
rect 5365 2965 5395 2995
rect 5395 2965 5396 2995
rect 5364 2964 5396 2965
rect 5364 2915 5396 2916
rect 5364 2885 5365 2915
rect 5365 2885 5395 2915
rect 5395 2885 5396 2915
rect 5364 2884 5396 2885
rect 5364 2835 5396 2836
rect 5364 2805 5365 2835
rect 5365 2805 5395 2835
rect 5395 2805 5396 2835
rect 5364 2804 5396 2805
rect 5364 2755 5396 2756
rect 5364 2725 5365 2755
rect 5365 2725 5395 2755
rect 5395 2725 5396 2755
rect 5364 2724 5396 2725
rect 5364 2675 5396 2676
rect 5364 2645 5365 2675
rect 5365 2645 5395 2675
rect 5395 2645 5396 2675
rect 5364 2644 5396 2645
rect 5364 2595 5396 2596
rect 5364 2565 5365 2595
rect 5365 2565 5395 2595
rect 5395 2565 5396 2595
rect 5364 2564 5396 2565
rect 5364 2515 5396 2516
rect 5364 2485 5365 2515
rect 5365 2485 5395 2515
rect 5395 2485 5396 2515
rect 5364 2484 5396 2485
rect 5364 2435 5396 2436
rect 5364 2405 5365 2435
rect 5365 2405 5395 2435
rect 5395 2405 5396 2435
rect 5364 2404 5396 2405
rect 5364 2355 5396 2356
rect 5364 2325 5365 2355
rect 5365 2325 5395 2355
rect 5395 2325 5396 2355
rect 5364 2324 5396 2325
rect 5364 2275 5396 2276
rect 5364 2245 5365 2275
rect 5365 2245 5395 2275
rect 5395 2245 5396 2275
rect 5364 2244 5396 2245
rect 5364 2195 5396 2196
rect 5364 2165 5365 2195
rect 5365 2165 5395 2195
rect 5395 2165 5396 2195
rect 5364 2164 5396 2165
rect 5364 2115 5396 2116
rect 5364 2085 5365 2115
rect 5365 2085 5395 2115
rect 5395 2085 5396 2115
rect 5364 2084 5396 2085
rect 5364 2035 5396 2036
rect 5364 2005 5365 2035
rect 5365 2005 5395 2035
rect 5395 2005 5396 2035
rect 5364 2004 5396 2005
rect 5364 1955 5396 1956
rect 5364 1925 5365 1955
rect 5365 1925 5395 1955
rect 5395 1925 5396 1955
rect 5364 1924 5396 1925
rect 5364 1844 5396 1876
rect 5364 1764 5396 1796
rect 5364 1715 5396 1716
rect 5364 1685 5365 1715
rect 5365 1685 5395 1715
rect 5395 1685 5396 1715
rect 5364 1684 5396 1685
rect 5364 1635 5396 1636
rect 5364 1605 5365 1635
rect 5365 1605 5395 1635
rect 5395 1605 5396 1635
rect 5364 1604 5396 1605
rect 5364 1555 5396 1556
rect 5364 1525 5365 1555
rect 5365 1525 5395 1555
rect 5395 1525 5396 1555
rect 5364 1524 5396 1525
rect 5364 1475 5396 1476
rect 5364 1445 5365 1475
rect 5365 1445 5395 1475
rect 5395 1445 5396 1475
rect 5364 1444 5396 1445
rect 5364 1395 5396 1396
rect 5364 1365 5365 1395
rect 5365 1365 5395 1395
rect 5395 1365 5396 1395
rect 5364 1364 5396 1365
rect 5364 1315 5396 1316
rect 5364 1285 5365 1315
rect 5365 1285 5395 1315
rect 5395 1285 5396 1315
rect 5364 1284 5396 1285
rect 5364 1235 5396 1236
rect 5364 1205 5365 1235
rect 5365 1205 5395 1235
rect 5395 1205 5396 1235
rect 5364 1204 5396 1205
rect 5364 1155 5396 1156
rect 5364 1125 5365 1155
rect 5365 1125 5395 1155
rect 5395 1125 5396 1155
rect 5364 1124 5396 1125
rect 5364 1075 5396 1076
rect 5364 1045 5365 1075
rect 5365 1045 5395 1075
rect 5395 1045 5396 1075
rect 5364 1044 5396 1045
rect 5364 995 5396 996
rect 5364 965 5365 995
rect 5365 965 5395 995
rect 5395 965 5396 995
rect 5364 964 5396 965
rect 5364 884 5396 916
rect 5364 835 5396 836
rect 5364 805 5365 835
rect 5365 805 5395 835
rect 5395 805 5396 835
rect 5364 804 5396 805
rect 5364 755 5396 756
rect 5364 725 5365 755
rect 5365 725 5395 755
rect 5395 725 5396 755
rect 5364 724 5396 725
rect 5364 675 5396 676
rect 5364 645 5365 675
rect 5365 645 5395 675
rect 5395 645 5396 675
rect 5364 644 5396 645
rect 5364 595 5396 596
rect 5364 565 5365 595
rect 5365 565 5395 595
rect 5395 565 5396 595
rect 5364 564 5396 565
rect 5364 515 5396 516
rect 5364 485 5365 515
rect 5365 485 5395 515
rect 5395 485 5396 515
rect 5364 484 5396 485
rect 5364 404 5396 436
rect 5364 324 5396 356
rect 5364 275 5396 276
rect 5364 245 5365 275
rect 5365 245 5395 275
rect 5395 245 5396 275
rect 5364 244 5396 245
rect 5364 195 5396 196
rect 5364 165 5365 195
rect 5365 165 5395 195
rect 5395 165 5396 195
rect 5364 164 5396 165
rect 5364 115 5396 116
rect 5364 85 5365 115
rect 5365 85 5395 115
rect 5395 85 5396 115
rect 5364 84 5396 85
rect 5364 35 5396 36
rect 5364 5 5365 35
rect 5365 5 5395 35
rect 5395 5 5396 35
rect 5364 4 5396 5
rect 5204 -716 5236 -524
rect 5524 15715 5556 15716
rect 5524 15685 5525 15715
rect 5525 15685 5555 15715
rect 5555 15685 5556 15715
rect 5524 15684 5556 15685
rect 5524 15635 5556 15636
rect 5524 15605 5525 15635
rect 5525 15605 5555 15635
rect 5555 15605 5556 15635
rect 5524 15604 5556 15605
rect 5524 15555 5556 15556
rect 5524 15525 5525 15555
rect 5525 15525 5555 15555
rect 5555 15525 5556 15555
rect 5524 15524 5556 15525
rect 5524 15475 5556 15476
rect 5524 15445 5525 15475
rect 5525 15445 5555 15475
rect 5555 15445 5556 15475
rect 5524 15444 5556 15445
rect 5524 15395 5556 15396
rect 5524 15365 5525 15395
rect 5525 15365 5555 15395
rect 5555 15365 5556 15395
rect 5524 15364 5556 15365
rect 5524 15315 5556 15316
rect 5524 15285 5525 15315
rect 5525 15285 5555 15315
rect 5555 15285 5556 15315
rect 5524 15284 5556 15285
rect 5524 15235 5556 15236
rect 5524 15205 5525 15235
rect 5525 15205 5555 15235
rect 5555 15205 5556 15235
rect 5524 15204 5556 15205
rect 5524 15155 5556 15156
rect 5524 15125 5525 15155
rect 5525 15125 5555 15155
rect 5555 15125 5556 15155
rect 5524 15124 5556 15125
rect 5524 15044 5556 15076
rect 5524 14995 5556 14996
rect 5524 14965 5525 14995
rect 5525 14965 5555 14995
rect 5555 14965 5556 14995
rect 5524 14964 5556 14965
rect 5524 14915 5556 14916
rect 5524 14885 5525 14915
rect 5525 14885 5555 14915
rect 5555 14885 5556 14915
rect 5524 14884 5556 14885
rect 5524 14835 5556 14836
rect 5524 14805 5525 14835
rect 5525 14805 5555 14835
rect 5555 14805 5556 14835
rect 5524 14804 5556 14805
rect 5524 14755 5556 14756
rect 5524 14725 5525 14755
rect 5525 14725 5555 14755
rect 5555 14725 5556 14755
rect 5524 14724 5556 14725
rect 5524 14675 5556 14676
rect 5524 14645 5525 14675
rect 5525 14645 5555 14675
rect 5555 14645 5556 14675
rect 5524 14644 5556 14645
rect 5524 14595 5556 14596
rect 5524 14565 5525 14595
rect 5525 14565 5555 14595
rect 5555 14565 5556 14595
rect 5524 14564 5556 14565
rect 5524 14515 5556 14516
rect 5524 14485 5525 14515
rect 5525 14485 5555 14515
rect 5555 14485 5556 14515
rect 5524 14484 5556 14485
rect 5524 14435 5556 14436
rect 5524 14405 5525 14435
rect 5525 14405 5555 14435
rect 5555 14405 5556 14435
rect 5524 14404 5556 14405
rect 5524 14324 5556 14356
rect 5524 14244 5556 14276
rect 5524 14164 5556 14196
rect 5524 14084 5556 14116
rect 5524 14035 5556 14036
rect 5524 14005 5525 14035
rect 5525 14005 5555 14035
rect 5555 14005 5556 14035
rect 5524 14004 5556 14005
rect 5524 13955 5556 13956
rect 5524 13925 5525 13955
rect 5525 13925 5555 13955
rect 5555 13925 5556 13955
rect 5524 13924 5556 13925
rect 5524 13875 5556 13876
rect 5524 13845 5525 13875
rect 5525 13845 5555 13875
rect 5555 13845 5556 13875
rect 5524 13844 5556 13845
rect 5524 13795 5556 13796
rect 5524 13765 5525 13795
rect 5525 13765 5555 13795
rect 5555 13765 5556 13795
rect 5524 13764 5556 13765
rect 5524 13715 5556 13716
rect 5524 13685 5525 13715
rect 5525 13685 5555 13715
rect 5555 13685 5556 13715
rect 5524 13684 5556 13685
rect 5524 13635 5556 13636
rect 5524 13605 5525 13635
rect 5525 13605 5555 13635
rect 5555 13605 5556 13635
rect 5524 13604 5556 13605
rect 5524 13555 5556 13556
rect 5524 13525 5525 13555
rect 5525 13525 5555 13555
rect 5555 13525 5556 13555
rect 5524 13524 5556 13525
rect 5524 13475 5556 13476
rect 5524 13445 5525 13475
rect 5525 13445 5555 13475
rect 5555 13445 5556 13475
rect 5524 13444 5556 13445
rect 5524 13364 5556 13396
rect 5524 13284 5556 13316
rect 5524 13204 5556 13236
rect 5524 13124 5556 13156
rect 5524 13075 5556 13076
rect 5524 13045 5525 13075
rect 5525 13045 5555 13075
rect 5555 13045 5556 13075
rect 5524 13044 5556 13045
rect 5524 12995 5556 12996
rect 5524 12965 5525 12995
rect 5525 12965 5555 12995
rect 5555 12965 5556 12995
rect 5524 12964 5556 12965
rect 5524 12915 5556 12916
rect 5524 12885 5525 12915
rect 5525 12885 5555 12915
rect 5555 12885 5556 12915
rect 5524 12884 5556 12885
rect 5524 12835 5556 12836
rect 5524 12805 5525 12835
rect 5525 12805 5555 12835
rect 5555 12805 5556 12835
rect 5524 12804 5556 12805
rect 5524 12755 5556 12756
rect 5524 12725 5525 12755
rect 5525 12725 5555 12755
rect 5555 12725 5556 12755
rect 5524 12724 5556 12725
rect 5524 12675 5556 12676
rect 5524 12645 5525 12675
rect 5525 12645 5555 12675
rect 5555 12645 5556 12675
rect 5524 12644 5556 12645
rect 5524 12595 5556 12596
rect 5524 12565 5525 12595
rect 5525 12565 5555 12595
rect 5555 12565 5556 12595
rect 5524 12564 5556 12565
rect 5524 12515 5556 12516
rect 5524 12485 5525 12515
rect 5525 12485 5555 12515
rect 5555 12485 5556 12515
rect 5524 12484 5556 12485
rect 5524 12404 5556 12436
rect 5524 12355 5556 12356
rect 5524 12325 5525 12355
rect 5525 12325 5555 12355
rect 5555 12325 5556 12355
rect 5524 12324 5556 12325
rect 5524 12275 5556 12276
rect 5524 12245 5525 12275
rect 5525 12245 5555 12275
rect 5555 12245 5556 12275
rect 5524 12244 5556 12245
rect 5524 12195 5556 12196
rect 5524 12165 5525 12195
rect 5525 12165 5555 12195
rect 5555 12165 5556 12195
rect 5524 12164 5556 12165
rect 5524 12115 5556 12116
rect 5524 12085 5525 12115
rect 5525 12085 5555 12115
rect 5555 12085 5556 12115
rect 5524 12084 5556 12085
rect 5524 12035 5556 12036
rect 5524 12005 5525 12035
rect 5525 12005 5555 12035
rect 5555 12005 5556 12035
rect 5524 12004 5556 12005
rect 5524 11955 5556 11956
rect 5524 11925 5525 11955
rect 5525 11925 5555 11955
rect 5555 11925 5556 11955
rect 5524 11924 5556 11925
rect 5524 11875 5556 11876
rect 5524 11845 5525 11875
rect 5525 11845 5555 11875
rect 5555 11845 5556 11875
rect 5524 11844 5556 11845
rect 5524 11795 5556 11796
rect 5524 11765 5525 11795
rect 5525 11765 5555 11795
rect 5555 11765 5556 11795
rect 5524 11764 5556 11765
rect 5524 11715 5556 11716
rect 5524 11685 5525 11715
rect 5525 11685 5555 11715
rect 5555 11685 5556 11715
rect 5524 11684 5556 11685
rect 5524 11635 5556 11636
rect 5524 11605 5525 11635
rect 5525 11605 5555 11635
rect 5555 11605 5556 11635
rect 5524 11604 5556 11605
rect 5524 11555 5556 11556
rect 5524 11525 5525 11555
rect 5525 11525 5555 11555
rect 5555 11525 5556 11555
rect 5524 11524 5556 11525
rect 5524 11475 5556 11476
rect 5524 11445 5525 11475
rect 5525 11445 5555 11475
rect 5555 11445 5556 11475
rect 5524 11444 5556 11445
rect 5524 11395 5556 11396
rect 5524 11365 5525 11395
rect 5525 11365 5555 11395
rect 5555 11365 5556 11395
rect 5524 11364 5556 11365
rect 5524 11315 5556 11316
rect 5524 11285 5525 11315
rect 5525 11285 5555 11315
rect 5555 11285 5556 11315
rect 5524 11284 5556 11285
rect 5524 11235 5556 11236
rect 5524 11205 5525 11235
rect 5525 11205 5555 11235
rect 5555 11205 5556 11235
rect 5524 11204 5556 11205
rect 5524 11155 5556 11156
rect 5524 11125 5525 11155
rect 5525 11125 5555 11155
rect 5555 11125 5556 11155
rect 5524 11124 5556 11125
rect 5524 11075 5556 11076
rect 5524 11045 5525 11075
rect 5525 11045 5555 11075
rect 5555 11045 5556 11075
rect 5524 11044 5556 11045
rect 5524 10964 5556 10996
rect 5524 10915 5556 10916
rect 5524 10885 5525 10915
rect 5525 10885 5555 10915
rect 5555 10885 5556 10915
rect 5524 10884 5556 10885
rect 5524 10835 5556 10836
rect 5524 10805 5525 10835
rect 5525 10805 5555 10835
rect 5555 10805 5556 10835
rect 5524 10804 5556 10805
rect 5524 10755 5556 10756
rect 5524 10725 5525 10755
rect 5525 10725 5555 10755
rect 5555 10725 5556 10755
rect 5524 10724 5556 10725
rect 5524 10675 5556 10676
rect 5524 10645 5525 10675
rect 5525 10645 5555 10675
rect 5555 10645 5556 10675
rect 5524 10644 5556 10645
rect 5524 10595 5556 10596
rect 5524 10565 5525 10595
rect 5525 10565 5555 10595
rect 5555 10565 5556 10595
rect 5524 10564 5556 10565
rect 5524 10515 5556 10516
rect 5524 10485 5525 10515
rect 5525 10485 5555 10515
rect 5555 10485 5556 10515
rect 5524 10484 5556 10485
rect 5524 10435 5556 10436
rect 5524 10405 5525 10435
rect 5525 10405 5555 10435
rect 5555 10405 5556 10435
rect 5524 10404 5556 10405
rect 5524 10355 5556 10356
rect 5524 10325 5525 10355
rect 5525 10325 5555 10355
rect 5555 10325 5556 10355
rect 5524 10324 5556 10325
rect 5524 10244 5556 10276
rect 5524 10164 5556 10196
rect 5524 10084 5556 10116
rect 5524 10004 5556 10036
rect 5524 9955 5556 9956
rect 5524 9925 5525 9955
rect 5525 9925 5555 9955
rect 5555 9925 5556 9955
rect 5524 9924 5556 9925
rect 5524 9875 5556 9876
rect 5524 9845 5525 9875
rect 5525 9845 5555 9875
rect 5555 9845 5556 9875
rect 5524 9844 5556 9845
rect 5524 9795 5556 9796
rect 5524 9765 5525 9795
rect 5525 9765 5555 9795
rect 5555 9765 5556 9795
rect 5524 9764 5556 9765
rect 5524 9715 5556 9716
rect 5524 9685 5525 9715
rect 5525 9685 5555 9715
rect 5555 9685 5556 9715
rect 5524 9684 5556 9685
rect 5524 9635 5556 9636
rect 5524 9605 5525 9635
rect 5525 9605 5555 9635
rect 5555 9605 5556 9635
rect 5524 9604 5556 9605
rect 5524 9555 5556 9556
rect 5524 9525 5525 9555
rect 5525 9525 5555 9555
rect 5555 9525 5556 9555
rect 5524 9524 5556 9525
rect 5524 9475 5556 9476
rect 5524 9445 5525 9475
rect 5525 9445 5555 9475
rect 5555 9445 5556 9475
rect 5524 9444 5556 9445
rect 5524 9395 5556 9396
rect 5524 9365 5525 9395
rect 5525 9365 5555 9395
rect 5555 9365 5556 9395
rect 5524 9364 5556 9365
rect 5524 9284 5556 9316
rect 5524 9204 5556 9236
rect 5524 9124 5556 9156
rect 5524 9044 5556 9076
rect 5524 8995 5556 8996
rect 5524 8965 5525 8995
rect 5525 8965 5555 8995
rect 5555 8965 5556 8995
rect 5524 8964 5556 8965
rect 5524 8915 5556 8916
rect 5524 8885 5525 8915
rect 5525 8885 5555 8915
rect 5555 8885 5556 8915
rect 5524 8884 5556 8885
rect 5524 8835 5556 8836
rect 5524 8805 5525 8835
rect 5525 8805 5555 8835
rect 5555 8805 5556 8835
rect 5524 8804 5556 8805
rect 5524 8755 5556 8756
rect 5524 8725 5525 8755
rect 5525 8725 5555 8755
rect 5555 8725 5556 8755
rect 5524 8724 5556 8725
rect 5524 8675 5556 8676
rect 5524 8645 5525 8675
rect 5525 8645 5555 8675
rect 5555 8645 5556 8675
rect 5524 8644 5556 8645
rect 5524 8595 5556 8596
rect 5524 8565 5525 8595
rect 5525 8565 5555 8595
rect 5555 8565 5556 8595
rect 5524 8564 5556 8565
rect 5524 8515 5556 8516
rect 5524 8485 5525 8515
rect 5525 8485 5555 8515
rect 5555 8485 5556 8515
rect 5524 8484 5556 8485
rect 5524 8435 5556 8436
rect 5524 8405 5525 8435
rect 5525 8405 5555 8435
rect 5555 8405 5556 8435
rect 5524 8404 5556 8405
rect 5524 8324 5556 8356
rect 5524 8275 5556 8276
rect 5524 8245 5525 8275
rect 5525 8245 5555 8275
rect 5555 8245 5556 8275
rect 5524 8244 5556 8245
rect 5524 8195 5556 8196
rect 5524 8165 5525 8195
rect 5525 8165 5555 8195
rect 5555 8165 5556 8195
rect 5524 8164 5556 8165
rect 5524 8115 5556 8116
rect 5524 8085 5525 8115
rect 5525 8085 5555 8115
rect 5555 8085 5556 8115
rect 5524 8084 5556 8085
rect 5524 8035 5556 8036
rect 5524 8005 5525 8035
rect 5525 8005 5555 8035
rect 5555 8005 5556 8035
rect 5524 8004 5556 8005
rect 5524 7955 5556 7956
rect 5524 7925 5525 7955
rect 5525 7925 5555 7955
rect 5555 7925 5556 7955
rect 5524 7924 5556 7925
rect 5524 7875 5556 7876
rect 5524 7845 5525 7875
rect 5525 7845 5555 7875
rect 5555 7845 5556 7875
rect 5524 7844 5556 7845
rect 5524 7795 5556 7796
rect 5524 7765 5525 7795
rect 5525 7765 5555 7795
rect 5555 7765 5556 7795
rect 5524 7764 5556 7765
rect 5524 7715 5556 7716
rect 5524 7685 5525 7715
rect 5525 7685 5555 7715
rect 5555 7685 5556 7715
rect 5524 7684 5556 7685
rect 5524 7635 5556 7636
rect 5524 7605 5525 7635
rect 5525 7605 5555 7635
rect 5555 7605 5556 7635
rect 5524 7604 5556 7605
rect 5524 7555 5556 7556
rect 5524 7525 5525 7555
rect 5525 7525 5555 7555
rect 5555 7525 5556 7555
rect 5524 7524 5556 7525
rect 5524 7475 5556 7476
rect 5524 7445 5525 7475
rect 5525 7445 5555 7475
rect 5555 7445 5556 7475
rect 5524 7444 5556 7445
rect 5524 7395 5556 7396
rect 5524 7365 5525 7395
rect 5525 7365 5555 7395
rect 5555 7365 5556 7395
rect 5524 7364 5556 7365
rect 5524 7315 5556 7316
rect 5524 7285 5525 7315
rect 5525 7285 5555 7315
rect 5555 7285 5556 7315
rect 5524 7284 5556 7285
rect 5524 7235 5556 7236
rect 5524 7205 5525 7235
rect 5525 7205 5555 7235
rect 5555 7205 5556 7235
rect 5524 7204 5556 7205
rect 5524 7155 5556 7156
rect 5524 7125 5525 7155
rect 5525 7125 5555 7155
rect 5555 7125 5556 7155
rect 5524 7124 5556 7125
rect 5524 7075 5556 7076
rect 5524 7045 5525 7075
rect 5525 7045 5555 7075
rect 5555 7045 5556 7075
rect 5524 7044 5556 7045
rect 5524 6995 5556 6996
rect 5524 6965 5525 6995
rect 5525 6965 5555 6995
rect 5555 6965 5556 6995
rect 5524 6964 5556 6965
rect 5524 6884 5556 6916
rect 5524 6835 5556 6836
rect 5524 6805 5525 6835
rect 5525 6805 5555 6835
rect 5555 6805 5556 6835
rect 5524 6804 5556 6805
rect 5524 6755 5556 6756
rect 5524 6725 5525 6755
rect 5525 6725 5555 6755
rect 5555 6725 5556 6755
rect 5524 6724 5556 6725
rect 5524 6675 5556 6676
rect 5524 6645 5525 6675
rect 5525 6645 5555 6675
rect 5555 6645 5556 6675
rect 5524 6644 5556 6645
rect 5524 6595 5556 6596
rect 5524 6565 5525 6595
rect 5525 6565 5555 6595
rect 5555 6565 5556 6595
rect 5524 6564 5556 6565
rect 5524 6515 5556 6516
rect 5524 6485 5525 6515
rect 5525 6485 5555 6515
rect 5555 6485 5556 6515
rect 5524 6484 5556 6485
rect 5524 6435 5556 6436
rect 5524 6405 5525 6435
rect 5525 6405 5555 6435
rect 5555 6405 5556 6435
rect 5524 6404 5556 6405
rect 5524 6355 5556 6356
rect 5524 6325 5525 6355
rect 5525 6325 5555 6355
rect 5555 6325 5556 6355
rect 5524 6324 5556 6325
rect 5524 6275 5556 6276
rect 5524 6245 5525 6275
rect 5525 6245 5555 6275
rect 5555 6245 5556 6275
rect 5524 6244 5556 6245
rect 5524 6164 5556 6196
rect 5524 6084 5556 6116
rect 5524 6004 5556 6036
rect 5524 5924 5556 5956
rect 5524 5875 5556 5876
rect 5524 5845 5525 5875
rect 5525 5845 5555 5875
rect 5555 5845 5556 5875
rect 5524 5844 5556 5845
rect 5524 5795 5556 5796
rect 5524 5765 5525 5795
rect 5525 5765 5555 5795
rect 5555 5765 5556 5795
rect 5524 5764 5556 5765
rect 5524 5715 5556 5716
rect 5524 5685 5525 5715
rect 5525 5685 5555 5715
rect 5555 5685 5556 5715
rect 5524 5684 5556 5685
rect 5524 5635 5556 5636
rect 5524 5605 5525 5635
rect 5525 5605 5555 5635
rect 5555 5605 5556 5635
rect 5524 5604 5556 5605
rect 5524 5555 5556 5556
rect 5524 5525 5525 5555
rect 5525 5525 5555 5555
rect 5555 5525 5556 5555
rect 5524 5524 5556 5525
rect 5524 5475 5556 5476
rect 5524 5445 5525 5475
rect 5525 5445 5555 5475
rect 5555 5445 5556 5475
rect 5524 5444 5556 5445
rect 5524 5395 5556 5396
rect 5524 5365 5525 5395
rect 5525 5365 5555 5395
rect 5555 5365 5556 5395
rect 5524 5364 5556 5365
rect 5524 5315 5556 5316
rect 5524 5285 5525 5315
rect 5525 5285 5555 5315
rect 5555 5285 5556 5315
rect 5524 5284 5556 5285
rect 5524 5235 5556 5236
rect 5524 5205 5525 5235
rect 5525 5205 5555 5235
rect 5555 5205 5556 5235
rect 5524 5204 5556 5205
rect 5524 5155 5556 5156
rect 5524 5125 5525 5155
rect 5525 5125 5555 5155
rect 5555 5125 5556 5155
rect 5524 5124 5556 5125
rect 5524 5075 5556 5076
rect 5524 5045 5525 5075
rect 5525 5045 5555 5075
rect 5555 5045 5556 5075
rect 5524 5044 5556 5045
rect 5524 4995 5556 4996
rect 5524 4965 5525 4995
rect 5525 4965 5555 4995
rect 5555 4965 5556 4995
rect 5524 4964 5556 4965
rect 5524 4915 5556 4916
rect 5524 4885 5525 4915
rect 5525 4885 5555 4915
rect 5555 4885 5556 4915
rect 5524 4884 5556 4885
rect 5524 4804 5556 4836
rect 5524 4755 5556 4756
rect 5524 4725 5525 4755
rect 5525 4725 5555 4755
rect 5555 4725 5556 4755
rect 5524 4724 5556 4725
rect 5524 4675 5556 4676
rect 5524 4645 5525 4675
rect 5525 4645 5555 4675
rect 5555 4645 5556 4675
rect 5524 4644 5556 4645
rect 5524 4564 5556 4596
rect 5524 4515 5556 4516
rect 5524 4485 5525 4515
rect 5525 4485 5555 4515
rect 5555 4485 5556 4515
rect 5524 4484 5556 4485
rect 5524 4435 5556 4436
rect 5524 4405 5525 4435
rect 5525 4405 5555 4435
rect 5555 4405 5556 4435
rect 5524 4404 5556 4405
rect 5524 4355 5556 4356
rect 5524 4325 5525 4355
rect 5525 4325 5555 4355
rect 5555 4325 5556 4355
rect 5524 4324 5556 4325
rect 5524 4275 5556 4276
rect 5524 4245 5525 4275
rect 5525 4245 5555 4275
rect 5555 4245 5556 4275
rect 5524 4244 5556 4245
rect 5524 4195 5556 4196
rect 5524 4165 5525 4195
rect 5525 4165 5555 4195
rect 5555 4165 5556 4195
rect 5524 4164 5556 4165
rect 5524 4115 5556 4116
rect 5524 4085 5525 4115
rect 5525 4085 5555 4115
rect 5555 4085 5556 4115
rect 5524 4084 5556 4085
rect 5524 4035 5556 4036
rect 5524 4005 5525 4035
rect 5525 4005 5555 4035
rect 5555 4005 5556 4035
rect 5524 4004 5556 4005
rect 5524 3955 5556 3956
rect 5524 3925 5525 3955
rect 5525 3925 5555 3955
rect 5555 3925 5556 3955
rect 5524 3924 5556 3925
rect 5524 3875 5556 3876
rect 5524 3845 5525 3875
rect 5525 3845 5555 3875
rect 5555 3845 5556 3875
rect 5524 3844 5556 3845
rect 5524 3764 5556 3796
rect 5524 3715 5556 3716
rect 5524 3685 5525 3715
rect 5525 3685 5555 3715
rect 5555 3685 5556 3715
rect 5524 3684 5556 3685
rect 5524 3635 5556 3636
rect 5524 3605 5525 3635
rect 5525 3605 5555 3635
rect 5555 3605 5556 3635
rect 5524 3604 5556 3605
rect 5524 3524 5556 3556
rect 5524 3475 5556 3476
rect 5524 3445 5525 3475
rect 5525 3445 5555 3475
rect 5555 3445 5556 3475
rect 5524 3444 5556 3445
rect 5524 3395 5556 3396
rect 5524 3365 5525 3395
rect 5525 3365 5555 3395
rect 5555 3365 5556 3395
rect 5524 3364 5556 3365
rect 5524 3284 5556 3316
rect 5524 3235 5556 3236
rect 5524 3205 5525 3235
rect 5525 3205 5555 3235
rect 5555 3205 5556 3235
rect 5524 3204 5556 3205
rect 5524 3155 5556 3156
rect 5524 3125 5525 3155
rect 5525 3125 5555 3155
rect 5555 3125 5556 3155
rect 5524 3124 5556 3125
rect 5524 3075 5556 3076
rect 5524 3045 5525 3075
rect 5525 3045 5555 3075
rect 5555 3045 5556 3075
rect 5524 3044 5556 3045
rect 5524 2995 5556 2996
rect 5524 2965 5525 2995
rect 5525 2965 5555 2995
rect 5555 2965 5556 2995
rect 5524 2964 5556 2965
rect 5524 2915 5556 2916
rect 5524 2885 5525 2915
rect 5525 2885 5555 2915
rect 5555 2885 5556 2915
rect 5524 2884 5556 2885
rect 5524 2835 5556 2836
rect 5524 2805 5525 2835
rect 5525 2805 5555 2835
rect 5555 2805 5556 2835
rect 5524 2804 5556 2805
rect 5524 2755 5556 2756
rect 5524 2725 5525 2755
rect 5525 2725 5555 2755
rect 5555 2725 5556 2755
rect 5524 2724 5556 2725
rect 5524 2675 5556 2676
rect 5524 2645 5525 2675
rect 5525 2645 5555 2675
rect 5555 2645 5556 2675
rect 5524 2644 5556 2645
rect 5524 2595 5556 2596
rect 5524 2565 5525 2595
rect 5525 2565 5555 2595
rect 5555 2565 5556 2595
rect 5524 2564 5556 2565
rect 5524 2515 5556 2516
rect 5524 2485 5525 2515
rect 5525 2485 5555 2515
rect 5555 2485 5556 2515
rect 5524 2484 5556 2485
rect 5524 2435 5556 2436
rect 5524 2405 5525 2435
rect 5525 2405 5555 2435
rect 5555 2405 5556 2435
rect 5524 2404 5556 2405
rect 5524 2355 5556 2356
rect 5524 2325 5525 2355
rect 5525 2325 5555 2355
rect 5555 2325 5556 2355
rect 5524 2324 5556 2325
rect 5524 2275 5556 2276
rect 5524 2245 5525 2275
rect 5525 2245 5555 2275
rect 5555 2245 5556 2275
rect 5524 2244 5556 2245
rect 5524 2195 5556 2196
rect 5524 2165 5525 2195
rect 5525 2165 5555 2195
rect 5555 2165 5556 2195
rect 5524 2164 5556 2165
rect 5524 2115 5556 2116
rect 5524 2085 5525 2115
rect 5525 2085 5555 2115
rect 5555 2085 5556 2115
rect 5524 2084 5556 2085
rect 5524 2035 5556 2036
rect 5524 2005 5525 2035
rect 5525 2005 5555 2035
rect 5555 2005 5556 2035
rect 5524 2004 5556 2005
rect 5524 1955 5556 1956
rect 5524 1925 5525 1955
rect 5525 1925 5555 1955
rect 5555 1925 5556 1955
rect 5524 1924 5556 1925
rect 5524 1844 5556 1876
rect 5524 1764 5556 1796
rect 5524 1715 5556 1716
rect 5524 1685 5525 1715
rect 5525 1685 5555 1715
rect 5555 1685 5556 1715
rect 5524 1684 5556 1685
rect 5524 1635 5556 1636
rect 5524 1605 5525 1635
rect 5525 1605 5555 1635
rect 5555 1605 5556 1635
rect 5524 1604 5556 1605
rect 5524 1555 5556 1556
rect 5524 1525 5525 1555
rect 5525 1525 5555 1555
rect 5555 1525 5556 1555
rect 5524 1524 5556 1525
rect 5524 1475 5556 1476
rect 5524 1445 5525 1475
rect 5525 1445 5555 1475
rect 5555 1445 5556 1475
rect 5524 1444 5556 1445
rect 5524 1395 5556 1396
rect 5524 1365 5525 1395
rect 5525 1365 5555 1395
rect 5555 1365 5556 1395
rect 5524 1364 5556 1365
rect 5524 1315 5556 1316
rect 5524 1285 5525 1315
rect 5525 1285 5555 1315
rect 5555 1285 5556 1315
rect 5524 1284 5556 1285
rect 5524 1235 5556 1236
rect 5524 1205 5525 1235
rect 5525 1205 5555 1235
rect 5555 1205 5556 1235
rect 5524 1204 5556 1205
rect 5524 1155 5556 1156
rect 5524 1125 5525 1155
rect 5525 1125 5555 1155
rect 5555 1125 5556 1155
rect 5524 1124 5556 1125
rect 5524 1075 5556 1076
rect 5524 1045 5525 1075
rect 5525 1045 5555 1075
rect 5555 1045 5556 1075
rect 5524 1044 5556 1045
rect 5524 995 5556 996
rect 5524 965 5525 995
rect 5525 965 5555 995
rect 5555 965 5556 995
rect 5524 964 5556 965
rect 5524 884 5556 916
rect 5524 835 5556 836
rect 5524 805 5525 835
rect 5525 805 5555 835
rect 5555 805 5556 835
rect 5524 804 5556 805
rect 5524 755 5556 756
rect 5524 725 5525 755
rect 5525 725 5555 755
rect 5555 725 5556 755
rect 5524 724 5556 725
rect 5524 675 5556 676
rect 5524 645 5525 675
rect 5525 645 5555 675
rect 5555 645 5556 675
rect 5524 644 5556 645
rect 5524 595 5556 596
rect 5524 565 5525 595
rect 5525 565 5555 595
rect 5555 565 5556 595
rect 5524 564 5556 565
rect 5524 515 5556 516
rect 5524 485 5525 515
rect 5525 485 5555 515
rect 5555 485 5556 515
rect 5524 484 5556 485
rect 5524 404 5556 436
rect 5524 324 5556 356
rect 5524 275 5556 276
rect 5524 245 5525 275
rect 5525 245 5555 275
rect 5555 245 5556 275
rect 5524 244 5556 245
rect 5524 195 5556 196
rect 5524 165 5525 195
rect 5525 165 5555 195
rect 5555 165 5556 195
rect 5524 164 5556 165
rect 5524 115 5556 116
rect 5524 85 5525 115
rect 5525 85 5555 115
rect 5555 85 5556 115
rect 5524 84 5556 85
rect 5524 35 5556 36
rect 5524 5 5525 35
rect 5525 5 5555 35
rect 5555 5 5556 35
rect 5524 4 5556 5
rect 5364 -716 5396 -524
rect 5684 15715 5716 15716
rect 5684 15685 5685 15715
rect 5685 15685 5715 15715
rect 5715 15685 5716 15715
rect 5684 15684 5716 15685
rect 5684 15635 5716 15636
rect 5684 15605 5685 15635
rect 5685 15605 5715 15635
rect 5715 15605 5716 15635
rect 5684 15604 5716 15605
rect 5684 15555 5716 15556
rect 5684 15525 5685 15555
rect 5685 15525 5715 15555
rect 5715 15525 5716 15555
rect 5684 15524 5716 15525
rect 5684 15475 5716 15476
rect 5684 15445 5685 15475
rect 5685 15445 5715 15475
rect 5715 15445 5716 15475
rect 5684 15444 5716 15445
rect 5684 15395 5716 15396
rect 5684 15365 5685 15395
rect 5685 15365 5715 15395
rect 5715 15365 5716 15395
rect 5684 15364 5716 15365
rect 5684 15315 5716 15316
rect 5684 15285 5685 15315
rect 5685 15285 5715 15315
rect 5715 15285 5716 15315
rect 5684 15284 5716 15285
rect 5684 15235 5716 15236
rect 5684 15205 5685 15235
rect 5685 15205 5715 15235
rect 5715 15205 5716 15235
rect 5684 15204 5716 15205
rect 5684 15155 5716 15156
rect 5684 15125 5685 15155
rect 5685 15125 5715 15155
rect 5715 15125 5716 15155
rect 5684 15124 5716 15125
rect 5684 15044 5716 15076
rect 5684 14995 5716 14996
rect 5684 14965 5685 14995
rect 5685 14965 5715 14995
rect 5715 14965 5716 14995
rect 5684 14964 5716 14965
rect 5684 14915 5716 14916
rect 5684 14885 5685 14915
rect 5685 14885 5715 14915
rect 5715 14885 5716 14915
rect 5684 14884 5716 14885
rect 5684 14835 5716 14836
rect 5684 14805 5685 14835
rect 5685 14805 5715 14835
rect 5715 14805 5716 14835
rect 5684 14804 5716 14805
rect 5684 14755 5716 14756
rect 5684 14725 5685 14755
rect 5685 14725 5715 14755
rect 5715 14725 5716 14755
rect 5684 14724 5716 14725
rect 5684 14675 5716 14676
rect 5684 14645 5685 14675
rect 5685 14645 5715 14675
rect 5715 14645 5716 14675
rect 5684 14644 5716 14645
rect 5684 14595 5716 14596
rect 5684 14565 5685 14595
rect 5685 14565 5715 14595
rect 5715 14565 5716 14595
rect 5684 14564 5716 14565
rect 5684 14515 5716 14516
rect 5684 14485 5685 14515
rect 5685 14485 5715 14515
rect 5715 14485 5716 14515
rect 5684 14484 5716 14485
rect 5684 14435 5716 14436
rect 5684 14405 5685 14435
rect 5685 14405 5715 14435
rect 5715 14405 5716 14435
rect 5684 14404 5716 14405
rect 5684 14324 5716 14356
rect 5684 14244 5716 14276
rect 5684 14164 5716 14196
rect 5684 14084 5716 14116
rect 5684 14035 5716 14036
rect 5684 14005 5685 14035
rect 5685 14005 5715 14035
rect 5715 14005 5716 14035
rect 5684 14004 5716 14005
rect 5684 13955 5716 13956
rect 5684 13925 5685 13955
rect 5685 13925 5715 13955
rect 5715 13925 5716 13955
rect 5684 13924 5716 13925
rect 5684 13875 5716 13876
rect 5684 13845 5685 13875
rect 5685 13845 5715 13875
rect 5715 13845 5716 13875
rect 5684 13844 5716 13845
rect 5684 13795 5716 13796
rect 5684 13765 5685 13795
rect 5685 13765 5715 13795
rect 5715 13765 5716 13795
rect 5684 13764 5716 13765
rect 5684 13715 5716 13716
rect 5684 13685 5685 13715
rect 5685 13685 5715 13715
rect 5715 13685 5716 13715
rect 5684 13684 5716 13685
rect 5684 13635 5716 13636
rect 5684 13605 5685 13635
rect 5685 13605 5715 13635
rect 5715 13605 5716 13635
rect 5684 13604 5716 13605
rect 5684 13555 5716 13556
rect 5684 13525 5685 13555
rect 5685 13525 5715 13555
rect 5715 13525 5716 13555
rect 5684 13524 5716 13525
rect 5684 13475 5716 13476
rect 5684 13445 5685 13475
rect 5685 13445 5715 13475
rect 5715 13445 5716 13475
rect 5684 13444 5716 13445
rect 5684 13364 5716 13396
rect 5684 13284 5716 13316
rect 5684 13204 5716 13236
rect 5684 13124 5716 13156
rect 5684 13075 5716 13076
rect 5684 13045 5685 13075
rect 5685 13045 5715 13075
rect 5715 13045 5716 13075
rect 5684 13044 5716 13045
rect 5684 12995 5716 12996
rect 5684 12965 5685 12995
rect 5685 12965 5715 12995
rect 5715 12965 5716 12995
rect 5684 12964 5716 12965
rect 5684 12915 5716 12916
rect 5684 12885 5685 12915
rect 5685 12885 5715 12915
rect 5715 12885 5716 12915
rect 5684 12884 5716 12885
rect 5684 12835 5716 12836
rect 5684 12805 5685 12835
rect 5685 12805 5715 12835
rect 5715 12805 5716 12835
rect 5684 12804 5716 12805
rect 5684 12755 5716 12756
rect 5684 12725 5685 12755
rect 5685 12725 5715 12755
rect 5715 12725 5716 12755
rect 5684 12724 5716 12725
rect 5684 12675 5716 12676
rect 5684 12645 5685 12675
rect 5685 12645 5715 12675
rect 5715 12645 5716 12675
rect 5684 12644 5716 12645
rect 5684 12595 5716 12596
rect 5684 12565 5685 12595
rect 5685 12565 5715 12595
rect 5715 12565 5716 12595
rect 5684 12564 5716 12565
rect 5684 12515 5716 12516
rect 5684 12485 5685 12515
rect 5685 12485 5715 12515
rect 5715 12485 5716 12515
rect 5684 12484 5716 12485
rect 5684 12404 5716 12436
rect 5684 12355 5716 12356
rect 5684 12325 5685 12355
rect 5685 12325 5715 12355
rect 5715 12325 5716 12355
rect 5684 12324 5716 12325
rect 5684 12275 5716 12276
rect 5684 12245 5685 12275
rect 5685 12245 5715 12275
rect 5715 12245 5716 12275
rect 5684 12244 5716 12245
rect 5684 12195 5716 12196
rect 5684 12165 5685 12195
rect 5685 12165 5715 12195
rect 5715 12165 5716 12195
rect 5684 12164 5716 12165
rect 5684 12115 5716 12116
rect 5684 12085 5685 12115
rect 5685 12085 5715 12115
rect 5715 12085 5716 12115
rect 5684 12084 5716 12085
rect 5684 12035 5716 12036
rect 5684 12005 5685 12035
rect 5685 12005 5715 12035
rect 5715 12005 5716 12035
rect 5684 12004 5716 12005
rect 5684 11955 5716 11956
rect 5684 11925 5685 11955
rect 5685 11925 5715 11955
rect 5715 11925 5716 11955
rect 5684 11924 5716 11925
rect 5684 11875 5716 11876
rect 5684 11845 5685 11875
rect 5685 11845 5715 11875
rect 5715 11845 5716 11875
rect 5684 11844 5716 11845
rect 5684 11795 5716 11796
rect 5684 11765 5685 11795
rect 5685 11765 5715 11795
rect 5715 11765 5716 11795
rect 5684 11764 5716 11765
rect 5684 11715 5716 11716
rect 5684 11685 5685 11715
rect 5685 11685 5715 11715
rect 5715 11685 5716 11715
rect 5684 11684 5716 11685
rect 5684 11635 5716 11636
rect 5684 11605 5685 11635
rect 5685 11605 5715 11635
rect 5715 11605 5716 11635
rect 5684 11604 5716 11605
rect 5684 11555 5716 11556
rect 5684 11525 5685 11555
rect 5685 11525 5715 11555
rect 5715 11525 5716 11555
rect 5684 11524 5716 11525
rect 5684 11475 5716 11476
rect 5684 11445 5685 11475
rect 5685 11445 5715 11475
rect 5715 11445 5716 11475
rect 5684 11444 5716 11445
rect 5684 11395 5716 11396
rect 5684 11365 5685 11395
rect 5685 11365 5715 11395
rect 5715 11365 5716 11395
rect 5684 11364 5716 11365
rect 5684 11315 5716 11316
rect 5684 11285 5685 11315
rect 5685 11285 5715 11315
rect 5715 11285 5716 11315
rect 5684 11284 5716 11285
rect 5684 11235 5716 11236
rect 5684 11205 5685 11235
rect 5685 11205 5715 11235
rect 5715 11205 5716 11235
rect 5684 11204 5716 11205
rect 5684 11155 5716 11156
rect 5684 11125 5685 11155
rect 5685 11125 5715 11155
rect 5715 11125 5716 11155
rect 5684 11124 5716 11125
rect 5684 11075 5716 11076
rect 5684 11045 5685 11075
rect 5685 11045 5715 11075
rect 5715 11045 5716 11075
rect 5684 11044 5716 11045
rect 5684 10964 5716 10996
rect 5684 10915 5716 10916
rect 5684 10885 5685 10915
rect 5685 10885 5715 10915
rect 5715 10885 5716 10915
rect 5684 10884 5716 10885
rect 5684 10835 5716 10836
rect 5684 10805 5685 10835
rect 5685 10805 5715 10835
rect 5715 10805 5716 10835
rect 5684 10804 5716 10805
rect 5684 10755 5716 10756
rect 5684 10725 5685 10755
rect 5685 10725 5715 10755
rect 5715 10725 5716 10755
rect 5684 10724 5716 10725
rect 5684 10675 5716 10676
rect 5684 10645 5685 10675
rect 5685 10645 5715 10675
rect 5715 10645 5716 10675
rect 5684 10644 5716 10645
rect 5684 10595 5716 10596
rect 5684 10565 5685 10595
rect 5685 10565 5715 10595
rect 5715 10565 5716 10595
rect 5684 10564 5716 10565
rect 5684 10515 5716 10516
rect 5684 10485 5685 10515
rect 5685 10485 5715 10515
rect 5715 10485 5716 10515
rect 5684 10484 5716 10485
rect 5684 10435 5716 10436
rect 5684 10405 5685 10435
rect 5685 10405 5715 10435
rect 5715 10405 5716 10435
rect 5684 10404 5716 10405
rect 5684 10355 5716 10356
rect 5684 10325 5685 10355
rect 5685 10325 5715 10355
rect 5715 10325 5716 10355
rect 5684 10324 5716 10325
rect 5684 10244 5716 10276
rect 5684 10164 5716 10196
rect 5684 10084 5716 10116
rect 5684 10004 5716 10036
rect 5684 9955 5716 9956
rect 5684 9925 5685 9955
rect 5685 9925 5715 9955
rect 5715 9925 5716 9955
rect 5684 9924 5716 9925
rect 5684 9875 5716 9876
rect 5684 9845 5685 9875
rect 5685 9845 5715 9875
rect 5715 9845 5716 9875
rect 5684 9844 5716 9845
rect 5684 9795 5716 9796
rect 5684 9765 5685 9795
rect 5685 9765 5715 9795
rect 5715 9765 5716 9795
rect 5684 9764 5716 9765
rect 5684 9715 5716 9716
rect 5684 9685 5685 9715
rect 5685 9685 5715 9715
rect 5715 9685 5716 9715
rect 5684 9684 5716 9685
rect 5684 9635 5716 9636
rect 5684 9605 5685 9635
rect 5685 9605 5715 9635
rect 5715 9605 5716 9635
rect 5684 9604 5716 9605
rect 5684 9555 5716 9556
rect 5684 9525 5685 9555
rect 5685 9525 5715 9555
rect 5715 9525 5716 9555
rect 5684 9524 5716 9525
rect 5684 9475 5716 9476
rect 5684 9445 5685 9475
rect 5685 9445 5715 9475
rect 5715 9445 5716 9475
rect 5684 9444 5716 9445
rect 5684 9395 5716 9396
rect 5684 9365 5685 9395
rect 5685 9365 5715 9395
rect 5715 9365 5716 9395
rect 5684 9364 5716 9365
rect 5684 9284 5716 9316
rect 5684 9204 5716 9236
rect 5684 9124 5716 9156
rect 5684 9044 5716 9076
rect 5684 8995 5716 8996
rect 5684 8965 5685 8995
rect 5685 8965 5715 8995
rect 5715 8965 5716 8995
rect 5684 8964 5716 8965
rect 5684 8915 5716 8916
rect 5684 8885 5685 8915
rect 5685 8885 5715 8915
rect 5715 8885 5716 8915
rect 5684 8884 5716 8885
rect 5684 8835 5716 8836
rect 5684 8805 5685 8835
rect 5685 8805 5715 8835
rect 5715 8805 5716 8835
rect 5684 8804 5716 8805
rect 5684 8755 5716 8756
rect 5684 8725 5685 8755
rect 5685 8725 5715 8755
rect 5715 8725 5716 8755
rect 5684 8724 5716 8725
rect 5684 8675 5716 8676
rect 5684 8645 5685 8675
rect 5685 8645 5715 8675
rect 5715 8645 5716 8675
rect 5684 8644 5716 8645
rect 5684 8595 5716 8596
rect 5684 8565 5685 8595
rect 5685 8565 5715 8595
rect 5715 8565 5716 8595
rect 5684 8564 5716 8565
rect 5684 8515 5716 8516
rect 5684 8485 5685 8515
rect 5685 8485 5715 8515
rect 5715 8485 5716 8515
rect 5684 8484 5716 8485
rect 5684 8435 5716 8436
rect 5684 8405 5685 8435
rect 5685 8405 5715 8435
rect 5715 8405 5716 8435
rect 5684 8404 5716 8405
rect 5684 8324 5716 8356
rect 5684 8275 5716 8276
rect 5684 8245 5685 8275
rect 5685 8245 5715 8275
rect 5715 8245 5716 8275
rect 5684 8244 5716 8245
rect 5684 8195 5716 8196
rect 5684 8165 5685 8195
rect 5685 8165 5715 8195
rect 5715 8165 5716 8195
rect 5684 8164 5716 8165
rect 5684 8115 5716 8116
rect 5684 8085 5685 8115
rect 5685 8085 5715 8115
rect 5715 8085 5716 8115
rect 5684 8084 5716 8085
rect 5684 8035 5716 8036
rect 5684 8005 5685 8035
rect 5685 8005 5715 8035
rect 5715 8005 5716 8035
rect 5684 8004 5716 8005
rect 5684 7955 5716 7956
rect 5684 7925 5685 7955
rect 5685 7925 5715 7955
rect 5715 7925 5716 7955
rect 5684 7924 5716 7925
rect 5684 7875 5716 7876
rect 5684 7845 5685 7875
rect 5685 7845 5715 7875
rect 5715 7845 5716 7875
rect 5684 7844 5716 7845
rect 5684 7795 5716 7796
rect 5684 7765 5685 7795
rect 5685 7765 5715 7795
rect 5715 7765 5716 7795
rect 5684 7764 5716 7765
rect 5684 7715 5716 7716
rect 5684 7685 5685 7715
rect 5685 7685 5715 7715
rect 5715 7685 5716 7715
rect 5684 7684 5716 7685
rect 5684 7635 5716 7636
rect 5684 7605 5685 7635
rect 5685 7605 5715 7635
rect 5715 7605 5716 7635
rect 5684 7604 5716 7605
rect 5684 7555 5716 7556
rect 5684 7525 5685 7555
rect 5685 7525 5715 7555
rect 5715 7525 5716 7555
rect 5684 7524 5716 7525
rect 5684 7475 5716 7476
rect 5684 7445 5685 7475
rect 5685 7445 5715 7475
rect 5715 7445 5716 7475
rect 5684 7444 5716 7445
rect 5684 7395 5716 7396
rect 5684 7365 5685 7395
rect 5685 7365 5715 7395
rect 5715 7365 5716 7395
rect 5684 7364 5716 7365
rect 5684 7315 5716 7316
rect 5684 7285 5685 7315
rect 5685 7285 5715 7315
rect 5715 7285 5716 7315
rect 5684 7284 5716 7285
rect 5684 7235 5716 7236
rect 5684 7205 5685 7235
rect 5685 7205 5715 7235
rect 5715 7205 5716 7235
rect 5684 7204 5716 7205
rect 5684 7155 5716 7156
rect 5684 7125 5685 7155
rect 5685 7125 5715 7155
rect 5715 7125 5716 7155
rect 5684 7124 5716 7125
rect 5684 7075 5716 7076
rect 5684 7045 5685 7075
rect 5685 7045 5715 7075
rect 5715 7045 5716 7075
rect 5684 7044 5716 7045
rect 5684 6995 5716 6996
rect 5684 6965 5685 6995
rect 5685 6965 5715 6995
rect 5715 6965 5716 6995
rect 5684 6964 5716 6965
rect 5684 6884 5716 6916
rect 5684 6835 5716 6836
rect 5684 6805 5685 6835
rect 5685 6805 5715 6835
rect 5715 6805 5716 6835
rect 5684 6804 5716 6805
rect 5684 6755 5716 6756
rect 5684 6725 5685 6755
rect 5685 6725 5715 6755
rect 5715 6725 5716 6755
rect 5684 6724 5716 6725
rect 5684 6675 5716 6676
rect 5684 6645 5685 6675
rect 5685 6645 5715 6675
rect 5715 6645 5716 6675
rect 5684 6644 5716 6645
rect 5684 6595 5716 6596
rect 5684 6565 5685 6595
rect 5685 6565 5715 6595
rect 5715 6565 5716 6595
rect 5684 6564 5716 6565
rect 5684 6515 5716 6516
rect 5684 6485 5685 6515
rect 5685 6485 5715 6515
rect 5715 6485 5716 6515
rect 5684 6484 5716 6485
rect 5684 6435 5716 6436
rect 5684 6405 5685 6435
rect 5685 6405 5715 6435
rect 5715 6405 5716 6435
rect 5684 6404 5716 6405
rect 5684 6355 5716 6356
rect 5684 6325 5685 6355
rect 5685 6325 5715 6355
rect 5715 6325 5716 6355
rect 5684 6324 5716 6325
rect 5684 6275 5716 6276
rect 5684 6245 5685 6275
rect 5685 6245 5715 6275
rect 5715 6245 5716 6275
rect 5684 6244 5716 6245
rect 5684 6164 5716 6196
rect 5684 6084 5716 6116
rect 5684 6004 5716 6036
rect 5684 5924 5716 5956
rect 5684 5875 5716 5876
rect 5684 5845 5685 5875
rect 5685 5845 5715 5875
rect 5715 5845 5716 5875
rect 5684 5844 5716 5845
rect 5684 5795 5716 5796
rect 5684 5765 5685 5795
rect 5685 5765 5715 5795
rect 5715 5765 5716 5795
rect 5684 5764 5716 5765
rect 5684 5715 5716 5716
rect 5684 5685 5685 5715
rect 5685 5685 5715 5715
rect 5715 5685 5716 5715
rect 5684 5684 5716 5685
rect 5684 5635 5716 5636
rect 5684 5605 5685 5635
rect 5685 5605 5715 5635
rect 5715 5605 5716 5635
rect 5684 5604 5716 5605
rect 5684 5555 5716 5556
rect 5684 5525 5685 5555
rect 5685 5525 5715 5555
rect 5715 5525 5716 5555
rect 5684 5524 5716 5525
rect 5684 5475 5716 5476
rect 5684 5445 5685 5475
rect 5685 5445 5715 5475
rect 5715 5445 5716 5475
rect 5684 5444 5716 5445
rect 5684 5395 5716 5396
rect 5684 5365 5685 5395
rect 5685 5365 5715 5395
rect 5715 5365 5716 5395
rect 5684 5364 5716 5365
rect 5684 5315 5716 5316
rect 5684 5285 5685 5315
rect 5685 5285 5715 5315
rect 5715 5285 5716 5315
rect 5684 5284 5716 5285
rect 5684 5235 5716 5236
rect 5684 5205 5685 5235
rect 5685 5205 5715 5235
rect 5715 5205 5716 5235
rect 5684 5204 5716 5205
rect 5684 5155 5716 5156
rect 5684 5125 5685 5155
rect 5685 5125 5715 5155
rect 5715 5125 5716 5155
rect 5684 5124 5716 5125
rect 5684 5075 5716 5076
rect 5684 5045 5685 5075
rect 5685 5045 5715 5075
rect 5715 5045 5716 5075
rect 5684 5044 5716 5045
rect 5684 4995 5716 4996
rect 5684 4965 5685 4995
rect 5685 4965 5715 4995
rect 5715 4965 5716 4995
rect 5684 4964 5716 4965
rect 5684 4915 5716 4916
rect 5684 4885 5685 4915
rect 5685 4885 5715 4915
rect 5715 4885 5716 4915
rect 5684 4884 5716 4885
rect 5684 4804 5716 4836
rect 5684 4755 5716 4756
rect 5684 4725 5685 4755
rect 5685 4725 5715 4755
rect 5715 4725 5716 4755
rect 5684 4724 5716 4725
rect 5684 4675 5716 4676
rect 5684 4645 5685 4675
rect 5685 4645 5715 4675
rect 5715 4645 5716 4675
rect 5684 4644 5716 4645
rect 5684 4564 5716 4596
rect 5684 4515 5716 4516
rect 5684 4485 5685 4515
rect 5685 4485 5715 4515
rect 5715 4485 5716 4515
rect 5684 4484 5716 4485
rect 5684 4435 5716 4436
rect 5684 4405 5685 4435
rect 5685 4405 5715 4435
rect 5715 4405 5716 4435
rect 5684 4404 5716 4405
rect 5684 4355 5716 4356
rect 5684 4325 5685 4355
rect 5685 4325 5715 4355
rect 5715 4325 5716 4355
rect 5684 4324 5716 4325
rect 5684 4275 5716 4276
rect 5684 4245 5685 4275
rect 5685 4245 5715 4275
rect 5715 4245 5716 4275
rect 5684 4244 5716 4245
rect 5684 4195 5716 4196
rect 5684 4165 5685 4195
rect 5685 4165 5715 4195
rect 5715 4165 5716 4195
rect 5684 4164 5716 4165
rect 5684 4115 5716 4116
rect 5684 4085 5685 4115
rect 5685 4085 5715 4115
rect 5715 4085 5716 4115
rect 5684 4084 5716 4085
rect 5684 4035 5716 4036
rect 5684 4005 5685 4035
rect 5685 4005 5715 4035
rect 5715 4005 5716 4035
rect 5684 4004 5716 4005
rect 5684 3955 5716 3956
rect 5684 3925 5685 3955
rect 5685 3925 5715 3955
rect 5715 3925 5716 3955
rect 5684 3924 5716 3925
rect 5684 3875 5716 3876
rect 5684 3845 5685 3875
rect 5685 3845 5715 3875
rect 5715 3845 5716 3875
rect 5684 3844 5716 3845
rect 5684 3764 5716 3796
rect 5684 3715 5716 3716
rect 5684 3685 5685 3715
rect 5685 3685 5715 3715
rect 5715 3685 5716 3715
rect 5684 3684 5716 3685
rect 5684 3635 5716 3636
rect 5684 3605 5685 3635
rect 5685 3605 5715 3635
rect 5715 3605 5716 3635
rect 5684 3604 5716 3605
rect 5684 3524 5716 3556
rect 5684 3475 5716 3476
rect 5684 3445 5685 3475
rect 5685 3445 5715 3475
rect 5715 3445 5716 3475
rect 5684 3444 5716 3445
rect 5684 3395 5716 3396
rect 5684 3365 5685 3395
rect 5685 3365 5715 3395
rect 5715 3365 5716 3395
rect 5684 3364 5716 3365
rect 5684 3284 5716 3316
rect 5684 3235 5716 3236
rect 5684 3205 5685 3235
rect 5685 3205 5715 3235
rect 5715 3205 5716 3235
rect 5684 3204 5716 3205
rect 5684 3155 5716 3156
rect 5684 3125 5685 3155
rect 5685 3125 5715 3155
rect 5715 3125 5716 3155
rect 5684 3124 5716 3125
rect 5684 3075 5716 3076
rect 5684 3045 5685 3075
rect 5685 3045 5715 3075
rect 5715 3045 5716 3075
rect 5684 3044 5716 3045
rect 5684 2995 5716 2996
rect 5684 2965 5685 2995
rect 5685 2965 5715 2995
rect 5715 2965 5716 2995
rect 5684 2964 5716 2965
rect 5684 2915 5716 2916
rect 5684 2885 5685 2915
rect 5685 2885 5715 2915
rect 5715 2885 5716 2915
rect 5684 2884 5716 2885
rect 5684 2835 5716 2836
rect 5684 2805 5685 2835
rect 5685 2805 5715 2835
rect 5715 2805 5716 2835
rect 5684 2804 5716 2805
rect 5684 2755 5716 2756
rect 5684 2725 5685 2755
rect 5685 2725 5715 2755
rect 5715 2725 5716 2755
rect 5684 2724 5716 2725
rect 5684 2675 5716 2676
rect 5684 2645 5685 2675
rect 5685 2645 5715 2675
rect 5715 2645 5716 2675
rect 5684 2644 5716 2645
rect 5684 2595 5716 2596
rect 5684 2565 5685 2595
rect 5685 2565 5715 2595
rect 5715 2565 5716 2595
rect 5684 2564 5716 2565
rect 5684 2515 5716 2516
rect 5684 2485 5685 2515
rect 5685 2485 5715 2515
rect 5715 2485 5716 2515
rect 5684 2484 5716 2485
rect 5684 2435 5716 2436
rect 5684 2405 5685 2435
rect 5685 2405 5715 2435
rect 5715 2405 5716 2435
rect 5684 2404 5716 2405
rect 5684 2355 5716 2356
rect 5684 2325 5685 2355
rect 5685 2325 5715 2355
rect 5715 2325 5716 2355
rect 5684 2324 5716 2325
rect 5684 2275 5716 2276
rect 5684 2245 5685 2275
rect 5685 2245 5715 2275
rect 5715 2245 5716 2275
rect 5684 2244 5716 2245
rect 5684 2195 5716 2196
rect 5684 2165 5685 2195
rect 5685 2165 5715 2195
rect 5715 2165 5716 2195
rect 5684 2164 5716 2165
rect 5684 2115 5716 2116
rect 5684 2085 5685 2115
rect 5685 2085 5715 2115
rect 5715 2085 5716 2115
rect 5684 2084 5716 2085
rect 5684 2035 5716 2036
rect 5684 2005 5685 2035
rect 5685 2005 5715 2035
rect 5715 2005 5716 2035
rect 5684 2004 5716 2005
rect 5684 1955 5716 1956
rect 5684 1925 5685 1955
rect 5685 1925 5715 1955
rect 5715 1925 5716 1955
rect 5684 1924 5716 1925
rect 5684 1844 5716 1876
rect 5684 1764 5716 1796
rect 5684 1715 5716 1716
rect 5684 1685 5685 1715
rect 5685 1685 5715 1715
rect 5715 1685 5716 1715
rect 5684 1684 5716 1685
rect 5684 1635 5716 1636
rect 5684 1605 5685 1635
rect 5685 1605 5715 1635
rect 5715 1605 5716 1635
rect 5684 1604 5716 1605
rect 5684 1555 5716 1556
rect 5684 1525 5685 1555
rect 5685 1525 5715 1555
rect 5715 1525 5716 1555
rect 5684 1524 5716 1525
rect 5684 1475 5716 1476
rect 5684 1445 5685 1475
rect 5685 1445 5715 1475
rect 5715 1445 5716 1475
rect 5684 1444 5716 1445
rect 5684 1395 5716 1396
rect 5684 1365 5685 1395
rect 5685 1365 5715 1395
rect 5715 1365 5716 1395
rect 5684 1364 5716 1365
rect 5684 1315 5716 1316
rect 5684 1285 5685 1315
rect 5685 1285 5715 1315
rect 5715 1285 5716 1315
rect 5684 1284 5716 1285
rect 5684 1235 5716 1236
rect 5684 1205 5685 1235
rect 5685 1205 5715 1235
rect 5715 1205 5716 1235
rect 5684 1204 5716 1205
rect 5684 1155 5716 1156
rect 5684 1125 5685 1155
rect 5685 1125 5715 1155
rect 5715 1125 5716 1155
rect 5684 1124 5716 1125
rect 5684 1075 5716 1076
rect 5684 1045 5685 1075
rect 5685 1045 5715 1075
rect 5715 1045 5716 1075
rect 5684 1044 5716 1045
rect 5684 995 5716 996
rect 5684 965 5685 995
rect 5685 965 5715 995
rect 5715 965 5716 995
rect 5684 964 5716 965
rect 5684 884 5716 916
rect 5684 835 5716 836
rect 5684 805 5685 835
rect 5685 805 5715 835
rect 5715 805 5716 835
rect 5684 804 5716 805
rect 5684 755 5716 756
rect 5684 725 5685 755
rect 5685 725 5715 755
rect 5715 725 5716 755
rect 5684 724 5716 725
rect 5684 675 5716 676
rect 5684 645 5685 675
rect 5685 645 5715 675
rect 5715 645 5716 675
rect 5684 644 5716 645
rect 5684 595 5716 596
rect 5684 565 5685 595
rect 5685 565 5715 595
rect 5715 565 5716 595
rect 5684 564 5716 565
rect 5684 515 5716 516
rect 5684 485 5685 515
rect 5685 485 5715 515
rect 5715 485 5716 515
rect 5684 484 5716 485
rect 5684 404 5716 436
rect 5684 324 5716 356
rect 5684 275 5716 276
rect 5684 245 5685 275
rect 5685 245 5715 275
rect 5715 245 5716 275
rect 5684 244 5716 245
rect 5684 195 5716 196
rect 5684 165 5685 195
rect 5685 165 5715 195
rect 5715 165 5716 195
rect 5684 164 5716 165
rect 5684 115 5716 116
rect 5684 85 5685 115
rect 5685 85 5715 115
rect 5715 85 5716 115
rect 5684 84 5716 85
rect 5684 35 5716 36
rect 5684 5 5685 35
rect 5685 5 5715 35
rect 5715 5 5716 35
rect 5684 4 5716 5
rect 5524 -716 5556 -524
rect 5684 -716 5716 -524
rect 5764 15715 5796 15716
rect 5764 15685 5765 15715
rect 5765 15685 5795 15715
rect 5795 15685 5796 15715
rect 5764 15684 5796 15685
rect 5764 15635 5796 15636
rect 5764 15605 5765 15635
rect 5765 15605 5795 15635
rect 5795 15605 5796 15635
rect 5764 15604 5796 15605
rect 5764 15555 5796 15556
rect 5764 15525 5765 15555
rect 5765 15525 5795 15555
rect 5795 15525 5796 15555
rect 5764 15524 5796 15525
rect 5764 15475 5796 15476
rect 5764 15445 5765 15475
rect 5765 15445 5795 15475
rect 5795 15445 5796 15475
rect 5764 15444 5796 15445
rect 5764 15395 5796 15396
rect 5764 15365 5765 15395
rect 5765 15365 5795 15395
rect 5795 15365 5796 15395
rect 5764 15364 5796 15365
rect 5764 15315 5796 15316
rect 5764 15285 5765 15315
rect 5765 15285 5795 15315
rect 5795 15285 5796 15315
rect 5764 15284 5796 15285
rect 5764 15235 5796 15236
rect 5764 15205 5765 15235
rect 5765 15205 5795 15235
rect 5795 15205 5796 15235
rect 5764 15204 5796 15205
rect 5764 15155 5796 15156
rect 5764 15125 5765 15155
rect 5765 15125 5795 15155
rect 5795 15125 5796 15155
rect 5764 15124 5796 15125
rect 5764 15044 5796 15076
rect 5764 14995 5796 14996
rect 5764 14965 5765 14995
rect 5765 14965 5795 14995
rect 5795 14965 5796 14995
rect 5764 14964 5796 14965
rect 5764 14915 5796 14916
rect 5764 14885 5765 14915
rect 5765 14885 5795 14915
rect 5795 14885 5796 14915
rect 5764 14884 5796 14885
rect 5764 14835 5796 14836
rect 5764 14805 5765 14835
rect 5765 14805 5795 14835
rect 5795 14805 5796 14835
rect 5764 14804 5796 14805
rect 5764 14755 5796 14756
rect 5764 14725 5765 14755
rect 5765 14725 5795 14755
rect 5795 14725 5796 14755
rect 5764 14724 5796 14725
rect 5764 14675 5796 14676
rect 5764 14645 5765 14675
rect 5765 14645 5795 14675
rect 5795 14645 5796 14675
rect 5764 14644 5796 14645
rect 5764 14595 5796 14596
rect 5764 14565 5765 14595
rect 5765 14565 5795 14595
rect 5795 14565 5796 14595
rect 5764 14564 5796 14565
rect 5764 14515 5796 14516
rect 5764 14485 5765 14515
rect 5765 14485 5795 14515
rect 5795 14485 5796 14515
rect 5764 14484 5796 14485
rect 5764 14435 5796 14436
rect 5764 14405 5765 14435
rect 5765 14405 5795 14435
rect 5795 14405 5796 14435
rect 5764 14404 5796 14405
rect 5764 14324 5796 14356
rect 5764 14244 5796 14276
rect 5764 14164 5796 14196
rect 5764 14084 5796 14116
rect 5764 14035 5796 14036
rect 5764 14005 5765 14035
rect 5765 14005 5795 14035
rect 5795 14005 5796 14035
rect 5764 14004 5796 14005
rect 5764 13955 5796 13956
rect 5764 13925 5765 13955
rect 5765 13925 5795 13955
rect 5795 13925 5796 13955
rect 5764 13924 5796 13925
rect 5764 13875 5796 13876
rect 5764 13845 5765 13875
rect 5765 13845 5795 13875
rect 5795 13845 5796 13875
rect 5764 13844 5796 13845
rect 5764 13795 5796 13796
rect 5764 13765 5765 13795
rect 5765 13765 5795 13795
rect 5795 13765 5796 13795
rect 5764 13764 5796 13765
rect 5764 13715 5796 13716
rect 5764 13685 5765 13715
rect 5765 13685 5795 13715
rect 5795 13685 5796 13715
rect 5764 13684 5796 13685
rect 5764 13635 5796 13636
rect 5764 13605 5765 13635
rect 5765 13605 5795 13635
rect 5795 13605 5796 13635
rect 5764 13604 5796 13605
rect 5764 13555 5796 13556
rect 5764 13525 5765 13555
rect 5765 13525 5795 13555
rect 5795 13525 5796 13555
rect 5764 13524 5796 13525
rect 5764 13475 5796 13476
rect 5764 13445 5765 13475
rect 5765 13445 5795 13475
rect 5795 13445 5796 13475
rect 5764 13444 5796 13445
rect 5764 13364 5796 13396
rect 5764 13284 5796 13316
rect 5764 13204 5796 13236
rect 5764 13124 5796 13156
rect 5764 13075 5796 13076
rect 5764 13045 5765 13075
rect 5765 13045 5795 13075
rect 5795 13045 5796 13075
rect 5764 13044 5796 13045
rect 5764 12995 5796 12996
rect 5764 12965 5765 12995
rect 5765 12965 5795 12995
rect 5795 12965 5796 12995
rect 5764 12964 5796 12965
rect 5764 12915 5796 12916
rect 5764 12885 5765 12915
rect 5765 12885 5795 12915
rect 5795 12885 5796 12915
rect 5764 12884 5796 12885
rect 5764 12835 5796 12836
rect 5764 12805 5765 12835
rect 5765 12805 5795 12835
rect 5795 12805 5796 12835
rect 5764 12804 5796 12805
rect 5764 12755 5796 12756
rect 5764 12725 5765 12755
rect 5765 12725 5795 12755
rect 5795 12725 5796 12755
rect 5764 12724 5796 12725
rect 5764 12675 5796 12676
rect 5764 12645 5765 12675
rect 5765 12645 5795 12675
rect 5795 12645 5796 12675
rect 5764 12644 5796 12645
rect 5764 12595 5796 12596
rect 5764 12565 5765 12595
rect 5765 12565 5795 12595
rect 5795 12565 5796 12595
rect 5764 12564 5796 12565
rect 5764 12515 5796 12516
rect 5764 12485 5765 12515
rect 5765 12485 5795 12515
rect 5795 12485 5796 12515
rect 5764 12484 5796 12485
rect 5764 12404 5796 12436
rect 5764 12355 5796 12356
rect 5764 12325 5765 12355
rect 5765 12325 5795 12355
rect 5795 12325 5796 12355
rect 5764 12324 5796 12325
rect 5764 12275 5796 12276
rect 5764 12245 5765 12275
rect 5765 12245 5795 12275
rect 5795 12245 5796 12275
rect 5764 12244 5796 12245
rect 5764 12195 5796 12196
rect 5764 12165 5765 12195
rect 5765 12165 5795 12195
rect 5795 12165 5796 12195
rect 5764 12164 5796 12165
rect 5764 12115 5796 12116
rect 5764 12085 5765 12115
rect 5765 12085 5795 12115
rect 5795 12085 5796 12115
rect 5764 12084 5796 12085
rect 5764 12035 5796 12036
rect 5764 12005 5765 12035
rect 5765 12005 5795 12035
rect 5795 12005 5796 12035
rect 5764 12004 5796 12005
rect 5764 11955 5796 11956
rect 5764 11925 5765 11955
rect 5765 11925 5795 11955
rect 5795 11925 5796 11955
rect 5764 11924 5796 11925
rect 5764 11875 5796 11876
rect 5764 11845 5765 11875
rect 5765 11845 5795 11875
rect 5795 11845 5796 11875
rect 5764 11844 5796 11845
rect 5764 11795 5796 11796
rect 5764 11765 5765 11795
rect 5765 11765 5795 11795
rect 5795 11765 5796 11795
rect 5764 11764 5796 11765
rect 5764 11715 5796 11716
rect 5764 11685 5765 11715
rect 5765 11685 5795 11715
rect 5795 11685 5796 11715
rect 5764 11684 5796 11685
rect 5764 11635 5796 11636
rect 5764 11605 5765 11635
rect 5765 11605 5795 11635
rect 5795 11605 5796 11635
rect 5764 11604 5796 11605
rect 5764 11555 5796 11556
rect 5764 11525 5765 11555
rect 5765 11525 5795 11555
rect 5795 11525 5796 11555
rect 5764 11524 5796 11525
rect 5764 11475 5796 11476
rect 5764 11445 5765 11475
rect 5765 11445 5795 11475
rect 5795 11445 5796 11475
rect 5764 11444 5796 11445
rect 5764 11395 5796 11396
rect 5764 11365 5765 11395
rect 5765 11365 5795 11395
rect 5795 11365 5796 11395
rect 5764 11364 5796 11365
rect 5764 11315 5796 11316
rect 5764 11285 5765 11315
rect 5765 11285 5795 11315
rect 5795 11285 5796 11315
rect 5764 11284 5796 11285
rect 5764 11235 5796 11236
rect 5764 11205 5765 11235
rect 5765 11205 5795 11235
rect 5795 11205 5796 11235
rect 5764 11204 5796 11205
rect 5764 11155 5796 11156
rect 5764 11125 5765 11155
rect 5765 11125 5795 11155
rect 5795 11125 5796 11155
rect 5764 11124 5796 11125
rect 5764 11075 5796 11076
rect 5764 11045 5765 11075
rect 5765 11045 5795 11075
rect 5795 11045 5796 11075
rect 5764 11044 5796 11045
rect 5764 10964 5796 10996
rect 5764 10915 5796 10916
rect 5764 10885 5765 10915
rect 5765 10885 5795 10915
rect 5795 10885 5796 10915
rect 5764 10884 5796 10885
rect 5764 10835 5796 10836
rect 5764 10805 5765 10835
rect 5765 10805 5795 10835
rect 5795 10805 5796 10835
rect 5764 10804 5796 10805
rect 5764 10755 5796 10756
rect 5764 10725 5765 10755
rect 5765 10725 5795 10755
rect 5795 10725 5796 10755
rect 5764 10724 5796 10725
rect 5764 10675 5796 10676
rect 5764 10645 5765 10675
rect 5765 10645 5795 10675
rect 5795 10645 5796 10675
rect 5764 10644 5796 10645
rect 5764 10595 5796 10596
rect 5764 10565 5765 10595
rect 5765 10565 5795 10595
rect 5795 10565 5796 10595
rect 5764 10564 5796 10565
rect 5764 10515 5796 10516
rect 5764 10485 5765 10515
rect 5765 10485 5795 10515
rect 5795 10485 5796 10515
rect 5764 10484 5796 10485
rect 5764 10435 5796 10436
rect 5764 10405 5765 10435
rect 5765 10405 5795 10435
rect 5795 10405 5796 10435
rect 5764 10404 5796 10405
rect 5764 10355 5796 10356
rect 5764 10325 5765 10355
rect 5765 10325 5795 10355
rect 5795 10325 5796 10355
rect 5764 10324 5796 10325
rect 5764 10244 5796 10276
rect 5764 10164 5796 10196
rect 5764 10084 5796 10116
rect 5764 10004 5796 10036
rect 5764 9955 5796 9956
rect 5764 9925 5765 9955
rect 5765 9925 5795 9955
rect 5795 9925 5796 9955
rect 5764 9924 5796 9925
rect 5764 9875 5796 9876
rect 5764 9845 5765 9875
rect 5765 9845 5795 9875
rect 5795 9845 5796 9875
rect 5764 9844 5796 9845
rect 5764 9795 5796 9796
rect 5764 9765 5765 9795
rect 5765 9765 5795 9795
rect 5795 9765 5796 9795
rect 5764 9764 5796 9765
rect 5764 9715 5796 9716
rect 5764 9685 5765 9715
rect 5765 9685 5795 9715
rect 5795 9685 5796 9715
rect 5764 9684 5796 9685
rect 5764 9635 5796 9636
rect 5764 9605 5765 9635
rect 5765 9605 5795 9635
rect 5795 9605 5796 9635
rect 5764 9604 5796 9605
rect 5764 9555 5796 9556
rect 5764 9525 5765 9555
rect 5765 9525 5795 9555
rect 5795 9525 5796 9555
rect 5764 9524 5796 9525
rect 5764 9475 5796 9476
rect 5764 9445 5765 9475
rect 5765 9445 5795 9475
rect 5795 9445 5796 9475
rect 5764 9444 5796 9445
rect 5764 9395 5796 9396
rect 5764 9365 5765 9395
rect 5765 9365 5795 9395
rect 5795 9365 5796 9395
rect 5764 9364 5796 9365
rect 5764 9284 5796 9316
rect 5764 9204 5796 9236
rect 5764 9124 5796 9156
rect 5764 9044 5796 9076
rect 5764 8995 5796 8996
rect 5764 8965 5765 8995
rect 5765 8965 5795 8995
rect 5795 8965 5796 8995
rect 5764 8964 5796 8965
rect 5764 8915 5796 8916
rect 5764 8885 5765 8915
rect 5765 8885 5795 8915
rect 5795 8885 5796 8915
rect 5764 8884 5796 8885
rect 5764 8835 5796 8836
rect 5764 8805 5765 8835
rect 5765 8805 5795 8835
rect 5795 8805 5796 8835
rect 5764 8804 5796 8805
rect 5764 8755 5796 8756
rect 5764 8725 5765 8755
rect 5765 8725 5795 8755
rect 5795 8725 5796 8755
rect 5764 8724 5796 8725
rect 5764 8675 5796 8676
rect 5764 8645 5765 8675
rect 5765 8645 5795 8675
rect 5795 8645 5796 8675
rect 5764 8644 5796 8645
rect 5764 8595 5796 8596
rect 5764 8565 5765 8595
rect 5765 8565 5795 8595
rect 5795 8565 5796 8595
rect 5764 8564 5796 8565
rect 5764 8515 5796 8516
rect 5764 8485 5765 8515
rect 5765 8485 5795 8515
rect 5795 8485 5796 8515
rect 5764 8484 5796 8485
rect 5764 8435 5796 8436
rect 5764 8405 5765 8435
rect 5765 8405 5795 8435
rect 5795 8405 5796 8435
rect 5764 8404 5796 8405
rect 5764 8324 5796 8356
rect 5764 8275 5796 8276
rect 5764 8245 5765 8275
rect 5765 8245 5795 8275
rect 5795 8245 5796 8275
rect 5764 8244 5796 8245
rect 5764 8195 5796 8196
rect 5764 8165 5765 8195
rect 5765 8165 5795 8195
rect 5795 8165 5796 8195
rect 5764 8164 5796 8165
rect 5764 8115 5796 8116
rect 5764 8085 5765 8115
rect 5765 8085 5795 8115
rect 5795 8085 5796 8115
rect 5764 8084 5796 8085
rect 5764 8035 5796 8036
rect 5764 8005 5765 8035
rect 5765 8005 5795 8035
rect 5795 8005 5796 8035
rect 5764 8004 5796 8005
rect 5764 7955 5796 7956
rect 5764 7925 5765 7955
rect 5765 7925 5795 7955
rect 5795 7925 5796 7955
rect 5764 7924 5796 7925
rect 5764 7875 5796 7876
rect 5764 7845 5765 7875
rect 5765 7845 5795 7875
rect 5795 7845 5796 7875
rect 5764 7844 5796 7845
rect 5764 7795 5796 7796
rect 5764 7765 5765 7795
rect 5765 7765 5795 7795
rect 5795 7765 5796 7795
rect 5764 7764 5796 7765
rect 5764 7715 5796 7716
rect 5764 7685 5765 7715
rect 5765 7685 5795 7715
rect 5795 7685 5796 7715
rect 5764 7684 5796 7685
rect 5764 7635 5796 7636
rect 5764 7605 5765 7635
rect 5765 7605 5795 7635
rect 5795 7605 5796 7635
rect 5764 7604 5796 7605
rect 5764 7555 5796 7556
rect 5764 7525 5765 7555
rect 5765 7525 5795 7555
rect 5795 7525 5796 7555
rect 5764 7524 5796 7525
rect 5764 7475 5796 7476
rect 5764 7445 5765 7475
rect 5765 7445 5795 7475
rect 5795 7445 5796 7475
rect 5764 7444 5796 7445
rect 5764 7395 5796 7396
rect 5764 7365 5765 7395
rect 5765 7365 5795 7395
rect 5795 7365 5796 7395
rect 5764 7364 5796 7365
rect 5764 7315 5796 7316
rect 5764 7285 5765 7315
rect 5765 7285 5795 7315
rect 5795 7285 5796 7315
rect 5764 7284 5796 7285
rect 5764 7235 5796 7236
rect 5764 7205 5765 7235
rect 5765 7205 5795 7235
rect 5795 7205 5796 7235
rect 5764 7204 5796 7205
rect 5764 7155 5796 7156
rect 5764 7125 5765 7155
rect 5765 7125 5795 7155
rect 5795 7125 5796 7155
rect 5764 7124 5796 7125
rect 5764 7075 5796 7076
rect 5764 7045 5765 7075
rect 5765 7045 5795 7075
rect 5795 7045 5796 7075
rect 5764 7044 5796 7045
rect 5764 6995 5796 6996
rect 5764 6965 5765 6995
rect 5765 6965 5795 6995
rect 5795 6965 5796 6995
rect 5764 6964 5796 6965
rect 5764 6884 5796 6916
rect 5764 6835 5796 6836
rect 5764 6805 5765 6835
rect 5765 6805 5795 6835
rect 5795 6805 5796 6835
rect 5764 6804 5796 6805
rect 5764 6755 5796 6756
rect 5764 6725 5765 6755
rect 5765 6725 5795 6755
rect 5795 6725 5796 6755
rect 5764 6724 5796 6725
rect 5764 6675 5796 6676
rect 5764 6645 5765 6675
rect 5765 6645 5795 6675
rect 5795 6645 5796 6675
rect 5764 6644 5796 6645
rect 5764 6595 5796 6596
rect 5764 6565 5765 6595
rect 5765 6565 5795 6595
rect 5795 6565 5796 6595
rect 5764 6564 5796 6565
rect 5764 6515 5796 6516
rect 5764 6485 5765 6515
rect 5765 6485 5795 6515
rect 5795 6485 5796 6515
rect 5764 6484 5796 6485
rect 5764 6435 5796 6436
rect 5764 6405 5765 6435
rect 5765 6405 5795 6435
rect 5795 6405 5796 6435
rect 5764 6404 5796 6405
rect 5764 6355 5796 6356
rect 5764 6325 5765 6355
rect 5765 6325 5795 6355
rect 5795 6325 5796 6355
rect 5764 6324 5796 6325
rect 5764 6275 5796 6276
rect 5764 6245 5765 6275
rect 5765 6245 5795 6275
rect 5795 6245 5796 6275
rect 5764 6244 5796 6245
rect 5764 6164 5796 6196
rect 5764 6084 5796 6116
rect 5764 6004 5796 6036
rect 5764 5924 5796 5956
rect 5764 5875 5796 5876
rect 5764 5845 5765 5875
rect 5765 5845 5795 5875
rect 5795 5845 5796 5875
rect 5764 5844 5796 5845
rect 5764 5795 5796 5796
rect 5764 5765 5765 5795
rect 5765 5765 5795 5795
rect 5795 5765 5796 5795
rect 5764 5764 5796 5765
rect 5764 5715 5796 5716
rect 5764 5685 5765 5715
rect 5765 5685 5795 5715
rect 5795 5685 5796 5715
rect 5764 5684 5796 5685
rect 5764 5635 5796 5636
rect 5764 5605 5765 5635
rect 5765 5605 5795 5635
rect 5795 5605 5796 5635
rect 5764 5604 5796 5605
rect 5764 5555 5796 5556
rect 5764 5525 5765 5555
rect 5765 5525 5795 5555
rect 5795 5525 5796 5555
rect 5764 5524 5796 5525
rect 5764 5475 5796 5476
rect 5764 5445 5765 5475
rect 5765 5445 5795 5475
rect 5795 5445 5796 5475
rect 5764 5444 5796 5445
rect 5764 5395 5796 5396
rect 5764 5365 5765 5395
rect 5765 5365 5795 5395
rect 5795 5365 5796 5395
rect 5764 5364 5796 5365
rect 5764 5315 5796 5316
rect 5764 5285 5765 5315
rect 5765 5285 5795 5315
rect 5795 5285 5796 5315
rect 5764 5284 5796 5285
rect 5764 5235 5796 5236
rect 5764 5205 5765 5235
rect 5765 5205 5795 5235
rect 5795 5205 5796 5235
rect 5764 5204 5796 5205
rect 5764 5155 5796 5156
rect 5764 5125 5765 5155
rect 5765 5125 5795 5155
rect 5795 5125 5796 5155
rect 5764 5124 5796 5125
rect 5764 5075 5796 5076
rect 5764 5045 5765 5075
rect 5765 5045 5795 5075
rect 5795 5045 5796 5075
rect 5764 5044 5796 5045
rect 5764 4995 5796 4996
rect 5764 4965 5765 4995
rect 5765 4965 5795 4995
rect 5795 4965 5796 4995
rect 5764 4964 5796 4965
rect 5764 4915 5796 4916
rect 5764 4885 5765 4915
rect 5765 4885 5795 4915
rect 5795 4885 5796 4915
rect 5764 4884 5796 4885
rect 5764 4804 5796 4836
rect 5764 4755 5796 4756
rect 5764 4725 5765 4755
rect 5765 4725 5795 4755
rect 5795 4725 5796 4755
rect 5764 4724 5796 4725
rect 5764 4675 5796 4676
rect 5764 4645 5765 4675
rect 5765 4645 5795 4675
rect 5795 4645 5796 4675
rect 5764 4644 5796 4645
rect 5764 4564 5796 4596
rect 5764 4515 5796 4516
rect 5764 4485 5765 4515
rect 5765 4485 5795 4515
rect 5795 4485 5796 4515
rect 5764 4484 5796 4485
rect 5764 4435 5796 4436
rect 5764 4405 5765 4435
rect 5765 4405 5795 4435
rect 5795 4405 5796 4435
rect 5764 4404 5796 4405
rect 5764 4355 5796 4356
rect 5764 4325 5765 4355
rect 5765 4325 5795 4355
rect 5795 4325 5796 4355
rect 5764 4324 5796 4325
rect 5764 4275 5796 4276
rect 5764 4245 5765 4275
rect 5765 4245 5795 4275
rect 5795 4245 5796 4275
rect 5764 4244 5796 4245
rect 5764 4195 5796 4196
rect 5764 4165 5765 4195
rect 5765 4165 5795 4195
rect 5795 4165 5796 4195
rect 5764 4164 5796 4165
rect 5764 4115 5796 4116
rect 5764 4085 5765 4115
rect 5765 4085 5795 4115
rect 5795 4085 5796 4115
rect 5764 4084 5796 4085
rect 5764 4035 5796 4036
rect 5764 4005 5765 4035
rect 5765 4005 5795 4035
rect 5795 4005 5796 4035
rect 5764 4004 5796 4005
rect 5764 3955 5796 3956
rect 5764 3925 5765 3955
rect 5765 3925 5795 3955
rect 5795 3925 5796 3955
rect 5764 3924 5796 3925
rect 5764 3875 5796 3876
rect 5764 3845 5765 3875
rect 5765 3845 5795 3875
rect 5795 3845 5796 3875
rect 5764 3844 5796 3845
rect 5764 3764 5796 3796
rect 5764 3715 5796 3716
rect 5764 3685 5765 3715
rect 5765 3685 5795 3715
rect 5795 3685 5796 3715
rect 5764 3684 5796 3685
rect 5764 3635 5796 3636
rect 5764 3605 5765 3635
rect 5765 3605 5795 3635
rect 5795 3605 5796 3635
rect 5764 3604 5796 3605
rect 5764 3524 5796 3556
rect 5764 3475 5796 3476
rect 5764 3445 5765 3475
rect 5765 3445 5795 3475
rect 5795 3445 5796 3475
rect 5764 3444 5796 3445
rect 5764 3395 5796 3396
rect 5764 3365 5765 3395
rect 5765 3365 5795 3395
rect 5795 3365 5796 3395
rect 5764 3364 5796 3365
rect 5764 3284 5796 3316
rect 5764 3235 5796 3236
rect 5764 3205 5765 3235
rect 5765 3205 5795 3235
rect 5795 3205 5796 3235
rect 5764 3204 5796 3205
rect 5764 3155 5796 3156
rect 5764 3125 5765 3155
rect 5765 3125 5795 3155
rect 5795 3125 5796 3155
rect 5764 3124 5796 3125
rect 5764 3075 5796 3076
rect 5764 3045 5765 3075
rect 5765 3045 5795 3075
rect 5795 3045 5796 3075
rect 5764 3044 5796 3045
rect 5764 2995 5796 2996
rect 5764 2965 5765 2995
rect 5765 2965 5795 2995
rect 5795 2965 5796 2995
rect 5764 2964 5796 2965
rect 5764 2915 5796 2916
rect 5764 2885 5765 2915
rect 5765 2885 5795 2915
rect 5795 2885 5796 2915
rect 5764 2884 5796 2885
rect 5764 2835 5796 2836
rect 5764 2805 5765 2835
rect 5765 2805 5795 2835
rect 5795 2805 5796 2835
rect 5764 2804 5796 2805
rect 5764 2755 5796 2756
rect 5764 2725 5765 2755
rect 5765 2725 5795 2755
rect 5795 2725 5796 2755
rect 5764 2724 5796 2725
rect 5764 2675 5796 2676
rect 5764 2645 5765 2675
rect 5765 2645 5795 2675
rect 5795 2645 5796 2675
rect 5764 2644 5796 2645
rect 5764 2595 5796 2596
rect 5764 2565 5765 2595
rect 5765 2565 5795 2595
rect 5795 2565 5796 2595
rect 5764 2564 5796 2565
rect 5764 2515 5796 2516
rect 5764 2485 5765 2515
rect 5765 2485 5795 2515
rect 5795 2485 5796 2515
rect 5764 2484 5796 2485
rect 5764 2435 5796 2436
rect 5764 2405 5765 2435
rect 5765 2405 5795 2435
rect 5795 2405 5796 2435
rect 5764 2404 5796 2405
rect 5764 2355 5796 2356
rect 5764 2325 5765 2355
rect 5765 2325 5795 2355
rect 5795 2325 5796 2355
rect 5764 2324 5796 2325
rect 5764 2275 5796 2276
rect 5764 2245 5765 2275
rect 5765 2245 5795 2275
rect 5795 2245 5796 2275
rect 5764 2244 5796 2245
rect 5764 2195 5796 2196
rect 5764 2165 5765 2195
rect 5765 2165 5795 2195
rect 5795 2165 5796 2195
rect 5764 2164 5796 2165
rect 5764 2115 5796 2116
rect 5764 2085 5765 2115
rect 5765 2085 5795 2115
rect 5795 2085 5796 2115
rect 5764 2084 5796 2085
rect 5764 2035 5796 2036
rect 5764 2005 5765 2035
rect 5765 2005 5795 2035
rect 5795 2005 5796 2035
rect 5764 2004 5796 2005
rect 5764 1955 5796 1956
rect 5764 1925 5765 1955
rect 5765 1925 5795 1955
rect 5795 1925 5796 1955
rect 5764 1924 5796 1925
rect 5764 1844 5796 1876
rect 5764 1764 5796 1796
rect 5764 1715 5796 1716
rect 5764 1685 5765 1715
rect 5765 1685 5795 1715
rect 5795 1685 5796 1715
rect 5764 1684 5796 1685
rect 5764 1635 5796 1636
rect 5764 1605 5765 1635
rect 5765 1605 5795 1635
rect 5795 1605 5796 1635
rect 5764 1604 5796 1605
rect 5764 1555 5796 1556
rect 5764 1525 5765 1555
rect 5765 1525 5795 1555
rect 5795 1525 5796 1555
rect 5764 1524 5796 1525
rect 5764 1475 5796 1476
rect 5764 1445 5765 1475
rect 5765 1445 5795 1475
rect 5795 1445 5796 1475
rect 5764 1444 5796 1445
rect 5764 1395 5796 1396
rect 5764 1365 5765 1395
rect 5765 1365 5795 1395
rect 5795 1365 5796 1395
rect 5764 1364 5796 1365
rect 5764 1315 5796 1316
rect 5764 1285 5765 1315
rect 5765 1285 5795 1315
rect 5795 1285 5796 1315
rect 5764 1284 5796 1285
rect 5764 1235 5796 1236
rect 5764 1205 5765 1235
rect 5765 1205 5795 1235
rect 5795 1205 5796 1235
rect 5764 1204 5796 1205
rect 5764 1155 5796 1156
rect 5764 1125 5765 1155
rect 5765 1125 5795 1155
rect 5795 1125 5796 1155
rect 5764 1124 5796 1125
rect 5764 1075 5796 1076
rect 5764 1045 5765 1075
rect 5765 1045 5795 1075
rect 5795 1045 5796 1075
rect 5764 1044 5796 1045
rect 5764 995 5796 996
rect 5764 965 5765 995
rect 5765 965 5795 995
rect 5795 965 5796 995
rect 5764 964 5796 965
rect 5764 884 5796 916
rect 5764 835 5796 836
rect 5764 805 5765 835
rect 5765 805 5795 835
rect 5795 805 5796 835
rect 5764 804 5796 805
rect 5764 755 5796 756
rect 5764 725 5765 755
rect 5765 725 5795 755
rect 5795 725 5796 755
rect 5764 724 5796 725
rect 5764 675 5796 676
rect 5764 645 5765 675
rect 5765 645 5795 675
rect 5795 645 5796 675
rect 5764 644 5796 645
rect 5764 595 5796 596
rect 5764 565 5765 595
rect 5765 565 5795 595
rect 5795 565 5796 595
rect 5764 564 5796 565
rect 5764 515 5796 516
rect 5764 485 5765 515
rect 5765 485 5795 515
rect 5795 485 5796 515
rect 5764 484 5796 485
rect 5764 404 5796 436
rect 5764 324 5796 356
rect 5764 275 5796 276
rect 5764 245 5765 275
rect 5765 245 5795 275
rect 5795 245 5796 275
rect 5764 244 5796 245
rect 5764 195 5796 196
rect 5764 165 5765 195
rect 5765 165 5795 195
rect 5795 165 5796 195
rect 5764 164 5796 165
rect 5764 115 5796 116
rect 5764 85 5765 115
rect 5765 85 5795 115
rect 5795 85 5796 115
rect 5764 84 5796 85
rect 5764 35 5796 36
rect 5764 5 5765 35
rect 5765 5 5795 35
rect 5795 5 5796 35
rect 5764 4 5796 5
rect 5924 15715 5956 15716
rect 5924 15685 5925 15715
rect 5925 15685 5955 15715
rect 5955 15685 5956 15715
rect 5924 15684 5956 15685
rect 5924 15635 5956 15636
rect 5924 15605 5925 15635
rect 5925 15605 5955 15635
rect 5955 15605 5956 15635
rect 5924 15604 5956 15605
rect 5924 15555 5956 15556
rect 5924 15525 5925 15555
rect 5925 15525 5955 15555
rect 5955 15525 5956 15555
rect 5924 15524 5956 15525
rect 5924 15475 5956 15476
rect 5924 15445 5925 15475
rect 5925 15445 5955 15475
rect 5955 15445 5956 15475
rect 5924 15444 5956 15445
rect 5924 15395 5956 15396
rect 5924 15365 5925 15395
rect 5925 15365 5955 15395
rect 5955 15365 5956 15395
rect 5924 15364 5956 15365
rect 5924 15315 5956 15316
rect 5924 15285 5925 15315
rect 5925 15285 5955 15315
rect 5955 15285 5956 15315
rect 5924 15284 5956 15285
rect 5924 15235 5956 15236
rect 5924 15205 5925 15235
rect 5925 15205 5955 15235
rect 5955 15205 5956 15235
rect 5924 15204 5956 15205
rect 5924 15155 5956 15156
rect 5924 15125 5925 15155
rect 5925 15125 5955 15155
rect 5955 15125 5956 15155
rect 5924 15124 5956 15125
rect 5924 15044 5956 15076
rect 5924 14995 5956 14996
rect 5924 14965 5925 14995
rect 5925 14965 5955 14995
rect 5955 14965 5956 14995
rect 5924 14964 5956 14965
rect 5924 14915 5956 14916
rect 5924 14885 5925 14915
rect 5925 14885 5955 14915
rect 5955 14885 5956 14915
rect 5924 14884 5956 14885
rect 5924 14835 5956 14836
rect 5924 14805 5925 14835
rect 5925 14805 5955 14835
rect 5955 14805 5956 14835
rect 5924 14804 5956 14805
rect 5924 14755 5956 14756
rect 5924 14725 5925 14755
rect 5925 14725 5955 14755
rect 5955 14725 5956 14755
rect 5924 14724 5956 14725
rect 5924 14675 5956 14676
rect 5924 14645 5925 14675
rect 5925 14645 5955 14675
rect 5955 14645 5956 14675
rect 5924 14644 5956 14645
rect 5924 14595 5956 14596
rect 5924 14565 5925 14595
rect 5925 14565 5955 14595
rect 5955 14565 5956 14595
rect 5924 14564 5956 14565
rect 5924 14515 5956 14516
rect 5924 14485 5925 14515
rect 5925 14485 5955 14515
rect 5955 14485 5956 14515
rect 5924 14484 5956 14485
rect 5924 14435 5956 14436
rect 5924 14405 5925 14435
rect 5925 14405 5955 14435
rect 5955 14405 5956 14435
rect 5924 14404 5956 14405
rect 5924 14324 5956 14356
rect 5924 14244 5956 14276
rect 5924 14164 5956 14196
rect 5924 14084 5956 14116
rect 5924 14035 5956 14036
rect 5924 14005 5925 14035
rect 5925 14005 5955 14035
rect 5955 14005 5956 14035
rect 5924 14004 5956 14005
rect 5924 13955 5956 13956
rect 5924 13925 5925 13955
rect 5925 13925 5955 13955
rect 5955 13925 5956 13955
rect 5924 13924 5956 13925
rect 5924 13875 5956 13876
rect 5924 13845 5925 13875
rect 5925 13845 5955 13875
rect 5955 13845 5956 13875
rect 5924 13844 5956 13845
rect 5924 13795 5956 13796
rect 5924 13765 5925 13795
rect 5925 13765 5955 13795
rect 5955 13765 5956 13795
rect 5924 13764 5956 13765
rect 5924 13715 5956 13716
rect 5924 13685 5925 13715
rect 5925 13685 5955 13715
rect 5955 13685 5956 13715
rect 5924 13684 5956 13685
rect 5924 13635 5956 13636
rect 5924 13605 5925 13635
rect 5925 13605 5955 13635
rect 5955 13605 5956 13635
rect 5924 13604 5956 13605
rect 5924 13555 5956 13556
rect 5924 13525 5925 13555
rect 5925 13525 5955 13555
rect 5955 13525 5956 13555
rect 5924 13524 5956 13525
rect 5924 13475 5956 13476
rect 5924 13445 5925 13475
rect 5925 13445 5955 13475
rect 5955 13445 5956 13475
rect 5924 13444 5956 13445
rect 5924 13364 5956 13396
rect 5924 13284 5956 13316
rect 5924 13204 5956 13236
rect 5924 13124 5956 13156
rect 5924 13075 5956 13076
rect 5924 13045 5925 13075
rect 5925 13045 5955 13075
rect 5955 13045 5956 13075
rect 5924 13044 5956 13045
rect 5924 12995 5956 12996
rect 5924 12965 5925 12995
rect 5925 12965 5955 12995
rect 5955 12965 5956 12995
rect 5924 12964 5956 12965
rect 5924 12915 5956 12916
rect 5924 12885 5925 12915
rect 5925 12885 5955 12915
rect 5955 12885 5956 12915
rect 5924 12884 5956 12885
rect 5924 12835 5956 12836
rect 5924 12805 5925 12835
rect 5925 12805 5955 12835
rect 5955 12805 5956 12835
rect 5924 12804 5956 12805
rect 5924 12755 5956 12756
rect 5924 12725 5925 12755
rect 5925 12725 5955 12755
rect 5955 12725 5956 12755
rect 5924 12724 5956 12725
rect 5924 12675 5956 12676
rect 5924 12645 5925 12675
rect 5925 12645 5955 12675
rect 5955 12645 5956 12675
rect 5924 12644 5956 12645
rect 5924 12595 5956 12596
rect 5924 12565 5925 12595
rect 5925 12565 5955 12595
rect 5955 12565 5956 12595
rect 5924 12564 5956 12565
rect 5924 12515 5956 12516
rect 5924 12485 5925 12515
rect 5925 12485 5955 12515
rect 5955 12485 5956 12515
rect 5924 12484 5956 12485
rect 5924 12404 5956 12436
rect 5924 12355 5956 12356
rect 5924 12325 5925 12355
rect 5925 12325 5955 12355
rect 5955 12325 5956 12355
rect 5924 12324 5956 12325
rect 5924 12275 5956 12276
rect 5924 12245 5925 12275
rect 5925 12245 5955 12275
rect 5955 12245 5956 12275
rect 5924 12244 5956 12245
rect 5924 12195 5956 12196
rect 5924 12165 5925 12195
rect 5925 12165 5955 12195
rect 5955 12165 5956 12195
rect 5924 12164 5956 12165
rect 5924 12115 5956 12116
rect 5924 12085 5925 12115
rect 5925 12085 5955 12115
rect 5955 12085 5956 12115
rect 5924 12084 5956 12085
rect 5924 12035 5956 12036
rect 5924 12005 5925 12035
rect 5925 12005 5955 12035
rect 5955 12005 5956 12035
rect 5924 12004 5956 12005
rect 5924 11955 5956 11956
rect 5924 11925 5925 11955
rect 5925 11925 5955 11955
rect 5955 11925 5956 11955
rect 5924 11924 5956 11925
rect 5924 11875 5956 11876
rect 5924 11845 5925 11875
rect 5925 11845 5955 11875
rect 5955 11845 5956 11875
rect 5924 11844 5956 11845
rect 5924 11795 5956 11796
rect 5924 11765 5925 11795
rect 5925 11765 5955 11795
rect 5955 11765 5956 11795
rect 5924 11764 5956 11765
rect 5924 11715 5956 11716
rect 5924 11685 5925 11715
rect 5925 11685 5955 11715
rect 5955 11685 5956 11715
rect 5924 11684 5956 11685
rect 5924 11635 5956 11636
rect 5924 11605 5925 11635
rect 5925 11605 5955 11635
rect 5955 11605 5956 11635
rect 5924 11604 5956 11605
rect 5924 11555 5956 11556
rect 5924 11525 5925 11555
rect 5925 11525 5955 11555
rect 5955 11525 5956 11555
rect 5924 11524 5956 11525
rect 5924 11475 5956 11476
rect 5924 11445 5925 11475
rect 5925 11445 5955 11475
rect 5955 11445 5956 11475
rect 5924 11444 5956 11445
rect 5924 11395 5956 11396
rect 5924 11365 5925 11395
rect 5925 11365 5955 11395
rect 5955 11365 5956 11395
rect 5924 11364 5956 11365
rect 5924 11315 5956 11316
rect 5924 11285 5925 11315
rect 5925 11285 5955 11315
rect 5955 11285 5956 11315
rect 5924 11284 5956 11285
rect 5924 11235 5956 11236
rect 5924 11205 5925 11235
rect 5925 11205 5955 11235
rect 5955 11205 5956 11235
rect 5924 11204 5956 11205
rect 5924 11155 5956 11156
rect 5924 11125 5925 11155
rect 5925 11125 5955 11155
rect 5955 11125 5956 11155
rect 5924 11124 5956 11125
rect 5924 11075 5956 11076
rect 5924 11045 5925 11075
rect 5925 11045 5955 11075
rect 5955 11045 5956 11075
rect 5924 11044 5956 11045
rect 5924 10964 5956 10996
rect 5924 10915 5956 10916
rect 5924 10885 5925 10915
rect 5925 10885 5955 10915
rect 5955 10885 5956 10915
rect 5924 10884 5956 10885
rect 5924 10835 5956 10836
rect 5924 10805 5925 10835
rect 5925 10805 5955 10835
rect 5955 10805 5956 10835
rect 5924 10804 5956 10805
rect 5924 10755 5956 10756
rect 5924 10725 5925 10755
rect 5925 10725 5955 10755
rect 5955 10725 5956 10755
rect 5924 10724 5956 10725
rect 5924 10675 5956 10676
rect 5924 10645 5925 10675
rect 5925 10645 5955 10675
rect 5955 10645 5956 10675
rect 5924 10644 5956 10645
rect 5924 10595 5956 10596
rect 5924 10565 5925 10595
rect 5925 10565 5955 10595
rect 5955 10565 5956 10595
rect 5924 10564 5956 10565
rect 5924 10515 5956 10516
rect 5924 10485 5925 10515
rect 5925 10485 5955 10515
rect 5955 10485 5956 10515
rect 5924 10484 5956 10485
rect 5924 10435 5956 10436
rect 5924 10405 5925 10435
rect 5925 10405 5955 10435
rect 5955 10405 5956 10435
rect 5924 10404 5956 10405
rect 5924 10355 5956 10356
rect 5924 10325 5925 10355
rect 5925 10325 5955 10355
rect 5955 10325 5956 10355
rect 5924 10324 5956 10325
rect 5924 10244 5956 10276
rect 5924 10164 5956 10196
rect 5924 10084 5956 10116
rect 5924 10004 5956 10036
rect 5924 9955 5956 9956
rect 5924 9925 5925 9955
rect 5925 9925 5955 9955
rect 5955 9925 5956 9955
rect 5924 9924 5956 9925
rect 5924 9875 5956 9876
rect 5924 9845 5925 9875
rect 5925 9845 5955 9875
rect 5955 9845 5956 9875
rect 5924 9844 5956 9845
rect 5924 9795 5956 9796
rect 5924 9765 5925 9795
rect 5925 9765 5955 9795
rect 5955 9765 5956 9795
rect 5924 9764 5956 9765
rect 5924 9715 5956 9716
rect 5924 9685 5925 9715
rect 5925 9685 5955 9715
rect 5955 9685 5956 9715
rect 5924 9684 5956 9685
rect 5924 9635 5956 9636
rect 5924 9605 5925 9635
rect 5925 9605 5955 9635
rect 5955 9605 5956 9635
rect 5924 9604 5956 9605
rect 5924 9555 5956 9556
rect 5924 9525 5925 9555
rect 5925 9525 5955 9555
rect 5955 9525 5956 9555
rect 5924 9524 5956 9525
rect 5924 9475 5956 9476
rect 5924 9445 5925 9475
rect 5925 9445 5955 9475
rect 5955 9445 5956 9475
rect 5924 9444 5956 9445
rect 5924 9395 5956 9396
rect 5924 9365 5925 9395
rect 5925 9365 5955 9395
rect 5955 9365 5956 9395
rect 5924 9364 5956 9365
rect 5924 9284 5956 9316
rect 5924 9204 5956 9236
rect 5924 9124 5956 9156
rect 5924 9044 5956 9076
rect 5924 8995 5956 8996
rect 5924 8965 5925 8995
rect 5925 8965 5955 8995
rect 5955 8965 5956 8995
rect 5924 8964 5956 8965
rect 5924 8915 5956 8916
rect 5924 8885 5925 8915
rect 5925 8885 5955 8915
rect 5955 8885 5956 8915
rect 5924 8884 5956 8885
rect 5924 8835 5956 8836
rect 5924 8805 5925 8835
rect 5925 8805 5955 8835
rect 5955 8805 5956 8835
rect 5924 8804 5956 8805
rect 5924 8755 5956 8756
rect 5924 8725 5925 8755
rect 5925 8725 5955 8755
rect 5955 8725 5956 8755
rect 5924 8724 5956 8725
rect 5924 8675 5956 8676
rect 5924 8645 5925 8675
rect 5925 8645 5955 8675
rect 5955 8645 5956 8675
rect 5924 8644 5956 8645
rect 5924 8595 5956 8596
rect 5924 8565 5925 8595
rect 5925 8565 5955 8595
rect 5955 8565 5956 8595
rect 5924 8564 5956 8565
rect 5924 8515 5956 8516
rect 5924 8485 5925 8515
rect 5925 8485 5955 8515
rect 5955 8485 5956 8515
rect 5924 8484 5956 8485
rect 5924 8435 5956 8436
rect 5924 8405 5925 8435
rect 5925 8405 5955 8435
rect 5955 8405 5956 8435
rect 5924 8404 5956 8405
rect 5924 8324 5956 8356
rect 5924 8275 5956 8276
rect 5924 8245 5925 8275
rect 5925 8245 5955 8275
rect 5955 8245 5956 8275
rect 5924 8244 5956 8245
rect 5924 8195 5956 8196
rect 5924 8165 5925 8195
rect 5925 8165 5955 8195
rect 5955 8165 5956 8195
rect 5924 8164 5956 8165
rect 5924 8115 5956 8116
rect 5924 8085 5925 8115
rect 5925 8085 5955 8115
rect 5955 8085 5956 8115
rect 5924 8084 5956 8085
rect 5924 8035 5956 8036
rect 5924 8005 5925 8035
rect 5925 8005 5955 8035
rect 5955 8005 5956 8035
rect 5924 8004 5956 8005
rect 5924 7955 5956 7956
rect 5924 7925 5925 7955
rect 5925 7925 5955 7955
rect 5955 7925 5956 7955
rect 5924 7924 5956 7925
rect 5924 7875 5956 7876
rect 5924 7845 5925 7875
rect 5925 7845 5955 7875
rect 5955 7845 5956 7875
rect 5924 7844 5956 7845
rect 5924 7795 5956 7796
rect 5924 7765 5925 7795
rect 5925 7765 5955 7795
rect 5955 7765 5956 7795
rect 5924 7764 5956 7765
rect 5924 7715 5956 7716
rect 5924 7685 5925 7715
rect 5925 7685 5955 7715
rect 5955 7685 5956 7715
rect 5924 7684 5956 7685
rect 5924 7635 5956 7636
rect 5924 7605 5925 7635
rect 5925 7605 5955 7635
rect 5955 7605 5956 7635
rect 5924 7604 5956 7605
rect 5924 7555 5956 7556
rect 5924 7525 5925 7555
rect 5925 7525 5955 7555
rect 5955 7525 5956 7555
rect 5924 7524 5956 7525
rect 5924 7475 5956 7476
rect 5924 7445 5925 7475
rect 5925 7445 5955 7475
rect 5955 7445 5956 7475
rect 5924 7444 5956 7445
rect 5924 7395 5956 7396
rect 5924 7365 5925 7395
rect 5925 7365 5955 7395
rect 5955 7365 5956 7395
rect 5924 7364 5956 7365
rect 5924 7315 5956 7316
rect 5924 7285 5925 7315
rect 5925 7285 5955 7315
rect 5955 7285 5956 7315
rect 5924 7284 5956 7285
rect 5924 7235 5956 7236
rect 5924 7205 5925 7235
rect 5925 7205 5955 7235
rect 5955 7205 5956 7235
rect 5924 7204 5956 7205
rect 5924 7155 5956 7156
rect 5924 7125 5925 7155
rect 5925 7125 5955 7155
rect 5955 7125 5956 7155
rect 5924 7124 5956 7125
rect 5924 7075 5956 7076
rect 5924 7045 5925 7075
rect 5925 7045 5955 7075
rect 5955 7045 5956 7075
rect 5924 7044 5956 7045
rect 5924 6995 5956 6996
rect 5924 6965 5925 6995
rect 5925 6965 5955 6995
rect 5955 6965 5956 6995
rect 5924 6964 5956 6965
rect 5924 6884 5956 6916
rect 5924 6835 5956 6836
rect 5924 6805 5925 6835
rect 5925 6805 5955 6835
rect 5955 6805 5956 6835
rect 5924 6804 5956 6805
rect 5924 6755 5956 6756
rect 5924 6725 5925 6755
rect 5925 6725 5955 6755
rect 5955 6725 5956 6755
rect 5924 6724 5956 6725
rect 5924 6675 5956 6676
rect 5924 6645 5925 6675
rect 5925 6645 5955 6675
rect 5955 6645 5956 6675
rect 5924 6644 5956 6645
rect 5924 6595 5956 6596
rect 5924 6565 5925 6595
rect 5925 6565 5955 6595
rect 5955 6565 5956 6595
rect 5924 6564 5956 6565
rect 5924 6515 5956 6516
rect 5924 6485 5925 6515
rect 5925 6485 5955 6515
rect 5955 6485 5956 6515
rect 5924 6484 5956 6485
rect 5924 6435 5956 6436
rect 5924 6405 5925 6435
rect 5925 6405 5955 6435
rect 5955 6405 5956 6435
rect 5924 6404 5956 6405
rect 5924 6355 5956 6356
rect 5924 6325 5925 6355
rect 5925 6325 5955 6355
rect 5955 6325 5956 6355
rect 5924 6324 5956 6325
rect 5924 6275 5956 6276
rect 5924 6245 5925 6275
rect 5925 6245 5955 6275
rect 5955 6245 5956 6275
rect 5924 6244 5956 6245
rect 5924 6164 5956 6196
rect 5924 6084 5956 6116
rect 5924 6004 5956 6036
rect 5924 5924 5956 5956
rect 5924 5875 5956 5876
rect 5924 5845 5925 5875
rect 5925 5845 5955 5875
rect 5955 5845 5956 5875
rect 5924 5844 5956 5845
rect 5924 5795 5956 5796
rect 5924 5765 5925 5795
rect 5925 5765 5955 5795
rect 5955 5765 5956 5795
rect 5924 5764 5956 5765
rect 5924 5715 5956 5716
rect 5924 5685 5925 5715
rect 5925 5685 5955 5715
rect 5955 5685 5956 5715
rect 5924 5684 5956 5685
rect 5924 5635 5956 5636
rect 5924 5605 5925 5635
rect 5925 5605 5955 5635
rect 5955 5605 5956 5635
rect 5924 5604 5956 5605
rect 5924 5555 5956 5556
rect 5924 5525 5925 5555
rect 5925 5525 5955 5555
rect 5955 5525 5956 5555
rect 5924 5524 5956 5525
rect 5924 5475 5956 5476
rect 5924 5445 5925 5475
rect 5925 5445 5955 5475
rect 5955 5445 5956 5475
rect 5924 5444 5956 5445
rect 5924 5395 5956 5396
rect 5924 5365 5925 5395
rect 5925 5365 5955 5395
rect 5955 5365 5956 5395
rect 5924 5364 5956 5365
rect 5924 5315 5956 5316
rect 5924 5285 5925 5315
rect 5925 5285 5955 5315
rect 5955 5285 5956 5315
rect 5924 5284 5956 5285
rect 5924 5235 5956 5236
rect 5924 5205 5925 5235
rect 5925 5205 5955 5235
rect 5955 5205 5956 5235
rect 5924 5204 5956 5205
rect 5924 5155 5956 5156
rect 5924 5125 5925 5155
rect 5925 5125 5955 5155
rect 5955 5125 5956 5155
rect 5924 5124 5956 5125
rect 5924 5075 5956 5076
rect 5924 5045 5925 5075
rect 5925 5045 5955 5075
rect 5955 5045 5956 5075
rect 5924 5044 5956 5045
rect 5924 4995 5956 4996
rect 5924 4965 5925 4995
rect 5925 4965 5955 4995
rect 5955 4965 5956 4995
rect 5924 4964 5956 4965
rect 5924 4915 5956 4916
rect 5924 4885 5925 4915
rect 5925 4885 5955 4915
rect 5955 4885 5956 4915
rect 5924 4884 5956 4885
rect 5924 4804 5956 4836
rect 5924 4755 5956 4756
rect 5924 4725 5925 4755
rect 5925 4725 5955 4755
rect 5955 4725 5956 4755
rect 5924 4724 5956 4725
rect 5924 4675 5956 4676
rect 5924 4645 5925 4675
rect 5925 4645 5955 4675
rect 5955 4645 5956 4675
rect 5924 4644 5956 4645
rect 5924 4564 5956 4596
rect 5924 4515 5956 4516
rect 5924 4485 5925 4515
rect 5925 4485 5955 4515
rect 5955 4485 5956 4515
rect 5924 4484 5956 4485
rect 5924 4435 5956 4436
rect 5924 4405 5925 4435
rect 5925 4405 5955 4435
rect 5955 4405 5956 4435
rect 5924 4404 5956 4405
rect 5924 4355 5956 4356
rect 5924 4325 5925 4355
rect 5925 4325 5955 4355
rect 5955 4325 5956 4355
rect 5924 4324 5956 4325
rect 5924 4275 5956 4276
rect 5924 4245 5925 4275
rect 5925 4245 5955 4275
rect 5955 4245 5956 4275
rect 5924 4244 5956 4245
rect 5924 4195 5956 4196
rect 5924 4165 5925 4195
rect 5925 4165 5955 4195
rect 5955 4165 5956 4195
rect 5924 4164 5956 4165
rect 5924 4115 5956 4116
rect 5924 4085 5925 4115
rect 5925 4085 5955 4115
rect 5955 4085 5956 4115
rect 5924 4084 5956 4085
rect 5924 4035 5956 4036
rect 5924 4005 5925 4035
rect 5925 4005 5955 4035
rect 5955 4005 5956 4035
rect 5924 4004 5956 4005
rect 5924 3955 5956 3956
rect 5924 3925 5925 3955
rect 5925 3925 5955 3955
rect 5955 3925 5956 3955
rect 5924 3924 5956 3925
rect 5924 3875 5956 3876
rect 5924 3845 5925 3875
rect 5925 3845 5955 3875
rect 5955 3845 5956 3875
rect 5924 3844 5956 3845
rect 5924 3764 5956 3796
rect 5924 3715 5956 3716
rect 5924 3685 5925 3715
rect 5925 3685 5955 3715
rect 5955 3685 5956 3715
rect 5924 3684 5956 3685
rect 5924 3635 5956 3636
rect 5924 3605 5925 3635
rect 5925 3605 5955 3635
rect 5955 3605 5956 3635
rect 5924 3604 5956 3605
rect 5924 3524 5956 3556
rect 5924 3475 5956 3476
rect 5924 3445 5925 3475
rect 5925 3445 5955 3475
rect 5955 3445 5956 3475
rect 5924 3444 5956 3445
rect 5924 3395 5956 3396
rect 5924 3365 5925 3395
rect 5925 3365 5955 3395
rect 5955 3365 5956 3395
rect 5924 3364 5956 3365
rect 5924 3284 5956 3316
rect 5924 3235 5956 3236
rect 5924 3205 5925 3235
rect 5925 3205 5955 3235
rect 5955 3205 5956 3235
rect 5924 3204 5956 3205
rect 5924 3155 5956 3156
rect 5924 3125 5925 3155
rect 5925 3125 5955 3155
rect 5955 3125 5956 3155
rect 5924 3124 5956 3125
rect 5924 3075 5956 3076
rect 5924 3045 5925 3075
rect 5925 3045 5955 3075
rect 5955 3045 5956 3075
rect 5924 3044 5956 3045
rect 5924 2995 5956 2996
rect 5924 2965 5925 2995
rect 5925 2965 5955 2995
rect 5955 2965 5956 2995
rect 5924 2964 5956 2965
rect 5924 2915 5956 2916
rect 5924 2885 5925 2915
rect 5925 2885 5955 2915
rect 5955 2885 5956 2915
rect 5924 2884 5956 2885
rect 5924 2835 5956 2836
rect 5924 2805 5925 2835
rect 5925 2805 5955 2835
rect 5955 2805 5956 2835
rect 5924 2804 5956 2805
rect 5924 2755 5956 2756
rect 5924 2725 5925 2755
rect 5925 2725 5955 2755
rect 5955 2725 5956 2755
rect 5924 2724 5956 2725
rect 5924 2675 5956 2676
rect 5924 2645 5925 2675
rect 5925 2645 5955 2675
rect 5955 2645 5956 2675
rect 5924 2644 5956 2645
rect 5924 2595 5956 2596
rect 5924 2565 5925 2595
rect 5925 2565 5955 2595
rect 5955 2565 5956 2595
rect 5924 2564 5956 2565
rect 5924 2515 5956 2516
rect 5924 2485 5925 2515
rect 5925 2485 5955 2515
rect 5955 2485 5956 2515
rect 5924 2484 5956 2485
rect 5924 2435 5956 2436
rect 5924 2405 5925 2435
rect 5925 2405 5955 2435
rect 5955 2405 5956 2435
rect 5924 2404 5956 2405
rect 5924 2355 5956 2356
rect 5924 2325 5925 2355
rect 5925 2325 5955 2355
rect 5955 2325 5956 2355
rect 5924 2324 5956 2325
rect 5924 2275 5956 2276
rect 5924 2245 5925 2275
rect 5925 2245 5955 2275
rect 5955 2245 5956 2275
rect 5924 2244 5956 2245
rect 5924 2195 5956 2196
rect 5924 2165 5925 2195
rect 5925 2165 5955 2195
rect 5955 2165 5956 2195
rect 5924 2164 5956 2165
rect 5924 2115 5956 2116
rect 5924 2085 5925 2115
rect 5925 2085 5955 2115
rect 5955 2085 5956 2115
rect 5924 2084 5956 2085
rect 5924 2035 5956 2036
rect 5924 2005 5925 2035
rect 5925 2005 5955 2035
rect 5955 2005 5956 2035
rect 5924 2004 5956 2005
rect 5924 1955 5956 1956
rect 5924 1925 5925 1955
rect 5925 1925 5955 1955
rect 5955 1925 5956 1955
rect 5924 1924 5956 1925
rect 5924 1844 5956 1876
rect 5924 1764 5956 1796
rect 5924 1715 5956 1716
rect 5924 1685 5925 1715
rect 5925 1685 5955 1715
rect 5955 1685 5956 1715
rect 5924 1684 5956 1685
rect 5924 1635 5956 1636
rect 5924 1605 5925 1635
rect 5925 1605 5955 1635
rect 5955 1605 5956 1635
rect 5924 1604 5956 1605
rect 5924 1555 5956 1556
rect 5924 1525 5925 1555
rect 5925 1525 5955 1555
rect 5955 1525 5956 1555
rect 5924 1524 5956 1525
rect 5924 1475 5956 1476
rect 5924 1445 5925 1475
rect 5925 1445 5955 1475
rect 5955 1445 5956 1475
rect 5924 1444 5956 1445
rect 5924 1395 5956 1396
rect 5924 1365 5925 1395
rect 5925 1365 5955 1395
rect 5955 1365 5956 1395
rect 5924 1364 5956 1365
rect 5924 1315 5956 1316
rect 5924 1285 5925 1315
rect 5925 1285 5955 1315
rect 5955 1285 5956 1315
rect 5924 1284 5956 1285
rect 5924 1235 5956 1236
rect 5924 1205 5925 1235
rect 5925 1205 5955 1235
rect 5955 1205 5956 1235
rect 5924 1204 5956 1205
rect 5924 1155 5956 1156
rect 5924 1125 5925 1155
rect 5925 1125 5955 1155
rect 5955 1125 5956 1155
rect 5924 1124 5956 1125
rect 5924 1075 5956 1076
rect 5924 1045 5925 1075
rect 5925 1045 5955 1075
rect 5955 1045 5956 1075
rect 5924 1044 5956 1045
rect 5924 995 5956 996
rect 5924 965 5925 995
rect 5925 965 5955 995
rect 5955 965 5956 995
rect 5924 964 5956 965
rect 5924 884 5956 916
rect 5924 835 5956 836
rect 5924 805 5925 835
rect 5925 805 5955 835
rect 5955 805 5956 835
rect 5924 804 5956 805
rect 5924 755 5956 756
rect 5924 725 5925 755
rect 5925 725 5955 755
rect 5955 725 5956 755
rect 5924 724 5956 725
rect 5924 675 5956 676
rect 5924 645 5925 675
rect 5925 645 5955 675
rect 5955 645 5956 675
rect 5924 644 5956 645
rect 5924 595 5956 596
rect 5924 565 5925 595
rect 5925 565 5955 595
rect 5955 565 5956 595
rect 5924 564 5956 565
rect 5924 515 5956 516
rect 5924 485 5925 515
rect 5925 485 5955 515
rect 5955 485 5956 515
rect 5924 484 5956 485
rect 5924 404 5956 436
rect 5924 324 5956 356
rect 5924 275 5956 276
rect 5924 245 5925 275
rect 5925 245 5955 275
rect 5955 245 5956 275
rect 5924 244 5956 245
rect 5924 195 5956 196
rect 5924 165 5925 195
rect 5925 165 5955 195
rect 5955 165 5956 195
rect 5924 164 5956 165
rect 5924 115 5956 116
rect 5924 85 5925 115
rect 5925 85 5955 115
rect 5955 85 5956 115
rect 5924 84 5956 85
rect 5924 35 5956 36
rect 5924 5 5925 35
rect 5925 5 5955 35
rect 5955 5 5956 35
rect 5924 4 5956 5
rect 5764 -236 5796 -44
rect 5924 -236 5956 -44
rect 6004 15715 6036 15716
rect 6004 15685 6005 15715
rect 6005 15685 6035 15715
rect 6035 15685 6036 15715
rect 6004 15684 6036 15685
rect 6004 15635 6036 15636
rect 6004 15605 6005 15635
rect 6005 15605 6035 15635
rect 6035 15605 6036 15635
rect 6004 15604 6036 15605
rect 6004 15555 6036 15556
rect 6004 15525 6005 15555
rect 6005 15525 6035 15555
rect 6035 15525 6036 15555
rect 6004 15524 6036 15525
rect 6004 15475 6036 15476
rect 6004 15445 6005 15475
rect 6005 15445 6035 15475
rect 6035 15445 6036 15475
rect 6004 15444 6036 15445
rect 6004 15395 6036 15396
rect 6004 15365 6005 15395
rect 6005 15365 6035 15395
rect 6035 15365 6036 15395
rect 6004 15364 6036 15365
rect 6004 15315 6036 15316
rect 6004 15285 6005 15315
rect 6005 15285 6035 15315
rect 6035 15285 6036 15315
rect 6004 15284 6036 15285
rect 6004 15235 6036 15236
rect 6004 15205 6005 15235
rect 6005 15205 6035 15235
rect 6035 15205 6036 15235
rect 6004 15204 6036 15205
rect 6004 15155 6036 15156
rect 6004 15125 6005 15155
rect 6005 15125 6035 15155
rect 6035 15125 6036 15155
rect 6004 15124 6036 15125
rect 6004 15044 6036 15076
rect 6004 14995 6036 14996
rect 6004 14965 6005 14995
rect 6005 14965 6035 14995
rect 6035 14965 6036 14995
rect 6004 14964 6036 14965
rect 6004 14915 6036 14916
rect 6004 14885 6005 14915
rect 6005 14885 6035 14915
rect 6035 14885 6036 14915
rect 6004 14884 6036 14885
rect 6004 14835 6036 14836
rect 6004 14805 6005 14835
rect 6005 14805 6035 14835
rect 6035 14805 6036 14835
rect 6004 14804 6036 14805
rect 6004 14755 6036 14756
rect 6004 14725 6005 14755
rect 6005 14725 6035 14755
rect 6035 14725 6036 14755
rect 6004 14724 6036 14725
rect 6004 14675 6036 14676
rect 6004 14645 6005 14675
rect 6005 14645 6035 14675
rect 6035 14645 6036 14675
rect 6004 14644 6036 14645
rect 6004 14595 6036 14596
rect 6004 14565 6005 14595
rect 6005 14565 6035 14595
rect 6035 14565 6036 14595
rect 6004 14564 6036 14565
rect 6004 14515 6036 14516
rect 6004 14485 6005 14515
rect 6005 14485 6035 14515
rect 6035 14485 6036 14515
rect 6004 14484 6036 14485
rect 6004 14435 6036 14436
rect 6004 14405 6005 14435
rect 6005 14405 6035 14435
rect 6035 14405 6036 14435
rect 6004 14404 6036 14405
rect 6004 14324 6036 14356
rect 6004 14244 6036 14276
rect 6004 14164 6036 14196
rect 6004 14084 6036 14116
rect 6004 14035 6036 14036
rect 6004 14005 6005 14035
rect 6005 14005 6035 14035
rect 6035 14005 6036 14035
rect 6004 14004 6036 14005
rect 6004 13955 6036 13956
rect 6004 13925 6005 13955
rect 6005 13925 6035 13955
rect 6035 13925 6036 13955
rect 6004 13924 6036 13925
rect 6004 13875 6036 13876
rect 6004 13845 6005 13875
rect 6005 13845 6035 13875
rect 6035 13845 6036 13875
rect 6004 13844 6036 13845
rect 6004 13795 6036 13796
rect 6004 13765 6005 13795
rect 6005 13765 6035 13795
rect 6035 13765 6036 13795
rect 6004 13764 6036 13765
rect 6004 13715 6036 13716
rect 6004 13685 6005 13715
rect 6005 13685 6035 13715
rect 6035 13685 6036 13715
rect 6004 13684 6036 13685
rect 6004 13635 6036 13636
rect 6004 13605 6005 13635
rect 6005 13605 6035 13635
rect 6035 13605 6036 13635
rect 6004 13604 6036 13605
rect 6004 13555 6036 13556
rect 6004 13525 6005 13555
rect 6005 13525 6035 13555
rect 6035 13525 6036 13555
rect 6004 13524 6036 13525
rect 6004 13475 6036 13476
rect 6004 13445 6005 13475
rect 6005 13445 6035 13475
rect 6035 13445 6036 13475
rect 6004 13444 6036 13445
rect 6004 13364 6036 13396
rect 6004 13284 6036 13316
rect 6004 13204 6036 13236
rect 6004 13124 6036 13156
rect 6004 13075 6036 13076
rect 6004 13045 6005 13075
rect 6005 13045 6035 13075
rect 6035 13045 6036 13075
rect 6004 13044 6036 13045
rect 6004 12995 6036 12996
rect 6004 12965 6005 12995
rect 6005 12965 6035 12995
rect 6035 12965 6036 12995
rect 6004 12964 6036 12965
rect 6004 12915 6036 12916
rect 6004 12885 6005 12915
rect 6005 12885 6035 12915
rect 6035 12885 6036 12915
rect 6004 12884 6036 12885
rect 6004 12835 6036 12836
rect 6004 12805 6005 12835
rect 6005 12805 6035 12835
rect 6035 12805 6036 12835
rect 6004 12804 6036 12805
rect 6004 12755 6036 12756
rect 6004 12725 6005 12755
rect 6005 12725 6035 12755
rect 6035 12725 6036 12755
rect 6004 12724 6036 12725
rect 6004 12675 6036 12676
rect 6004 12645 6005 12675
rect 6005 12645 6035 12675
rect 6035 12645 6036 12675
rect 6004 12644 6036 12645
rect 6004 12595 6036 12596
rect 6004 12565 6005 12595
rect 6005 12565 6035 12595
rect 6035 12565 6036 12595
rect 6004 12564 6036 12565
rect 6004 12515 6036 12516
rect 6004 12485 6005 12515
rect 6005 12485 6035 12515
rect 6035 12485 6036 12515
rect 6004 12484 6036 12485
rect 6004 12404 6036 12436
rect 6004 12355 6036 12356
rect 6004 12325 6005 12355
rect 6005 12325 6035 12355
rect 6035 12325 6036 12355
rect 6004 12324 6036 12325
rect 6004 12275 6036 12276
rect 6004 12245 6005 12275
rect 6005 12245 6035 12275
rect 6035 12245 6036 12275
rect 6004 12244 6036 12245
rect 6004 12195 6036 12196
rect 6004 12165 6005 12195
rect 6005 12165 6035 12195
rect 6035 12165 6036 12195
rect 6004 12164 6036 12165
rect 6004 12115 6036 12116
rect 6004 12085 6005 12115
rect 6005 12085 6035 12115
rect 6035 12085 6036 12115
rect 6004 12084 6036 12085
rect 6004 12035 6036 12036
rect 6004 12005 6005 12035
rect 6005 12005 6035 12035
rect 6035 12005 6036 12035
rect 6004 12004 6036 12005
rect 6004 11955 6036 11956
rect 6004 11925 6005 11955
rect 6005 11925 6035 11955
rect 6035 11925 6036 11955
rect 6004 11924 6036 11925
rect 6004 11875 6036 11876
rect 6004 11845 6005 11875
rect 6005 11845 6035 11875
rect 6035 11845 6036 11875
rect 6004 11844 6036 11845
rect 6004 11795 6036 11796
rect 6004 11765 6005 11795
rect 6005 11765 6035 11795
rect 6035 11765 6036 11795
rect 6004 11764 6036 11765
rect 6004 11715 6036 11716
rect 6004 11685 6005 11715
rect 6005 11685 6035 11715
rect 6035 11685 6036 11715
rect 6004 11684 6036 11685
rect 6004 11635 6036 11636
rect 6004 11605 6005 11635
rect 6005 11605 6035 11635
rect 6035 11605 6036 11635
rect 6004 11604 6036 11605
rect 6004 11555 6036 11556
rect 6004 11525 6005 11555
rect 6005 11525 6035 11555
rect 6035 11525 6036 11555
rect 6004 11524 6036 11525
rect 6004 11475 6036 11476
rect 6004 11445 6005 11475
rect 6005 11445 6035 11475
rect 6035 11445 6036 11475
rect 6004 11444 6036 11445
rect 6004 11395 6036 11396
rect 6004 11365 6005 11395
rect 6005 11365 6035 11395
rect 6035 11365 6036 11395
rect 6004 11364 6036 11365
rect 6004 11315 6036 11316
rect 6004 11285 6005 11315
rect 6005 11285 6035 11315
rect 6035 11285 6036 11315
rect 6004 11284 6036 11285
rect 6004 11235 6036 11236
rect 6004 11205 6005 11235
rect 6005 11205 6035 11235
rect 6035 11205 6036 11235
rect 6004 11204 6036 11205
rect 6004 11155 6036 11156
rect 6004 11125 6005 11155
rect 6005 11125 6035 11155
rect 6035 11125 6036 11155
rect 6004 11124 6036 11125
rect 6004 11075 6036 11076
rect 6004 11045 6005 11075
rect 6005 11045 6035 11075
rect 6035 11045 6036 11075
rect 6004 11044 6036 11045
rect 6004 10964 6036 10996
rect 6004 10915 6036 10916
rect 6004 10885 6005 10915
rect 6005 10885 6035 10915
rect 6035 10885 6036 10915
rect 6004 10884 6036 10885
rect 6004 10835 6036 10836
rect 6004 10805 6005 10835
rect 6005 10805 6035 10835
rect 6035 10805 6036 10835
rect 6004 10804 6036 10805
rect 6004 10755 6036 10756
rect 6004 10725 6005 10755
rect 6005 10725 6035 10755
rect 6035 10725 6036 10755
rect 6004 10724 6036 10725
rect 6004 10675 6036 10676
rect 6004 10645 6005 10675
rect 6005 10645 6035 10675
rect 6035 10645 6036 10675
rect 6004 10644 6036 10645
rect 6004 10595 6036 10596
rect 6004 10565 6005 10595
rect 6005 10565 6035 10595
rect 6035 10565 6036 10595
rect 6004 10564 6036 10565
rect 6004 10515 6036 10516
rect 6004 10485 6005 10515
rect 6005 10485 6035 10515
rect 6035 10485 6036 10515
rect 6004 10484 6036 10485
rect 6004 10435 6036 10436
rect 6004 10405 6005 10435
rect 6005 10405 6035 10435
rect 6035 10405 6036 10435
rect 6004 10404 6036 10405
rect 6004 10355 6036 10356
rect 6004 10325 6005 10355
rect 6005 10325 6035 10355
rect 6035 10325 6036 10355
rect 6004 10324 6036 10325
rect 6004 10244 6036 10276
rect 6004 10164 6036 10196
rect 6004 10084 6036 10116
rect 6004 10004 6036 10036
rect 6004 9955 6036 9956
rect 6004 9925 6005 9955
rect 6005 9925 6035 9955
rect 6035 9925 6036 9955
rect 6004 9924 6036 9925
rect 6004 9875 6036 9876
rect 6004 9845 6005 9875
rect 6005 9845 6035 9875
rect 6035 9845 6036 9875
rect 6004 9844 6036 9845
rect 6004 9795 6036 9796
rect 6004 9765 6005 9795
rect 6005 9765 6035 9795
rect 6035 9765 6036 9795
rect 6004 9764 6036 9765
rect 6004 9715 6036 9716
rect 6004 9685 6005 9715
rect 6005 9685 6035 9715
rect 6035 9685 6036 9715
rect 6004 9684 6036 9685
rect 6004 9635 6036 9636
rect 6004 9605 6005 9635
rect 6005 9605 6035 9635
rect 6035 9605 6036 9635
rect 6004 9604 6036 9605
rect 6004 9555 6036 9556
rect 6004 9525 6005 9555
rect 6005 9525 6035 9555
rect 6035 9525 6036 9555
rect 6004 9524 6036 9525
rect 6004 9475 6036 9476
rect 6004 9445 6005 9475
rect 6005 9445 6035 9475
rect 6035 9445 6036 9475
rect 6004 9444 6036 9445
rect 6004 9395 6036 9396
rect 6004 9365 6005 9395
rect 6005 9365 6035 9395
rect 6035 9365 6036 9395
rect 6004 9364 6036 9365
rect 6004 9284 6036 9316
rect 6004 9204 6036 9236
rect 6004 9124 6036 9156
rect 6004 9044 6036 9076
rect 6004 8995 6036 8996
rect 6004 8965 6005 8995
rect 6005 8965 6035 8995
rect 6035 8965 6036 8995
rect 6004 8964 6036 8965
rect 6004 8915 6036 8916
rect 6004 8885 6005 8915
rect 6005 8885 6035 8915
rect 6035 8885 6036 8915
rect 6004 8884 6036 8885
rect 6004 8835 6036 8836
rect 6004 8805 6005 8835
rect 6005 8805 6035 8835
rect 6035 8805 6036 8835
rect 6004 8804 6036 8805
rect 6004 8755 6036 8756
rect 6004 8725 6005 8755
rect 6005 8725 6035 8755
rect 6035 8725 6036 8755
rect 6004 8724 6036 8725
rect 6004 8675 6036 8676
rect 6004 8645 6005 8675
rect 6005 8645 6035 8675
rect 6035 8645 6036 8675
rect 6004 8644 6036 8645
rect 6004 8595 6036 8596
rect 6004 8565 6005 8595
rect 6005 8565 6035 8595
rect 6035 8565 6036 8595
rect 6004 8564 6036 8565
rect 6004 8515 6036 8516
rect 6004 8485 6005 8515
rect 6005 8485 6035 8515
rect 6035 8485 6036 8515
rect 6004 8484 6036 8485
rect 6004 8435 6036 8436
rect 6004 8405 6005 8435
rect 6005 8405 6035 8435
rect 6035 8405 6036 8435
rect 6004 8404 6036 8405
rect 6004 8324 6036 8356
rect 6004 8275 6036 8276
rect 6004 8245 6005 8275
rect 6005 8245 6035 8275
rect 6035 8245 6036 8275
rect 6004 8244 6036 8245
rect 6004 8195 6036 8196
rect 6004 8165 6005 8195
rect 6005 8165 6035 8195
rect 6035 8165 6036 8195
rect 6004 8164 6036 8165
rect 6004 8115 6036 8116
rect 6004 8085 6005 8115
rect 6005 8085 6035 8115
rect 6035 8085 6036 8115
rect 6004 8084 6036 8085
rect 6004 8035 6036 8036
rect 6004 8005 6005 8035
rect 6005 8005 6035 8035
rect 6035 8005 6036 8035
rect 6004 8004 6036 8005
rect 6004 7955 6036 7956
rect 6004 7925 6005 7955
rect 6005 7925 6035 7955
rect 6035 7925 6036 7955
rect 6004 7924 6036 7925
rect 6004 7875 6036 7876
rect 6004 7845 6005 7875
rect 6005 7845 6035 7875
rect 6035 7845 6036 7875
rect 6004 7844 6036 7845
rect 6004 7795 6036 7796
rect 6004 7765 6005 7795
rect 6005 7765 6035 7795
rect 6035 7765 6036 7795
rect 6004 7764 6036 7765
rect 6004 7715 6036 7716
rect 6004 7685 6005 7715
rect 6005 7685 6035 7715
rect 6035 7685 6036 7715
rect 6004 7684 6036 7685
rect 6004 7635 6036 7636
rect 6004 7605 6005 7635
rect 6005 7605 6035 7635
rect 6035 7605 6036 7635
rect 6004 7604 6036 7605
rect 6004 7555 6036 7556
rect 6004 7525 6005 7555
rect 6005 7525 6035 7555
rect 6035 7525 6036 7555
rect 6004 7524 6036 7525
rect 6004 7475 6036 7476
rect 6004 7445 6005 7475
rect 6005 7445 6035 7475
rect 6035 7445 6036 7475
rect 6004 7444 6036 7445
rect 6004 7395 6036 7396
rect 6004 7365 6005 7395
rect 6005 7365 6035 7395
rect 6035 7365 6036 7395
rect 6004 7364 6036 7365
rect 6004 7315 6036 7316
rect 6004 7285 6005 7315
rect 6005 7285 6035 7315
rect 6035 7285 6036 7315
rect 6004 7284 6036 7285
rect 6004 7235 6036 7236
rect 6004 7205 6005 7235
rect 6005 7205 6035 7235
rect 6035 7205 6036 7235
rect 6004 7204 6036 7205
rect 6004 7155 6036 7156
rect 6004 7125 6005 7155
rect 6005 7125 6035 7155
rect 6035 7125 6036 7155
rect 6004 7124 6036 7125
rect 6004 7075 6036 7076
rect 6004 7045 6005 7075
rect 6005 7045 6035 7075
rect 6035 7045 6036 7075
rect 6004 7044 6036 7045
rect 6004 6995 6036 6996
rect 6004 6965 6005 6995
rect 6005 6965 6035 6995
rect 6035 6965 6036 6995
rect 6004 6964 6036 6965
rect 6004 6884 6036 6916
rect 6004 6835 6036 6836
rect 6004 6805 6005 6835
rect 6005 6805 6035 6835
rect 6035 6805 6036 6835
rect 6004 6804 6036 6805
rect 6004 6755 6036 6756
rect 6004 6725 6005 6755
rect 6005 6725 6035 6755
rect 6035 6725 6036 6755
rect 6004 6724 6036 6725
rect 6004 6675 6036 6676
rect 6004 6645 6005 6675
rect 6005 6645 6035 6675
rect 6035 6645 6036 6675
rect 6004 6644 6036 6645
rect 6004 6595 6036 6596
rect 6004 6565 6005 6595
rect 6005 6565 6035 6595
rect 6035 6565 6036 6595
rect 6004 6564 6036 6565
rect 6004 6515 6036 6516
rect 6004 6485 6005 6515
rect 6005 6485 6035 6515
rect 6035 6485 6036 6515
rect 6004 6484 6036 6485
rect 6004 6435 6036 6436
rect 6004 6405 6005 6435
rect 6005 6405 6035 6435
rect 6035 6405 6036 6435
rect 6004 6404 6036 6405
rect 6004 6355 6036 6356
rect 6004 6325 6005 6355
rect 6005 6325 6035 6355
rect 6035 6325 6036 6355
rect 6004 6324 6036 6325
rect 6004 6275 6036 6276
rect 6004 6245 6005 6275
rect 6005 6245 6035 6275
rect 6035 6245 6036 6275
rect 6004 6244 6036 6245
rect 6004 6164 6036 6196
rect 6004 6084 6036 6116
rect 6004 6004 6036 6036
rect 6004 5924 6036 5956
rect 6004 5875 6036 5876
rect 6004 5845 6005 5875
rect 6005 5845 6035 5875
rect 6035 5845 6036 5875
rect 6004 5844 6036 5845
rect 6004 5795 6036 5796
rect 6004 5765 6005 5795
rect 6005 5765 6035 5795
rect 6035 5765 6036 5795
rect 6004 5764 6036 5765
rect 6004 5715 6036 5716
rect 6004 5685 6005 5715
rect 6005 5685 6035 5715
rect 6035 5685 6036 5715
rect 6004 5684 6036 5685
rect 6004 5635 6036 5636
rect 6004 5605 6005 5635
rect 6005 5605 6035 5635
rect 6035 5605 6036 5635
rect 6004 5604 6036 5605
rect 6004 5555 6036 5556
rect 6004 5525 6005 5555
rect 6005 5525 6035 5555
rect 6035 5525 6036 5555
rect 6004 5524 6036 5525
rect 6004 5475 6036 5476
rect 6004 5445 6005 5475
rect 6005 5445 6035 5475
rect 6035 5445 6036 5475
rect 6004 5444 6036 5445
rect 6004 5395 6036 5396
rect 6004 5365 6005 5395
rect 6005 5365 6035 5395
rect 6035 5365 6036 5395
rect 6004 5364 6036 5365
rect 6004 5315 6036 5316
rect 6004 5285 6005 5315
rect 6005 5285 6035 5315
rect 6035 5285 6036 5315
rect 6004 5284 6036 5285
rect 6004 5235 6036 5236
rect 6004 5205 6005 5235
rect 6005 5205 6035 5235
rect 6035 5205 6036 5235
rect 6004 5204 6036 5205
rect 6004 5155 6036 5156
rect 6004 5125 6005 5155
rect 6005 5125 6035 5155
rect 6035 5125 6036 5155
rect 6004 5124 6036 5125
rect 6004 5075 6036 5076
rect 6004 5045 6005 5075
rect 6005 5045 6035 5075
rect 6035 5045 6036 5075
rect 6004 5044 6036 5045
rect 6004 4995 6036 4996
rect 6004 4965 6005 4995
rect 6005 4965 6035 4995
rect 6035 4965 6036 4995
rect 6004 4964 6036 4965
rect 6004 4915 6036 4916
rect 6004 4885 6005 4915
rect 6005 4885 6035 4915
rect 6035 4885 6036 4915
rect 6004 4884 6036 4885
rect 6004 4804 6036 4836
rect 6004 4755 6036 4756
rect 6004 4725 6005 4755
rect 6005 4725 6035 4755
rect 6035 4725 6036 4755
rect 6004 4724 6036 4725
rect 6004 4675 6036 4676
rect 6004 4645 6005 4675
rect 6005 4645 6035 4675
rect 6035 4645 6036 4675
rect 6004 4644 6036 4645
rect 6004 4564 6036 4596
rect 6004 4515 6036 4516
rect 6004 4485 6005 4515
rect 6005 4485 6035 4515
rect 6035 4485 6036 4515
rect 6004 4484 6036 4485
rect 6004 4435 6036 4436
rect 6004 4405 6005 4435
rect 6005 4405 6035 4435
rect 6035 4405 6036 4435
rect 6004 4404 6036 4405
rect 6004 4355 6036 4356
rect 6004 4325 6005 4355
rect 6005 4325 6035 4355
rect 6035 4325 6036 4355
rect 6004 4324 6036 4325
rect 6004 4275 6036 4276
rect 6004 4245 6005 4275
rect 6005 4245 6035 4275
rect 6035 4245 6036 4275
rect 6004 4244 6036 4245
rect 6004 4195 6036 4196
rect 6004 4165 6005 4195
rect 6005 4165 6035 4195
rect 6035 4165 6036 4195
rect 6004 4164 6036 4165
rect 6004 4115 6036 4116
rect 6004 4085 6005 4115
rect 6005 4085 6035 4115
rect 6035 4085 6036 4115
rect 6004 4084 6036 4085
rect 6004 4035 6036 4036
rect 6004 4005 6005 4035
rect 6005 4005 6035 4035
rect 6035 4005 6036 4035
rect 6004 4004 6036 4005
rect 6004 3955 6036 3956
rect 6004 3925 6005 3955
rect 6005 3925 6035 3955
rect 6035 3925 6036 3955
rect 6004 3924 6036 3925
rect 6004 3875 6036 3876
rect 6004 3845 6005 3875
rect 6005 3845 6035 3875
rect 6035 3845 6036 3875
rect 6004 3844 6036 3845
rect 6004 3764 6036 3796
rect 6004 3715 6036 3716
rect 6004 3685 6005 3715
rect 6005 3685 6035 3715
rect 6035 3685 6036 3715
rect 6004 3684 6036 3685
rect 6004 3635 6036 3636
rect 6004 3605 6005 3635
rect 6005 3605 6035 3635
rect 6035 3605 6036 3635
rect 6004 3604 6036 3605
rect 6004 3524 6036 3556
rect 6004 3475 6036 3476
rect 6004 3445 6005 3475
rect 6005 3445 6035 3475
rect 6035 3445 6036 3475
rect 6004 3444 6036 3445
rect 6004 3395 6036 3396
rect 6004 3365 6005 3395
rect 6005 3365 6035 3395
rect 6035 3365 6036 3395
rect 6004 3364 6036 3365
rect 6004 3284 6036 3316
rect 6004 3235 6036 3236
rect 6004 3205 6005 3235
rect 6005 3205 6035 3235
rect 6035 3205 6036 3235
rect 6004 3204 6036 3205
rect 6004 3155 6036 3156
rect 6004 3125 6005 3155
rect 6005 3125 6035 3155
rect 6035 3125 6036 3155
rect 6004 3124 6036 3125
rect 6004 3075 6036 3076
rect 6004 3045 6005 3075
rect 6005 3045 6035 3075
rect 6035 3045 6036 3075
rect 6004 3044 6036 3045
rect 6004 2995 6036 2996
rect 6004 2965 6005 2995
rect 6005 2965 6035 2995
rect 6035 2965 6036 2995
rect 6004 2964 6036 2965
rect 6004 2915 6036 2916
rect 6004 2885 6005 2915
rect 6005 2885 6035 2915
rect 6035 2885 6036 2915
rect 6004 2884 6036 2885
rect 6004 2835 6036 2836
rect 6004 2805 6005 2835
rect 6005 2805 6035 2835
rect 6035 2805 6036 2835
rect 6004 2804 6036 2805
rect 6004 2755 6036 2756
rect 6004 2725 6005 2755
rect 6005 2725 6035 2755
rect 6035 2725 6036 2755
rect 6004 2724 6036 2725
rect 6004 2675 6036 2676
rect 6004 2645 6005 2675
rect 6005 2645 6035 2675
rect 6035 2645 6036 2675
rect 6004 2644 6036 2645
rect 6004 2595 6036 2596
rect 6004 2565 6005 2595
rect 6005 2565 6035 2595
rect 6035 2565 6036 2595
rect 6004 2564 6036 2565
rect 6004 2515 6036 2516
rect 6004 2485 6005 2515
rect 6005 2485 6035 2515
rect 6035 2485 6036 2515
rect 6004 2484 6036 2485
rect 6004 2435 6036 2436
rect 6004 2405 6005 2435
rect 6005 2405 6035 2435
rect 6035 2405 6036 2435
rect 6004 2404 6036 2405
rect 6004 2355 6036 2356
rect 6004 2325 6005 2355
rect 6005 2325 6035 2355
rect 6035 2325 6036 2355
rect 6004 2324 6036 2325
rect 6004 2275 6036 2276
rect 6004 2245 6005 2275
rect 6005 2245 6035 2275
rect 6035 2245 6036 2275
rect 6004 2244 6036 2245
rect 6004 2195 6036 2196
rect 6004 2165 6005 2195
rect 6005 2165 6035 2195
rect 6035 2165 6036 2195
rect 6004 2164 6036 2165
rect 6004 2115 6036 2116
rect 6004 2085 6005 2115
rect 6005 2085 6035 2115
rect 6035 2085 6036 2115
rect 6004 2084 6036 2085
rect 6004 2035 6036 2036
rect 6004 2005 6005 2035
rect 6005 2005 6035 2035
rect 6035 2005 6036 2035
rect 6004 2004 6036 2005
rect 6004 1955 6036 1956
rect 6004 1925 6005 1955
rect 6005 1925 6035 1955
rect 6035 1925 6036 1955
rect 6004 1924 6036 1925
rect 6004 1844 6036 1876
rect 6004 1764 6036 1796
rect 6004 1715 6036 1716
rect 6004 1685 6005 1715
rect 6005 1685 6035 1715
rect 6035 1685 6036 1715
rect 6004 1684 6036 1685
rect 6004 1635 6036 1636
rect 6004 1605 6005 1635
rect 6005 1605 6035 1635
rect 6035 1605 6036 1635
rect 6004 1604 6036 1605
rect 6004 1555 6036 1556
rect 6004 1525 6005 1555
rect 6005 1525 6035 1555
rect 6035 1525 6036 1555
rect 6004 1524 6036 1525
rect 6004 1475 6036 1476
rect 6004 1445 6005 1475
rect 6005 1445 6035 1475
rect 6035 1445 6036 1475
rect 6004 1444 6036 1445
rect 6004 1395 6036 1396
rect 6004 1365 6005 1395
rect 6005 1365 6035 1395
rect 6035 1365 6036 1395
rect 6004 1364 6036 1365
rect 6004 1315 6036 1316
rect 6004 1285 6005 1315
rect 6005 1285 6035 1315
rect 6035 1285 6036 1315
rect 6004 1284 6036 1285
rect 6004 1235 6036 1236
rect 6004 1205 6005 1235
rect 6005 1205 6035 1235
rect 6035 1205 6036 1235
rect 6004 1204 6036 1205
rect 6004 1155 6036 1156
rect 6004 1125 6005 1155
rect 6005 1125 6035 1155
rect 6035 1125 6036 1155
rect 6004 1124 6036 1125
rect 6004 1075 6036 1076
rect 6004 1045 6005 1075
rect 6005 1045 6035 1075
rect 6035 1045 6036 1075
rect 6004 1044 6036 1045
rect 6004 995 6036 996
rect 6004 965 6005 995
rect 6005 965 6035 995
rect 6035 965 6036 995
rect 6004 964 6036 965
rect 6004 884 6036 916
rect 6004 835 6036 836
rect 6004 805 6005 835
rect 6005 805 6035 835
rect 6035 805 6036 835
rect 6004 804 6036 805
rect 6004 755 6036 756
rect 6004 725 6005 755
rect 6005 725 6035 755
rect 6035 725 6036 755
rect 6004 724 6036 725
rect 6004 675 6036 676
rect 6004 645 6005 675
rect 6005 645 6035 675
rect 6035 645 6036 675
rect 6004 644 6036 645
rect 6004 595 6036 596
rect 6004 565 6005 595
rect 6005 565 6035 595
rect 6035 565 6036 595
rect 6004 564 6036 565
rect 6004 515 6036 516
rect 6004 485 6005 515
rect 6005 485 6035 515
rect 6035 485 6036 515
rect 6004 484 6036 485
rect 6004 404 6036 436
rect 6004 324 6036 356
rect 6004 275 6036 276
rect 6004 245 6005 275
rect 6005 245 6035 275
rect 6035 245 6036 275
rect 6004 244 6036 245
rect 6004 195 6036 196
rect 6004 165 6005 195
rect 6005 165 6035 195
rect 6035 165 6036 195
rect 6004 164 6036 165
rect 6004 115 6036 116
rect 6004 85 6005 115
rect 6005 85 6035 115
rect 6035 85 6036 115
rect 6004 84 6036 85
rect 6004 35 6036 36
rect 6004 5 6005 35
rect 6005 5 6035 35
rect 6035 5 6036 35
rect 6004 4 6036 5
rect 6164 15715 6196 15716
rect 6164 15685 6165 15715
rect 6165 15685 6195 15715
rect 6195 15685 6196 15715
rect 6164 15684 6196 15685
rect 6164 15635 6196 15636
rect 6164 15605 6165 15635
rect 6165 15605 6195 15635
rect 6195 15605 6196 15635
rect 6164 15604 6196 15605
rect 6164 15555 6196 15556
rect 6164 15525 6165 15555
rect 6165 15525 6195 15555
rect 6195 15525 6196 15555
rect 6164 15524 6196 15525
rect 6164 15475 6196 15476
rect 6164 15445 6165 15475
rect 6165 15445 6195 15475
rect 6195 15445 6196 15475
rect 6164 15444 6196 15445
rect 6164 15395 6196 15396
rect 6164 15365 6165 15395
rect 6165 15365 6195 15395
rect 6195 15365 6196 15395
rect 6164 15364 6196 15365
rect 6164 15315 6196 15316
rect 6164 15285 6165 15315
rect 6165 15285 6195 15315
rect 6195 15285 6196 15315
rect 6164 15284 6196 15285
rect 6164 15235 6196 15236
rect 6164 15205 6165 15235
rect 6165 15205 6195 15235
rect 6195 15205 6196 15235
rect 6164 15204 6196 15205
rect 6164 15155 6196 15156
rect 6164 15125 6165 15155
rect 6165 15125 6195 15155
rect 6195 15125 6196 15155
rect 6164 15124 6196 15125
rect 6164 15044 6196 15076
rect 6164 14995 6196 14996
rect 6164 14965 6165 14995
rect 6165 14965 6195 14995
rect 6195 14965 6196 14995
rect 6164 14964 6196 14965
rect 6164 14915 6196 14916
rect 6164 14885 6165 14915
rect 6165 14885 6195 14915
rect 6195 14885 6196 14915
rect 6164 14884 6196 14885
rect 6164 14835 6196 14836
rect 6164 14805 6165 14835
rect 6165 14805 6195 14835
rect 6195 14805 6196 14835
rect 6164 14804 6196 14805
rect 6164 14755 6196 14756
rect 6164 14725 6165 14755
rect 6165 14725 6195 14755
rect 6195 14725 6196 14755
rect 6164 14724 6196 14725
rect 6164 14675 6196 14676
rect 6164 14645 6165 14675
rect 6165 14645 6195 14675
rect 6195 14645 6196 14675
rect 6164 14644 6196 14645
rect 6164 14595 6196 14596
rect 6164 14565 6165 14595
rect 6165 14565 6195 14595
rect 6195 14565 6196 14595
rect 6164 14564 6196 14565
rect 6164 14515 6196 14516
rect 6164 14485 6165 14515
rect 6165 14485 6195 14515
rect 6195 14485 6196 14515
rect 6164 14484 6196 14485
rect 6164 14435 6196 14436
rect 6164 14405 6165 14435
rect 6165 14405 6195 14435
rect 6195 14405 6196 14435
rect 6164 14404 6196 14405
rect 6164 14324 6196 14356
rect 6164 14244 6196 14276
rect 6164 14164 6196 14196
rect 6164 14084 6196 14116
rect 6164 14035 6196 14036
rect 6164 14005 6165 14035
rect 6165 14005 6195 14035
rect 6195 14005 6196 14035
rect 6164 14004 6196 14005
rect 6164 13955 6196 13956
rect 6164 13925 6165 13955
rect 6165 13925 6195 13955
rect 6195 13925 6196 13955
rect 6164 13924 6196 13925
rect 6164 13875 6196 13876
rect 6164 13845 6165 13875
rect 6165 13845 6195 13875
rect 6195 13845 6196 13875
rect 6164 13844 6196 13845
rect 6164 13795 6196 13796
rect 6164 13765 6165 13795
rect 6165 13765 6195 13795
rect 6195 13765 6196 13795
rect 6164 13764 6196 13765
rect 6164 13715 6196 13716
rect 6164 13685 6165 13715
rect 6165 13685 6195 13715
rect 6195 13685 6196 13715
rect 6164 13684 6196 13685
rect 6164 13635 6196 13636
rect 6164 13605 6165 13635
rect 6165 13605 6195 13635
rect 6195 13605 6196 13635
rect 6164 13604 6196 13605
rect 6164 13555 6196 13556
rect 6164 13525 6165 13555
rect 6165 13525 6195 13555
rect 6195 13525 6196 13555
rect 6164 13524 6196 13525
rect 6164 13475 6196 13476
rect 6164 13445 6165 13475
rect 6165 13445 6195 13475
rect 6195 13445 6196 13475
rect 6164 13444 6196 13445
rect 6164 13364 6196 13396
rect 6164 13284 6196 13316
rect 6164 13204 6196 13236
rect 6164 13124 6196 13156
rect 6164 13075 6196 13076
rect 6164 13045 6165 13075
rect 6165 13045 6195 13075
rect 6195 13045 6196 13075
rect 6164 13044 6196 13045
rect 6164 12995 6196 12996
rect 6164 12965 6165 12995
rect 6165 12965 6195 12995
rect 6195 12965 6196 12995
rect 6164 12964 6196 12965
rect 6164 12915 6196 12916
rect 6164 12885 6165 12915
rect 6165 12885 6195 12915
rect 6195 12885 6196 12915
rect 6164 12884 6196 12885
rect 6164 12835 6196 12836
rect 6164 12805 6165 12835
rect 6165 12805 6195 12835
rect 6195 12805 6196 12835
rect 6164 12804 6196 12805
rect 6164 12755 6196 12756
rect 6164 12725 6165 12755
rect 6165 12725 6195 12755
rect 6195 12725 6196 12755
rect 6164 12724 6196 12725
rect 6164 12675 6196 12676
rect 6164 12645 6165 12675
rect 6165 12645 6195 12675
rect 6195 12645 6196 12675
rect 6164 12644 6196 12645
rect 6164 12595 6196 12596
rect 6164 12565 6165 12595
rect 6165 12565 6195 12595
rect 6195 12565 6196 12595
rect 6164 12564 6196 12565
rect 6164 12515 6196 12516
rect 6164 12485 6165 12515
rect 6165 12485 6195 12515
rect 6195 12485 6196 12515
rect 6164 12484 6196 12485
rect 6164 12404 6196 12436
rect 6164 12355 6196 12356
rect 6164 12325 6165 12355
rect 6165 12325 6195 12355
rect 6195 12325 6196 12355
rect 6164 12324 6196 12325
rect 6164 12275 6196 12276
rect 6164 12245 6165 12275
rect 6165 12245 6195 12275
rect 6195 12245 6196 12275
rect 6164 12244 6196 12245
rect 6164 12195 6196 12196
rect 6164 12165 6165 12195
rect 6165 12165 6195 12195
rect 6195 12165 6196 12195
rect 6164 12164 6196 12165
rect 6164 12115 6196 12116
rect 6164 12085 6165 12115
rect 6165 12085 6195 12115
rect 6195 12085 6196 12115
rect 6164 12084 6196 12085
rect 6164 12035 6196 12036
rect 6164 12005 6165 12035
rect 6165 12005 6195 12035
rect 6195 12005 6196 12035
rect 6164 12004 6196 12005
rect 6164 11955 6196 11956
rect 6164 11925 6165 11955
rect 6165 11925 6195 11955
rect 6195 11925 6196 11955
rect 6164 11924 6196 11925
rect 6164 11875 6196 11876
rect 6164 11845 6165 11875
rect 6165 11845 6195 11875
rect 6195 11845 6196 11875
rect 6164 11844 6196 11845
rect 6164 11795 6196 11796
rect 6164 11765 6165 11795
rect 6165 11765 6195 11795
rect 6195 11765 6196 11795
rect 6164 11764 6196 11765
rect 6164 11715 6196 11716
rect 6164 11685 6165 11715
rect 6165 11685 6195 11715
rect 6195 11685 6196 11715
rect 6164 11684 6196 11685
rect 6164 11635 6196 11636
rect 6164 11605 6165 11635
rect 6165 11605 6195 11635
rect 6195 11605 6196 11635
rect 6164 11604 6196 11605
rect 6164 11555 6196 11556
rect 6164 11525 6165 11555
rect 6165 11525 6195 11555
rect 6195 11525 6196 11555
rect 6164 11524 6196 11525
rect 6164 11475 6196 11476
rect 6164 11445 6165 11475
rect 6165 11445 6195 11475
rect 6195 11445 6196 11475
rect 6164 11444 6196 11445
rect 6164 11395 6196 11396
rect 6164 11365 6165 11395
rect 6165 11365 6195 11395
rect 6195 11365 6196 11395
rect 6164 11364 6196 11365
rect 6164 11315 6196 11316
rect 6164 11285 6165 11315
rect 6165 11285 6195 11315
rect 6195 11285 6196 11315
rect 6164 11284 6196 11285
rect 6164 11235 6196 11236
rect 6164 11205 6165 11235
rect 6165 11205 6195 11235
rect 6195 11205 6196 11235
rect 6164 11204 6196 11205
rect 6164 11155 6196 11156
rect 6164 11125 6165 11155
rect 6165 11125 6195 11155
rect 6195 11125 6196 11155
rect 6164 11124 6196 11125
rect 6164 11075 6196 11076
rect 6164 11045 6165 11075
rect 6165 11045 6195 11075
rect 6195 11045 6196 11075
rect 6164 11044 6196 11045
rect 6164 10964 6196 10996
rect 6164 10915 6196 10916
rect 6164 10885 6165 10915
rect 6165 10885 6195 10915
rect 6195 10885 6196 10915
rect 6164 10884 6196 10885
rect 6164 10835 6196 10836
rect 6164 10805 6165 10835
rect 6165 10805 6195 10835
rect 6195 10805 6196 10835
rect 6164 10804 6196 10805
rect 6164 10755 6196 10756
rect 6164 10725 6165 10755
rect 6165 10725 6195 10755
rect 6195 10725 6196 10755
rect 6164 10724 6196 10725
rect 6164 10675 6196 10676
rect 6164 10645 6165 10675
rect 6165 10645 6195 10675
rect 6195 10645 6196 10675
rect 6164 10644 6196 10645
rect 6164 10595 6196 10596
rect 6164 10565 6165 10595
rect 6165 10565 6195 10595
rect 6195 10565 6196 10595
rect 6164 10564 6196 10565
rect 6164 10515 6196 10516
rect 6164 10485 6165 10515
rect 6165 10485 6195 10515
rect 6195 10485 6196 10515
rect 6164 10484 6196 10485
rect 6164 10435 6196 10436
rect 6164 10405 6165 10435
rect 6165 10405 6195 10435
rect 6195 10405 6196 10435
rect 6164 10404 6196 10405
rect 6164 10355 6196 10356
rect 6164 10325 6165 10355
rect 6165 10325 6195 10355
rect 6195 10325 6196 10355
rect 6164 10324 6196 10325
rect 6164 10244 6196 10276
rect 6164 10164 6196 10196
rect 6164 10084 6196 10116
rect 6164 10004 6196 10036
rect 6164 9955 6196 9956
rect 6164 9925 6165 9955
rect 6165 9925 6195 9955
rect 6195 9925 6196 9955
rect 6164 9924 6196 9925
rect 6164 9875 6196 9876
rect 6164 9845 6165 9875
rect 6165 9845 6195 9875
rect 6195 9845 6196 9875
rect 6164 9844 6196 9845
rect 6164 9795 6196 9796
rect 6164 9765 6165 9795
rect 6165 9765 6195 9795
rect 6195 9765 6196 9795
rect 6164 9764 6196 9765
rect 6164 9715 6196 9716
rect 6164 9685 6165 9715
rect 6165 9685 6195 9715
rect 6195 9685 6196 9715
rect 6164 9684 6196 9685
rect 6164 9635 6196 9636
rect 6164 9605 6165 9635
rect 6165 9605 6195 9635
rect 6195 9605 6196 9635
rect 6164 9604 6196 9605
rect 6164 9555 6196 9556
rect 6164 9525 6165 9555
rect 6165 9525 6195 9555
rect 6195 9525 6196 9555
rect 6164 9524 6196 9525
rect 6164 9475 6196 9476
rect 6164 9445 6165 9475
rect 6165 9445 6195 9475
rect 6195 9445 6196 9475
rect 6164 9444 6196 9445
rect 6164 9395 6196 9396
rect 6164 9365 6165 9395
rect 6165 9365 6195 9395
rect 6195 9365 6196 9395
rect 6164 9364 6196 9365
rect 6164 9284 6196 9316
rect 6164 9204 6196 9236
rect 6164 9124 6196 9156
rect 6164 9044 6196 9076
rect 6164 8995 6196 8996
rect 6164 8965 6165 8995
rect 6165 8965 6195 8995
rect 6195 8965 6196 8995
rect 6164 8964 6196 8965
rect 6164 8915 6196 8916
rect 6164 8885 6165 8915
rect 6165 8885 6195 8915
rect 6195 8885 6196 8915
rect 6164 8884 6196 8885
rect 6164 8835 6196 8836
rect 6164 8805 6165 8835
rect 6165 8805 6195 8835
rect 6195 8805 6196 8835
rect 6164 8804 6196 8805
rect 6164 8755 6196 8756
rect 6164 8725 6165 8755
rect 6165 8725 6195 8755
rect 6195 8725 6196 8755
rect 6164 8724 6196 8725
rect 6164 8675 6196 8676
rect 6164 8645 6165 8675
rect 6165 8645 6195 8675
rect 6195 8645 6196 8675
rect 6164 8644 6196 8645
rect 6164 8595 6196 8596
rect 6164 8565 6165 8595
rect 6165 8565 6195 8595
rect 6195 8565 6196 8595
rect 6164 8564 6196 8565
rect 6164 8515 6196 8516
rect 6164 8485 6165 8515
rect 6165 8485 6195 8515
rect 6195 8485 6196 8515
rect 6164 8484 6196 8485
rect 6164 8435 6196 8436
rect 6164 8405 6165 8435
rect 6165 8405 6195 8435
rect 6195 8405 6196 8435
rect 6164 8404 6196 8405
rect 6164 8324 6196 8356
rect 6164 8275 6196 8276
rect 6164 8245 6165 8275
rect 6165 8245 6195 8275
rect 6195 8245 6196 8275
rect 6164 8244 6196 8245
rect 6164 8195 6196 8196
rect 6164 8165 6165 8195
rect 6165 8165 6195 8195
rect 6195 8165 6196 8195
rect 6164 8164 6196 8165
rect 6164 8115 6196 8116
rect 6164 8085 6165 8115
rect 6165 8085 6195 8115
rect 6195 8085 6196 8115
rect 6164 8084 6196 8085
rect 6164 8035 6196 8036
rect 6164 8005 6165 8035
rect 6165 8005 6195 8035
rect 6195 8005 6196 8035
rect 6164 8004 6196 8005
rect 6164 7955 6196 7956
rect 6164 7925 6165 7955
rect 6165 7925 6195 7955
rect 6195 7925 6196 7955
rect 6164 7924 6196 7925
rect 6164 7875 6196 7876
rect 6164 7845 6165 7875
rect 6165 7845 6195 7875
rect 6195 7845 6196 7875
rect 6164 7844 6196 7845
rect 6164 7795 6196 7796
rect 6164 7765 6165 7795
rect 6165 7765 6195 7795
rect 6195 7765 6196 7795
rect 6164 7764 6196 7765
rect 6164 7715 6196 7716
rect 6164 7685 6165 7715
rect 6165 7685 6195 7715
rect 6195 7685 6196 7715
rect 6164 7684 6196 7685
rect 6164 7635 6196 7636
rect 6164 7605 6165 7635
rect 6165 7605 6195 7635
rect 6195 7605 6196 7635
rect 6164 7604 6196 7605
rect 6164 7555 6196 7556
rect 6164 7525 6165 7555
rect 6165 7525 6195 7555
rect 6195 7525 6196 7555
rect 6164 7524 6196 7525
rect 6164 7475 6196 7476
rect 6164 7445 6165 7475
rect 6165 7445 6195 7475
rect 6195 7445 6196 7475
rect 6164 7444 6196 7445
rect 6164 7395 6196 7396
rect 6164 7365 6165 7395
rect 6165 7365 6195 7395
rect 6195 7365 6196 7395
rect 6164 7364 6196 7365
rect 6164 7315 6196 7316
rect 6164 7285 6165 7315
rect 6165 7285 6195 7315
rect 6195 7285 6196 7315
rect 6164 7284 6196 7285
rect 6164 7235 6196 7236
rect 6164 7205 6165 7235
rect 6165 7205 6195 7235
rect 6195 7205 6196 7235
rect 6164 7204 6196 7205
rect 6164 7155 6196 7156
rect 6164 7125 6165 7155
rect 6165 7125 6195 7155
rect 6195 7125 6196 7155
rect 6164 7124 6196 7125
rect 6164 7075 6196 7076
rect 6164 7045 6165 7075
rect 6165 7045 6195 7075
rect 6195 7045 6196 7075
rect 6164 7044 6196 7045
rect 6164 6995 6196 6996
rect 6164 6965 6165 6995
rect 6165 6965 6195 6995
rect 6195 6965 6196 6995
rect 6164 6964 6196 6965
rect 6164 6884 6196 6916
rect 6164 6835 6196 6836
rect 6164 6805 6165 6835
rect 6165 6805 6195 6835
rect 6195 6805 6196 6835
rect 6164 6804 6196 6805
rect 6164 6755 6196 6756
rect 6164 6725 6165 6755
rect 6165 6725 6195 6755
rect 6195 6725 6196 6755
rect 6164 6724 6196 6725
rect 6164 6675 6196 6676
rect 6164 6645 6165 6675
rect 6165 6645 6195 6675
rect 6195 6645 6196 6675
rect 6164 6644 6196 6645
rect 6164 6595 6196 6596
rect 6164 6565 6165 6595
rect 6165 6565 6195 6595
rect 6195 6565 6196 6595
rect 6164 6564 6196 6565
rect 6164 6515 6196 6516
rect 6164 6485 6165 6515
rect 6165 6485 6195 6515
rect 6195 6485 6196 6515
rect 6164 6484 6196 6485
rect 6164 6435 6196 6436
rect 6164 6405 6165 6435
rect 6165 6405 6195 6435
rect 6195 6405 6196 6435
rect 6164 6404 6196 6405
rect 6164 6355 6196 6356
rect 6164 6325 6165 6355
rect 6165 6325 6195 6355
rect 6195 6325 6196 6355
rect 6164 6324 6196 6325
rect 6164 6275 6196 6276
rect 6164 6245 6165 6275
rect 6165 6245 6195 6275
rect 6195 6245 6196 6275
rect 6164 6244 6196 6245
rect 6164 6164 6196 6196
rect 6164 6084 6196 6116
rect 6164 6004 6196 6036
rect 6164 5924 6196 5956
rect 6164 5875 6196 5876
rect 6164 5845 6165 5875
rect 6165 5845 6195 5875
rect 6195 5845 6196 5875
rect 6164 5844 6196 5845
rect 6164 5795 6196 5796
rect 6164 5765 6165 5795
rect 6165 5765 6195 5795
rect 6195 5765 6196 5795
rect 6164 5764 6196 5765
rect 6164 5715 6196 5716
rect 6164 5685 6165 5715
rect 6165 5685 6195 5715
rect 6195 5685 6196 5715
rect 6164 5684 6196 5685
rect 6164 5635 6196 5636
rect 6164 5605 6165 5635
rect 6165 5605 6195 5635
rect 6195 5605 6196 5635
rect 6164 5604 6196 5605
rect 6164 5555 6196 5556
rect 6164 5525 6165 5555
rect 6165 5525 6195 5555
rect 6195 5525 6196 5555
rect 6164 5524 6196 5525
rect 6164 5475 6196 5476
rect 6164 5445 6165 5475
rect 6165 5445 6195 5475
rect 6195 5445 6196 5475
rect 6164 5444 6196 5445
rect 6164 5395 6196 5396
rect 6164 5365 6165 5395
rect 6165 5365 6195 5395
rect 6195 5365 6196 5395
rect 6164 5364 6196 5365
rect 6164 5315 6196 5316
rect 6164 5285 6165 5315
rect 6165 5285 6195 5315
rect 6195 5285 6196 5315
rect 6164 5284 6196 5285
rect 6164 5235 6196 5236
rect 6164 5205 6165 5235
rect 6165 5205 6195 5235
rect 6195 5205 6196 5235
rect 6164 5204 6196 5205
rect 6164 5155 6196 5156
rect 6164 5125 6165 5155
rect 6165 5125 6195 5155
rect 6195 5125 6196 5155
rect 6164 5124 6196 5125
rect 6164 5075 6196 5076
rect 6164 5045 6165 5075
rect 6165 5045 6195 5075
rect 6195 5045 6196 5075
rect 6164 5044 6196 5045
rect 6164 4995 6196 4996
rect 6164 4965 6165 4995
rect 6165 4965 6195 4995
rect 6195 4965 6196 4995
rect 6164 4964 6196 4965
rect 6164 4915 6196 4916
rect 6164 4885 6165 4915
rect 6165 4885 6195 4915
rect 6195 4885 6196 4915
rect 6164 4884 6196 4885
rect 6164 4804 6196 4836
rect 6164 4755 6196 4756
rect 6164 4725 6165 4755
rect 6165 4725 6195 4755
rect 6195 4725 6196 4755
rect 6164 4724 6196 4725
rect 6164 4675 6196 4676
rect 6164 4645 6165 4675
rect 6165 4645 6195 4675
rect 6195 4645 6196 4675
rect 6164 4644 6196 4645
rect 6164 4564 6196 4596
rect 6164 4515 6196 4516
rect 6164 4485 6165 4515
rect 6165 4485 6195 4515
rect 6195 4485 6196 4515
rect 6164 4484 6196 4485
rect 6164 4435 6196 4436
rect 6164 4405 6165 4435
rect 6165 4405 6195 4435
rect 6195 4405 6196 4435
rect 6164 4404 6196 4405
rect 6164 4355 6196 4356
rect 6164 4325 6165 4355
rect 6165 4325 6195 4355
rect 6195 4325 6196 4355
rect 6164 4324 6196 4325
rect 6164 4275 6196 4276
rect 6164 4245 6165 4275
rect 6165 4245 6195 4275
rect 6195 4245 6196 4275
rect 6164 4244 6196 4245
rect 6164 4195 6196 4196
rect 6164 4165 6165 4195
rect 6165 4165 6195 4195
rect 6195 4165 6196 4195
rect 6164 4164 6196 4165
rect 6164 4115 6196 4116
rect 6164 4085 6165 4115
rect 6165 4085 6195 4115
rect 6195 4085 6196 4115
rect 6164 4084 6196 4085
rect 6164 4035 6196 4036
rect 6164 4005 6165 4035
rect 6165 4005 6195 4035
rect 6195 4005 6196 4035
rect 6164 4004 6196 4005
rect 6164 3955 6196 3956
rect 6164 3925 6165 3955
rect 6165 3925 6195 3955
rect 6195 3925 6196 3955
rect 6164 3924 6196 3925
rect 6164 3875 6196 3876
rect 6164 3845 6165 3875
rect 6165 3845 6195 3875
rect 6195 3845 6196 3875
rect 6164 3844 6196 3845
rect 6164 3764 6196 3796
rect 6164 3715 6196 3716
rect 6164 3685 6165 3715
rect 6165 3685 6195 3715
rect 6195 3685 6196 3715
rect 6164 3684 6196 3685
rect 6164 3635 6196 3636
rect 6164 3605 6165 3635
rect 6165 3605 6195 3635
rect 6195 3605 6196 3635
rect 6164 3604 6196 3605
rect 6164 3524 6196 3556
rect 6164 3475 6196 3476
rect 6164 3445 6165 3475
rect 6165 3445 6195 3475
rect 6195 3445 6196 3475
rect 6164 3444 6196 3445
rect 6164 3395 6196 3396
rect 6164 3365 6165 3395
rect 6165 3365 6195 3395
rect 6195 3365 6196 3395
rect 6164 3364 6196 3365
rect 6164 3284 6196 3316
rect 6164 3235 6196 3236
rect 6164 3205 6165 3235
rect 6165 3205 6195 3235
rect 6195 3205 6196 3235
rect 6164 3204 6196 3205
rect 6164 3155 6196 3156
rect 6164 3125 6165 3155
rect 6165 3125 6195 3155
rect 6195 3125 6196 3155
rect 6164 3124 6196 3125
rect 6164 3075 6196 3076
rect 6164 3045 6165 3075
rect 6165 3045 6195 3075
rect 6195 3045 6196 3075
rect 6164 3044 6196 3045
rect 6164 2995 6196 2996
rect 6164 2965 6165 2995
rect 6165 2965 6195 2995
rect 6195 2965 6196 2995
rect 6164 2964 6196 2965
rect 6164 2915 6196 2916
rect 6164 2885 6165 2915
rect 6165 2885 6195 2915
rect 6195 2885 6196 2915
rect 6164 2884 6196 2885
rect 6164 2835 6196 2836
rect 6164 2805 6165 2835
rect 6165 2805 6195 2835
rect 6195 2805 6196 2835
rect 6164 2804 6196 2805
rect 6164 2755 6196 2756
rect 6164 2725 6165 2755
rect 6165 2725 6195 2755
rect 6195 2725 6196 2755
rect 6164 2724 6196 2725
rect 6164 2675 6196 2676
rect 6164 2645 6165 2675
rect 6165 2645 6195 2675
rect 6195 2645 6196 2675
rect 6164 2644 6196 2645
rect 6164 2595 6196 2596
rect 6164 2565 6165 2595
rect 6165 2565 6195 2595
rect 6195 2565 6196 2595
rect 6164 2564 6196 2565
rect 6164 2515 6196 2516
rect 6164 2485 6165 2515
rect 6165 2485 6195 2515
rect 6195 2485 6196 2515
rect 6164 2484 6196 2485
rect 6164 2435 6196 2436
rect 6164 2405 6165 2435
rect 6165 2405 6195 2435
rect 6195 2405 6196 2435
rect 6164 2404 6196 2405
rect 6164 2355 6196 2356
rect 6164 2325 6165 2355
rect 6165 2325 6195 2355
rect 6195 2325 6196 2355
rect 6164 2324 6196 2325
rect 6164 2275 6196 2276
rect 6164 2245 6165 2275
rect 6165 2245 6195 2275
rect 6195 2245 6196 2275
rect 6164 2244 6196 2245
rect 6164 2195 6196 2196
rect 6164 2165 6165 2195
rect 6165 2165 6195 2195
rect 6195 2165 6196 2195
rect 6164 2164 6196 2165
rect 6164 2115 6196 2116
rect 6164 2085 6165 2115
rect 6165 2085 6195 2115
rect 6195 2085 6196 2115
rect 6164 2084 6196 2085
rect 6164 2035 6196 2036
rect 6164 2005 6165 2035
rect 6165 2005 6195 2035
rect 6195 2005 6196 2035
rect 6164 2004 6196 2005
rect 6164 1955 6196 1956
rect 6164 1925 6165 1955
rect 6165 1925 6195 1955
rect 6195 1925 6196 1955
rect 6164 1924 6196 1925
rect 6164 1844 6196 1876
rect 6164 1764 6196 1796
rect 6164 1715 6196 1716
rect 6164 1685 6165 1715
rect 6165 1685 6195 1715
rect 6195 1685 6196 1715
rect 6164 1684 6196 1685
rect 6164 1635 6196 1636
rect 6164 1605 6165 1635
rect 6165 1605 6195 1635
rect 6195 1605 6196 1635
rect 6164 1604 6196 1605
rect 6164 1555 6196 1556
rect 6164 1525 6165 1555
rect 6165 1525 6195 1555
rect 6195 1525 6196 1555
rect 6164 1524 6196 1525
rect 6164 1475 6196 1476
rect 6164 1445 6165 1475
rect 6165 1445 6195 1475
rect 6195 1445 6196 1475
rect 6164 1444 6196 1445
rect 6164 1395 6196 1396
rect 6164 1365 6165 1395
rect 6165 1365 6195 1395
rect 6195 1365 6196 1395
rect 6164 1364 6196 1365
rect 6164 1315 6196 1316
rect 6164 1285 6165 1315
rect 6165 1285 6195 1315
rect 6195 1285 6196 1315
rect 6164 1284 6196 1285
rect 6164 1235 6196 1236
rect 6164 1205 6165 1235
rect 6165 1205 6195 1235
rect 6195 1205 6196 1235
rect 6164 1204 6196 1205
rect 6164 1155 6196 1156
rect 6164 1125 6165 1155
rect 6165 1125 6195 1155
rect 6195 1125 6196 1155
rect 6164 1124 6196 1125
rect 6164 1075 6196 1076
rect 6164 1045 6165 1075
rect 6165 1045 6195 1075
rect 6195 1045 6196 1075
rect 6164 1044 6196 1045
rect 6164 995 6196 996
rect 6164 965 6165 995
rect 6165 965 6195 995
rect 6195 965 6196 995
rect 6164 964 6196 965
rect 6164 884 6196 916
rect 6164 835 6196 836
rect 6164 805 6165 835
rect 6165 805 6195 835
rect 6195 805 6196 835
rect 6164 804 6196 805
rect 6164 755 6196 756
rect 6164 725 6165 755
rect 6165 725 6195 755
rect 6195 725 6196 755
rect 6164 724 6196 725
rect 6164 675 6196 676
rect 6164 645 6165 675
rect 6165 645 6195 675
rect 6195 645 6196 675
rect 6164 644 6196 645
rect 6164 595 6196 596
rect 6164 565 6165 595
rect 6165 565 6195 595
rect 6195 565 6196 595
rect 6164 564 6196 565
rect 6164 515 6196 516
rect 6164 485 6165 515
rect 6165 485 6195 515
rect 6195 485 6196 515
rect 6164 484 6196 485
rect 6164 404 6196 436
rect 6164 324 6196 356
rect 6164 275 6196 276
rect 6164 245 6165 275
rect 6165 245 6195 275
rect 6195 245 6196 275
rect 6164 244 6196 245
rect 6164 195 6196 196
rect 6164 165 6165 195
rect 6165 165 6195 195
rect 6195 165 6196 195
rect 6164 164 6196 165
rect 6164 115 6196 116
rect 6164 85 6165 115
rect 6165 85 6195 115
rect 6195 85 6196 115
rect 6164 84 6196 85
rect 6164 35 6196 36
rect 6164 5 6165 35
rect 6165 5 6195 35
rect 6195 5 6196 35
rect 6164 4 6196 5
rect 6004 -716 6036 -524
rect 6164 -716 6196 -524
rect 4644 -1036 4676 -1004
rect 10284 -1036 10316 -1004
rect 244 -1116 276 -1084
rect 1204 -1116 1236 -1084
rect 1364 -1116 1396 -1084
rect 2324 -1116 2356 -1084
rect 2484 -1116 2516 -1084
rect 3444 -1116 3476 -1084
rect 3604 -1116 3636 -1084
rect 4564 -1116 4596 -1084
rect 4724 -1116 4756 -1084
rect 5684 -1116 5716 -1084
rect 5844 -1116 5876 -1084
rect 6804 -1116 6836 -1084
rect 6964 -1116 6996 -1084
rect 7924 -1116 7956 -1084
rect 8084 -1116 8116 -1084
rect 9044 -1116 9076 -1084
rect 9204 -1116 9236 -1084
rect 10164 -1116 10196 -1084
rect 124 -2316 156 -2284
rect 10284 -2316 10316 -2284
<< mimcap >>
rect 280 -1240 1200 -1200
rect 280 -2160 320 -1240
rect 1160 -2160 1200 -1240
rect 280 -2200 1200 -2160
rect 1400 -1240 2320 -1200
rect 1400 -2160 1440 -1240
rect 2280 -2160 2320 -1240
rect 1400 -2200 2320 -2160
rect 2520 -1240 3440 -1200
rect 2520 -2160 2560 -1240
rect 3400 -2160 3440 -1240
rect 2520 -2200 3440 -2160
rect 3640 -1240 4560 -1200
rect 3640 -2160 3680 -1240
rect 4520 -2160 4560 -1240
rect 3640 -2200 4560 -2160
rect 4760 -1240 5680 -1200
rect 4760 -2160 4800 -1240
rect 5640 -2160 5680 -1240
rect 4760 -2200 5680 -2160
rect 5880 -1240 6800 -1200
rect 5880 -2160 5920 -1240
rect 6760 -2160 6800 -1240
rect 5880 -2200 6800 -2160
rect 7000 -1240 7920 -1200
rect 7000 -2160 7040 -1240
rect 7880 -2160 7920 -1240
rect 7000 -2200 7920 -2160
rect 8120 -1240 9040 -1200
rect 8120 -2160 8160 -1240
rect 9000 -2160 9040 -1240
rect 8120 -2200 9040 -2160
rect 9240 -1240 10160 -1200
rect 9240 -2160 9280 -1240
rect 10120 -2160 10160 -1240
rect 9240 -2200 10160 -2160
<< mimcapcontact >>
rect 320 -2160 1160 -1240
rect 1440 -2160 2280 -1240
rect 2560 -2160 3400 -1240
rect 3680 -2160 4520 -1240
rect 4800 -2160 5640 -1240
rect 5920 -2160 6760 -1240
rect 7040 -2160 7880 -1240
rect 8160 -2160 9000 -1240
rect 9280 -2160 10120 -1240
<< metal4 >>
rect 4240 15716 4440 15720
rect 4240 15684 4244 15716
rect 4276 15684 4404 15716
rect 4436 15684 4440 15716
rect 4240 15680 4440 15684
rect 4480 15716 4680 15720
rect 4480 15684 4484 15716
rect 4516 15684 4644 15716
rect 4676 15684 4680 15716
rect 4480 15680 4680 15684
rect 4720 15716 5720 15720
rect 4720 15684 4724 15716
rect 4756 15684 4884 15716
rect 4916 15684 5044 15716
rect 5076 15684 5204 15716
rect 5236 15684 5364 15716
rect 5396 15684 5524 15716
rect 5556 15684 5684 15716
rect 5716 15684 5720 15716
rect 4720 15680 5720 15684
rect 5760 15716 5960 15720
rect 5760 15684 5764 15716
rect 5796 15684 5924 15716
rect 5956 15684 5960 15716
rect 5760 15680 5960 15684
rect 6000 15716 6200 15720
rect 6000 15684 6004 15716
rect 6036 15684 6164 15716
rect 6196 15684 6200 15716
rect 6000 15680 6200 15684
rect 4240 15636 4440 15640
rect 4240 15604 4244 15636
rect 4276 15604 4404 15636
rect 4436 15604 4440 15636
rect 4240 15600 4440 15604
rect 4480 15636 4680 15640
rect 4480 15604 4484 15636
rect 4516 15604 4644 15636
rect 4676 15604 4680 15636
rect 4480 15600 4680 15604
rect 4720 15636 5720 15640
rect 4720 15604 4724 15636
rect 4756 15604 4884 15636
rect 4916 15604 5044 15636
rect 5076 15604 5204 15636
rect 5236 15604 5364 15636
rect 5396 15604 5524 15636
rect 5556 15604 5684 15636
rect 5716 15604 5720 15636
rect 4720 15600 5720 15604
rect 5760 15636 5960 15640
rect 5760 15604 5764 15636
rect 5796 15604 5924 15636
rect 5956 15604 5960 15636
rect 5760 15600 5960 15604
rect 6000 15636 6200 15640
rect 6000 15604 6004 15636
rect 6036 15604 6164 15636
rect 6196 15604 6200 15636
rect 6000 15600 6200 15604
rect 4240 15556 4440 15560
rect 4240 15524 4244 15556
rect 4276 15524 4404 15556
rect 4436 15524 4440 15556
rect 4240 15520 4440 15524
rect 4480 15556 4680 15560
rect 4480 15524 4484 15556
rect 4516 15524 4644 15556
rect 4676 15524 4680 15556
rect 4480 15520 4680 15524
rect 4720 15556 5720 15560
rect 4720 15524 4724 15556
rect 4756 15524 4884 15556
rect 4916 15524 5044 15556
rect 5076 15524 5204 15556
rect 5236 15524 5364 15556
rect 5396 15524 5524 15556
rect 5556 15524 5684 15556
rect 5716 15524 5720 15556
rect 4720 15520 5720 15524
rect 5760 15556 5960 15560
rect 5760 15524 5764 15556
rect 5796 15524 5924 15556
rect 5956 15524 5960 15556
rect 5760 15520 5960 15524
rect 6000 15556 6200 15560
rect 6000 15524 6004 15556
rect 6036 15524 6164 15556
rect 6196 15524 6200 15556
rect 6000 15520 6200 15524
rect 4240 15476 4440 15480
rect 4240 15444 4244 15476
rect 4276 15444 4404 15476
rect 4436 15444 4440 15476
rect 4240 15440 4440 15444
rect 4480 15476 4680 15480
rect 4480 15444 4484 15476
rect 4516 15444 4644 15476
rect 4676 15444 4680 15476
rect 4480 15440 4680 15444
rect 4720 15476 5720 15480
rect 4720 15444 4724 15476
rect 4756 15444 4884 15476
rect 4916 15444 5044 15476
rect 5076 15444 5204 15476
rect 5236 15444 5364 15476
rect 5396 15444 5524 15476
rect 5556 15444 5684 15476
rect 5716 15444 5720 15476
rect 4720 15440 5720 15444
rect 5760 15476 5960 15480
rect 5760 15444 5764 15476
rect 5796 15444 5924 15476
rect 5956 15444 5960 15476
rect 5760 15440 5960 15444
rect 6000 15476 6200 15480
rect 6000 15444 6004 15476
rect 6036 15444 6164 15476
rect 6196 15444 6200 15476
rect 6000 15440 6200 15444
rect 4240 15396 4440 15400
rect 4240 15364 4244 15396
rect 4276 15364 4404 15396
rect 4436 15364 4440 15396
rect 4240 15360 4440 15364
rect 4480 15396 4680 15400
rect 4480 15364 4484 15396
rect 4516 15364 4644 15396
rect 4676 15364 4680 15396
rect 4480 15360 4680 15364
rect 4720 15396 5720 15400
rect 4720 15364 4724 15396
rect 4756 15364 4884 15396
rect 4916 15364 5044 15396
rect 5076 15364 5204 15396
rect 5236 15364 5364 15396
rect 5396 15364 5524 15396
rect 5556 15364 5684 15396
rect 5716 15364 5720 15396
rect 4720 15360 5720 15364
rect 5760 15396 5960 15400
rect 5760 15364 5764 15396
rect 5796 15364 5924 15396
rect 5956 15364 5960 15396
rect 5760 15360 5960 15364
rect 6000 15396 6200 15400
rect 6000 15364 6004 15396
rect 6036 15364 6164 15396
rect 6196 15364 6200 15396
rect 6000 15360 6200 15364
rect 4240 15316 4440 15320
rect 4240 15284 4244 15316
rect 4276 15284 4404 15316
rect 4436 15284 4440 15316
rect 4240 15280 4440 15284
rect 4480 15316 4680 15320
rect 4480 15284 4484 15316
rect 4516 15284 4644 15316
rect 4676 15284 4680 15316
rect 4480 15280 4680 15284
rect 4720 15316 5720 15320
rect 4720 15284 4724 15316
rect 4756 15284 4884 15316
rect 4916 15284 5044 15316
rect 5076 15284 5204 15316
rect 5236 15284 5364 15316
rect 5396 15284 5524 15316
rect 5556 15284 5684 15316
rect 5716 15284 5720 15316
rect 4720 15280 5720 15284
rect 5760 15316 5960 15320
rect 5760 15284 5764 15316
rect 5796 15284 5924 15316
rect 5956 15284 5960 15316
rect 5760 15280 5960 15284
rect 6000 15316 6200 15320
rect 6000 15284 6004 15316
rect 6036 15284 6164 15316
rect 6196 15284 6200 15316
rect 6000 15280 6200 15284
rect 4240 15236 4440 15240
rect 4240 15204 4244 15236
rect 4276 15204 4404 15236
rect 4436 15204 4440 15236
rect 4240 15200 4440 15204
rect 4480 15236 4680 15240
rect 4480 15204 4484 15236
rect 4516 15204 4644 15236
rect 4676 15204 4680 15236
rect 4480 15200 4680 15204
rect 4720 15236 5720 15240
rect 4720 15204 4724 15236
rect 4756 15204 4884 15236
rect 4916 15204 5044 15236
rect 5076 15204 5204 15236
rect 5236 15204 5364 15236
rect 5396 15204 5524 15236
rect 5556 15204 5684 15236
rect 5716 15204 5720 15236
rect 4720 15200 5720 15204
rect 5760 15236 5960 15240
rect 5760 15204 5764 15236
rect 5796 15204 5924 15236
rect 5956 15204 5960 15236
rect 5760 15200 5960 15204
rect 6000 15236 6200 15240
rect 6000 15204 6004 15236
rect 6036 15204 6164 15236
rect 6196 15204 6200 15236
rect 6000 15200 6200 15204
rect 4240 15156 4440 15160
rect 4240 15124 4244 15156
rect 4276 15124 4404 15156
rect 4436 15124 4440 15156
rect 4240 15120 4440 15124
rect 4480 15156 4680 15160
rect 4480 15124 4484 15156
rect 4516 15124 4644 15156
rect 4676 15124 4680 15156
rect 4480 15120 4680 15124
rect 4720 15156 5720 15160
rect 4720 15124 4724 15156
rect 4756 15124 4884 15156
rect 4916 15124 5044 15156
rect 5076 15124 5204 15156
rect 5236 15124 5364 15156
rect 5396 15124 5524 15156
rect 5556 15124 5684 15156
rect 5716 15124 5720 15156
rect 4720 15120 5720 15124
rect 5760 15156 5960 15160
rect 5760 15124 5764 15156
rect 5796 15124 5924 15156
rect 5956 15124 5960 15156
rect 5760 15120 5960 15124
rect 6000 15156 6200 15160
rect 6000 15124 6004 15156
rect 6036 15124 6164 15156
rect 6196 15124 6200 15156
rect 6000 15120 6200 15124
rect 4240 15076 4440 15080
rect 4240 15044 4244 15076
rect 4276 15044 4404 15076
rect 4436 15044 4440 15076
rect 4240 15040 4440 15044
rect 4480 15076 4680 15080
rect 4480 15044 4484 15076
rect 4516 15044 4644 15076
rect 4676 15044 4680 15076
rect 4480 15040 4680 15044
rect 4720 15076 5720 15080
rect 4720 15044 4724 15076
rect 4756 15044 4884 15076
rect 4916 15044 5044 15076
rect 5076 15044 5204 15076
rect 5236 15044 5364 15076
rect 5396 15044 5524 15076
rect 5556 15044 5684 15076
rect 5716 15044 5720 15076
rect 4720 15040 5720 15044
rect 5760 15076 5960 15080
rect 5760 15044 5764 15076
rect 5796 15044 5924 15076
rect 5956 15044 5960 15076
rect 5760 15040 5960 15044
rect 6000 15076 6200 15080
rect 6000 15044 6004 15076
rect 6036 15044 6164 15076
rect 6196 15044 6200 15076
rect 6000 15040 6200 15044
rect 4240 14996 4440 15000
rect 4240 14964 4244 14996
rect 4276 14964 4404 14996
rect 4436 14964 4440 14996
rect 4240 14960 4440 14964
rect 4480 14996 4680 15000
rect 4480 14964 4484 14996
rect 4516 14964 4644 14996
rect 4676 14964 4680 14996
rect 4480 14960 4680 14964
rect 4720 14996 5720 15000
rect 4720 14964 4724 14996
rect 4756 14964 4884 14996
rect 4916 14964 5044 14996
rect 5076 14964 5204 14996
rect 5236 14964 5364 14996
rect 5396 14964 5524 14996
rect 5556 14964 5684 14996
rect 5716 14964 5720 14996
rect 4720 14960 5720 14964
rect 5760 14996 5960 15000
rect 5760 14964 5764 14996
rect 5796 14964 5924 14996
rect 5956 14964 5960 14996
rect 5760 14960 5960 14964
rect 6000 14996 6200 15000
rect 6000 14964 6004 14996
rect 6036 14964 6164 14996
rect 6196 14964 6200 14996
rect 6000 14960 6200 14964
rect 4240 14916 4440 14920
rect 4240 14884 4244 14916
rect 4276 14884 4404 14916
rect 4436 14884 4440 14916
rect 4240 14880 4440 14884
rect 4480 14916 4680 14920
rect 4480 14884 4484 14916
rect 4516 14884 4644 14916
rect 4676 14884 4680 14916
rect 4480 14880 4680 14884
rect 4720 14916 5720 14920
rect 4720 14884 4724 14916
rect 4756 14884 4884 14916
rect 4916 14884 5044 14916
rect 5076 14884 5204 14916
rect 5236 14884 5364 14916
rect 5396 14884 5524 14916
rect 5556 14884 5684 14916
rect 5716 14884 5720 14916
rect 4720 14880 5720 14884
rect 5760 14916 5960 14920
rect 5760 14884 5764 14916
rect 5796 14884 5924 14916
rect 5956 14884 5960 14916
rect 5760 14880 5960 14884
rect 6000 14916 6200 14920
rect 6000 14884 6004 14916
rect 6036 14884 6164 14916
rect 6196 14884 6200 14916
rect 6000 14880 6200 14884
rect 4240 14836 4440 14840
rect 4240 14804 4244 14836
rect 4276 14804 4404 14836
rect 4436 14804 4440 14836
rect 4240 14800 4440 14804
rect 4480 14836 4680 14840
rect 4480 14804 4484 14836
rect 4516 14804 4644 14836
rect 4676 14804 4680 14836
rect 4480 14800 4680 14804
rect 4720 14836 5720 14840
rect 4720 14804 4724 14836
rect 4756 14804 4884 14836
rect 4916 14804 5044 14836
rect 5076 14804 5204 14836
rect 5236 14804 5364 14836
rect 5396 14804 5524 14836
rect 5556 14804 5684 14836
rect 5716 14804 5720 14836
rect 4720 14800 5720 14804
rect 5760 14836 5960 14840
rect 5760 14804 5764 14836
rect 5796 14804 5924 14836
rect 5956 14804 5960 14836
rect 5760 14800 5960 14804
rect 6000 14836 6200 14840
rect 6000 14804 6004 14836
rect 6036 14804 6164 14836
rect 6196 14804 6200 14836
rect 6000 14800 6200 14804
rect 4240 14756 4440 14760
rect 4240 14724 4244 14756
rect 4276 14724 4404 14756
rect 4436 14724 4440 14756
rect 4240 14720 4440 14724
rect 4480 14756 4680 14760
rect 4480 14724 4484 14756
rect 4516 14724 4644 14756
rect 4676 14724 4680 14756
rect 4480 14720 4680 14724
rect 4720 14756 5720 14760
rect 4720 14724 4724 14756
rect 4756 14724 4884 14756
rect 4916 14724 5044 14756
rect 5076 14724 5204 14756
rect 5236 14724 5364 14756
rect 5396 14724 5524 14756
rect 5556 14724 5684 14756
rect 5716 14724 5720 14756
rect 4720 14720 5720 14724
rect 5760 14756 5960 14760
rect 5760 14724 5764 14756
rect 5796 14724 5924 14756
rect 5956 14724 5960 14756
rect 5760 14720 5960 14724
rect 6000 14756 6200 14760
rect 6000 14724 6004 14756
rect 6036 14724 6164 14756
rect 6196 14724 6200 14756
rect 6000 14720 6200 14724
rect 4240 14676 4440 14680
rect 4240 14644 4244 14676
rect 4276 14644 4404 14676
rect 4436 14644 4440 14676
rect 4240 14640 4440 14644
rect 4480 14676 4680 14680
rect 4480 14644 4484 14676
rect 4516 14644 4644 14676
rect 4676 14644 4680 14676
rect 4480 14640 4680 14644
rect 4720 14676 5720 14680
rect 4720 14644 4724 14676
rect 4756 14644 4884 14676
rect 4916 14644 5044 14676
rect 5076 14644 5204 14676
rect 5236 14644 5364 14676
rect 5396 14644 5524 14676
rect 5556 14644 5684 14676
rect 5716 14644 5720 14676
rect 4720 14640 5720 14644
rect 5760 14676 5960 14680
rect 5760 14644 5764 14676
rect 5796 14644 5924 14676
rect 5956 14644 5960 14676
rect 5760 14640 5960 14644
rect 6000 14676 6200 14680
rect 6000 14644 6004 14676
rect 6036 14644 6164 14676
rect 6196 14644 6200 14676
rect 6000 14640 6200 14644
rect 4240 14596 4440 14600
rect 4240 14564 4244 14596
rect 4276 14564 4404 14596
rect 4436 14564 4440 14596
rect 4240 14560 4440 14564
rect 4480 14596 4680 14600
rect 4480 14564 4484 14596
rect 4516 14564 4644 14596
rect 4676 14564 4680 14596
rect 4480 14560 4680 14564
rect 4720 14596 5720 14600
rect 4720 14564 4724 14596
rect 4756 14564 4884 14596
rect 4916 14564 5044 14596
rect 5076 14564 5204 14596
rect 5236 14564 5364 14596
rect 5396 14564 5524 14596
rect 5556 14564 5684 14596
rect 5716 14564 5720 14596
rect 4720 14560 5720 14564
rect 5760 14596 5960 14600
rect 5760 14564 5764 14596
rect 5796 14564 5924 14596
rect 5956 14564 5960 14596
rect 5760 14560 5960 14564
rect 6000 14596 6200 14600
rect 6000 14564 6004 14596
rect 6036 14564 6164 14596
rect 6196 14564 6200 14596
rect 6000 14560 6200 14564
rect 4240 14516 4440 14520
rect 4240 14484 4244 14516
rect 4276 14484 4404 14516
rect 4436 14484 4440 14516
rect 4240 14480 4440 14484
rect 4480 14516 4680 14520
rect 4480 14484 4484 14516
rect 4516 14484 4644 14516
rect 4676 14484 4680 14516
rect 4480 14480 4680 14484
rect 4720 14516 5720 14520
rect 4720 14484 4724 14516
rect 4756 14484 4884 14516
rect 4916 14484 5044 14516
rect 5076 14484 5204 14516
rect 5236 14484 5364 14516
rect 5396 14484 5524 14516
rect 5556 14484 5684 14516
rect 5716 14484 5720 14516
rect 4720 14480 5720 14484
rect 5760 14516 5960 14520
rect 5760 14484 5764 14516
rect 5796 14484 5924 14516
rect 5956 14484 5960 14516
rect 5760 14480 5960 14484
rect 6000 14516 6200 14520
rect 6000 14484 6004 14516
rect 6036 14484 6164 14516
rect 6196 14484 6200 14516
rect 6000 14480 6200 14484
rect 4240 14436 4440 14440
rect 4240 14404 4244 14436
rect 4276 14404 4404 14436
rect 4436 14404 4440 14436
rect 4240 14400 4440 14404
rect 4480 14436 4680 14440
rect 4480 14404 4484 14436
rect 4516 14404 4644 14436
rect 4676 14404 4680 14436
rect 4480 14400 4680 14404
rect 4720 14436 5720 14440
rect 4720 14404 4724 14436
rect 4756 14404 4884 14436
rect 4916 14404 5044 14436
rect 5076 14404 5204 14436
rect 5236 14404 5364 14436
rect 5396 14404 5524 14436
rect 5556 14404 5684 14436
rect 5716 14404 5720 14436
rect 4720 14400 5720 14404
rect 5760 14436 5960 14440
rect 5760 14404 5764 14436
rect 5796 14404 5924 14436
rect 5956 14404 5960 14436
rect 5760 14400 5960 14404
rect 6000 14436 6200 14440
rect 6000 14404 6004 14436
rect 6036 14404 6164 14436
rect 6196 14404 6200 14436
rect 6000 14400 6200 14404
rect 4240 14356 4440 14360
rect 4240 14324 4244 14356
rect 4276 14324 4404 14356
rect 4436 14324 4440 14356
rect 4240 14320 4440 14324
rect 4480 14356 4680 14360
rect 4480 14324 4484 14356
rect 4516 14324 4644 14356
rect 4676 14324 4680 14356
rect 4480 14320 4680 14324
rect 4720 14356 5720 14360
rect 4720 14324 4724 14356
rect 4756 14324 4884 14356
rect 4916 14324 5044 14356
rect 5076 14324 5204 14356
rect 5236 14324 5364 14356
rect 5396 14324 5524 14356
rect 5556 14324 5684 14356
rect 5716 14324 5720 14356
rect 4720 14320 5720 14324
rect 5760 14356 5960 14360
rect 5760 14324 5764 14356
rect 5796 14324 5924 14356
rect 5956 14324 5960 14356
rect 5760 14320 5960 14324
rect 6000 14356 6200 14360
rect 6000 14324 6004 14356
rect 6036 14324 6164 14356
rect 6196 14324 6200 14356
rect 6000 14320 6200 14324
rect 4240 14276 4440 14280
rect 4240 14244 4244 14276
rect 4276 14244 4404 14276
rect 4436 14244 4440 14276
rect 4240 14240 4440 14244
rect 4480 14276 4680 14280
rect 4480 14244 4484 14276
rect 4516 14244 4644 14276
rect 4676 14244 4680 14276
rect 4480 14240 4680 14244
rect 4720 14276 5720 14280
rect 4720 14244 4724 14276
rect 4756 14244 4884 14276
rect 4916 14244 5044 14276
rect 5076 14244 5204 14276
rect 5236 14244 5364 14276
rect 5396 14244 5524 14276
rect 5556 14244 5684 14276
rect 5716 14244 5720 14276
rect 4720 14240 5720 14244
rect 5760 14276 5960 14280
rect 5760 14244 5764 14276
rect 5796 14244 5924 14276
rect 5956 14244 5960 14276
rect 5760 14240 5960 14244
rect 6000 14276 6200 14280
rect 6000 14244 6004 14276
rect 6036 14244 6164 14276
rect 6196 14244 6200 14276
rect 6000 14240 6200 14244
rect 4240 14196 4440 14200
rect 4240 14164 4244 14196
rect 4276 14164 4404 14196
rect 4436 14164 4440 14196
rect 4240 14160 4440 14164
rect 4480 14196 4680 14200
rect 4480 14164 4484 14196
rect 4516 14164 4644 14196
rect 4676 14164 4680 14196
rect 4480 14160 4680 14164
rect 4720 14196 5720 14200
rect 4720 14164 4724 14196
rect 4756 14164 4884 14196
rect 4916 14164 5044 14196
rect 5076 14164 5204 14196
rect 5236 14164 5364 14196
rect 5396 14164 5524 14196
rect 5556 14164 5684 14196
rect 5716 14164 5720 14196
rect 4720 14160 5720 14164
rect 5760 14196 5960 14200
rect 5760 14164 5764 14196
rect 5796 14164 5924 14196
rect 5956 14164 5960 14196
rect 5760 14160 5960 14164
rect 6000 14196 6200 14200
rect 6000 14164 6004 14196
rect 6036 14164 6164 14196
rect 6196 14164 6200 14196
rect 6000 14160 6200 14164
rect 4240 14116 4440 14120
rect 4240 14084 4244 14116
rect 4276 14084 4404 14116
rect 4436 14084 4440 14116
rect 4240 14080 4440 14084
rect 4480 14116 4680 14120
rect 4480 14084 4484 14116
rect 4516 14084 4644 14116
rect 4676 14084 4680 14116
rect 4480 14080 4680 14084
rect 4720 14116 5720 14120
rect 4720 14084 4724 14116
rect 4756 14084 4884 14116
rect 4916 14084 5044 14116
rect 5076 14084 5204 14116
rect 5236 14084 5364 14116
rect 5396 14084 5524 14116
rect 5556 14084 5684 14116
rect 5716 14084 5720 14116
rect 4720 14080 5720 14084
rect 5760 14116 5960 14120
rect 5760 14084 5764 14116
rect 5796 14084 5924 14116
rect 5956 14084 5960 14116
rect 5760 14080 5960 14084
rect 6000 14116 6200 14120
rect 6000 14084 6004 14116
rect 6036 14084 6164 14116
rect 6196 14084 6200 14116
rect 6000 14080 6200 14084
rect 4240 14036 4440 14040
rect 4240 14004 4244 14036
rect 4276 14004 4404 14036
rect 4436 14004 4440 14036
rect 4240 14000 4440 14004
rect 4480 14036 4680 14040
rect 4480 14004 4484 14036
rect 4516 14004 4644 14036
rect 4676 14004 4680 14036
rect 4480 14000 4680 14004
rect 4720 14036 5720 14040
rect 4720 14004 4724 14036
rect 4756 14004 4884 14036
rect 4916 14004 5044 14036
rect 5076 14004 5204 14036
rect 5236 14004 5364 14036
rect 5396 14004 5524 14036
rect 5556 14004 5684 14036
rect 5716 14004 5720 14036
rect 4720 14000 5720 14004
rect 5760 14036 5960 14040
rect 5760 14004 5764 14036
rect 5796 14004 5924 14036
rect 5956 14004 5960 14036
rect 5760 14000 5960 14004
rect 6000 14036 6200 14040
rect 6000 14004 6004 14036
rect 6036 14004 6164 14036
rect 6196 14004 6200 14036
rect 6000 14000 6200 14004
rect 4240 13956 4440 13960
rect 4240 13924 4244 13956
rect 4276 13924 4404 13956
rect 4436 13924 4440 13956
rect 4240 13920 4440 13924
rect 4480 13956 4680 13960
rect 4480 13924 4484 13956
rect 4516 13924 4644 13956
rect 4676 13924 4680 13956
rect 4480 13920 4680 13924
rect 4720 13956 5720 13960
rect 4720 13924 4724 13956
rect 4756 13924 4884 13956
rect 4916 13924 5044 13956
rect 5076 13924 5204 13956
rect 5236 13924 5364 13956
rect 5396 13924 5524 13956
rect 5556 13924 5684 13956
rect 5716 13924 5720 13956
rect 4720 13920 5720 13924
rect 5760 13956 5960 13960
rect 5760 13924 5764 13956
rect 5796 13924 5924 13956
rect 5956 13924 5960 13956
rect 5760 13920 5960 13924
rect 6000 13956 6200 13960
rect 6000 13924 6004 13956
rect 6036 13924 6164 13956
rect 6196 13924 6200 13956
rect 6000 13920 6200 13924
rect 4240 13876 4440 13880
rect 4240 13844 4244 13876
rect 4276 13844 4404 13876
rect 4436 13844 4440 13876
rect 4240 13840 4440 13844
rect 4480 13876 4680 13880
rect 4480 13844 4484 13876
rect 4516 13844 4644 13876
rect 4676 13844 4680 13876
rect 4480 13840 4680 13844
rect 4720 13876 5720 13880
rect 4720 13844 4724 13876
rect 4756 13844 4884 13876
rect 4916 13844 5044 13876
rect 5076 13844 5204 13876
rect 5236 13844 5364 13876
rect 5396 13844 5524 13876
rect 5556 13844 5684 13876
rect 5716 13844 5720 13876
rect 4720 13840 5720 13844
rect 5760 13876 5960 13880
rect 5760 13844 5764 13876
rect 5796 13844 5924 13876
rect 5956 13844 5960 13876
rect 5760 13840 5960 13844
rect 6000 13876 6200 13880
rect 6000 13844 6004 13876
rect 6036 13844 6164 13876
rect 6196 13844 6200 13876
rect 6000 13840 6200 13844
rect 4240 13796 4440 13800
rect 4240 13764 4244 13796
rect 4276 13764 4404 13796
rect 4436 13764 4440 13796
rect 4240 13760 4440 13764
rect 4480 13796 4680 13800
rect 4480 13764 4484 13796
rect 4516 13764 4644 13796
rect 4676 13764 4680 13796
rect 4480 13760 4680 13764
rect 4720 13796 5720 13800
rect 4720 13764 4724 13796
rect 4756 13764 4884 13796
rect 4916 13764 5044 13796
rect 5076 13764 5204 13796
rect 5236 13764 5364 13796
rect 5396 13764 5524 13796
rect 5556 13764 5684 13796
rect 5716 13764 5720 13796
rect 4720 13760 5720 13764
rect 5760 13796 5960 13800
rect 5760 13764 5764 13796
rect 5796 13764 5924 13796
rect 5956 13764 5960 13796
rect 5760 13760 5960 13764
rect 6000 13796 6200 13800
rect 6000 13764 6004 13796
rect 6036 13764 6164 13796
rect 6196 13764 6200 13796
rect 6000 13760 6200 13764
rect 4240 13716 4440 13720
rect 4240 13684 4244 13716
rect 4276 13684 4404 13716
rect 4436 13684 4440 13716
rect 4240 13680 4440 13684
rect 4480 13716 4680 13720
rect 4480 13684 4484 13716
rect 4516 13684 4644 13716
rect 4676 13684 4680 13716
rect 4480 13680 4680 13684
rect 4720 13716 5720 13720
rect 4720 13684 4724 13716
rect 4756 13684 4884 13716
rect 4916 13684 5044 13716
rect 5076 13684 5204 13716
rect 5236 13684 5364 13716
rect 5396 13684 5524 13716
rect 5556 13684 5684 13716
rect 5716 13684 5720 13716
rect 4720 13680 5720 13684
rect 5760 13716 5960 13720
rect 5760 13684 5764 13716
rect 5796 13684 5924 13716
rect 5956 13684 5960 13716
rect 5760 13680 5960 13684
rect 6000 13716 6200 13720
rect 6000 13684 6004 13716
rect 6036 13684 6164 13716
rect 6196 13684 6200 13716
rect 6000 13680 6200 13684
rect 4240 13636 4440 13640
rect 4240 13604 4244 13636
rect 4276 13604 4404 13636
rect 4436 13604 4440 13636
rect 4240 13600 4440 13604
rect 4480 13636 4680 13640
rect 4480 13604 4484 13636
rect 4516 13604 4644 13636
rect 4676 13604 4680 13636
rect 4480 13600 4680 13604
rect 4720 13636 5720 13640
rect 4720 13604 4724 13636
rect 4756 13604 4884 13636
rect 4916 13604 5044 13636
rect 5076 13604 5204 13636
rect 5236 13604 5364 13636
rect 5396 13604 5524 13636
rect 5556 13604 5684 13636
rect 5716 13604 5720 13636
rect 4720 13600 5720 13604
rect 5760 13636 5960 13640
rect 5760 13604 5764 13636
rect 5796 13604 5924 13636
rect 5956 13604 5960 13636
rect 5760 13600 5960 13604
rect 6000 13636 6200 13640
rect 6000 13604 6004 13636
rect 6036 13604 6164 13636
rect 6196 13604 6200 13636
rect 6000 13600 6200 13604
rect 4240 13556 4440 13560
rect 4240 13524 4244 13556
rect 4276 13524 4404 13556
rect 4436 13524 4440 13556
rect 4240 13520 4440 13524
rect 4480 13556 4680 13560
rect 4480 13524 4484 13556
rect 4516 13524 4644 13556
rect 4676 13524 4680 13556
rect 4480 13520 4680 13524
rect 4720 13556 5720 13560
rect 4720 13524 4724 13556
rect 4756 13524 4884 13556
rect 4916 13524 5044 13556
rect 5076 13524 5204 13556
rect 5236 13524 5364 13556
rect 5396 13524 5524 13556
rect 5556 13524 5684 13556
rect 5716 13524 5720 13556
rect 4720 13520 5720 13524
rect 5760 13556 5960 13560
rect 5760 13524 5764 13556
rect 5796 13524 5924 13556
rect 5956 13524 5960 13556
rect 5760 13520 5960 13524
rect 6000 13556 6200 13560
rect 6000 13524 6004 13556
rect 6036 13524 6164 13556
rect 6196 13524 6200 13556
rect 6000 13520 6200 13524
rect 4240 13476 4440 13480
rect 4240 13444 4244 13476
rect 4276 13444 4404 13476
rect 4436 13444 4440 13476
rect 4240 13440 4440 13444
rect 4480 13476 4680 13480
rect 4480 13444 4484 13476
rect 4516 13444 4644 13476
rect 4676 13444 4680 13476
rect 4480 13440 4680 13444
rect 4720 13476 5720 13480
rect 4720 13444 4724 13476
rect 4756 13444 4884 13476
rect 4916 13444 5044 13476
rect 5076 13444 5204 13476
rect 5236 13444 5364 13476
rect 5396 13444 5524 13476
rect 5556 13444 5684 13476
rect 5716 13444 5720 13476
rect 4720 13440 5720 13444
rect 5760 13476 5960 13480
rect 5760 13444 5764 13476
rect 5796 13444 5924 13476
rect 5956 13444 5960 13476
rect 5760 13440 5960 13444
rect 6000 13476 6200 13480
rect 6000 13444 6004 13476
rect 6036 13444 6164 13476
rect 6196 13444 6200 13476
rect 6000 13440 6200 13444
rect 4240 13396 4440 13400
rect 4240 13364 4244 13396
rect 4276 13364 4404 13396
rect 4436 13364 4440 13396
rect 4240 13360 4440 13364
rect 4480 13396 4680 13400
rect 4480 13364 4484 13396
rect 4516 13364 4644 13396
rect 4676 13364 4680 13396
rect 4480 13360 4680 13364
rect 4720 13396 5720 13400
rect 4720 13364 4724 13396
rect 4756 13364 4884 13396
rect 4916 13364 5044 13396
rect 5076 13364 5204 13396
rect 5236 13364 5364 13396
rect 5396 13364 5524 13396
rect 5556 13364 5684 13396
rect 5716 13364 5720 13396
rect 4720 13360 5720 13364
rect 5760 13396 5960 13400
rect 5760 13364 5764 13396
rect 5796 13364 5924 13396
rect 5956 13364 5960 13396
rect 5760 13360 5960 13364
rect 6000 13396 6200 13400
rect 6000 13364 6004 13396
rect 6036 13364 6164 13396
rect 6196 13364 6200 13396
rect 6000 13360 6200 13364
rect 4240 13316 4440 13320
rect 4240 13284 4244 13316
rect 4276 13284 4404 13316
rect 4436 13284 4440 13316
rect 4240 13280 4440 13284
rect 4480 13316 4680 13320
rect 4480 13284 4484 13316
rect 4516 13284 4644 13316
rect 4676 13284 4680 13316
rect 4480 13280 4680 13284
rect 4720 13316 5720 13320
rect 4720 13284 4724 13316
rect 4756 13284 4884 13316
rect 4916 13284 5044 13316
rect 5076 13284 5204 13316
rect 5236 13284 5364 13316
rect 5396 13284 5524 13316
rect 5556 13284 5684 13316
rect 5716 13284 5720 13316
rect 4720 13280 5720 13284
rect 5760 13316 5960 13320
rect 5760 13284 5764 13316
rect 5796 13284 5924 13316
rect 5956 13284 5960 13316
rect 5760 13280 5960 13284
rect 6000 13316 6200 13320
rect 6000 13284 6004 13316
rect 6036 13284 6164 13316
rect 6196 13284 6200 13316
rect 6000 13280 6200 13284
rect 4240 13236 4440 13240
rect 4240 13204 4244 13236
rect 4276 13204 4404 13236
rect 4436 13204 4440 13236
rect 4240 13200 4440 13204
rect 4480 13236 4680 13240
rect 4480 13204 4484 13236
rect 4516 13204 4644 13236
rect 4676 13204 4680 13236
rect 4480 13200 4680 13204
rect 4720 13236 5720 13240
rect 4720 13204 4724 13236
rect 4756 13204 4884 13236
rect 4916 13204 5044 13236
rect 5076 13204 5204 13236
rect 5236 13204 5364 13236
rect 5396 13204 5524 13236
rect 5556 13204 5684 13236
rect 5716 13204 5720 13236
rect 4720 13200 5720 13204
rect 5760 13236 5960 13240
rect 5760 13204 5764 13236
rect 5796 13204 5924 13236
rect 5956 13204 5960 13236
rect 5760 13200 5960 13204
rect 6000 13236 6200 13240
rect 6000 13204 6004 13236
rect 6036 13204 6164 13236
rect 6196 13204 6200 13236
rect 6000 13200 6200 13204
rect 4240 13156 4440 13160
rect 4240 13124 4244 13156
rect 4276 13124 4404 13156
rect 4436 13124 4440 13156
rect 4240 13120 4440 13124
rect 4480 13156 4680 13160
rect 4480 13124 4484 13156
rect 4516 13124 4644 13156
rect 4676 13124 4680 13156
rect 4480 13120 4680 13124
rect 4720 13156 5720 13160
rect 4720 13124 4724 13156
rect 4756 13124 4884 13156
rect 4916 13124 5044 13156
rect 5076 13124 5204 13156
rect 5236 13124 5364 13156
rect 5396 13124 5524 13156
rect 5556 13124 5684 13156
rect 5716 13124 5720 13156
rect 4720 13120 5720 13124
rect 5760 13156 5960 13160
rect 5760 13124 5764 13156
rect 5796 13124 5924 13156
rect 5956 13124 5960 13156
rect 5760 13120 5960 13124
rect 6000 13156 6200 13160
rect 6000 13124 6004 13156
rect 6036 13124 6164 13156
rect 6196 13124 6200 13156
rect 6000 13120 6200 13124
rect 4240 13076 4440 13080
rect 4240 13044 4244 13076
rect 4276 13044 4404 13076
rect 4436 13044 4440 13076
rect 4240 13040 4440 13044
rect 4480 13076 4680 13080
rect 4480 13044 4484 13076
rect 4516 13044 4644 13076
rect 4676 13044 4680 13076
rect 4480 13040 4680 13044
rect 4720 13076 5720 13080
rect 4720 13044 4724 13076
rect 4756 13044 4884 13076
rect 4916 13044 5044 13076
rect 5076 13044 5204 13076
rect 5236 13044 5364 13076
rect 5396 13044 5524 13076
rect 5556 13044 5684 13076
rect 5716 13044 5720 13076
rect 4720 13040 5720 13044
rect 5760 13076 5960 13080
rect 5760 13044 5764 13076
rect 5796 13044 5924 13076
rect 5956 13044 5960 13076
rect 5760 13040 5960 13044
rect 6000 13076 6200 13080
rect 6000 13044 6004 13076
rect 6036 13044 6164 13076
rect 6196 13044 6200 13076
rect 6000 13040 6200 13044
rect 4240 12996 4440 13000
rect 4240 12964 4244 12996
rect 4276 12964 4404 12996
rect 4436 12964 4440 12996
rect 4240 12960 4440 12964
rect 4480 12996 4680 13000
rect 4480 12964 4484 12996
rect 4516 12964 4644 12996
rect 4676 12964 4680 12996
rect 4480 12960 4680 12964
rect 4720 12996 5720 13000
rect 4720 12964 4724 12996
rect 4756 12964 4884 12996
rect 4916 12964 5044 12996
rect 5076 12964 5204 12996
rect 5236 12964 5364 12996
rect 5396 12964 5524 12996
rect 5556 12964 5684 12996
rect 5716 12964 5720 12996
rect 4720 12960 5720 12964
rect 5760 12996 5960 13000
rect 5760 12964 5764 12996
rect 5796 12964 5924 12996
rect 5956 12964 5960 12996
rect 5760 12960 5960 12964
rect 6000 12996 6200 13000
rect 6000 12964 6004 12996
rect 6036 12964 6164 12996
rect 6196 12964 6200 12996
rect 6000 12960 6200 12964
rect 4240 12916 4440 12920
rect 4240 12884 4244 12916
rect 4276 12884 4404 12916
rect 4436 12884 4440 12916
rect 4240 12880 4440 12884
rect 4480 12916 4680 12920
rect 4480 12884 4484 12916
rect 4516 12884 4644 12916
rect 4676 12884 4680 12916
rect 4480 12880 4680 12884
rect 4720 12916 5720 12920
rect 4720 12884 4724 12916
rect 4756 12884 4884 12916
rect 4916 12884 5044 12916
rect 5076 12884 5204 12916
rect 5236 12884 5364 12916
rect 5396 12884 5524 12916
rect 5556 12884 5684 12916
rect 5716 12884 5720 12916
rect 4720 12880 5720 12884
rect 5760 12916 5960 12920
rect 5760 12884 5764 12916
rect 5796 12884 5924 12916
rect 5956 12884 5960 12916
rect 5760 12880 5960 12884
rect 6000 12916 6200 12920
rect 6000 12884 6004 12916
rect 6036 12884 6164 12916
rect 6196 12884 6200 12916
rect 6000 12880 6200 12884
rect 4240 12836 4440 12840
rect 4240 12804 4244 12836
rect 4276 12804 4404 12836
rect 4436 12804 4440 12836
rect 4240 12800 4440 12804
rect 4480 12836 4680 12840
rect 4480 12804 4484 12836
rect 4516 12804 4644 12836
rect 4676 12804 4680 12836
rect 4480 12800 4680 12804
rect 4720 12836 5720 12840
rect 4720 12804 4724 12836
rect 4756 12804 4884 12836
rect 4916 12804 5044 12836
rect 5076 12804 5204 12836
rect 5236 12804 5364 12836
rect 5396 12804 5524 12836
rect 5556 12804 5684 12836
rect 5716 12804 5720 12836
rect 4720 12800 5720 12804
rect 5760 12836 5960 12840
rect 5760 12804 5764 12836
rect 5796 12804 5924 12836
rect 5956 12804 5960 12836
rect 5760 12800 5960 12804
rect 6000 12836 6200 12840
rect 6000 12804 6004 12836
rect 6036 12804 6164 12836
rect 6196 12804 6200 12836
rect 6000 12800 6200 12804
rect 4240 12756 4440 12760
rect 4240 12724 4244 12756
rect 4276 12724 4404 12756
rect 4436 12724 4440 12756
rect 4240 12720 4440 12724
rect 4480 12756 4680 12760
rect 4480 12724 4484 12756
rect 4516 12724 4644 12756
rect 4676 12724 4680 12756
rect 4480 12720 4680 12724
rect 4720 12756 5720 12760
rect 4720 12724 4724 12756
rect 4756 12724 4884 12756
rect 4916 12724 5044 12756
rect 5076 12724 5204 12756
rect 5236 12724 5364 12756
rect 5396 12724 5524 12756
rect 5556 12724 5684 12756
rect 5716 12724 5720 12756
rect 4720 12720 5720 12724
rect 5760 12756 5960 12760
rect 5760 12724 5764 12756
rect 5796 12724 5924 12756
rect 5956 12724 5960 12756
rect 5760 12720 5960 12724
rect 6000 12756 6200 12760
rect 6000 12724 6004 12756
rect 6036 12724 6164 12756
rect 6196 12724 6200 12756
rect 6000 12720 6200 12724
rect 4240 12676 4440 12680
rect 4240 12644 4244 12676
rect 4276 12644 4404 12676
rect 4436 12644 4440 12676
rect 4240 12640 4440 12644
rect 4480 12676 4680 12680
rect 4480 12644 4484 12676
rect 4516 12644 4644 12676
rect 4676 12644 4680 12676
rect 4480 12640 4680 12644
rect 4720 12676 5720 12680
rect 4720 12644 4724 12676
rect 4756 12644 4884 12676
rect 4916 12644 5044 12676
rect 5076 12644 5204 12676
rect 5236 12644 5364 12676
rect 5396 12644 5524 12676
rect 5556 12644 5684 12676
rect 5716 12644 5720 12676
rect 4720 12640 5720 12644
rect 5760 12676 5960 12680
rect 5760 12644 5764 12676
rect 5796 12644 5924 12676
rect 5956 12644 5960 12676
rect 5760 12640 5960 12644
rect 6000 12676 6200 12680
rect 6000 12644 6004 12676
rect 6036 12644 6164 12676
rect 6196 12644 6200 12676
rect 6000 12640 6200 12644
rect 4240 12596 4440 12600
rect 4240 12564 4244 12596
rect 4276 12564 4404 12596
rect 4436 12564 4440 12596
rect 4240 12560 4440 12564
rect 4480 12596 4680 12600
rect 4480 12564 4484 12596
rect 4516 12564 4644 12596
rect 4676 12564 4680 12596
rect 4480 12560 4680 12564
rect 4720 12596 5720 12600
rect 4720 12564 4724 12596
rect 4756 12564 4884 12596
rect 4916 12564 5044 12596
rect 5076 12564 5204 12596
rect 5236 12564 5364 12596
rect 5396 12564 5524 12596
rect 5556 12564 5684 12596
rect 5716 12564 5720 12596
rect 4720 12560 5720 12564
rect 5760 12596 5960 12600
rect 5760 12564 5764 12596
rect 5796 12564 5924 12596
rect 5956 12564 5960 12596
rect 5760 12560 5960 12564
rect 6000 12596 6200 12600
rect 6000 12564 6004 12596
rect 6036 12564 6164 12596
rect 6196 12564 6200 12596
rect 6000 12560 6200 12564
rect 4240 12516 4440 12520
rect 4240 12484 4244 12516
rect 4276 12484 4404 12516
rect 4436 12484 4440 12516
rect 4240 12480 4440 12484
rect 4480 12516 4680 12520
rect 4480 12484 4484 12516
rect 4516 12484 4644 12516
rect 4676 12484 4680 12516
rect 4480 12480 4680 12484
rect 4720 12516 5720 12520
rect 4720 12484 4724 12516
rect 4756 12484 4884 12516
rect 4916 12484 5044 12516
rect 5076 12484 5204 12516
rect 5236 12484 5364 12516
rect 5396 12484 5524 12516
rect 5556 12484 5684 12516
rect 5716 12484 5720 12516
rect 4720 12480 5720 12484
rect 5760 12516 5960 12520
rect 5760 12484 5764 12516
rect 5796 12484 5924 12516
rect 5956 12484 5960 12516
rect 5760 12480 5960 12484
rect 6000 12516 6200 12520
rect 6000 12484 6004 12516
rect 6036 12484 6164 12516
rect 6196 12484 6200 12516
rect 6000 12480 6200 12484
rect 4240 12436 4440 12440
rect 4240 12404 4244 12436
rect 4276 12404 4404 12436
rect 4436 12404 4440 12436
rect 4240 12400 4440 12404
rect 4480 12436 4680 12440
rect 4480 12404 4484 12436
rect 4516 12404 4644 12436
rect 4676 12404 4680 12436
rect 4480 12400 4680 12404
rect 4720 12436 5720 12440
rect 4720 12404 4724 12436
rect 4756 12404 4884 12436
rect 4916 12404 5044 12436
rect 5076 12404 5204 12436
rect 5236 12404 5364 12436
rect 5396 12404 5524 12436
rect 5556 12404 5684 12436
rect 5716 12404 5720 12436
rect 4720 12400 5720 12404
rect 5760 12436 5960 12440
rect 5760 12404 5764 12436
rect 5796 12404 5924 12436
rect 5956 12404 5960 12436
rect 5760 12400 5960 12404
rect 6000 12436 6200 12440
rect 6000 12404 6004 12436
rect 6036 12404 6164 12436
rect 6196 12404 6200 12436
rect 6000 12400 6200 12404
rect 4240 12356 4440 12360
rect 4240 12324 4244 12356
rect 4276 12324 4404 12356
rect 4436 12324 4440 12356
rect 4240 12320 4440 12324
rect 4480 12356 4680 12360
rect 4480 12324 4484 12356
rect 4516 12324 4644 12356
rect 4676 12324 4680 12356
rect 4480 12320 4680 12324
rect 4720 12356 5720 12360
rect 4720 12324 4724 12356
rect 4756 12324 4884 12356
rect 4916 12324 5044 12356
rect 5076 12324 5204 12356
rect 5236 12324 5364 12356
rect 5396 12324 5524 12356
rect 5556 12324 5684 12356
rect 5716 12324 5720 12356
rect 4720 12320 5720 12324
rect 5760 12356 5960 12360
rect 5760 12324 5764 12356
rect 5796 12324 5924 12356
rect 5956 12324 5960 12356
rect 5760 12320 5960 12324
rect 6000 12356 6200 12360
rect 6000 12324 6004 12356
rect 6036 12324 6164 12356
rect 6196 12324 6200 12356
rect 6000 12320 6200 12324
rect 4240 12276 4440 12280
rect 4240 12244 4244 12276
rect 4276 12244 4404 12276
rect 4436 12244 4440 12276
rect 4240 12240 4440 12244
rect 4480 12276 4680 12280
rect 4480 12244 4484 12276
rect 4516 12244 4644 12276
rect 4676 12244 4680 12276
rect 4480 12240 4680 12244
rect 4720 12276 5720 12280
rect 4720 12244 4724 12276
rect 4756 12244 4884 12276
rect 4916 12244 5044 12276
rect 5076 12244 5204 12276
rect 5236 12244 5364 12276
rect 5396 12244 5524 12276
rect 5556 12244 5684 12276
rect 5716 12244 5720 12276
rect 4720 12240 5720 12244
rect 5760 12276 5960 12280
rect 5760 12244 5764 12276
rect 5796 12244 5924 12276
rect 5956 12244 5960 12276
rect 5760 12240 5960 12244
rect 6000 12276 6200 12280
rect 6000 12244 6004 12276
rect 6036 12244 6164 12276
rect 6196 12244 6200 12276
rect 6000 12240 6200 12244
rect 4240 12196 4440 12200
rect 4240 12164 4244 12196
rect 4276 12164 4404 12196
rect 4436 12164 4440 12196
rect 4240 12160 4440 12164
rect 4480 12196 4680 12200
rect 4480 12164 4484 12196
rect 4516 12164 4644 12196
rect 4676 12164 4680 12196
rect 4480 12160 4680 12164
rect 4720 12196 5720 12200
rect 4720 12164 4724 12196
rect 4756 12164 4884 12196
rect 4916 12164 5044 12196
rect 5076 12164 5204 12196
rect 5236 12164 5364 12196
rect 5396 12164 5524 12196
rect 5556 12164 5684 12196
rect 5716 12164 5720 12196
rect 4720 12160 5720 12164
rect 5760 12196 5960 12200
rect 5760 12164 5764 12196
rect 5796 12164 5924 12196
rect 5956 12164 5960 12196
rect 5760 12160 5960 12164
rect 6000 12196 6200 12200
rect 6000 12164 6004 12196
rect 6036 12164 6164 12196
rect 6196 12164 6200 12196
rect 6000 12160 6200 12164
rect 4240 12116 4440 12120
rect 4240 12084 4244 12116
rect 4276 12084 4404 12116
rect 4436 12084 4440 12116
rect 4240 12080 4440 12084
rect 4480 12116 4680 12120
rect 4480 12084 4484 12116
rect 4516 12084 4644 12116
rect 4676 12084 4680 12116
rect 4480 12080 4680 12084
rect 4720 12116 5720 12120
rect 4720 12084 4724 12116
rect 4756 12084 4884 12116
rect 4916 12084 5044 12116
rect 5076 12084 5204 12116
rect 5236 12084 5364 12116
rect 5396 12084 5524 12116
rect 5556 12084 5684 12116
rect 5716 12084 5720 12116
rect 4720 12080 5720 12084
rect 5760 12116 5960 12120
rect 5760 12084 5764 12116
rect 5796 12084 5924 12116
rect 5956 12084 5960 12116
rect 5760 12080 5960 12084
rect 6000 12116 6200 12120
rect 6000 12084 6004 12116
rect 6036 12084 6164 12116
rect 6196 12084 6200 12116
rect 6000 12080 6200 12084
rect 4240 12036 4440 12040
rect 4240 12004 4244 12036
rect 4276 12004 4404 12036
rect 4436 12004 4440 12036
rect 4240 12000 4440 12004
rect 4480 12036 4680 12040
rect 4480 12004 4484 12036
rect 4516 12004 4644 12036
rect 4676 12004 4680 12036
rect 4480 12000 4680 12004
rect 4720 12036 5720 12040
rect 4720 12004 4724 12036
rect 4756 12004 4884 12036
rect 4916 12004 5044 12036
rect 5076 12004 5204 12036
rect 5236 12004 5364 12036
rect 5396 12004 5524 12036
rect 5556 12004 5684 12036
rect 5716 12004 5720 12036
rect 4720 12000 5720 12004
rect 5760 12036 5960 12040
rect 5760 12004 5764 12036
rect 5796 12004 5924 12036
rect 5956 12004 5960 12036
rect 5760 12000 5960 12004
rect 6000 12036 6200 12040
rect 6000 12004 6004 12036
rect 6036 12004 6164 12036
rect 6196 12004 6200 12036
rect 6000 12000 6200 12004
rect 4240 11956 4440 11960
rect 4240 11924 4244 11956
rect 4276 11924 4404 11956
rect 4436 11924 4440 11956
rect 4240 11920 4440 11924
rect 4480 11956 4680 11960
rect 4480 11924 4484 11956
rect 4516 11924 4644 11956
rect 4676 11924 4680 11956
rect 4480 11920 4680 11924
rect 4720 11956 5720 11960
rect 4720 11924 4724 11956
rect 4756 11924 4884 11956
rect 4916 11924 5044 11956
rect 5076 11924 5204 11956
rect 5236 11924 5364 11956
rect 5396 11924 5524 11956
rect 5556 11924 5684 11956
rect 5716 11924 5720 11956
rect 4720 11920 5720 11924
rect 5760 11956 5960 11960
rect 5760 11924 5764 11956
rect 5796 11924 5924 11956
rect 5956 11924 5960 11956
rect 5760 11920 5960 11924
rect 6000 11956 6200 11960
rect 6000 11924 6004 11956
rect 6036 11924 6164 11956
rect 6196 11924 6200 11956
rect 6000 11920 6200 11924
rect 4240 11876 4440 11880
rect 4240 11844 4244 11876
rect 4276 11844 4404 11876
rect 4436 11844 4440 11876
rect 4240 11840 4440 11844
rect 4480 11876 4680 11880
rect 4480 11844 4484 11876
rect 4516 11844 4644 11876
rect 4676 11844 4680 11876
rect 4480 11840 4680 11844
rect 4720 11876 5720 11880
rect 4720 11844 4724 11876
rect 4756 11844 4884 11876
rect 4916 11844 5044 11876
rect 5076 11844 5204 11876
rect 5236 11844 5364 11876
rect 5396 11844 5524 11876
rect 5556 11844 5684 11876
rect 5716 11844 5720 11876
rect 4720 11840 5720 11844
rect 5760 11876 5960 11880
rect 5760 11844 5764 11876
rect 5796 11844 5924 11876
rect 5956 11844 5960 11876
rect 5760 11840 5960 11844
rect 6000 11876 6200 11880
rect 6000 11844 6004 11876
rect 6036 11844 6164 11876
rect 6196 11844 6200 11876
rect 6000 11840 6200 11844
rect 4240 11796 4440 11800
rect 4240 11764 4244 11796
rect 4276 11764 4404 11796
rect 4436 11764 4440 11796
rect 4240 11760 4440 11764
rect 4480 11796 4680 11800
rect 4480 11764 4484 11796
rect 4516 11764 4644 11796
rect 4676 11764 4680 11796
rect 4480 11760 4680 11764
rect 4720 11796 5720 11800
rect 4720 11764 4724 11796
rect 4756 11764 4884 11796
rect 4916 11764 5044 11796
rect 5076 11764 5204 11796
rect 5236 11764 5364 11796
rect 5396 11764 5524 11796
rect 5556 11764 5684 11796
rect 5716 11764 5720 11796
rect 4720 11760 5720 11764
rect 5760 11796 5960 11800
rect 5760 11764 5764 11796
rect 5796 11764 5924 11796
rect 5956 11764 5960 11796
rect 5760 11760 5960 11764
rect 6000 11796 6200 11800
rect 6000 11764 6004 11796
rect 6036 11764 6164 11796
rect 6196 11764 6200 11796
rect 6000 11760 6200 11764
rect 4240 11716 4440 11720
rect 4240 11684 4244 11716
rect 4276 11684 4404 11716
rect 4436 11684 4440 11716
rect 4240 11680 4440 11684
rect 4480 11716 4680 11720
rect 4480 11684 4484 11716
rect 4516 11684 4644 11716
rect 4676 11684 4680 11716
rect 4480 11680 4680 11684
rect 4720 11716 5720 11720
rect 4720 11684 4724 11716
rect 4756 11684 4884 11716
rect 4916 11684 5044 11716
rect 5076 11684 5204 11716
rect 5236 11684 5364 11716
rect 5396 11684 5524 11716
rect 5556 11684 5684 11716
rect 5716 11684 5720 11716
rect 4720 11680 5720 11684
rect 5760 11716 5960 11720
rect 5760 11684 5764 11716
rect 5796 11684 5924 11716
rect 5956 11684 5960 11716
rect 5760 11680 5960 11684
rect 6000 11716 6200 11720
rect 6000 11684 6004 11716
rect 6036 11684 6164 11716
rect 6196 11684 6200 11716
rect 6000 11680 6200 11684
rect 4240 11636 4440 11640
rect 4240 11604 4244 11636
rect 4276 11604 4404 11636
rect 4436 11604 4440 11636
rect 4240 11600 4440 11604
rect 4480 11636 4680 11640
rect 4480 11604 4484 11636
rect 4516 11604 4644 11636
rect 4676 11604 4680 11636
rect 4480 11600 4680 11604
rect 4720 11636 5720 11640
rect 4720 11604 4724 11636
rect 4756 11604 4884 11636
rect 4916 11604 5044 11636
rect 5076 11604 5204 11636
rect 5236 11604 5364 11636
rect 5396 11604 5524 11636
rect 5556 11604 5684 11636
rect 5716 11604 5720 11636
rect 4720 11600 5720 11604
rect 5760 11636 5960 11640
rect 5760 11604 5764 11636
rect 5796 11604 5924 11636
rect 5956 11604 5960 11636
rect 5760 11600 5960 11604
rect 6000 11636 6200 11640
rect 6000 11604 6004 11636
rect 6036 11604 6164 11636
rect 6196 11604 6200 11636
rect 6000 11600 6200 11604
rect 4240 11556 4440 11560
rect 4240 11524 4244 11556
rect 4276 11524 4404 11556
rect 4436 11524 4440 11556
rect 4240 11520 4440 11524
rect 4480 11556 4680 11560
rect 4480 11524 4484 11556
rect 4516 11524 4644 11556
rect 4676 11524 4680 11556
rect 4480 11520 4680 11524
rect 4720 11556 5720 11560
rect 4720 11524 4724 11556
rect 4756 11524 4884 11556
rect 4916 11524 5044 11556
rect 5076 11524 5204 11556
rect 5236 11524 5364 11556
rect 5396 11524 5524 11556
rect 5556 11524 5684 11556
rect 5716 11524 5720 11556
rect 4720 11520 5720 11524
rect 5760 11556 5960 11560
rect 5760 11524 5764 11556
rect 5796 11524 5924 11556
rect 5956 11524 5960 11556
rect 5760 11520 5960 11524
rect 6000 11556 6200 11560
rect 6000 11524 6004 11556
rect 6036 11524 6164 11556
rect 6196 11524 6200 11556
rect 6000 11520 6200 11524
rect 4240 11476 4440 11480
rect 4240 11444 4244 11476
rect 4276 11444 4404 11476
rect 4436 11444 4440 11476
rect 4240 11440 4440 11444
rect 4480 11476 4680 11480
rect 4480 11444 4484 11476
rect 4516 11444 4644 11476
rect 4676 11444 4680 11476
rect 4480 11440 4680 11444
rect 4720 11476 5720 11480
rect 4720 11444 4724 11476
rect 4756 11444 4884 11476
rect 4916 11444 5044 11476
rect 5076 11444 5204 11476
rect 5236 11444 5364 11476
rect 5396 11444 5524 11476
rect 5556 11444 5684 11476
rect 5716 11444 5720 11476
rect 4720 11440 5720 11444
rect 5760 11476 5960 11480
rect 5760 11444 5764 11476
rect 5796 11444 5924 11476
rect 5956 11444 5960 11476
rect 5760 11440 5960 11444
rect 6000 11476 6200 11480
rect 6000 11444 6004 11476
rect 6036 11444 6164 11476
rect 6196 11444 6200 11476
rect 6000 11440 6200 11444
rect 4240 11396 4440 11400
rect 4240 11364 4244 11396
rect 4276 11364 4404 11396
rect 4436 11364 4440 11396
rect 4240 11360 4440 11364
rect 4480 11396 4680 11400
rect 4480 11364 4484 11396
rect 4516 11364 4644 11396
rect 4676 11364 4680 11396
rect 4480 11360 4680 11364
rect 4720 11396 5720 11400
rect 4720 11364 4724 11396
rect 4756 11364 4884 11396
rect 4916 11364 5044 11396
rect 5076 11364 5204 11396
rect 5236 11364 5364 11396
rect 5396 11364 5524 11396
rect 5556 11364 5684 11396
rect 5716 11364 5720 11396
rect 4720 11360 5720 11364
rect 5760 11396 5960 11400
rect 5760 11364 5764 11396
rect 5796 11364 5924 11396
rect 5956 11364 5960 11396
rect 5760 11360 5960 11364
rect 6000 11396 6200 11400
rect 6000 11364 6004 11396
rect 6036 11364 6164 11396
rect 6196 11364 6200 11396
rect 6000 11360 6200 11364
rect 4240 11316 4440 11320
rect 4240 11284 4244 11316
rect 4276 11284 4404 11316
rect 4436 11284 4440 11316
rect 4240 11280 4440 11284
rect 4480 11316 4680 11320
rect 4480 11284 4484 11316
rect 4516 11284 4644 11316
rect 4676 11284 4680 11316
rect 4480 11280 4680 11284
rect 4720 11316 5720 11320
rect 4720 11284 4724 11316
rect 4756 11284 4884 11316
rect 4916 11284 5044 11316
rect 5076 11284 5204 11316
rect 5236 11284 5364 11316
rect 5396 11284 5524 11316
rect 5556 11284 5684 11316
rect 5716 11284 5720 11316
rect 4720 11280 5720 11284
rect 5760 11316 5960 11320
rect 5760 11284 5764 11316
rect 5796 11284 5924 11316
rect 5956 11284 5960 11316
rect 5760 11280 5960 11284
rect 6000 11316 6200 11320
rect 6000 11284 6004 11316
rect 6036 11284 6164 11316
rect 6196 11284 6200 11316
rect 6000 11280 6200 11284
rect 4240 11236 4440 11240
rect 4240 11204 4244 11236
rect 4276 11204 4404 11236
rect 4436 11204 4440 11236
rect 4240 11200 4440 11204
rect 4480 11236 4680 11240
rect 4480 11204 4484 11236
rect 4516 11204 4644 11236
rect 4676 11204 4680 11236
rect 4480 11200 4680 11204
rect 4720 11236 5720 11240
rect 4720 11204 4724 11236
rect 4756 11204 4884 11236
rect 4916 11204 5044 11236
rect 5076 11204 5204 11236
rect 5236 11204 5364 11236
rect 5396 11204 5524 11236
rect 5556 11204 5684 11236
rect 5716 11204 5720 11236
rect 4720 11200 5720 11204
rect 5760 11236 5960 11240
rect 5760 11204 5764 11236
rect 5796 11204 5924 11236
rect 5956 11204 5960 11236
rect 5760 11200 5960 11204
rect 6000 11236 6200 11240
rect 6000 11204 6004 11236
rect 6036 11204 6164 11236
rect 6196 11204 6200 11236
rect 6000 11200 6200 11204
rect 4240 11156 4440 11160
rect 4240 11124 4244 11156
rect 4276 11124 4404 11156
rect 4436 11124 4440 11156
rect 4240 11120 4440 11124
rect 4480 11156 4680 11160
rect 4480 11124 4484 11156
rect 4516 11124 4644 11156
rect 4676 11124 4680 11156
rect 4480 11120 4680 11124
rect 4720 11156 5720 11160
rect 4720 11124 4724 11156
rect 4756 11124 4884 11156
rect 4916 11124 5044 11156
rect 5076 11124 5204 11156
rect 5236 11124 5364 11156
rect 5396 11124 5524 11156
rect 5556 11124 5684 11156
rect 5716 11124 5720 11156
rect 4720 11120 5720 11124
rect 5760 11156 5960 11160
rect 5760 11124 5764 11156
rect 5796 11124 5924 11156
rect 5956 11124 5960 11156
rect 5760 11120 5960 11124
rect 6000 11156 6200 11160
rect 6000 11124 6004 11156
rect 6036 11124 6164 11156
rect 6196 11124 6200 11156
rect 6000 11120 6200 11124
rect 4240 11076 4440 11080
rect 4240 11044 4244 11076
rect 4276 11044 4404 11076
rect 4436 11044 4440 11076
rect 4240 11040 4440 11044
rect 4480 11076 4680 11080
rect 4480 11044 4484 11076
rect 4516 11044 4644 11076
rect 4676 11044 4680 11076
rect 4480 11040 4680 11044
rect 4720 11076 5720 11080
rect 4720 11044 4724 11076
rect 4756 11044 4884 11076
rect 4916 11044 5044 11076
rect 5076 11044 5204 11076
rect 5236 11044 5364 11076
rect 5396 11044 5524 11076
rect 5556 11044 5684 11076
rect 5716 11044 5720 11076
rect 4720 11040 5720 11044
rect 5760 11076 5960 11080
rect 5760 11044 5764 11076
rect 5796 11044 5924 11076
rect 5956 11044 5960 11076
rect 5760 11040 5960 11044
rect 6000 11076 6200 11080
rect 6000 11044 6004 11076
rect 6036 11044 6164 11076
rect 6196 11044 6200 11076
rect 6000 11040 6200 11044
rect 4240 10996 4440 11000
rect 4240 10964 4244 10996
rect 4276 10964 4404 10996
rect 4436 10964 4440 10996
rect 4240 10960 4440 10964
rect 4480 10996 4680 11000
rect 4480 10964 4484 10996
rect 4516 10964 4644 10996
rect 4676 10964 4680 10996
rect 4480 10960 4680 10964
rect 4720 10996 5720 11000
rect 4720 10964 4724 10996
rect 4756 10964 4884 10996
rect 4916 10964 5044 10996
rect 5076 10964 5204 10996
rect 5236 10964 5364 10996
rect 5396 10964 5524 10996
rect 5556 10964 5684 10996
rect 5716 10964 5720 10996
rect 4720 10960 5720 10964
rect 5760 10996 5960 11000
rect 5760 10964 5764 10996
rect 5796 10964 5924 10996
rect 5956 10964 5960 10996
rect 5760 10960 5960 10964
rect 6000 10996 6200 11000
rect 6000 10964 6004 10996
rect 6036 10964 6164 10996
rect 6196 10964 6200 10996
rect 6000 10960 6200 10964
rect 4240 10916 4440 10920
rect 4240 10884 4244 10916
rect 4276 10884 4404 10916
rect 4436 10884 4440 10916
rect 4240 10880 4440 10884
rect 4480 10916 4680 10920
rect 4480 10884 4484 10916
rect 4516 10884 4644 10916
rect 4676 10884 4680 10916
rect 4480 10880 4680 10884
rect 4720 10916 5720 10920
rect 4720 10884 4724 10916
rect 4756 10884 4884 10916
rect 4916 10884 5044 10916
rect 5076 10884 5204 10916
rect 5236 10884 5364 10916
rect 5396 10884 5524 10916
rect 5556 10884 5684 10916
rect 5716 10884 5720 10916
rect 4720 10880 5720 10884
rect 5760 10916 5960 10920
rect 5760 10884 5764 10916
rect 5796 10884 5924 10916
rect 5956 10884 5960 10916
rect 5760 10880 5960 10884
rect 6000 10916 6200 10920
rect 6000 10884 6004 10916
rect 6036 10884 6164 10916
rect 6196 10884 6200 10916
rect 6000 10880 6200 10884
rect 4240 10836 4440 10840
rect 4240 10804 4244 10836
rect 4276 10804 4404 10836
rect 4436 10804 4440 10836
rect 4240 10800 4440 10804
rect 4480 10836 4680 10840
rect 4480 10804 4484 10836
rect 4516 10804 4644 10836
rect 4676 10804 4680 10836
rect 4480 10800 4680 10804
rect 4720 10836 5720 10840
rect 4720 10804 4724 10836
rect 4756 10804 4884 10836
rect 4916 10804 5044 10836
rect 5076 10804 5204 10836
rect 5236 10804 5364 10836
rect 5396 10804 5524 10836
rect 5556 10804 5684 10836
rect 5716 10804 5720 10836
rect 4720 10800 5720 10804
rect 5760 10836 5960 10840
rect 5760 10804 5764 10836
rect 5796 10804 5924 10836
rect 5956 10804 5960 10836
rect 5760 10800 5960 10804
rect 6000 10836 6200 10840
rect 6000 10804 6004 10836
rect 6036 10804 6164 10836
rect 6196 10804 6200 10836
rect 6000 10800 6200 10804
rect 4240 10756 4440 10760
rect 4240 10724 4244 10756
rect 4276 10724 4404 10756
rect 4436 10724 4440 10756
rect 4240 10720 4440 10724
rect 4480 10756 4680 10760
rect 4480 10724 4484 10756
rect 4516 10724 4644 10756
rect 4676 10724 4680 10756
rect 4480 10720 4680 10724
rect 4720 10756 5720 10760
rect 4720 10724 4724 10756
rect 4756 10724 4884 10756
rect 4916 10724 5044 10756
rect 5076 10724 5204 10756
rect 5236 10724 5364 10756
rect 5396 10724 5524 10756
rect 5556 10724 5684 10756
rect 5716 10724 5720 10756
rect 4720 10720 5720 10724
rect 5760 10756 5960 10760
rect 5760 10724 5764 10756
rect 5796 10724 5924 10756
rect 5956 10724 5960 10756
rect 5760 10720 5960 10724
rect 6000 10756 6200 10760
rect 6000 10724 6004 10756
rect 6036 10724 6164 10756
rect 6196 10724 6200 10756
rect 6000 10720 6200 10724
rect 4240 10676 4440 10680
rect 4240 10644 4244 10676
rect 4276 10644 4404 10676
rect 4436 10644 4440 10676
rect 4240 10640 4440 10644
rect 4480 10676 4680 10680
rect 4480 10644 4484 10676
rect 4516 10644 4644 10676
rect 4676 10644 4680 10676
rect 4480 10640 4680 10644
rect 4720 10676 5720 10680
rect 4720 10644 4724 10676
rect 4756 10644 4884 10676
rect 4916 10644 5044 10676
rect 5076 10644 5204 10676
rect 5236 10644 5364 10676
rect 5396 10644 5524 10676
rect 5556 10644 5684 10676
rect 5716 10644 5720 10676
rect 4720 10640 5720 10644
rect 5760 10676 5960 10680
rect 5760 10644 5764 10676
rect 5796 10644 5924 10676
rect 5956 10644 5960 10676
rect 5760 10640 5960 10644
rect 6000 10676 6200 10680
rect 6000 10644 6004 10676
rect 6036 10644 6164 10676
rect 6196 10644 6200 10676
rect 6000 10640 6200 10644
rect 4240 10596 4440 10600
rect 4240 10564 4244 10596
rect 4276 10564 4404 10596
rect 4436 10564 4440 10596
rect 4240 10560 4440 10564
rect 4480 10596 4680 10600
rect 4480 10564 4484 10596
rect 4516 10564 4644 10596
rect 4676 10564 4680 10596
rect 4480 10560 4680 10564
rect 4720 10596 5720 10600
rect 4720 10564 4724 10596
rect 4756 10564 4884 10596
rect 4916 10564 5044 10596
rect 5076 10564 5204 10596
rect 5236 10564 5364 10596
rect 5396 10564 5524 10596
rect 5556 10564 5684 10596
rect 5716 10564 5720 10596
rect 4720 10560 5720 10564
rect 5760 10596 5960 10600
rect 5760 10564 5764 10596
rect 5796 10564 5924 10596
rect 5956 10564 5960 10596
rect 5760 10560 5960 10564
rect 6000 10596 6200 10600
rect 6000 10564 6004 10596
rect 6036 10564 6164 10596
rect 6196 10564 6200 10596
rect 6000 10560 6200 10564
rect 4240 10516 4440 10520
rect 4240 10484 4244 10516
rect 4276 10484 4404 10516
rect 4436 10484 4440 10516
rect 4240 10480 4440 10484
rect 4480 10516 4680 10520
rect 4480 10484 4484 10516
rect 4516 10484 4644 10516
rect 4676 10484 4680 10516
rect 4480 10480 4680 10484
rect 4720 10516 5720 10520
rect 4720 10484 4724 10516
rect 4756 10484 4884 10516
rect 4916 10484 5044 10516
rect 5076 10484 5204 10516
rect 5236 10484 5364 10516
rect 5396 10484 5524 10516
rect 5556 10484 5684 10516
rect 5716 10484 5720 10516
rect 4720 10480 5720 10484
rect 5760 10516 5960 10520
rect 5760 10484 5764 10516
rect 5796 10484 5924 10516
rect 5956 10484 5960 10516
rect 5760 10480 5960 10484
rect 6000 10516 6200 10520
rect 6000 10484 6004 10516
rect 6036 10484 6164 10516
rect 6196 10484 6200 10516
rect 6000 10480 6200 10484
rect 4240 10436 4440 10440
rect 4240 10404 4244 10436
rect 4276 10404 4404 10436
rect 4436 10404 4440 10436
rect 4240 10400 4440 10404
rect 4480 10436 4680 10440
rect 4480 10404 4484 10436
rect 4516 10404 4644 10436
rect 4676 10404 4680 10436
rect 4480 10400 4680 10404
rect 4720 10436 5720 10440
rect 4720 10404 4724 10436
rect 4756 10404 4884 10436
rect 4916 10404 5044 10436
rect 5076 10404 5204 10436
rect 5236 10404 5364 10436
rect 5396 10404 5524 10436
rect 5556 10404 5684 10436
rect 5716 10404 5720 10436
rect 4720 10400 5720 10404
rect 5760 10436 5960 10440
rect 5760 10404 5764 10436
rect 5796 10404 5924 10436
rect 5956 10404 5960 10436
rect 5760 10400 5960 10404
rect 6000 10436 6200 10440
rect 6000 10404 6004 10436
rect 6036 10404 6164 10436
rect 6196 10404 6200 10436
rect 6000 10400 6200 10404
rect 4240 10356 4440 10360
rect 4240 10324 4244 10356
rect 4276 10324 4404 10356
rect 4436 10324 4440 10356
rect 4240 10320 4440 10324
rect 4480 10356 4680 10360
rect 4480 10324 4484 10356
rect 4516 10324 4644 10356
rect 4676 10324 4680 10356
rect 4480 10320 4680 10324
rect 4720 10356 5720 10360
rect 4720 10324 4724 10356
rect 4756 10324 4884 10356
rect 4916 10324 5044 10356
rect 5076 10324 5204 10356
rect 5236 10324 5364 10356
rect 5396 10324 5524 10356
rect 5556 10324 5684 10356
rect 5716 10324 5720 10356
rect 4720 10320 5720 10324
rect 5760 10356 5960 10360
rect 5760 10324 5764 10356
rect 5796 10324 5924 10356
rect 5956 10324 5960 10356
rect 5760 10320 5960 10324
rect 6000 10356 6200 10360
rect 6000 10324 6004 10356
rect 6036 10324 6164 10356
rect 6196 10324 6200 10356
rect 6000 10320 6200 10324
rect 4240 10276 4440 10280
rect 4240 10244 4244 10276
rect 4276 10244 4404 10276
rect 4436 10244 4440 10276
rect 4240 10240 4440 10244
rect 4480 10276 4680 10280
rect 4480 10244 4484 10276
rect 4516 10244 4644 10276
rect 4676 10244 4680 10276
rect 4480 10240 4680 10244
rect 4720 10276 5720 10280
rect 4720 10244 4724 10276
rect 4756 10244 4884 10276
rect 4916 10244 5044 10276
rect 5076 10244 5204 10276
rect 5236 10244 5364 10276
rect 5396 10244 5524 10276
rect 5556 10244 5684 10276
rect 5716 10244 5720 10276
rect 4720 10240 5720 10244
rect 5760 10276 5960 10280
rect 5760 10244 5764 10276
rect 5796 10244 5924 10276
rect 5956 10244 5960 10276
rect 5760 10240 5960 10244
rect 6000 10276 6200 10280
rect 6000 10244 6004 10276
rect 6036 10244 6164 10276
rect 6196 10244 6200 10276
rect 6000 10240 6200 10244
rect 4240 10196 4440 10200
rect 4240 10164 4244 10196
rect 4276 10164 4404 10196
rect 4436 10164 4440 10196
rect 4240 10160 4440 10164
rect 4480 10196 4680 10200
rect 4480 10164 4484 10196
rect 4516 10164 4644 10196
rect 4676 10164 4680 10196
rect 4480 10160 4680 10164
rect 4720 10196 5720 10200
rect 4720 10164 4724 10196
rect 4756 10164 4884 10196
rect 4916 10164 5044 10196
rect 5076 10164 5204 10196
rect 5236 10164 5364 10196
rect 5396 10164 5524 10196
rect 5556 10164 5684 10196
rect 5716 10164 5720 10196
rect 4720 10160 5720 10164
rect 5760 10196 5960 10200
rect 5760 10164 5764 10196
rect 5796 10164 5924 10196
rect 5956 10164 5960 10196
rect 5760 10160 5960 10164
rect 6000 10196 6200 10200
rect 6000 10164 6004 10196
rect 6036 10164 6164 10196
rect 6196 10164 6200 10196
rect 6000 10160 6200 10164
rect 4240 10116 4440 10120
rect 4240 10084 4244 10116
rect 4276 10084 4404 10116
rect 4436 10084 4440 10116
rect 4240 10080 4440 10084
rect 4480 10116 4680 10120
rect 4480 10084 4484 10116
rect 4516 10084 4644 10116
rect 4676 10084 4680 10116
rect 4480 10080 4680 10084
rect 4720 10116 5720 10120
rect 4720 10084 4724 10116
rect 4756 10084 4884 10116
rect 4916 10084 5044 10116
rect 5076 10084 5204 10116
rect 5236 10084 5364 10116
rect 5396 10084 5524 10116
rect 5556 10084 5684 10116
rect 5716 10084 5720 10116
rect 4720 10080 5720 10084
rect 5760 10116 5960 10120
rect 5760 10084 5764 10116
rect 5796 10084 5924 10116
rect 5956 10084 5960 10116
rect 5760 10080 5960 10084
rect 6000 10116 6200 10120
rect 6000 10084 6004 10116
rect 6036 10084 6164 10116
rect 6196 10084 6200 10116
rect 6000 10080 6200 10084
rect 4240 10036 4440 10040
rect 4240 10004 4244 10036
rect 4276 10004 4404 10036
rect 4436 10004 4440 10036
rect 4240 10000 4440 10004
rect 4480 10036 4680 10040
rect 4480 10004 4484 10036
rect 4516 10004 4644 10036
rect 4676 10004 4680 10036
rect 4480 10000 4680 10004
rect 4720 10036 5720 10040
rect 4720 10004 4724 10036
rect 4756 10004 4884 10036
rect 4916 10004 5044 10036
rect 5076 10004 5204 10036
rect 5236 10004 5364 10036
rect 5396 10004 5524 10036
rect 5556 10004 5684 10036
rect 5716 10004 5720 10036
rect 4720 10000 5720 10004
rect 5760 10036 5960 10040
rect 5760 10004 5764 10036
rect 5796 10004 5924 10036
rect 5956 10004 5960 10036
rect 5760 10000 5960 10004
rect 6000 10036 6200 10040
rect 6000 10004 6004 10036
rect 6036 10004 6164 10036
rect 6196 10004 6200 10036
rect 6000 10000 6200 10004
rect 4240 9956 4440 9960
rect 4240 9924 4244 9956
rect 4276 9924 4404 9956
rect 4436 9924 4440 9956
rect 4240 9920 4440 9924
rect 4480 9956 4680 9960
rect 4480 9924 4484 9956
rect 4516 9924 4644 9956
rect 4676 9924 4680 9956
rect 4480 9920 4680 9924
rect 4720 9956 5720 9960
rect 4720 9924 4724 9956
rect 4756 9924 4884 9956
rect 4916 9924 5044 9956
rect 5076 9924 5204 9956
rect 5236 9924 5364 9956
rect 5396 9924 5524 9956
rect 5556 9924 5684 9956
rect 5716 9924 5720 9956
rect 4720 9920 5720 9924
rect 5760 9956 5960 9960
rect 5760 9924 5764 9956
rect 5796 9924 5924 9956
rect 5956 9924 5960 9956
rect 5760 9920 5960 9924
rect 6000 9956 6200 9960
rect 6000 9924 6004 9956
rect 6036 9924 6164 9956
rect 6196 9924 6200 9956
rect 6000 9920 6200 9924
rect 4240 9876 4440 9880
rect 4240 9844 4244 9876
rect 4276 9844 4404 9876
rect 4436 9844 4440 9876
rect 4240 9840 4440 9844
rect 4480 9876 4680 9880
rect 4480 9844 4484 9876
rect 4516 9844 4644 9876
rect 4676 9844 4680 9876
rect 4480 9840 4680 9844
rect 4720 9876 5720 9880
rect 4720 9844 4724 9876
rect 4756 9844 4884 9876
rect 4916 9844 5044 9876
rect 5076 9844 5204 9876
rect 5236 9844 5364 9876
rect 5396 9844 5524 9876
rect 5556 9844 5684 9876
rect 5716 9844 5720 9876
rect 4720 9840 5720 9844
rect 5760 9876 5960 9880
rect 5760 9844 5764 9876
rect 5796 9844 5924 9876
rect 5956 9844 5960 9876
rect 5760 9840 5960 9844
rect 6000 9876 6200 9880
rect 6000 9844 6004 9876
rect 6036 9844 6164 9876
rect 6196 9844 6200 9876
rect 6000 9840 6200 9844
rect 4240 9796 4440 9800
rect 4240 9764 4244 9796
rect 4276 9764 4404 9796
rect 4436 9764 4440 9796
rect 4240 9760 4440 9764
rect 4480 9796 4680 9800
rect 4480 9764 4484 9796
rect 4516 9764 4644 9796
rect 4676 9764 4680 9796
rect 4480 9760 4680 9764
rect 4720 9796 5720 9800
rect 4720 9764 4724 9796
rect 4756 9764 4884 9796
rect 4916 9764 5044 9796
rect 5076 9764 5204 9796
rect 5236 9764 5364 9796
rect 5396 9764 5524 9796
rect 5556 9764 5684 9796
rect 5716 9764 5720 9796
rect 4720 9760 5720 9764
rect 5760 9796 5960 9800
rect 5760 9764 5764 9796
rect 5796 9764 5924 9796
rect 5956 9764 5960 9796
rect 5760 9760 5960 9764
rect 6000 9796 6200 9800
rect 6000 9764 6004 9796
rect 6036 9764 6164 9796
rect 6196 9764 6200 9796
rect 6000 9760 6200 9764
rect 4240 9716 4440 9720
rect 4240 9684 4244 9716
rect 4276 9684 4404 9716
rect 4436 9684 4440 9716
rect 4240 9680 4440 9684
rect 4480 9716 4680 9720
rect 4480 9684 4484 9716
rect 4516 9684 4644 9716
rect 4676 9684 4680 9716
rect 4480 9680 4680 9684
rect 4720 9716 5720 9720
rect 4720 9684 4724 9716
rect 4756 9684 4884 9716
rect 4916 9684 5044 9716
rect 5076 9684 5204 9716
rect 5236 9684 5364 9716
rect 5396 9684 5524 9716
rect 5556 9684 5684 9716
rect 5716 9684 5720 9716
rect 4720 9680 5720 9684
rect 5760 9716 5960 9720
rect 5760 9684 5764 9716
rect 5796 9684 5924 9716
rect 5956 9684 5960 9716
rect 5760 9680 5960 9684
rect 6000 9716 6200 9720
rect 6000 9684 6004 9716
rect 6036 9684 6164 9716
rect 6196 9684 6200 9716
rect 6000 9680 6200 9684
rect 4240 9636 4440 9640
rect 4240 9604 4244 9636
rect 4276 9604 4404 9636
rect 4436 9604 4440 9636
rect 4240 9600 4440 9604
rect 4480 9636 4680 9640
rect 4480 9604 4484 9636
rect 4516 9604 4644 9636
rect 4676 9604 4680 9636
rect 4480 9600 4680 9604
rect 4720 9636 5720 9640
rect 4720 9604 4724 9636
rect 4756 9604 4884 9636
rect 4916 9604 5044 9636
rect 5076 9604 5204 9636
rect 5236 9604 5364 9636
rect 5396 9604 5524 9636
rect 5556 9604 5684 9636
rect 5716 9604 5720 9636
rect 4720 9600 5720 9604
rect 5760 9636 5960 9640
rect 5760 9604 5764 9636
rect 5796 9604 5924 9636
rect 5956 9604 5960 9636
rect 5760 9600 5960 9604
rect 6000 9636 6200 9640
rect 6000 9604 6004 9636
rect 6036 9604 6164 9636
rect 6196 9604 6200 9636
rect 6000 9600 6200 9604
rect 4240 9556 4440 9560
rect 4240 9524 4244 9556
rect 4276 9524 4404 9556
rect 4436 9524 4440 9556
rect 4240 9520 4440 9524
rect 4480 9556 4680 9560
rect 4480 9524 4484 9556
rect 4516 9524 4644 9556
rect 4676 9524 4680 9556
rect 4480 9520 4680 9524
rect 4720 9556 5720 9560
rect 4720 9524 4724 9556
rect 4756 9524 4884 9556
rect 4916 9524 5044 9556
rect 5076 9524 5204 9556
rect 5236 9524 5364 9556
rect 5396 9524 5524 9556
rect 5556 9524 5684 9556
rect 5716 9524 5720 9556
rect 4720 9520 5720 9524
rect 5760 9556 5960 9560
rect 5760 9524 5764 9556
rect 5796 9524 5924 9556
rect 5956 9524 5960 9556
rect 5760 9520 5960 9524
rect 6000 9556 6200 9560
rect 6000 9524 6004 9556
rect 6036 9524 6164 9556
rect 6196 9524 6200 9556
rect 6000 9520 6200 9524
rect 4240 9476 4440 9480
rect 4240 9444 4244 9476
rect 4276 9444 4404 9476
rect 4436 9444 4440 9476
rect 4240 9440 4440 9444
rect 4480 9476 4680 9480
rect 4480 9444 4484 9476
rect 4516 9444 4644 9476
rect 4676 9444 4680 9476
rect 4480 9440 4680 9444
rect 4720 9476 5720 9480
rect 4720 9444 4724 9476
rect 4756 9444 4884 9476
rect 4916 9444 5044 9476
rect 5076 9444 5204 9476
rect 5236 9444 5364 9476
rect 5396 9444 5524 9476
rect 5556 9444 5684 9476
rect 5716 9444 5720 9476
rect 4720 9440 5720 9444
rect 5760 9476 5960 9480
rect 5760 9444 5764 9476
rect 5796 9444 5924 9476
rect 5956 9444 5960 9476
rect 5760 9440 5960 9444
rect 6000 9476 6200 9480
rect 6000 9444 6004 9476
rect 6036 9444 6164 9476
rect 6196 9444 6200 9476
rect 6000 9440 6200 9444
rect 4240 9396 4440 9400
rect 4240 9364 4244 9396
rect 4276 9364 4404 9396
rect 4436 9364 4440 9396
rect 4240 9360 4440 9364
rect 4480 9396 4680 9400
rect 4480 9364 4484 9396
rect 4516 9364 4644 9396
rect 4676 9364 4680 9396
rect 4480 9360 4680 9364
rect 4720 9396 5720 9400
rect 4720 9364 4724 9396
rect 4756 9364 4884 9396
rect 4916 9364 5044 9396
rect 5076 9364 5204 9396
rect 5236 9364 5364 9396
rect 5396 9364 5524 9396
rect 5556 9364 5684 9396
rect 5716 9364 5720 9396
rect 4720 9360 5720 9364
rect 5760 9396 5960 9400
rect 5760 9364 5764 9396
rect 5796 9364 5924 9396
rect 5956 9364 5960 9396
rect 5760 9360 5960 9364
rect 6000 9396 6200 9400
rect 6000 9364 6004 9396
rect 6036 9364 6164 9396
rect 6196 9364 6200 9396
rect 6000 9360 6200 9364
rect 4240 9316 4440 9320
rect 4240 9284 4244 9316
rect 4276 9284 4404 9316
rect 4436 9284 4440 9316
rect 4240 9280 4440 9284
rect 4480 9316 4680 9320
rect 4480 9284 4484 9316
rect 4516 9284 4644 9316
rect 4676 9284 4680 9316
rect 4480 9280 4680 9284
rect 4720 9316 5720 9320
rect 4720 9284 4724 9316
rect 4756 9284 4884 9316
rect 4916 9284 5044 9316
rect 5076 9284 5204 9316
rect 5236 9284 5364 9316
rect 5396 9284 5524 9316
rect 5556 9284 5684 9316
rect 5716 9284 5720 9316
rect 4720 9280 5720 9284
rect 5760 9316 5960 9320
rect 5760 9284 5764 9316
rect 5796 9284 5924 9316
rect 5956 9284 5960 9316
rect 5760 9280 5960 9284
rect 6000 9316 6200 9320
rect 6000 9284 6004 9316
rect 6036 9284 6164 9316
rect 6196 9284 6200 9316
rect 6000 9280 6200 9284
rect 4240 9236 4440 9240
rect 4240 9204 4244 9236
rect 4276 9204 4404 9236
rect 4436 9204 4440 9236
rect 4240 9200 4440 9204
rect 4480 9236 4680 9240
rect 4480 9204 4484 9236
rect 4516 9204 4644 9236
rect 4676 9204 4680 9236
rect 4480 9200 4680 9204
rect 4720 9236 5720 9240
rect 4720 9204 4724 9236
rect 4756 9204 4884 9236
rect 4916 9204 5044 9236
rect 5076 9204 5204 9236
rect 5236 9204 5364 9236
rect 5396 9204 5524 9236
rect 5556 9204 5684 9236
rect 5716 9204 5720 9236
rect 4720 9200 5720 9204
rect 5760 9236 5960 9240
rect 5760 9204 5764 9236
rect 5796 9204 5924 9236
rect 5956 9204 5960 9236
rect 5760 9200 5960 9204
rect 6000 9236 6200 9240
rect 6000 9204 6004 9236
rect 6036 9204 6164 9236
rect 6196 9204 6200 9236
rect 6000 9200 6200 9204
rect 4240 9156 4440 9160
rect 4240 9124 4244 9156
rect 4276 9124 4404 9156
rect 4436 9124 4440 9156
rect 4240 9120 4440 9124
rect 4480 9156 4680 9160
rect 4480 9124 4484 9156
rect 4516 9124 4644 9156
rect 4676 9124 4680 9156
rect 4480 9120 4680 9124
rect 4720 9156 5720 9160
rect 4720 9124 4724 9156
rect 4756 9124 4884 9156
rect 4916 9124 5044 9156
rect 5076 9124 5204 9156
rect 5236 9124 5364 9156
rect 5396 9124 5524 9156
rect 5556 9124 5684 9156
rect 5716 9124 5720 9156
rect 4720 9120 5720 9124
rect 5760 9156 5960 9160
rect 5760 9124 5764 9156
rect 5796 9124 5924 9156
rect 5956 9124 5960 9156
rect 5760 9120 5960 9124
rect 6000 9156 6200 9160
rect 6000 9124 6004 9156
rect 6036 9124 6164 9156
rect 6196 9124 6200 9156
rect 6000 9120 6200 9124
rect 4240 9076 4440 9080
rect 4240 9044 4244 9076
rect 4276 9044 4404 9076
rect 4436 9044 4440 9076
rect 4240 9040 4440 9044
rect 4480 9076 4680 9080
rect 4480 9044 4484 9076
rect 4516 9044 4644 9076
rect 4676 9044 4680 9076
rect 4480 9040 4680 9044
rect 4720 9076 5720 9080
rect 4720 9044 4724 9076
rect 4756 9044 4884 9076
rect 4916 9044 5044 9076
rect 5076 9044 5204 9076
rect 5236 9044 5364 9076
rect 5396 9044 5524 9076
rect 5556 9044 5684 9076
rect 5716 9044 5720 9076
rect 4720 9040 5720 9044
rect 5760 9076 5960 9080
rect 5760 9044 5764 9076
rect 5796 9044 5924 9076
rect 5956 9044 5960 9076
rect 5760 9040 5960 9044
rect 6000 9076 6200 9080
rect 6000 9044 6004 9076
rect 6036 9044 6164 9076
rect 6196 9044 6200 9076
rect 6000 9040 6200 9044
rect 4240 8996 4440 9000
rect 4240 8964 4244 8996
rect 4276 8964 4404 8996
rect 4436 8964 4440 8996
rect 4240 8960 4440 8964
rect 4480 8996 4680 9000
rect 4480 8964 4484 8996
rect 4516 8964 4644 8996
rect 4676 8964 4680 8996
rect 4480 8960 4680 8964
rect 4720 8996 5720 9000
rect 4720 8964 4724 8996
rect 4756 8964 4884 8996
rect 4916 8964 5044 8996
rect 5076 8964 5204 8996
rect 5236 8964 5364 8996
rect 5396 8964 5524 8996
rect 5556 8964 5684 8996
rect 5716 8964 5720 8996
rect 4720 8960 5720 8964
rect 5760 8996 5960 9000
rect 5760 8964 5764 8996
rect 5796 8964 5924 8996
rect 5956 8964 5960 8996
rect 5760 8960 5960 8964
rect 6000 8996 6200 9000
rect 6000 8964 6004 8996
rect 6036 8964 6164 8996
rect 6196 8964 6200 8996
rect 6000 8960 6200 8964
rect 4240 8916 4440 8920
rect 4240 8884 4244 8916
rect 4276 8884 4404 8916
rect 4436 8884 4440 8916
rect 4240 8880 4440 8884
rect 4480 8916 4680 8920
rect 4480 8884 4484 8916
rect 4516 8884 4644 8916
rect 4676 8884 4680 8916
rect 4480 8880 4680 8884
rect 4720 8916 5720 8920
rect 4720 8884 4724 8916
rect 4756 8884 4884 8916
rect 4916 8884 5044 8916
rect 5076 8884 5204 8916
rect 5236 8884 5364 8916
rect 5396 8884 5524 8916
rect 5556 8884 5684 8916
rect 5716 8884 5720 8916
rect 4720 8880 5720 8884
rect 5760 8916 5960 8920
rect 5760 8884 5764 8916
rect 5796 8884 5924 8916
rect 5956 8884 5960 8916
rect 5760 8880 5960 8884
rect 6000 8916 6200 8920
rect 6000 8884 6004 8916
rect 6036 8884 6164 8916
rect 6196 8884 6200 8916
rect 6000 8880 6200 8884
rect 4240 8836 4440 8840
rect 4240 8804 4244 8836
rect 4276 8804 4404 8836
rect 4436 8804 4440 8836
rect 4240 8800 4440 8804
rect 4480 8836 4680 8840
rect 4480 8804 4484 8836
rect 4516 8804 4644 8836
rect 4676 8804 4680 8836
rect 4480 8800 4680 8804
rect 4720 8836 5720 8840
rect 4720 8804 4724 8836
rect 4756 8804 4884 8836
rect 4916 8804 5044 8836
rect 5076 8804 5204 8836
rect 5236 8804 5364 8836
rect 5396 8804 5524 8836
rect 5556 8804 5684 8836
rect 5716 8804 5720 8836
rect 4720 8800 5720 8804
rect 5760 8836 5960 8840
rect 5760 8804 5764 8836
rect 5796 8804 5924 8836
rect 5956 8804 5960 8836
rect 5760 8800 5960 8804
rect 6000 8836 6200 8840
rect 6000 8804 6004 8836
rect 6036 8804 6164 8836
rect 6196 8804 6200 8836
rect 6000 8800 6200 8804
rect 4240 8756 4440 8760
rect 4240 8724 4244 8756
rect 4276 8724 4404 8756
rect 4436 8724 4440 8756
rect 4240 8720 4440 8724
rect 4480 8756 4680 8760
rect 4480 8724 4484 8756
rect 4516 8724 4644 8756
rect 4676 8724 4680 8756
rect 4480 8720 4680 8724
rect 4720 8756 5720 8760
rect 4720 8724 4724 8756
rect 4756 8724 4884 8756
rect 4916 8724 5044 8756
rect 5076 8724 5204 8756
rect 5236 8724 5364 8756
rect 5396 8724 5524 8756
rect 5556 8724 5684 8756
rect 5716 8724 5720 8756
rect 4720 8720 5720 8724
rect 5760 8756 5960 8760
rect 5760 8724 5764 8756
rect 5796 8724 5924 8756
rect 5956 8724 5960 8756
rect 5760 8720 5960 8724
rect 6000 8756 6200 8760
rect 6000 8724 6004 8756
rect 6036 8724 6164 8756
rect 6196 8724 6200 8756
rect 6000 8720 6200 8724
rect 4240 8676 4440 8680
rect 4240 8644 4244 8676
rect 4276 8644 4404 8676
rect 4436 8644 4440 8676
rect 4240 8640 4440 8644
rect 4480 8676 4680 8680
rect 4480 8644 4484 8676
rect 4516 8644 4644 8676
rect 4676 8644 4680 8676
rect 4480 8640 4680 8644
rect 4720 8676 5720 8680
rect 4720 8644 4724 8676
rect 4756 8644 4884 8676
rect 4916 8644 5044 8676
rect 5076 8644 5204 8676
rect 5236 8644 5364 8676
rect 5396 8644 5524 8676
rect 5556 8644 5684 8676
rect 5716 8644 5720 8676
rect 4720 8640 5720 8644
rect 5760 8676 5960 8680
rect 5760 8644 5764 8676
rect 5796 8644 5924 8676
rect 5956 8644 5960 8676
rect 5760 8640 5960 8644
rect 6000 8676 6200 8680
rect 6000 8644 6004 8676
rect 6036 8644 6164 8676
rect 6196 8644 6200 8676
rect 6000 8640 6200 8644
rect 4240 8596 4440 8600
rect 4240 8564 4244 8596
rect 4276 8564 4404 8596
rect 4436 8564 4440 8596
rect 4240 8560 4440 8564
rect 4480 8596 4680 8600
rect 4480 8564 4484 8596
rect 4516 8564 4644 8596
rect 4676 8564 4680 8596
rect 4480 8560 4680 8564
rect 4720 8596 5720 8600
rect 4720 8564 4724 8596
rect 4756 8564 4884 8596
rect 4916 8564 5044 8596
rect 5076 8564 5204 8596
rect 5236 8564 5364 8596
rect 5396 8564 5524 8596
rect 5556 8564 5684 8596
rect 5716 8564 5720 8596
rect 4720 8560 5720 8564
rect 5760 8596 5960 8600
rect 5760 8564 5764 8596
rect 5796 8564 5924 8596
rect 5956 8564 5960 8596
rect 5760 8560 5960 8564
rect 6000 8596 6200 8600
rect 6000 8564 6004 8596
rect 6036 8564 6164 8596
rect 6196 8564 6200 8596
rect 6000 8560 6200 8564
rect 4240 8516 4440 8520
rect 4240 8484 4244 8516
rect 4276 8484 4404 8516
rect 4436 8484 4440 8516
rect 4240 8480 4440 8484
rect 4480 8516 4680 8520
rect 4480 8484 4484 8516
rect 4516 8484 4644 8516
rect 4676 8484 4680 8516
rect 4480 8480 4680 8484
rect 4720 8516 5720 8520
rect 4720 8484 4724 8516
rect 4756 8484 4884 8516
rect 4916 8484 5044 8516
rect 5076 8484 5204 8516
rect 5236 8484 5364 8516
rect 5396 8484 5524 8516
rect 5556 8484 5684 8516
rect 5716 8484 5720 8516
rect 4720 8480 5720 8484
rect 5760 8516 5960 8520
rect 5760 8484 5764 8516
rect 5796 8484 5924 8516
rect 5956 8484 5960 8516
rect 5760 8480 5960 8484
rect 6000 8516 6200 8520
rect 6000 8484 6004 8516
rect 6036 8484 6164 8516
rect 6196 8484 6200 8516
rect 6000 8480 6200 8484
rect 4240 8436 4440 8440
rect 4240 8404 4244 8436
rect 4276 8404 4404 8436
rect 4436 8404 4440 8436
rect 4240 8400 4440 8404
rect 4480 8436 4680 8440
rect 4480 8404 4484 8436
rect 4516 8404 4644 8436
rect 4676 8404 4680 8436
rect 4480 8400 4680 8404
rect 4720 8436 5720 8440
rect 4720 8404 4724 8436
rect 4756 8404 4884 8436
rect 4916 8404 5044 8436
rect 5076 8404 5204 8436
rect 5236 8404 5364 8436
rect 5396 8404 5524 8436
rect 5556 8404 5684 8436
rect 5716 8404 5720 8436
rect 4720 8400 5720 8404
rect 5760 8436 5960 8440
rect 5760 8404 5764 8436
rect 5796 8404 5924 8436
rect 5956 8404 5960 8436
rect 5760 8400 5960 8404
rect 6000 8436 6200 8440
rect 6000 8404 6004 8436
rect 6036 8404 6164 8436
rect 6196 8404 6200 8436
rect 6000 8400 6200 8404
rect 4240 8356 4440 8360
rect 4240 8324 4244 8356
rect 4276 8324 4404 8356
rect 4436 8324 4440 8356
rect 4240 8320 4440 8324
rect 4480 8356 4680 8360
rect 4480 8324 4484 8356
rect 4516 8324 4644 8356
rect 4676 8324 4680 8356
rect 4480 8320 4680 8324
rect 4720 8356 5720 8360
rect 4720 8324 4724 8356
rect 4756 8324 4884 8356
rect 4916 8324 5044 8356
rect 5076 8324 5204 8356
rect 5236 8324 5364 8356
rect 5396 8324 5524 8356
rect 5556 8324 5684 8356
rect 5716 8324 5720 8356
rect 4720 8320 5720 8324
rect 5760 8356 5960 8360
rect 5760 8324 5764 8356
rect 5796 8324 5924 8356
rect 5956 8324 5960 8356
rect 5760 8320 5960 8324
rect 6000 8356 6200 8360
rect 6000 8324 6004 8356
rect 6036 8324 6164 8356
rect 6196 8324 6200 8356
rect 6000 8320 6200 8324
rect 4240 8276 4440 8280
rect 4240 8244 4244 8276
rect 4276 8244 4404 8276
rect 4436 8244 4440 8276
rect 4240 8240 4440 8244
rect 4480 8276 4680 8280
rect 4480 8244 4484 8276
rect 4516 8244 4644 8276
rect 4676 8244 4680 8276
rect 4480 8240 4680 8244
rect 4720 8276 5720 8280
rect 4720 8244 4724 8276
rect 4756 8244 4884 8276
rect 4916 8244 5044 8276
rect 5076 8244 5204 8276
rect 5236 8244 5364 8276
rect 5396 8244 5524 8276
rect 5556 8244 5684 8276
rect 5716 8244 5720 8276
rect 4720 8240 5720 8244
rect 5760 8276 5960 8280
rect 5760 8244 5764 8276
rect 5796 8244 5924 8276
rect 5956 8244 5960 8276
rect 5760 8240 5960 8244
rect 6000 8276 6200 8280
rect 6000 8244 6004 8276
rect 6036 8244 6164 8276
rect 6196 8244 6200 8276
rect 6000 8240 6200 8244
rect 4240 8196 4440 8200
rect 4240 8164 4244 8196
rect 4276 8164 4404 8196
rect 4436 8164 4440 8196
rect 4240 8160 4440 8164
rect 4480 8196 4680 8200
rect 4480 8164 4484 8196
rect 4516 8164 4644 8196
rect 4676 8164 4680 8196
rect 4480 8160 4680 8164
rect 4720 8196 5720 8200
rect 4720 8164 4724 8196
rect 4756 8164 4884 8196
rect 4916 8164 5044 8196
rect 5076 8164 5204 8196
rect 5236 8164 5364 8196
rect 5396 8164 5524 8196
rect 5556 8164 5684 8196
rect 5716 8164 5720 8196
rect 4720 8160 5720 8164
rect 5760 8196 5960 8200
rect 5760 8164 5764 8196
rect 5796 8164 5924 8196
rect 5956 8164 5960 8196
rect 5760 8160 5960 8164
rect 6000 8196 6200 8200
rect 6000 8164 6004 8196
rect 6036 8164 6164 8196
rect 6196 8164 6200 8196
rect 6000 8160 6200 8164
rect 4240 8116 4440 8120
rect 4240 8084 4244 8116
rect 4276 8084 4404 8116
rect 4436 8084 4440 8116
rect 4240 8080 4440 8084
rect 4480 8116 4680 8120
rect 4480 8084 4484 8116
rect 4516 8084 4644 8116
rect 4676 8084 4680 8116
rect 4480 8080 4680 8084
rect 4720 8116 5720 8120
rect 4720 8084 4724 8116
rect 4756 8084 4884 8116
rect 4916 8084 5044 8116
rect 5076 8084 5204 8116
rect 5236 8084 5364 8116
rect 5396 8084 5524 8116
rect 5556 8084 5684 8116
rect 5716 8084 5720 8116
rect 4720 8080 5720 8084
rect 5760 8116 5960 8120
rect 5760 8084 5764 8116
rect 5796 8084 5924 8116
rect 5956 8084 5960 8116
rect 5760 8080 5960 8084
rect 6000 8116 6200 8120
rect 6000 8084 6004 8116
rect 6036 8084 6164 8116
rect 6196 8084 6200 8116
rect 6000 8080 6200 8084
rect 4240 8036 4440 8040
rect 4240 8004 4244 8036
rect 4276 8004 4404 8036
rect 4436 8004 4440 8036
rect 4240 8000 4440 8004
rect 4480 8036 4680 8040
rect 4480 8004 4484 8036
rect 4516 8004 4644 8036
rect 4676 8004 4680 8036
rect 4480 8000 4680 8004
rect 4720 8036 5720 8040
rect 4720 8004 4724 8036
rect 4756 8004 4884 8036
rect 4916 8004 5044 8036
rect 5076 8004 5204 8036
rect 5236 8004 5364 8036
rect 5396 8004 5524 8036
rect 5556 8004 5684 8036
rect 5716 8004 5720 8036
rect 4720 8000 5720 8004
rect 5760 8036 5960 8040
rect 5760 8004 5764 8036
rect 5796 8004 5924 8036
rect 5956 8004 5960 8036
rect 5760 8000 5960 8004
rect 6000 8036 6200 8040
rect 6000 8004 6004 8036
rect 6036 8004 6164 8036
rect 6196 8004 6200 8036
rect 6000 8000 6200 8004
rect 4240 7956 4440 7960
rect 4240 7924 4244 7956
rect 4276 7924 4404 7956
rect 4436 7924 4440 7956
rect 4240 7920 4440 7924
rect 4480 7956 4680 7960
rect 4480 7924 4484 7956
rect 4516 7924 4644 7956
rect 4676 7924 4680 7956
rect 4480 7920 4680 7924
rect 4720 7956 5720 7960
rect 4720 7924 4724 7956
rect 4756 7924 4884 7956
rect 4916 7924 5044 7956
rect 5076 7924 5204 7956
rect 5236 7924 5364 7956
rect 5396 7924 5524 7956
rect 5556 7924 5684 7956
rect 5716 7924 5720 7956
rect 4720 7920 5720 7924
rect 5760 7956 5960 7960
rect 5760 7924 5764 7956
rect 5796 7924 5924 7956
rect 5956 7924 5960 7956
rect 5760 7920 5960 7924
rect 6000 7956 6200 7960
rect 6000 7924 6004 7956
rect 6036 7924 6164 7956
rect 6196 7924 6200 7956
rect 6000 7920 6200 7924
rect 4240 7876 4440 7880
rect 4240 7844 4244 7876
rect 4276 7844 4404 7876
rect 4436 7844 4440 7876
rect 4240 7840 4440 7844
rect 4480 7876 4680 7880
rect 4480 7844 4484 7876
rect 4516 7844 4644 7876
rect 4676 7844 4680 7876
rect 4480 7840 4680 7844
rect 4720 7876 5720 7880
rect 4720 7844 4724 7876
rect 4756 7844 4884 7876
rect 4916 7844 5044 7876
rect 5076 7844 5204 7876
rect 5236 7844 5364 7876
rect 5396 7844 5524 7876
rect 5556 7844 5684 7876
rect 5716 7844 5720 7876
rect 4720 7840 5720 7844
rect 5760 7876 5960 7880
rect 5760 7844 5764 7876
rect 5796 7844 5924 7876
rect 5956 7844 5960 7876
rect 5760 7840 5960 7844
rect 6000 7876 6200 7880
rect 6000 7844 6004 7876
rect 6036 7844 6164 7876
rect 6196 7844 6200 7876
rect 6000 7840 6200 7844
rect 4240 7796 4440 7800
rect 4240 7764 4244 7796
rect 4276 7764 4404 7796
rect 4436 7764 4440 7796
rect 4240 7760 4440 7764
rect 4480 7796 4680 7800
rect 4480 7764 4484 7796
rect 4516 7764 4644 7796
rect 4676 7764 4680 7796
rect 4480 7760 4680 7764
rect 4720 7796 5720 7800
rect 4720 7764 4724 7796
rect 4756 7764 4884 7796
rect 4916 7764 5044 7796
rect 5076 7764 5204 7796
rect 5236 7764 5364 7796
rect 5396 7764 5524 7796
rect 5556 7764 5684 7796
rect 5716 7764 5720 7796
rect 4720 7760 5720 7764
rect 5760 7796 5960 7800
rect 5760 7764 5764 7796
rect 5796 7764 5924 7796
rect 5956 7764 5960 7796
rect 5760 7760 5960 7764
rect 6000 7796 6200 7800
rect 6000 7764 6004 7796
rect 6036 7764 6164 7796
rect 6196 7764 6200 7796
rect 6000 7760 6200 7764
rect 4240 7716 4440 7720
rect 4240 7684 4244 7716
rect 4276 7684 4404 7716
rect 4436 7684 4440 7716
rect 4240 7680 4440 7684
rect 4480 7716 4680 7720
rect 4480 7684 4484 7716
rect 4516 7684 4644 7716
rect 4676 7684 4680 7716
rect 4480 7680 4680 7684
rect 4720 7716 5720 7720
rect 4720 7684 4724 7716
rect 4756 7684 4884 7716
rect 4916 7684 5044 7716
rect 5076 7684 5204 7716
rect 5236 7684 5364 7716
rect 5396 7684 5524 7716
rect 5556 7684 5684 7716
rect 5716 7684 5720 7716
rect 4720 7680 5720 7684
rect 5760 7716 5960 7720
rect 5760 7684 5764 7716
rect 5796 7684 5924 7716
rect 5956 7684 5960 7716
rect 5760 7680 5960 7684
rect 6000 7716 6200 7720
rect 6000 7684 6004 7716
rect 6036 7684 6164 7716
rect 6196 7684 6200 7716
rect 6000 7680 6200 7684
rect 4240 7636 4440 7640
rect 4240 7604 4244 7636
rect 4276 7604 4404 7636
rect 4436 7604 4440 7636
rect 4240 7600 4440 7604
rect 4480 7636 4680 7640
rect 4480 7604 4484 7636
rect 4516 7604 4644 7636
rect 4676 7604 4680 7636
rect 4480 7600 4680 7604
rect 4720 7636 5720 7640
rect 4720 7604 4724 7636
rect 4756 7604 4884 7636
rect 4916 7604 5044 7636
rect 5076 7604 5204 7636
rect 5236 7604 5364 7636
rect 5396 7604 5524 7636
rect 5556 7604 5684 7636
rect 5716 7604 5720 7636
rect 4720 7600 5720 7604
rect 5760 7636 5960 7640
rect 5760 7604 5764 7636
rect 5796 7604 5924 7636
rect 5956 7604 5960 7636
rect 5760 7600 5960 7604
rect 6000 7636 6200 7640
rect 6000 7604 6004 7636
rect 6036 7604 6164 7636
rect 6196 7604 6200 7636
rect 6000 7600 6200 7604
rect 4240 7556 4440 7560
rect 4240 7524 4244 7556
rect 4276 7524 4404 7556
rect 4436 7524 4440 7556
rect 4240 7520 4440 7524
rect 4480 7556 4680 7560
rect 4480 7524 4484 7556
rect 4516 7524 4644 7556
rect 4676 7524 4680 7556
rect 4480 7520 4680 7524
rect 4720 7556 5720 7560
rect 4720 7524 4724 7556
rect 4756 7524 4884 7556
rect 4916 7524 5044 7556
rect 5076 7524 5204 7556
rect 5236 7524 5364 7556
rect 5396 7524 5524 7556
rect 5556 7524 5684 7556
rect 5716 7524 5720 7556
rect 4720 7520 5720 7524
rect 5760 7556 5960 7560
rect 5760 7524 5764 7556
rect 5796 7524 5924 7556
rect 5956 7524 5960 7556
rect 5760 7520 5960 7524
rect 6000 7556 6200 7560
rect 6000 7524 6004 7556
rect 6036 7524 6164 7556
rect 6196 7524 6200 7556
rect 6000 7520 6200 7524
rect 4240 7476 4440 7480
rect 4240 7444 4244 7476
rect 4276 7444 4404 7476
rect 4436 7444 4440 7476
rect 4240 7440 4440 7444
rect 4480 7476 4680 7480
rect 4480 7444 4484 7476
rect 4516 7444 4644 7476
rect 4676 7444 4680 7476
rect 4480 7440 4680 7444
rect 4720 7476 5720 7480
rect 4720 7444 4724 7476
rect 4756 7444 4884 7476
rect 4916 7444 5044 7476
rect 5076 7444 5204 7476
rect 5236 7444 5364 7476
rect 5396 7444 5524 7476
rect 5556 7444 5684 7476
rect 5716 7444 5720 7476
rect 4720 7440 5720 7444
rect 5760 7476 5960 7480
rect 5760 7444 5764 7476
rect 5796 7444 5924 7476
rect 5956 7444 5960 7476
rect 5760 7440 5960 7444
rect 6000 7476 6200 7480
rect 6000 7444 6004 7476
rect 6036 7444 6164 7476
rect 6196 7444 6200 7476
rect 6000 7440 6200 7444
rect 4240 7396 4440 7400
rect 4240 7364 4244 7396
rect 4276 7364 4404 7396
rect 4436 7364 4440 7396
rect 4240 7360 4440 7364
rect 4480 7396 4680 7400
rect 4480 7364 4484 7396
rect 4516 7364 4644 7396
rect 4676 7364 4680 7396
rect 4480 7360 4680 7364
rect 4720 7396 5720 7400
rect 4720 7364 4724 7396
rect 4756 7364 4884 7396
rect 4916 7364 5044 7396
rect 5076 7364 5204 7396
rect 5236 7364 5364 7396
rect 5396 7364 5524 7396
rect 5556 7364 5684 7396
rect 5716 7364 5720 7396
rect 4720 7360 5720 7364
rect 5760 7396 5960 7400
rect 5760 7364 5764 7396
rect 5796 7364 5924 7396
rect 5956 7364 5960 7396
rect 5760 7360 5960 7364
rect 6000 7396 6200 7400
rect 6000 7364 6004 7396
rect 6036 7364 6164 7396
rect 6196 7364 6200 7396
rect 6000 7360 6200 7364
rect 4240 7316 4440 7320
rect 4240 7284 4244 7316
rect 4276 7284 4404 7316
rect 4436 7284 4440 7316
rect 4240 7280 4440 7284
rect 4480 7316 4680 7320
rect 4480 7284 4484 7316
rect 4516 7284 4644 7316
rect 4676 7284 4680 7316
rect 4480 7280 4680 7284
rect 4720 7316 5720 7320
rect 4720 7284 4724 7316
rect 4756 7284 4884 7316
rect 4916 7284 5044 7316
rect 5076 7284 5204 7316
rect 5236 7284 5364 7316
rect 5396 7284 5524 7316
rect 5556 7284 5684 7316
rect 5716 7284 5720 7316
rect 4720 7280 5720 7284
rect 5760 7316 5960 7320
rect 5760 7284 5764 7316
rect 5796 7284 5924 7316
rect 5956 7284 5960 7316
rect 5760 7280 5960 7284
rect 6000 7316 6200 7320
rect 6000 7284 6004 7316
rect 6036 7284 6164 7316
rect 6196 7284 6200 7316
rect 6000 7280 6200 7284
rect 4240 7236 4440 7240
rect 4240 7204 4244 7236
rect 4276 7204 4404 7236
rect 4436 7204 4440 7236
rect 4240 7200 4440 7204
rect 4480 7236 4680 7240
rect 4480 7204 4484 7236
rect 4516 7204 4644 7236
rect 4676 7204 4680 7236
rect 4480 7200 4680 7204
rect 4720 7236 5720 7240
rect 4720 7204 4724 7236
rect 4756 7204 4884 7236
rect 4916 7204 5044 7236
rect 5076 7204 5204 7236
rect 5236 7204 5364 7236
rect 5396 7204 5524 7236
rect 5556 7204 5684 7236
rect 5716 7204 5720 7236
rect 4720 7200 5720 7204
rect 5760 7236 5960 7240
rect 5760 7204 5764 7236
rect 5796 7204 5924 7236
rect 5956 7204 5960 7236
rect 5760 7200 5960 7204
rect 6000 7236 6200 7240
rect 6000 7204 6004 7236
rect 6036 7204 6164 7236
rect 6196 7204 6200 7236
rect 6000 7200 6200 7204
rect 4240 7156 4440 7160
rect 4240 7124 4244 7156
rect 4276 7124 4404 7156
rect 4436 7124 4440 7156
rect 4240 7120 4440 7124
rect 4480 7156 4680 7160
rect 4480 7124 4484 7156
rect 4516 7124 4644 7156
rect 4676 7124 4680 7156
rect 4480 7120 4680 7124
rect 4720 7156 5720 7160
rect 4720 7124 4724 7156
rect 4756 7124 4884 7156
rect 4916 7124 5044 7156
rect 5076 7124 5204 7156
rect 5236 7124 5364 7156
rect 5396 7124 5524 7156
rect 5556 7124 5684 7156
rect 5716 7124 5720 7156
rect 4720 7120 5720 7124
rect 5760 7156 5960 7160
rect 5760 7124 5764 7156
rect 5796 7124 5924 7156
rect 5956 7124 5960 7156
rect 5760 7120 5960 7124
rect 6000 7156 6200 7160
rect 6000 7124 6004 7156
rect 6036 7124 6164 7156
rect 6196 7124 6200 7156
rect 6000 7120 6200 7124
rect 4240 7076 4440 7080
rect 4240 7044 4244 7076
rect 4276 7044 4404 7076
rect 4436 7044 4440 7076
rect 4240 7040 4440 7044
rect 4480 7076 4680 7080
rect 4480 7044 4484 7076
rect 4516 7044 4644 7076
rect 4676 7044 4680 7076
rect 4480 7040 4680 7044
rect 4720 7076 5720 7080
rect 4720 7044 4724 7076
rect 4756 7044 4884 7076
rect 4916 7044 5044 7076
rect 5076 7044 5204 7076
rect 5236 7044 5364 7076
rect 5396 7044 5524 7076
rect 5556 7044 5684 7076
rect 5716 7044 5720 7076
rect 4720 7040 5720 7044
rect 5760 7076 5960 7080
rect 5760 7044 5764 7076
rect 5796 7044 5924 7076
rect 5956 7044 5960 7076
rect 5760 7040 5960 7044
rect 6000 7076 6200 7080
rect 6000 7044 6004 7076
rect 6036 7044 6164 7076
rect 6196 7044 6200 7076
rect 6000 7040 6200 7044
rect 4240 6996 4440 7000
rect 4240 6964 4244 6996
rect 4276 6964 4404 6996
rect 4436 6964 4440 6996
rect 4240 6960 4440 6964
rect 4480 6996 4680 7000
rect 4480 6964 4484 6996
rect 4516 6964 4644 6996
rect 4676 6964 4680 6996
rect 4480 6960 4680 6964
rect 4720 6996 5720 7000
rect 4720 6964 4724 6996
rect 4756 6964 4884 6996
rect 4916 6964 5044 6996
rect 5076 6964 5204 6996
rect 5236 6964 5364 6996
rect 5396 6964 5524 6996
rect 5556 6964 5684 6996
rect 5716 6964 5720 6996
rect 4720 6960 5720 6964
rect 5760 6996 5960 7000
rect 5760 6964 5764 6996
rect 5796 6964 5924 6996
rect 5956 6964 5960 6996
rect 5760 6960 5960 6964
rect 6000 6996 6200 7000
rect 6000 6964 6004 6996
rect 6036 6964 6164 6996
rect 6196 6964 6200 6996
rect 6000 6960 6200 6964
rect 4240 6916 4440 6920
rect 4240 6884 4244 6916
rect 4276 6884 4404 6916
rect 4436 6884 4440 6916
rect 4240 6880 4440 6884
rect 4480 6916 4680 6920
rect 4480 6884 4484 6916
rect 4516 6884 4644 6916
rect 4676 6884 4680 6916
rect 4480 6880 4680 6884
rect 4720 6916 5720 6920
rect 4720 6884 4724 6916
rect 4756 6884 4884 6916
rect 4916 6884 5044 6916
rect 5076 6884 5204 6916
rect 5236 6884 5364 6916
rect 5396 6884 5524 6916
rect 5556 6884 5684 6916
rect 5716 6884 5720 6916
rect 4720 6880 5720 6884
rect 5760 6916 5960 6920
rect 5760 6884 5764 6916
rect 5796 6884 5924 6916
rect 5956 6884 5960 6916
rect 5760 6880 5960 6884
rect 6000 6916 6200 6920
rect 6000 6884 6004 6916
rect 6036 6884 6164 6916
rect 6196 6884 6200 6916
rect 6000 6880 6200 6884
rect 4240 6836 4440 6840
rect 4240 6804 4244 6836
rect 4276 6804 4404 6836
rect 4436 6804 4440 6836
rect 4240 6800 4440 6804
rect 4480 6836 4680 6840
rect 4480 6804 4484 6836
rect 4516 6804 4644 6836
rect 4676 6804 4680 6836
rect 4480 6800 4680 6804
rect 4720 6836 5720 6840
rect 4720 6804 4724 6836
rect 4756 6804 4884 6836
rect 4916 6804 5044 6836
rect 5076 6804 5204 6836
rect 5236 6804 5364 6836
rect 5396 6804 5524 6836
rect 5556 6804 5684 6836
rect 5716 6804 5720 6836
rect 4720 6800 5720 6804
rect 5760 6836 5960 6840
rect 5760 6804 5764 6836
rect 5796 6804 5924 6836
rect 5956 6804 5960 6836
rect 5760 6800 5960 6804
rect 6000 6836 6200 6840
rect 6000 6804 6004 6836
rect 6036 6804 6164 6836
rect 6196 6804 6200 6836
rect 6000 6800 6200 6804
rect 4240 6756 4440 6760
rect 4240 6724 4244 6756
rect 4276 6724 4404 6756
rect 4436 6724 4440 6756
rect 4240 6720 4440 6724
rect 4480 6756 4680 6760
rect 4480 6724 4484 6756
rect 4516 6724 4644 6756
rect 4676 6724 4680 6756
rect 4480 6720 4680 6724
rect 4720 6756 5720 6760
rect 4720 6724 4724 6756
rect 4756 6724 4884 6756
rect 4916 6724 5044 6756
rect 5076 6724 5204 6756
rect 5236 6724 5364 6756
rect 5396 6724 5524 6756
rect 5556 6724 5684 6756
rect 5716 6724 5720 6756
rect 4720 6720 5720 6724
rect 5760 6756 5960 6760
rect 5760 6724 5764 6756
rect 5796 6724 5924 6756
rect 5956 6724 5960 6756
rect 5760 6720 5960 6724
rect 6000 6756 6200 6760
rect 6000 6724 6004 6756
rect 6036 6724 6164 6756
rect 6196 6724 6200 6756
rect 6000 6720 6200 6724
rect 4240 6676 4440 6680
rect 4240 6644 4244 6676
rect 4276 6644 4404 6676
rect 4436 6644 4440 6676
rect 4240 6640 4440 6644
rect 4480 6676 4680 6680
rect 4480 6644 4484 6676
rect 4516 6644 4644 6676
rect 4676 6644 4680 6676
rect 4480 6640 4680 6644
rect 4720 6676 5720 6680
rect 4720 6644 4724 6676
rect 4756 6644 4884 6676
rect 4916 6644 5044 6676
rect 5076 6644 5204 6676
rect 5236 6644 5364 6676
rect 5396 6644 5524 6676
rect 5556 6644 5684 6676
rect 5716 6644 5720 6676
rect 4720 6640 5720 6644
rect 5760 6676 5960 6680
rect 5760 6644 5764 6676
rect 5796 6644 5924 6676
rect 5956 6644 5960 6676
rect 5760 6640 5960 6644
rect 6000 6676 6200 6680
rect 6000 6644 6004 6676
rect 6036 6644 6164 6676
rect 6196 6644 6200 6676
rect 6000 6640 6200 6644
rect 4240 6596 4440 6600
rect 4240 6564 4244 6596
rect 4276 6564 4404 6596
rect 4436 6564 4440 6596
rect 4240 6560 4440 6564
rect 4480 6596 4680 6600
rect 4480 6564 4484 6596
rect 4516 6564 4644 6596
rect 4676 6564 4680 6596
rect 4480 6560 4680 6564
rect 4720 6596 5720 6600
rect 4720 6564 4724 6596
rect 4756 6564 4884 6596
rect 4916 6564 5044 6596
rect 5076 6564 5204 6596
rect 5236 6564 5364 6596
rect 5396 6564 5524 6596
rect 5556 6564 5684 6596
rect 5716 6564 5720 6596
rect 4720 6560 5720 6564
rect 5760 6596 5960 6600
rect 5760 6564 5764 6596
rect 5796 6564 5924 6596
rect 5956 6564 5960 6596
rect 5760 6560 5960 6564
rect 6000 6596 6200 6600
rect 6000 6564 6004 6596
rect 6036 6564 6164 6596
rect 6196 6564 6200 6596
rect 6000 6560 6200 6564
rect 4240 6516 4440 6520
rect 4240 6484 4244 6516
rect 4276 6484 4404 6516
rect 4436 6484 4440 6516
rect 4240 6480 4440 6484
rect 4480 6516 4680 6520
rect 4480 6484 4484 6516
rect 4516 6484 4644 6516
rect 4676 6484 4680 6516
rect 4480 6480 4680 6484
rect 4720 6516 5720 6520
rect 4720 6484 4724 6516
rect 4756 6484 4884 6516
rect 4916 6484 5044 6516
rect 5076 6484 5204 6516
rect 5236 6484 5364 6516
rect 5396 6484 5524 6516
rect 5556 6484 5684 6516
rect 5716 6484 5720 6516
rect 4720 6480 5720 6484
rect 5760 6516 5960 6520
rect 5760 6484 5764 6516
rect 5796 6484 5924 6516
rect 5956 6484 5960 6516
rect 5760 6480 5960 6484
rect 6000 6516 6200 6520
rect 6000 6484 6004 6516
rect 6036 6484 6164 6516
rect 6196 6484 6200 6516
rect 6000 6480 6200 6484
rect 4240 6436 4440 6440
rect 4240 6404 4244 6436
rect 4276 6404 4404 6436
rect 4436 6404 4440 6436
rect 4240 6400 4440 6404
rect 4480 6436 4680 6440
rect 4480 6404 4484 6436
rect 4516 6404 4644 6436
rect 4676 6404 4680 6436
rect 4480 6400 4680 6404
rect 4720 6436 5720 6440
rect 4720 6404 4724 6436
rect 4756 6404 4884 6436
rect 4916 6404 5044 6436
rect 5076 6404 5204 6436
rect 5236 6404 5364 6436
rect 5396 6404 5524 6436
rect 5556 6404 5684 6436
rect 5716 6404 5720 6436
rect 4720 6400 5720 6404
rect 5760 6436 5960 6440
rect 5760 6404 5764 6436
rect 5796 6404 5924 6436
rect 5956 6404 5960 6436
rect 5760 6400 5960 6404
rect 6000 6436 6200 6440
rect 6000 6404 6004 6436
rect 6036 6404 6164 6436
rect 6196 6404 6200 6436
rect 6000 6400 6200 6404
rect 4240 6356 4440 6360
rect 4240 6324 4244 6356
rect 4276 6324 4404 6356
rect 4436 6324 4440 6356
rect 4240 6320 4440 6324
rect 4480 6356 4680 6360
rect 4480 6324 4484 6356
rect 4516 6324 4644 6356
rect 4676 6324 4680 6356
rect 4480 6320 4680 6324
rect 4720 6356 5720 6360
rect 4720 6324 4724 6356
rect 4756 6324 4884 6356
rect 4916 6324 5044 6356
rect 5076 6324 5204 6356
rect 5236 6324 5364 6356
rect 5396 6324 5524 6356
rect 5556 6324 5684 6356
rect 5716 6324 5720 6356
rect 4720 6320 5720 6324
rect 5760 6356 5960 6360
rect 5760 6324 5764 6356
rect 5796 6324 5924 6356
rect 5956 6324 5960 6356
rect 5760 6320 5960 6324
rect 6000 6356 6200 6360
rect 6000 6324 6004 6356
rect 6036 6324 6164 6356
rect 6196 6324 6200 6356
rect 6000 6320 6200 6324
rect 4240 6276 4440 6280
rect 4240 6244 4244 6276
rect 4276 6244 4404 6276
rect 4436 6244 4440 6276
rect 4240 6240 4440 6244
rect 4480 6276 4680 6280
rect 4480 6244 4484 6276
rect 4516 6244 4644 6276
rect 4676 6244 4680 6276
rect 4480 6240 4680 6244
rect 4720 6276 5720 6280
rect 4720 6244 4724 6276
rect 4756 6244 4884 6276
rect 4916 6244 5044 6276
rect 5076 6244 5204 6276
rect 5236 6244 5364 6276
rect 5396 6244 5524 6276
rect 5556 6244 5684 6276
rect 5716 6244 5720 6276
rect 4720 6240 5720 6244
rect 5760 6276 5960 6280
rect 5760 6244 5764 6276
rect 5796 6244 5924 6276
rect 5956 6244 5960 6276
rect 5760 6240 5960 6244
rect 6000 6276 6200 6280
rect 6000 6244 6004 6276
rect 6036 6244 6164 6276
rect 6196 6244 6200 6276
rect 6000 6240 6200 6244
rect 4240 6196 4440 6200
rect 4240 6164 4244 6196
rect 4276 6164 4404 6196
rect 4436 6164 4440 6196
rect 4240 6160 4440 6164
rect 4480 6196 4680 6200
rect 4480 6164 4484 6196
rect 4516 6164 4644 6196
rect 4676 6164 4680 6196
rect 4480 6160 4680 6164
rect 4720 6196 5720 6200
rect 4720 6164 4724 6196
rect 4756 6164 4884 6196
rect 4916 6164 5044 6196
rect 5076 6164 5204 6196
rect 5236 6164 5364 6196
rect 5396 6164 5524 6196
rect 5556 6164 5684 6196
rect 5716 6164 5720 6196
rect 4720 6160 5720 6164
rect 5760 6196 5960 6200
rect 5760 6164 5764 6196
rect 5796 6164 5924 6196
rect 5956 6164 5960 6196
rect 5760 6160 5960 6164
rect 6000 6196 6200 6200
rect 6000 6164 6004 6196
rect 6036 6164 6164 6196
rect 6196 6164 6200 6196
rect 6000 6160 6200 6164
rect 4240 6116 4440 6120
rect 4240 6084 4244 6116
rect 4276 6084 4404 6116
rect 4436 6084 4440 6116
rect 4240 6080 4440 6084
rect 4480 6116 4680 6120
rect 4480 6084 4484 6116
rect 4516 6084 4644 6116
rect 4676 6084 4680 6116
rect 4480 6080 4680 6084
rect 4720 6116 5720 6120
rect 4720 6084 4724 6116
rect 4756 6084 4884 6116
rect 4916 6084 5044 6116
rect 5076 6084 5204 6116
rect 5236 6084 5364 6116
rect 5396 6084 5524 6116
rect 5556 6084 5684 6116
rect 5716 6084 5720 6116
rect 4720 6080 5720 6084
rect 5760 6116 5960 6120
rect 5760 6084 5764 6116
rect 5796 6084 5924 6116
rect 5956 6084 5960 6116
rect 5760 6080 5960 6084
rect 6000 6116 6200 6120
rect 6000 6084 6004 6116
rect 6036 6084 6164 6116
rect 6196 6084 6200 6116
rect 6000 6080 6200 6084
rect 4240 6036 4440 6040
rect 4240 6004 4244 6036
rect 4276 6004 4404 6036
rect 4436 6004 4440 6036
rect 4240 6000 4440 6004
rect 4480 6036 4680 6040
rect 4480 6004 4484 6036
rect 4516 6004 4644 6036
rect 4676 6004 4680 6036
rect 4480 6000 4680 6004
rect 4720 6036 5720 6040
rect 4720 6004 4724 6036
rect 4756 6004 4884 6036
rect 4916 6004 5044 6036
rect 5076 6004 5204 6036
rect 5236 6004 5364 6036
rect 5396 6004 5524 6036
rect 5556 6004 5684 6036
rect 5716 6004 5720 6036
rect 4720 6000 5720 6004
rect 5760 6036 5960 6040
rect 5760 6004 5764 6036
rect 5796 6004 5924 6036
rect 5956 6004 5960 6036
rect 5760 6000 5960 6004
rect 6000 6036 6200 6040
rect 6000 6004 6004 6036
rect 6036 6004 6164 6036
rect 6196 6004 6200 6036
rect 6000 6000 6200 6004
rect 4240 5956 4440 5960
rect 4240 5924 4244 5956
rect 4276 5924 4404 5956
rect 4436 5924 4440 5956
rect 4240 5920 4440 5924
rect 4480 5956 4680 5960
rect 4480 5924 4484 5956
rect 4516 5924 4644 5956
rect 4676 5924 4680 5956
rect 4480 5920 4680 5924
rect 4720 5956 5720 5960
rect 4720 5924 4724 5956
rect 4756 5924 4884 5956
rect 4916 5924 5044 5956
rect 5076 5924 5204 5956
rect 5236 5924 5364 5956
rect 5396 5924 5524 5956
rect 5556 5924 5684 5956
rect 5716 5924 5720 5956
rect 4720 5920 5720 5924
rect 5760 5956 5960 5960
rect 5760 5924 5764 5956
rect 5796 5924 5924 5956
rect 5956 5924 5960 5956
rect 5760 5920 5960 5924
rect 6000 5956 6200 5960
rect 6000 5924 6004 5956
rect 6036 5924 6164 5956
rect 6196 5924 6200 5956
rect 6000 5920 6200 5924
rect 4240 5876 4440 5880
rect 4240 5844 4244 5876
rect 4276 5844 4404 5876
rect 4436 5844 4440 5876
rect 4240 5840 4440 5844
rect 4480 5876 4680 5880
rect 4480 5844 4484 5876
rect 4516 5844 4644 5876
rect 4676 5844 4680 5876
rect 4480 5840 4680 5844
rect 4720 5876 5720 5880
rect 4720 5844 4724 5876
rect 4756 5844 4884 5876
rect 4916 5844 5044 5876
rect 5076 5844 5204 5876
rect 5236 5844 5364 5876
rect 5396 5844 5524 5876
rect 5556 5844 5684 5876
rect 5716 5844 5720 5876
rect 4720 5840 5720 5844
rect 5760 5876 5960 5880
rect 5760 5844 5764 5876
rect 5796 5844 5924 5876
rect 5956 5844 5960 5876
rect 5760 5840 5960 5844
rect 6000 5876 6200 5880
rect 6000 5844 6004 5876
rect 6036 5844 6164 5876
rect 6196 5844 6200 5876
rect 6000 5840 6200 5844
rect 4240 5796 4440 5800
rect 4240 5764 4244 5796
rect 4276 5764 4404 5796
rect 4436 5764 4440 5796
rect 4240 5760 4440 5764
rect 4480 5796 4680 5800
rect 4480 5764 4484 5796
rect 4516 5764 4644 5796
rect 4676 5764 4680 5796
rect 4480 5760 4680 5764
rect 4720 5796 5720 5800
rect 4720 5764 4724 5796
rect 4756 5764 4884 5796
rect 4916 5764 5044 5796
rect 5076 5764 5204 5796
rect 5236 5764 5364 5796
rect 5396 5764 5524 5796
rect 5556 5764 5684 5796
rect 5716 5764 5720 5796
rect 4720 5760 5720 5764
rect 5760 5796 5960 5800
rect 5760 5764 5764 5796
rect 5796 5764 5924 5796
rect 5956 5764 5960 5796
rect 5760 5760 5960 5764
rect 6000 5796 6200 5800
rect 6000 5764 6004 5796
rect 6036 5764 6164 5796
rect 6196 5764 6200 5796
rect 6000 5760 6200 5764
rect 4240 5716 4440 5720
rect 4240 5684 4244 5716
rect 4276 5684 4404 5716
rect 4436 5684 4440 5716
rect 4240 5680 4440 5684
rect 4480 5716 4680 5720
rect 4480 5684 4484 5716
rect 4516 5684 4644 5716
rect 4676 5684 4680 5716
rect 4480 5680 4680 5684
rect 4720 5716 5720 5720
rect 4720 5684 4724 5716
rect 4756 5684 4884 5716
rect 4916 5684 5044 5716
rect 5076 5684 5204 5716
rect 5236 5684 5364 5716
rect 5396 5684 5524 5716
rect 5556 5684 5684 5716
rect 5716 5684 5720 5716
rect 4720 5680 5720 5684
rect 5760 5716 5960 5720
rect 5760 5684 5764 5716
rect 5796 5684 5924 5716
rect 5956 5684 5960 5716
rect 5760 5680 5960 5684
rect 6000 5716 6200 5720
rect 6000 5684 6004 5716
rect 6036 5684 6164 5716
rect 6196 5684 6200 5716
rect 6000 5680 6200 5684
rect 4240 5636 4440 5640
rect 4240 5604 4244 5636
rect 4276 5604 4404 5636
rect 4436 5604 4440 5636
rect 4240 5600 4440 5604
rect 4480 5636 4680 5640
rect 4480 5604 4484 5636
rect 4516 5604 4644 5636
rect 4676 5604 4680 5636
rect 4480 5600 4680 5604
rect 4720 5636 5720 5640
rect 4720 5604 4724 5636
rect 4756 5604 4884 5636
rect 4916 5604 5044 5636
rect 5076 5604 5204 5636
rect 5236 5604 5364 5636
rect 5396 5604 5524 5636
rect 5556 5604 5684 5636
rect 5716 5604 5720 5636
rect 4720 5600 5720 5604
rect 5760 5636 5960 5640
rect 5760 5604 5764 5636
rect 5796 5604 5924 5636
rect 5956 5604 5960 5636
rect 5760 5600 5960 5604
rect 6000 5636 6200 5640
rect 6000 5604 6004 5636
rect 6036 5604 6164 5636
rect 6196 5604 6200 5636
rect 6000 5600 6200 5604
rect 4240 5556 4440 5560
rect 4240 5524 4244 5556
rect 4276 5524 4404 5556
rect 4436 5524 4440 5556
rect 4240 5520 4440 5524
rect 4480 5556 4680 5560
rect 4480 5524 4484 5556
rect 4516 5524 4644 5556
rect 4676 5524 4680 5556
rect 4480 5520 4680 5524
rect 4720 5556 5720 5560
rect 4720 5524 4724 5556
rect 4756 5524 4884 5556
rect 4916 5524 5044 5556
rect 5076 5524 5204 5556
rect 5236 5524 5364 5556
rect 5396 5524 5524 5556
rect 5556 5524 5684 5556
rect 5716 5524 5720 5556
rect 4720 5520 5720 5524
rect 5760 5556 5960 5560
rect 5760 5524 5764 5556
rect 5796 5524 5924 5556
rect 5956 5524 5960 5556
rect 5760 5520 5960 5524
rect 6000 5556 6200 5560
rect 6000 5524 6004 5556
rect 6036 5524 6164 5556
rect 6196 5524 6200 5556
rect 6000 5520 6200 5524
rect 4240 5476 4440 5480
rect 4240 5444 4244 5476
rect 4276 5444 4404 5476
rect 4436 5444 4440 5476
rect 4240 5440 4440 5444
rect 4480 5476 4680 5480
rect 4480 5444 4484 5476
rect 4516 5444 4644 5476
rect 4676 5444 4680 5476
rect 4480 5440 4680 5444
rect 4720 5476 5720 5480
rect 4720 5444 4724 5476
rect 4756 5444 4884 5476
rect 4916 5444 5044 5476
rect 5076 5444 5204 5476
rect 5236 5444 5364 5476
rect 5396 5444 5524 5476
rect 5556 5444 5684 5476
rect 5716 5444 5720 5476
rect 4720 5440 5720 5444
rect 5760 5476 5960 5480
rect 5760 5444 5764 5476
rect 5796 5444 5924 5476
rect 5956 5444 5960 5476
rect 5760 5440 5960 5444
rect 6000 5476 6200 5480
rect 6000 5444 6004 5476
rect 6036 5444 6164 5476
rect 6196 5444 6200 5476
rect 6000 5440 6200 5444
rect 4240 5396 4440 5400
rect 4240 5364 4244 5396
rect 4276 5364 4404 5396
rect 4436 5364 4440 5396
rect 4240 5360 4440 5364
rect 4480 5396 4680 5400
rect 4480 5364 4484 5396
rect 4516 5364 4644 5396
rect 4676 5364 4680 5396
rect 4480 5360 4680 5364
rect 4720 5396 5720 5400
rect 4720 5364 4724 5396
rect 4756 5364 4884 5396
rect 4916 5364 5044 5396
rect 5076 5364 5204 5396
rect 5236 5364 5364 5396
rect 5396 5364 5524 5396
rect 5556 5364 5684 5396
rect 5716 5364 5720 5396
rect 4720 5360 5720 5364
rect 5760 5396 5960 5400
rect 5760 5364 5764 5396
rect 5796 5364 5924 5396
rect 5956 5364 5960 5396
rect 5760 5360 5960 5364
rect 6000 5396 6200 5400
rect 6000 5364 6004 5396
rect 6036 5364 6164 5396
rect 6196 5364 6200 5396
rect 6000 5360 6200 5364
rect 4240 5316 4440 5320
rect 4240 5284 4244 5316
rect 4276 5284 4404 5316
rect 4436 5284 4440 5316
rect 4240 5280 4440 5284
rect 4480 5316 4680 5320
rect 4480 5284 4484 5316
rect 4516 5284 4644 5316
rect 4676 5284 4680 5316
rect 4480 5280 4680 5284
rect 4720 5316 5720 5320
rect 4720 5284 4724 5316
rect 4756 5284 4884 5316
rect 4916 5284 5044 5316
rect 5076 5284 5204 5316
rect 5236 5284 5364 5316
rect 5396 5284 5524 5316
rect 5556 5284 5684 5316
rect 5716 5284 5720 5316
rect 4720 5280 5720 5284
rect 5760 5316 5960 5320
rect 5760 5284 5764 5316
rect 5796 5284 5924 5316
rect 5956 5284 5960 5316
rect 5760 5280 5960 5284
rect 6000 5316 6200 5320
rect 6000 5284 6004 5316
rect 6036 5284 6164 5316
rect 6196 5284 6200 5316
rect 6000 5280 6200 5284
rect 4240 5236 4440 5240
rect 4240 5204 4244 5236
rect 4276 5204 4404 5236
rect 4436 5204 4440 5236
rect 4240 5200 4440 5204
rect 4480 5236 4680 5240
rect 4480 5204 4484 5236
rect 4516 5204 4644 5236
rect 4676 5204 4680 5236
rect 4480 5200 4680 5204
rect 4720 5236 5720 5240
rect 4720 5204 4724 5236
rect 4756 5204 4884 5236
rect 4916 5204 5044 5236
rect 5076 5204 5204 5236
rect 5236 5204 5364 5236
rect 5396 5204 5524 5236
rect 5556 5204 5684 5236
rect 5716 5204 5720 5236
rect 4720 5200 5720 5204
rect 5760 5236 5960 5240
rect 5760 5204 5764 5236
rect 5796 5204 5924 5236
rect 5956 5204 5960 5236
rect 5760 5200 5960 5204
rect 6000 5236 6200 5240
rect 6000 5204 6004 5236
rect 6036 5204 6164 5236
rect 6196 5204 6200 5236
rect 6000 5200 6200 5204
rect 4240 5156 4440 5160
rect 4240 5124 4244 5156
rect 4276 5124 4404 5156
rect 4436 5124 4440 5156
rect 4240 5120 4440 5124
rect 4480 5156 4680 5160
rect 4480 5124 4484 5156
rect 4516 5124 4644 5156
rect 4676 5124 4680 5156
rect 4480 5120 4680 5124
rect 4720 5156 5720 5160
rect 4720 5124 4724 5156
rect 4756 5124 4884 5156
rect 4916 5124 5044 5156
rect 5076 5124 5204 5156
rect 5236 5124 5364 5156
rect 5396 5124 5524 5156
rect 5556 5124 5684 5156
rect 5716 5124 5720 5156
rect 4720 5120 5720 5124
rect 5760 5156 5960 5160
rect 5760 5124 5764 5156
rect 5796 5124 5924 5156
rect 5956 5124 5960 5156
rect 5760 5120 5960 5124
rect 6000 5156 6200 5160
rect 6000 5124 6004 5156
rect 6036 5124 6164 5156
rect 6196 5124 6200 5156
rect 6000 5120 6200 5124
rect 4240 5076 4440 5080
rect 4240 5044 4244 5076
rect 4276 5044 4404 5076
rect 4436 5044 4440 5076
rect 4240 5040 4440 5044
rect 4480 5076 4680 5080
rect 4480 5044 4484 5076
rect 4516 5044 4644 5076
rect 4676 5044 4680 5076
rect 4480 5040 4680 5044
rect 4720 5076 5720 5080
rect 4720 5044 4724 5076
rect 4756 5044 4884 5076
rect 4916 5044 5044 5076
rect 5076 5044 5204 5076
rect 5236 5044 5364 5076
rect 5396 5044 5524 5076
rect 5556 5044 5684 5076
rect 5716 5044 5720 5076
rect 4720 5040 5720 5044
rect 5760 5076 5960 5080
rect 5760 5044 5764 5076
rect 5796 5044 5924 5076
rect 5956 5044 5960 5076
rect 5760 5040 5960 5044
rect 6000 5076 6200 5080
rect 6000 5044 6004 5076
rect 6036 5044 6164 5076
rect 6196 5044 6200 5076
rect 6000 5040 6200 5044
rect 4240 4996 4440 5000
rect 4240 4964 4244 4996
rect 4276 4964 4404 4996
rect 4436 4964 4440 4996
rect 4240 4960 4440 4964
rect 4480 4996 4680 5000
rect 4480 4964 4484 4996
rect 4516 4964 4644 4996
rect 4676 4964 4680 4996
rect 4480 4960 4680 4964
rect 4720 4996 5720 5000
rect 4720 4964 4724 4996
rect 4756 4964 4884 4996
rect 4916 4964 5044 4996
rect 5076 4964 5204 4996
rect 5236 4964 5364 4996
rect 5396 4964 5524 4996
rect 5556 4964 5684 4996
rect 5716 4964 5720 4996
rect 4720 4960 5720 4964
rect 5760 4996 5960 5000
rect 5760 4964 5764 4996
rect 5796 4964 5924 4996
rect 5956 4964 5960 4996
rect 5760 4960 5960 4964
rect 6000 4996 6200 5000
rect 6000 4964 6004 4996
rect 6036 4964 6164 4996
rect 6196 4964 6200 4996
rect 6000 4960 6200 4964
rect 4240 4916 4440 4920
rect 4240 4884 4244 4916
rect 4276 4884 4404 4916
rect 4436 4884 4440 4916
rect 4240 4880 4440 4884
rect 4480 4916 4680 4920
rect 4480 4884 4484 4916
rect 4516 4884 4644 4916
rect 4676 4884 4680 4916
rect 4480 4880 4680 4884
rect 4720 4916 5720 4920
rect 4720 4884 4724 4916
rect 4756 4884 4884 4916
rect 4916 4884 5044 4916
rect 5076 4884 5204 4916
rect 5236 4884 5364 4916
rect 5396 4884 5524 4916
rect 5556 4884 5684 4916
rect 5716 4884 5720 4916
rect 4720 4880 5720 4884
rect 5760 4916 5960 4920
rect 5760 4884 5764 4916
rect 5796 4884 5924 4916
rect 5956 4884 5960 4916
rect 5760 4880 5960 4884
rect 6000 4916 6200 4920
rect 6000 4884 6004 4916
rect 6036 4884 6164 4916
rect 6196 4884 6200 4916
rect 6000 4880 6200 4884
rect 4240 4836 4440 4840
rect 4240 4804 4244 4836
rect 4276 4804 4404 4836
rect 4436 4804 4440 4836
rect 4240 4800 4440 4804
rect 4480 4836 4680 4840
rect 4480 4804 4484 4836
rect 4516 4804 4644 4836
rect 4676 4804 4680 4836
rect 4480 4800 4680 4804
rect 4720 4836 5720 4840
rect 4720 4804 4724 4836
rect 4756 4804 4884 4836
rect 4916 4804 5044 4836
rect 5076 4804 5204 4836
rect 5236 4804 5364 4836
rect 5396 4804 5524 4836
rect 5556 4804 5684 4836
rect 5716 4804 5720 4836
rect 4720 4800 5720 4804
rect 5760 4836 5960 4840
rect 5760 4804 5764 4836
rect 5796 4804 5924 4836
rect 5956 4804 5960 4836
rect 5760 4800 5960 4804
rect 6000 4836 6200 4840
rect 6000 4804 6004 4836
rect 6036 4804 6164 4836
rect 6196 4804 6200 4836
rect 6000 4800 6200 4804
rect 4240 4756 4440 4760
rect 4240 4724 4244 4756
rect 4276 4724 4404 4756
rect 4436 4724 4440 4756
rect 4240 4720 4440 4724
rect 4480 4756 4680 4760
rect 4480 4724 4484 4756
rect 4516 4724 4644 4756
rect 4676 4724 4680 4756
rect 4480 4720 4680 4724
rect 4720 4756 5720 4760
rect 4720 4724 4724 4756
rect 4756 4724 4884 4756
rect 4916 4724 5044 4756
rect 5076 4724 5204 4756
rect 5236 4724 5364 4756
rect 5396 4724 5524 4756
rect 5556 4724 5684 4756
rect 5716 4724 5720 4756
rect 4720 4720 5720 4724
rect 5760 4756 5960 4760
rect 5760 4724 5764 4756
rect 5796 4724 5924 4756
rect 5956 4724 5960 4756
rect 5760 4720 5960 4724
rect 6000 4756 6200 4760
rect 6000 4724 6004 4756
rect 6036 4724 6164 4756
rect 6196 4724 6200 4756
rect 6000 4720 6200 4724
rect 4240 4676 4440 4680
rect 4240 4644 4244 4676
rect 4276 4644 4404 4676
rect 4436 4644 4440 4676
rect 4240 4640 4440 4644
rect 4480 4676 4680 4680
rect 4480 4644 4484 4676
rect 4516 4644 4644 4676
rect 4676 4644 4680 4676
rect 4480 4640 4680 4644
rect 4720 4676 5720 4680
rect 4720 4644 4724 4676
rect 4756 4644 4884 4676
rect 4916 4644 5044 4676
rect 5076 4644 5204 4676
rect 5236 4644 5364 4676
rect 5396 4644 5524 4676
rect 5556 4644 5684 4676
rect 5716 4644 5720 4676
rect 4720 4640 5720 4644
rect 5760 4676 5960 4680
rect 5760 4644 5764 4676
rect 5796 4644 5924 4676
rect 5956 4644 5960 4676
rect 5760 4640 5960 4644
rect 6000 4676 6200 4680
rect 6000 4644 6004 4676
rect 6036 4644 6164 4676
rect 6196 4644 6200 4676
rect 6000 4640 6200 4644
rect 4240 4596 4440 4600
rect 4240 4564 4244 4596
rect 4276 4564 4404 4596
rect 4436 4564 4440 4596
rect 4240 4560 4440 4564
rect 4480 4596 4680 4600
rect 4480 4564 4484 4596
rect 4516 4564 4644 4596
rect 4676 4564 4680 4596
rect 4480 4560 4680 4564
rect 4720 4596 5720 4600
rect 4720 4564 4724 4596
rect 4756 4564 4884 4596
rect 4916 4564 5044 4596
rect 5076 4564 5204 4596
rect 5236 4564 5364 4596
rect 5396 4564 5524 4596
rect 5556 4564 5684 4596
rect 5716 4564 5720 4596
rect 4720 4560 5720 4564
rect 5760 4596 5960 4600
rect 5760 4564 5764 4596
rect 5796 4564 5924 4596
rect 5956 4564 5960 4596
rect 5760 4560 5960 4564
rect 6000 4596 6200 4600
rect 6000 4564 6004 4596
rect 6036 4564 6164 4596
rect 6196 4564 6200 4596
rect 6000 4560 6200 4564
rect 4240 4516 4440 4520
rect 4240 4484 4244 4516
rect 4276 4484 4404 4516
rect 4436 4484 4440 4516
rect 4240 4480 4440 4484
rect 4480 4516 4680 4520
rect 4480 4484 4484 4516
rect 4516 4484 4644 4516
rect 4676 4484 4680 4516
rect 4480 4480 4680 4484
rect 4720 4516 5720 4520
rect 4720 4484 4724 4516
rect 4756 4484 4884 4516
rect 4916 4484 5044 4516
rect 5076 4484 5204 4516
rect 5236 4484 5364 4516
rect 5396 4484 5524 4516
rect 5556 4484 5684 4516
rect 5716 4484 5720 4516
rect 4720 4480 5720 4484
rect 5760 4516 5960 4520
rect 5760 4484 5764 4516
rect 5796 4484 5924 4516
rect 5956 4484 5960 4516
rect 5760 4480 5960 4484
rect 6000 4516 6200 4520
rect 6000 4484 6004 4516
rect 6036 4484 6164 4516
rect 6196 4484 6200 4516
rect 6000 4480 6200 4484
rect 4240 4436 4440 4440
rect 4240 4404 4244 4436
rect 4276 4404 4404 4436
rect 4436 4404 4440 4436
rect 4240 4400 4440 4404
rect 4480 4436 4680 4440
rect 4480 4404 4484 4436
rect 4516 4404 4644 4436
rect 4676 4404 4680 4436
rect 4480 4400 4680 4404
rect 4720 4436 5720 4440
rect 4720 4404 4724 4436
rect 4756 4404 4884 4436
rect 4916 4404 5044 4436
rect 5076 4404 5204 4436
rect 5236 4404 5364 4436
rect 5396 4404 5524 4436
rect 5556 4404 5684 4436
rect 5716 4404 5720 4436
rect 4720 4400 5720 4404
rect 5760 4436 5960 4440
rect 5760 4404 5764 4436
rect 5796 4404 5924 4436
rect 5956 4404 5960 4436
rect 5760 4400 5960 4404
rect 6000 4436 6200 4440
rect 6000 4404 6004 4436
rect 6036 4404 6164 4436
rect 6196 4404 6200 4436
rect 6000 4400 6200 4404
rect 4240 4356 4440 4360
rect 4240 4324 4244 4356
rect 4276 4324 4404 4356
rect 4436 4324 4440 4356
rect 4240 4320 4440 4324
rect 4480 4356 4680 4360
rect 4480 4324 4484 4356
rect 4516 4324 4644 4356
rect 4676 4324 4680 4356
rect 4480 4320 4680 4324
rect 4720 4356 5720 4360
rect 4720 4324 4724 4356
rect 4756 4324 4884 4356
rect 4916 4324 5044 4356
rect 5076 4324 5204 4356
rect 5236 4324 5364 4356
rect 5396 4324 5524 4356
rect 5556 4324 5684 4356
rect 5716 4324 5720 4356
rect 4720 4320 5720 4324
rect 5760 4356 5960 4360
rect 5760 4324 5764 4356
rect 5796 4324 5924 4356
rect 5956 4324 5960 4356
rect 5760 4320 5960 4324
rect 6000 4356 6200 4360
rect 6000 4324 6004 4356
rect 6036 4324 6164 4356
rect 6196 4324 6200 4356
rect 6000 4320 6200 4324
rect 4240 4276 4440 4280
rect 4240 4244 4244 4276
rect 4276 4244 4404 4276
rect 4436 4244 4440 4276
rect 4240 4240 4440 4244
rect 4480 4276 4680 4280
rect 4480 4244 4484 4276
rect 4516 4244 4644 4276
rect 4676 4244 4680 4276
rect 4480 4240 4680 4244
rect 4720 4276 5720 4280
rect 4720 4244 4724 4276
rect 4756 4244 4884 4276
rect 4916 4244 5044 4276
rect 5076 4244 5204 4276
rect 5236 4244 5364 4276
rect 5396 4244 5524 4276
rect 5556 4244 5684 4276
rect 5716 4244 5720 4276
rect 4720 4240 5720 4244
rect 5760 4276 5960 4280
rect 5760 4244 5764 4276
rect 5796 4244 5924 4276
rect 5956 4244 5960 4276
rect 5760 4240 5960 4244
rect 6000 4276 6200 4280
rect 6000 4244 6004 4276
rect 6036 4244 6164 4276
rect 6196 4244 6200 4276
rect 6000 4240 6200 4244
rect 4240 4196 4440 4200
rect 4240 4164 4244 4196
rect 4276 4164 4404 4196
rect 4436 4164 4440 4196
rect 4240 4160 4440 4164
rect 4480 4196 4680 4200
rect 4480 4164 4484 4196
rect 4516 4164 4644 4196
rect 4676 4164 4680 4196
rect 4480 4160 4680 4164
rect 4720 4196 5720 4200
rect 4720 4164 4724 4196
rect 4756 4164 4884 4196
rect 4916 4164 5044 4196
rect 5076 4164 5204 4196
rect 5236 4164 5364 4196
rect 5396 4164 5524 4196
rect 5556 4164 5684 4196
rect 5716 4164 5720 4196
rect 4720 4160 5720 4164
rect 5760 4196 5960 4200
rect 5760 4164 5764 4196
rect 5796 4164 5924 4196
rect 5956 4164 5960 4196
rect 5760 4160 5960 4164
rect 6000 4196 6200 4200
rect 6000 4164 6004 4196
rect 6036 4164 6164 4196
rect 6196 4164 6200 4196
rect 6000 4160 6200 4164
rect 4240 4116 4440 4120
rect 4240 4084 4244 4116
rect 4276 4084 4404 4116
rect 4436 4084 4440 4116
rect 4240 4080 4440 4084
rect 4480 4116 4680 4120
rect 4480 4084 4484 4116
rect 4516 4084 4644 4116
rect 4676 4084 4680 4116
rect 4480 4080 4680 4084
rect 4720 4116 5720 4120
rect 4720 4084 4724 4116
rect 4756 4084 4884 4116
rect 4916 4084 5044 4116
rect 5076 4084 5204 4116
rect 5236 4084 5364 4116
rect 5396 4084 5524 4116
rect 5556 4084 5684 4116
rect 5716 4084 5720 4116
rect 4720 4080 5720 4084
rect 5760 4116 5960 4120
rect 5760 4084 5764 4116
rect 5796 4084 5924 4116
rect 5956 4084 5960 4116
rect 5760 4080 5960 4084
rect 6000 4116 6200 4120
rect 6000 4084 6004 4116
rect 6036 4084 6164 4116
rect 6196 4084 6200 4116
rect 6000 4080 6200 4084
rect 4240 4036 4440 4040
rect 4240 4004 4244 4036
rect 4276 4004 4404 4036
rect 4436 4004 4440 4036
rect 4240 4000 4440 4004
rect 4480 4036 4680 4040
rect 4480 4004 4484 4036
rect 4516 4004 4644 4036
rect 4676 4004 4680 4036
rect 4480 4000 4680 4004
rect 4720 4036 5720 4040
rect 4720 4004 4724 4036
rect 4756 4004 4884 4036
rect 4916 4004 5044 4036
rect 5076 4004 5204 4036
rect 5236 4004 5364 4036
rect 5396 4004 5524 4036
rect 5556 4004 5684 4036
rect 5716 4004 5720 4036
rect 4720 4000 5720 4004
rect 5760 4036 5960 4040
rect 5760 4004 5764 4036
rect 5796 4004 5924 4036
rect 5956 4004 5960 4036
rect 5760 4000 5960 4004
rect 6000 4036 6200 4040
rect 6000 4004 6004 4036
rect 6036 4004 6164 4036
rect 6196 4004 6200 4036
rect 6000 4000 6200 4004
rect 4240 3956 4440 3960
rect 4240 3924 4244 3956
rect 4276 3924 4404 3956
rect 4436 3924 4440 3956
rect 4240 3920 4440 3924
rect 4480 3956 4680 3960
rect 4480 3924 4484 3956
rect 4516 3924 4644 3956
rect 4676 3924 4680 3956
rect 4480 3920 4680 3924
rect 4720 3956 5720 3960
rect 4720 3924 4724 3956
rect 4756 3924 4884 3956
rect 4916 3924 5044 3956
rect 5076 3924 5204 3956
rect 5236 3924 5364 3956
rect 5396 3924 5524 3956
rect 5556 3924 5684 3956
rect 5716 3924 5720 3956
rect 4720 3920 5720 3924
rect 5760 3956 5960 3960
rect 5760 3924 5764 3956
rect 5796 3924 5924 3956
rect 5956 3924 5960 3956
rect 5760 3920 5960 3924
rect 6000 3956 6200 3960
rect 6000 3924 6004 3956
rect 6036 3924 6164 3956
rect 6196 3924 6200 3956
rect 6000 3920 6200 3924
rect 4240 3876 4440 3880
rect 4240 3844 4244 3876
rect 4276 3844 4404 3876
rect 4436 3844 4440 3876
rect 4240 3840 4440 3844
rect 4480 3876 4680 3880
rect 4480 3844 4484 3876
rect 4516 3844 4644 3876
rect 4676 3844 4680 3876
rect 4480 3840 4680 3844
rect 4720 3876 5720 3880
rect 4720 3844 4724 3876
rect 4756 3844 4884 3876
rect 4916 3844 5044 3876
rect 5076 3844 5204 3876
rect 5236 3844 5364 3876
rect 5396 3844 5524 3876
rect 5556 3844 5684 3876
rect 5716 3844 5720 3876
rect 4720 3840 5720 3844
rect 5760 3876 5960 3880
rect 5760 3844 5764 3876
rect 5796 3844 5924 3876
rect 5956 3844 5960 3876
rect 5760 3840 5960 3844
rect 6000 3876 6200 3880
rect 6000 3844 6004 3876
rect 6036 3844 6164 3876
rect 6196 3844 6200 3876
rect 6000 3840 6200 3844
rect 4240 3796 4440 3800
rect 4240 3764 4244 3796
rect 4276 3764 4404 3796
rect 4436 3764 4440 3796
rect 4240 3760 4440 3764
rect 4480 3796 4680 3800
rect 4480 3764 4484 3796
rect 4516 3764 4644 3796
rect 4676 3764 4680 3796
rect 4480 3760 4680 3764
rect 4720 3796 5720 3800
rect 4720 3764 4724 3796
rect 4756 3764 4884 3796
rect 4916 3764 5044 3796
rect 5076 3764 5204 3796
rect 5236 3764 5364 3796
rect 5396 3764 5524 3796
rect 5556 3764 5684 3796
rect 5716 3764 5720 3796
rect 4720 3760 5720 3764
rect 5760 3796 5960 3800
rect 5760 3764 5764 3796
rect 5796 3764 5924 3796
rect 5956 3764 5960 3796
rect 5760 3760 5960 3764
rect 6000 3796 6200 3800
rect 6000 3764 6004 3796
rect 6036 3764 6164 3796
rect 6196 3764 6200 3796
rect 6000 3760 6200 3764
rect 4240 3716 4440 3720
rect 4240 3684 4244 3716
rect 4276 3684 4404 3716
rect 4436 3684 4440 3716
rect 4240 3680 4440 3684
rect 4480 3716 4680 3720
rect 4480 3684 4484 3716
rect 4516 3684 4644 3716
rect 4676 3684 4680 3716
rect 4480 3680 4680 3684
rect 4720 3716 5720 3720
rect 4720 3684 4724 3716
rect 4756 3684 4884 3716
rect 4916 3684 5044 3716
rect 5076 3684 5204 3716
rect 5236 3684 5364 3716
rect 5396 3684 5524 3716
rect 5556 3684 5684 3716
rect 5716 3684 5720 3716
rect 4720 3680 5720 3684
rect 5760 3716 5960 3720
rect 5760 3684 5764 3716
rect 5796 3684 5924 3716
rect 5956 3684 5960 3716
rect 5760 3680 5960 3684
rect 6000 3716 6200 3720
rect 6000 3684 6004 3716
rect 6036 3684 6164 3716
rect 6196 3684 6200 3716
rect 6000 3680 6200 3684
rect 4240 3636 4440 3640
rect 4240 3604 4244 3636
rect 4276 3604 4404 3636
rect 4436 3604 4440 3636
rect 4240 3600 4440 3604
rect 4480 3636 4680 3640
rect 4480 3604 4484 3636
rect 4516 3604 4644 3636
rect 4676 3604 4680 3636
rect 4480 3600 4680 3604
rect 4720 3636 5720 3640
rect 4720 3604 4724 3636
rect 4756 3604 4884 3636
rect 4916 3604 5044 3636
rect 5076 3604 5204 3636
rect 5236 3604 5364 3636
rect 5396 3604 5524 3636
rect 5556 3604 5684 3636
rect 5716 3604 5720 3636
rect 4720 3600 5720 3604
rect 5760 3636 5960 3640
rect 5760 3604 5764 3636
rect 5796 3604 5924 3636
rect 5956 3604 5960 3636
rect 5760 3600 5960 3604
rect 6000 3636 6200 3640
rect 6000 3604 6004 3636
rect 6036 3604 6164 3636
rect 6196 3604 6200 3636
rect 6000 3600 6200 3604
rect 4240 3556 4440 3560
rect 4240 3524 4244 3556
rect 4276 3524 4404 3556
rect 4436 3524 4440 3556
rect 4240 3520 4440 3524
rect 4480 3556 4680 3560
rect 4480 3524 4484 3556
rect 4516 3524 4644 3556
rect 4676 3524 4680 3556
rect 4480 3520 4680 3524
rect 4720 3556 5720 3560
rect 4720 3524 4724 3556
rect 4756 3524 4884 3556
rect 4916 3524 5044 3556
rect 5076 3524 5204 3556
rect 5236 3524 5364 3556
rect 5396 3524 5524 3556
rect 5556 3524 5684 3556
rect 5716 3524 5720 3556
rect 4720 3520 5720 3524
rect 5760 3556 5960 3560
rect 5760 3524 5764 3556
rect 5796 3524 5924 3556
rect 5956 3524 5960 3556
rect 5760 3520 5960 3524
rect 6000 3556 6200 3560
rect 6000 3524 6004 3556
rect 6036 3524 6164 3556
rect 6196 3524 6200 3556
rect 6000 3520 6200 3524
rect 4240 3476 4440 3480
rect 4240 3444 4244 3476
rect 4276 3444 4404 3476
rect 4436 3444 4440 3476
rect 4240 3440 4440 3444
rect 4480 3476 4680 3480
rect 4480 3444 4484 3476
rect 4516 3444 4644 3476
rect 4676 3444 4680 3476
rect 4480 3440 4680 3444
rect 4720 3476 5720 3480
rect 4720 3444 4724 3476
rect 4756 3444 4884 3476
rect 4916 3444 5044 3476
rect 5076 3444 5204 3476
rect 5236 3444 5364 3476
rect 5396 3444 5524 3476
rect 5556 3444 5684 3476
rect 5716 3444 5720 3476
rect 4720 3440 5720 3444
rect 5760 3476 5960 3480
rect 5760 3444 5764 3476
rect 5796 3444 5924 3476
rect 5956 3444 5960 3476
rect 5760 3440 5960 3444
rect 6000 3476 6200 3480
rect 6000 3444 6004 3476
rect 6036 3444 6164 3476
rect 6196 3444 6200 3476
rect 6000 3440 6200 3444
rect 4240 3396 4440 3400
rect 4240 3364 4244 3396
rect 4276 3364 4404 3396
rect 4436 3364 4440 3396
rect 4240 3360 4440 3364
rect 4480 3396 4680 3400
rect 4480 3364 4484 3396
rect 4516 3364 4644 3396
rect 4676 3364 4680 3396
rect 4480 3360 4680 3364
rect 4720 3396 5720 3400
rect 4720 3364 4724 3396
rect 4756 3364 4884 3396
rect 4916 3364 5044 3396
rect 5076 3364 5204 3396
rect 5236 3364 5364 3396
rect 5396 3364 5524 3396
rect 5556 3364 5684 3396
rect 5716 3364 5720 3396
rect 4720 3360 5720 3364
rect 5760 3396 5960 3400
rect 5760 3364 5764 3396
rect 5796 3364 5924 3396
rect 5956 3364 5960 3396
rect 5760 3360 5960 3364
rect 6000 3396 6200 3400
rect 6000 3364 6004 3396
rect 6036 3364 6164 3396
rect 6196 3364 6200 3396
rect 6000 3360 6200 3364
rect 4240 3316 4440 3320
rect 4240 3284 4244 3316
rect 4276 3284 4404 3316
rect 4436 3284 4440 3316
rect 4240 3280 4440 3284
rect 4480 3316 4680 3320
rect 4480 3284 4484 3316
rect 4516 3284 4644 3316
rect 4676 3284 4680 3316
rect 4480 3280 4680 3284
rect 4720 3316 5720 3320
rect 4720 3284 4724 3316
rect 4756 3284 4884 3316
rect 4916 3284 5044 3316
rect 5076 3284 5204 3316
rect 5236 3284 5364 3316
rect 5396 3284 5524 3316
rect 5556 3284 5684 3316
rect 5716 3284 5720 3316
rect 4720 3280 5720 3284
rect 5760 3316 5960 3320
rect 5760 3284 5764 3316
rect 5796 3284 5924 3316
rect 5956 3284 5960 3316
rect 5760 3280 5960 3284
rect 6000 3316 6200 3320
rect 6000 3284 6004 3316
rect 6036 3284 6164 3316
rect 6196 3284 6200 3316
rect 6000 3280 6200 3284
rect 4240 3236 4440 3240
rect 4240 3204 4244 3236
rect 4276 3204 4404 3236
rect 4436 3204 4440 3236
rect 4240 3200 4440 3204
rect 4480 3236 4680 3240
rect 4480 3204 4484 3236
rect 4516 3204 4644 3236
rect 4676 3204 4680 3236
rect 4480 3200 4680 3204
rect 4720 3236 5720 3240
rect 4720 3204 4724 3236
rect 4756 3204 4884 3236
rect 4916 3204 5044 3236
rect 5076 3204 5204 3236
rect 5236 3204 5364 3236
rect 5396 3204 5524 3236
rect 5556 3204 5684 3236
rect 5716 3204 5720 3236
rect 4720 3200 5720 3204
rect 5760 3236 5960 3240
rect 5760 3204 5764 3236
rect 5796 3204 5924 3236
rect 5956 3204 5960 3236
rect 5760 3200 5960 3204
rect 6000 3236 6200 3240
rect 6000 3204 6004 3236
rect 6036 3204 6164 3236
rect 6196 3204 6200 3236
rect 6000 3200 6200 3204
rect 4240 3156 4440 3160
rect 4240 3124 4244 3156
rect 4276 3124 4404 3156
rect 4436 3124 4440 3156
rect 4240 3120 4440 3124
rect 4480 3156 4680 3160
rect 4480 3124 4484 3156
rect 4516 3124 4644 3156
rect 4676 3124 4680 3156
rect 4480 3120 4680 3124
rect 4720 3156 5720 3160
rect 4720 3124 4724 3156
rect 4756 3124 4884 3156
rect 4916 3124 5044 3156
rect 5076 3124 5204 3156
rect 5236 3124 5364 3156
rect 5396 3124 5524 3156
rect 5556 3124 5684 3156
rect 5716 3124 5720 3156
rect 4720 3120 5720 3124
rect 5760 3156 5960 3160
rect 5760 3124 5764 3156
rect 5796 3124 5924 3156
rect 5956 3124 5960 3156
rect 5760 3120 5960 3124
rect 6000 3156 6200 3160
rect 6000 3124 6004 3156
rect 6036 3124 6164 3156
rect 6196 3124 6200 3156
rect 6000 3120 6200 3124
rect 4240 3076 4440 3080
rect 4240 3044 4244 3076
rect 4276 3044 4404 3076
rect 4436 3044 4440 3076
rect 4240 3040 4440 3044
rect 4480 3076 4680 3080
rect 4480 3044 4484 3076
rect 4516 3044 4644 3076
rect 4676 3044 4680 3076
rect 4480 3040 4680 3044
rect 4720 3076 5720 3080
rect 4720 3044 4724 3076
rect 4756 3044 4884 3076
rect 4916 3044 5044 3076
rect 5076 3044 5204 3076
rect 5236 3044 5364 3076
rect 5396 3044 5524 3076
rect 5556 3044 5684 3076
rect 5716 3044 5720 3076
rect 4720 3040 5720 3044
rect 5760 3076 5960 3080
rect 5760 3044 5764 3076
rect 5796 3044 5924 3076
rect 5956 3044 5960 3076
rect 5760 3040 5960 3044
rect 6000 3076 6200 3080
rect 6000 3044 6004 3076
rect 6036 3044 6164 3076
rect 6196 3044 6200 3076
rect 6000 3040 6200 3044
rect 4240 2996 4440 3000
rect 4240 2964 4244 2996
rect 4276 2964 4404 2996
rect 4436 2964 4440 2996
rect 4240 2960 4440 2964
rect 4480 2996 4680 3000
rect 4480 2964 4484 2996
rect 4516 2964 4644 2996
rect 4676 2964 4680 2996
rect 4480 2960 4680 2964
rect 4720 2996 5720 3000
rect 4720 2964 4724 2996
rect 4756 2964 4884 2996
rect 4916 2964 5044 2996
rect 5076 2964 5204 2996
rect 5236 2964 5364 2996
rect 5396 2964 5524 2996
rect 5556 2964 5684 2996
rect 5716 2964 5720 2996
rect 4720 2960 5720 2964
rect 5760 2996 5960 3000
rect 5760 2964 5764 2996
rect 5796 2964 5924 2996
rect 5956 2964 5960 2996
rect 5760 2960 5960 2964
rect 6000 2996 6200 3000
rect 6000 2964 6004 2996
rect 6036 2964 6164 2996
rect 6196 2964 6200 2996
rect 6000 2960 6200 2964
rect 4240 2916 4440 2920
rect 4240 2884 4244 2916
rect 4276 2884 4404 2916
rect 4436 2884 4440 2916
rect 4240 2880 4440 2884
rect 4480 2916 4680 2920
rect 4480 2884 4484 2916
rect 4516 2884 4644 2916
rect 4676 2884 4680 2916
rect 4480 2880 4680 2884
rect 4720 2916 5720 2920
rect 4720 2884 4724 2916
rect 4756 2884 4884 2916
rect 4916 2884 5044 2916
rect 5076 2884 5204 2916
rect 5236 2884 5364 2916
rect 5396 2884 5524 2916
rect 5556 2884 5684 2916
rect 5716 2884 5720 2916
rect 4720 2880 5720 2884
rect 5760 2916 5960 2920
rect 5760 2884 5764 2916
rect 5796 2884 5924 2916
rect 5956 2884 5960 2916
rect 5760 2880 5960 2884
rect 6000 2916 6200 2920
rect 6000 2884 6004 2916
rect 6036 2884 6164 2916
rect 6196 2884 6200 2916
rect 6000 2880 6200 2884
rect 4240 2836 4440 2840
rect 4240 2804 4244 2836
rect 4276 2804 4404 2836
rect 4436 2804 4440 2836
rect 4240 2800 4440 2804
rect 4480 2836 4680 2840
rect 4480 2804 4484 2836
rect 4516 2804 4644 2836
rect 4676 2804 4680 2836
rect 4480 2800 4680 2804
rect 4720 2836 5720 2840
rect 4720 2804 4724 2836
rect 4756 2804 4884 2836
rect 4916 2804 5044 2836
rect 5076 2804 5204 2836
rect 5236 2804 5364 2836
rect 5396 2804 5524 2836
rect 5556 2804 5684 2836
rect 5716 2804 5720 2836
rect 4720 2800 5720 2804
rect 5760 2836 5960 2840
rect 5760 2804 5764 2836
rect 5796 2804 5924 2836
rect 5956 2804 5960 2836
rect 5760 2800 5960 2804
rect 6000 2836 6200 2840
rect 6000 2804 6004 2836
rect 6036 2804 6164 2836
rect 6196 2804 6200 2836
rect 6000 2800 6200 2804
rect 4240 2756 4440 2760
rect 4240 2724 4244 2756
rect 4276 2724 4404 2756
rect 4436 2724 4440 2756
rect 4240 2720 4440 2724
rect 4480 2756 4680 2760
rect 4480 2724 4484 2756
rect 4516 2724 4644 2756
rect 4676 2724 4680 2756
rect 4480 2720 4680 2724
rect 4720 2756 5720 2760
rect 4720 2724 4724 2756
rect 4756 2724 4884 2756
rect 4916 2724 5044 2756
rect 5076 2724 5204 2756
rect 5236 2724 5364 2756
rect 5396 2724 5524 2756
rect 5556 2724 5684 2756
rect 5716 2724 5720 2756
rect 4720 2720 5720 2724
rect 5760 2756 5960 2760
rect 5760 2724 5764 2756
rect 5796 2724 5924 2756
rect 5956 2724 5960 2756
rect 5760 2720 5960 2724
rect 6000 2756 6200 2760
rect 6000 2724 6004 2756
rect 6036 2724 6164 2756
rect 6196 2724 6200 2756
rect 6000 2720 6200 2724
rect 4240 2676 4440 2680
rect 4240 2644 4244 2676
rect 4276 2644 4404 2676
rect 4436 2644 4440 2676
rect 4240 2640 4440 2644
rect 4480 2676 4680 2680
rect 4480 2644 4484 2676
rect 4516 2644 4644 2676
rect 4676 2644 4680 2676
rect 4480 2640 4680 2644
rect 4720 2676 5720 2680
rect 4720 2644 4724 2676
rect 4756 2644 4884 2676
rect 4916 2644 5044 2676
rect 5076 2644 5204 2676
rect 5236 2644 5364 2676
rect 5396 2644 5524 2676
rect 5556 2644 5684 2676
rect 5716 2644 5720 2676
rect 4720 2640 5720 2644
rect 5760 2676 5960 2680
rect 5760 2644 5764 2676
rect 5796 2644 5924 2676
rect 5956 2644 5960 2676
rect 5760 2640 5960 2644
rect 6000 2676 6200 2680
rect 6000 2644 6004 2676
rect 6036 2644 6164 2676
rect 6196 2644 6200 2676
rect 6000 2640 6200 2644
rect 4240 2596 4440 2600
rect 4240 2564 4244 2596
rect 4276 2564 4404 2596
rect 4436 2564 4440 2596
rect 4240 2560 4440 2564
rect 4480 2596 4680 2600
rect 4480 2564 4484 2596
rect 4516 2564 4644 2596
rect 4676 2564 4680 2596
rect 4480 2560 4680 2564
rect 4720 2596 5720 2600
rect 4720 2564 4724 2596
rect 4756 2564 4884 2596
rect 4916 2564 5044 2596
rect 5076 2564 5204 2596
rect 5236 2564 5364 2596
rect 5396 2564 5524 2596
rect 5556 2564 5684 2596
rect 5716 2564 5720 2596
rect 4720 2560 5720 2564
rect 5760 2596 5960 2600
rect 5760 2564 5764 2596
rect 5796 2564 5924 2596
rect 5956 2564 5960 2596
rect 5760 2560 5960 2564
rect 6000 2596 6200 2600
rect 6000 2564 6004 2596
rect 6036 2564 6164 2596
rect 6196 2564 6200 2596
rect 6000 2560 6200 2564
rect 4240 2516 4440 2520
rect 4240 2484 4244 2516
rect 4276 2484 4404 2516
rect 4436 2484 4440 2516
rect 4240 2480 4440 2484
rect 4480 2516 4680 2520
rect 4480 2484 4484 2516
rect 4516 2484 4644 2516
rect 4676 2484 4680 2516
rect 4480 2480 4680 2484
rect 4720 2516 5720 2520
rect 4720 2484 4724 2516
rect 4756 2484 4884 2516
rect 4916 2484 5044 2516
rect 5076 2484 5204 2516
rect 5236 2484 5364 2516
rect 5396 2484 5524 2516
rect 5556 2484 5684 2516
rect 5716 2484 5720 2516
rect 4720 2480 5720 2484
rect 5760 2516 5960 2520
rect 5760 2484 5764 2516
rect 5796 2484 5924 2516
rect 5956 2484 5960 2516
rect 5760 2480 5960 2484
rect 6000 2516 6200 2520
rect 6000 2484 6004 2516
rect 6036 2484 6164 2516
rect 6196 2484 6200 2516
rect 6000 2480 6200 2484
rect 4240 2436 4440 2440
rect 4240 2404 4244 2436
rect 4276 2404 4404 2436
rect 4436 2404 4440 2436
rect 4240 2400 4440 2404
rect 4480 2436 4680 2440
rect 4480 2404 4484 2436
rect 4516 2404 4644 2436
rect 4676 2404 4680 2436
rect 4480 2400 4680 2404
rect 4720 2436 5720 2440
rect 4720 2404 4724 2436
rect 4756 2404 4884 2436
rect 4916 2404 5044 2436
rect 5076 2404 5204 2436
rect 5236 2404 5364 2436
rect 5396 2404 5524 2436
rect 5556 2404 5684 2436
rect 5716 2404 5720 2436
rect 4720 2400 5720 2404
rect 5760 2436 5960 2440
rect 5760 2404 5764 2436
rect 5796 2404 5924 2436
rect 5956 2404 5960 2436
rect 5760 2400 5960 2404
rect 6000 2436 6200 2440
rect 6000 2404 6004 2436
rect 6036 2404 6164 2436
rect 6196 2404 6200 2436
rect 6000 2400 6200 2404
rect 4240 2356 4440 2360
rect 4240 2324 4244 2356
rect 4276 2324 4404 2356
rect 4436 2324 4440 2356
rect 4240 2320 4440 2324
rect 4480 2356 4680 2360
rect 4480 2324 4484 2356
rect 4516 2324 4644 2356
rect 4676 2324 4680 2356
rect 4480 2320 4680 2324
rect 4720 2356 5720 2360
rect 4720 2324 4724 2356
rect 4756 2324 4884 2356
rect 4916 2324 5044 2356
rect 5076 2324 5204 2356
rect 5236 2324 5364 2356
rect 5396 2324 5524 2356
rect 5556 2324 5684 2356
rect 5716 2324 5720 2356
rect 4720 2320 5720 2324
rect 5760 2356 5960 2360
rect 5760 2324 5764 2356
rect 5796 2324 5924 2356
rect 5956 2324 5960 2356
rect 5760 2320 5960 2324
rect 6000 2356 6200 2360
rect 6000 2324 6004 2356
rect 6036 2324 6164 2356
rect 6196 2324 6200 2356
rect 6000 2320 6200 2324
rect 4240 2276 4440 2280
rect 4240 2244 4244 2276
rect 4276 2244 4404 2276
rect 4436 2244 4440 2276
rect 4240 2240 4440 2244
rect 4480 2276 4680 2280
rect 4480 2244 4484 2276
rect 4516 2244 4644 2276
rect 4676 2244 4680 2276
rect 4480 2240 4680 2244
rect 4720 2276 5720 2280
rect 4720 2244 4724 2276
rect 4756 2244 4884 2276
rect 4916 2244 5044 2276
rect 5076 2244 5204 2276
rect 5236 2244 5364 2276
rect 5396 2244 5524 2276
rect 5556 2244 5684 2276
rect 5716 2244 5720 2276
rect 4720 2240 5720 2244
rect 5760 2276 5960 2280
rect 5760 2244 5764 2276
rect 5796 2244 5924 2276
rect 5956 2244 5960 2276
rect 5760 2240 5960 2244
rect 6000 2276 6200 2280
rect 6000 2244 6004 2276
rect 6036 2244 6164 2276
rect 6196 2244 6200 2276
rect 6000 2240 6200 2244
rect 4240 2196 4440 2200
rect 4240 2164 4244 2196
rect 4276 2164 4404 2196
rect 4436 2164 4440 2196
rect 4240 2160 4440 2164
rect 4480 2196 4680 2200
rect 4480 2164 4484 2196
rect 4516 2164 4644 2196
rect 4676 2164 4680 2196
rect 4480 2160 4680 2164
rect 4720 2196 5720 2200
rect 4720 2164 4724 2196
rect 4756 2164 4884 2196
rect 4916 2164 5044 2196
rect 5076 2164 5204 2196
rect 5236 2164 5364 2196
rect 5396 2164 5524 2196
rect 5556 2164 5684 2196
rect 5716 2164 5720 2196
rect 4720 2160 5720 2164
rect 5760 2196 5960 2200
rect 5760 2164 5764 2196
rect 5796 2164 5924 2196
rect 5956 2164 5960 2196
rect 5760 2160 5960 2164
rect 6000 2196 6200 2200
rect 6000 2164 6004 2196
rect 6036 2164 6164 2196
rect 6196 2164 6200 2196
rect 6000 2160 6200 2164
rect 4240 2116 4440 2120
rect 4240 2084 4244 2116
rect 4276 2084 4404 2116
rect 4436 2084 4440 2116
rect 4240 2080 4440 2084
rect 4480 2116 4680 2120
rect 4480 2084 4484 2116
rect 4516 2084 4644 2116
rect 4676 2084 4680 2116
rect 4480 2080 4680 2084
rect 4720 2116 5720 2120
rect 4720 2084 4724 2116
rect 4756 2084 4884 2116
rect 4916 2084 5044 2116
rect 5076 2084 5204 2116
rect 5236 2084 5364 2116
rect 5396 2084 5524 2116
rect 5556 2084 5684 2116
rect 5716 2084 5720 2116
rect 4720 2080 5720 2084
rect 5760 2116 5960 2120
rect 5760 2084 5764 2116
rect 5796 2084 5924 2116
rect 5956 2084 5960 2116
rect 5760 2080 5960 2084
rect 6000 2116 6200 2120
rect 6000 2084 6004 2116
rect 6036 2084 6164 2116
rect 6196 2084 6200 2116
rect 6000 2080 6200 2084
rect 4240 2036 4440 2040
rect 4240 2004 4244 2036
rect 4276 2004 4404 2036
rect 4436 2004 4440 2036
rect 4240 2000 4440 2004
rect 4480 2036 4680 2040
rect 4480 2004 4484 2036
rect 4516 2004 4644 2036
rect 4676 2004 4680 2036
rect 4480 2000 4680 2004
rect 4720 2036 5720 2040
rect 4720 2004 4724 2036
rect 4756 2004 4884 2036
rect 4916 2004 5044 2036
rect 5076 2004 5204 2036
rect 5236 2004 5364 2036
rect 5396 2004 5524 2036
rect 5556 2004 5684 2036
rect 5716 2004 5720 2036
rect 4720 2000 5720 2004
rect 5760 2036 5960 2040
rect 5760 2004 5764 2036
rect 5796 2004 5924 2036
rect 5956 2004 5960 2036
rect 5760 2000 5960 2004
rect 6000 2036 6200 2040
rect 6000 2004 6004 2036
rect 6036 2004 6164 2036
rect 6196 2004 6200 2036
rect 6000 2000 6200 2004
rect 4240 1956 4440 1960
rect 4240 1924 4244 1956
rect 4276 1924 4404 1956
rect 4436 1924 4440 1956
rect 4240 1920 4440 1924
rect 4480 1956 4680 1960
rect 4480 1924 4484 1956
rect 4516 1924 4644 1956
rect 4676 1924 4680 1956
rect 4480 1920 4680 1924
rect 4720 1956 5720 1960
rect 4720 1924 4724 1956
rect 4756 1924 4884 1956
rect 4916 1924 5044 1956
rect 5076 1924 5204 1956
rect 5236 1924 5364 1956
rect 5396 1924 5524 1956
rect 5556 1924 5684 1956
rect 5716 1924 5720 1956
rect 4720 1920 5720 1924
rect 5760 1956 5960 1960
rect 5760 1924 5764 1956
rect 5796 1924 5924 1956
rect 5956 1924 5960 1956
rect 5760 1920 5960 1924
rect 6000 1956 6200 1960
rect 6000 1924 6004 1956
rect 6036 1924 6164 1956
rect 6196 1924 6200 1956
rect 6000 1920 6200 1924
rect 4240 1876 4440 1880
rect 4240 1844 4244 1876
rect 4276 1844 4404 1876
rect 4436 1844 4440 1876
rect 4240 1840 4440 1844
rect 4480 1876 4680 1880
rect 4480 1844 4484 1876
rect 4516 1844 4644 1876
rect 4676 1844 4680 1876
rect 4480 1840 4680 1844
rect 4720 1876 5720 1880
rect 4720 1844 4724 1876
rect 4756 1844 4884 1876
rect 4916 1844 5044 1876
rect 5076 1844 5204 1876
rect 5236 1844 5364 1876
rect 5396 1844 5524 1876
rect 5556 1844 5684 1876
rect 5716 1844 5720 1876
rect 4720 1840 5720 1844
rect 5760 1876 5960 1880
rect 5760 1844 5764 1876
rect 5796 1844 5924 1876
rect 5956 1844 5960 1876
rect 5760 1840 5960 1844
rect 6000 1876 6200 1880
rect 6000 1844 6004 1876
rect 6036 1844 6164 1876
rect 6196 1844 6200 1876
rect 6000 1840 6200 1844
rect 4240 1796 4440 1800
rect 4240 1764 4244 1796
rect 4276 1764 4404 1796
rect 4436 1764 4440 1796
rect 4240 1760 4440 1764
rect 4480 1796 4680 1800
rect 4480 1764 4484 1796
rect 4516 1764 4644 1796
rect 4676 1764 4680 1796
rect 4480 1760 4680 1764
rect 4720 1796 5720 1800
rect 4720 1764 4724 1796
rect 4756 1764 4884 1796
rect 4916 1764 5044 1796
rect 5076 1764 5204 1796
rect 5236 1764 5364 1796
rect 5396 1764 5524 1796
rect 5556 1764 5684 1796
rect 5716 1764 5720 1796
rect 4720 1760 5720 1764
rect 5760 1796 5960 1800
rect 5760 1764 5764 1796
rect 5796 1764 5924 1796
rect 5956 1764 5960 1796
rect 5760 1760 5960 1764
rect 6000 1796 6200 1800
rect 6000 1764 6004 1796
rect 6036 1764 6164 1796
rect 6196 1764 6200 1796
rect 6000 1760 6200 1764
rect 4240 1716 4440 1720
rect 4240 1684 4244 1716
rect 4276 1684 4404 1716
rect 4436 1684 4440 1716
rect 4240 1680 4440 1684
rect 4480 1716 4680 1720
rect 4480 1684 4484 1716
rect 4516 1684 4644 1716
rect 4676 1684 4680 1716
rect 4480 1680 4680 1684
rect 4720 1716 5720 1720
rect 4720 1684 4724 1716
rect 4756 1684 4884 1716
rect 4916 1684 5044 1716
rect 5076 1684 5204 1716
rect 5236 1684 5364 1716
rect 5396 1684 5524 1716
rect 5556 1684 5684 1716
rect 5716 1684 5720 1716
rect 4720 1680 5720 1684
rect 5760 1716 5960 1720
rect 5760 1684 5764 1716
rect 5796 1684 5924 1716
rect 5956 1684 5960 1716
rect 5760 1680 5960 1684
rect 6000 1716 6200 1720
rect 6000 1684 6004 1716
rect 6036 1684 6164 1716
rect 6196 1684 6200 1716
rect 6000 1680 6200 1684
rect 4240 1636 4440 1640
rect 4240 1604 4244 1636
rect 4276 1604 4404 1636
rect 4436 1604 4440 1636
rect 4240 1600 4440 1604
rect 4480 1636 4680 1640
rect 4480 1604 4484 1636
rect 4516 1604 4644 1636
rect 4676 1604 4680 1636
rect 4480 1600 4680 1604
rect 4720 1636 5720 1640
rect 4720 1604 4724 1636
rect 4756 1604 4884 1636
rect 4916 1604 5044 1636
rect 5076 1604 5204 1636
rect 5236 1604 5364 1636
rect 5396 1604 5524 1636
rect 5556 1604 5684 1636
rect 5716 1604 5720 1636
rect 4720 1600 5720 1604
rect 5760 1636 5960 1640
rect 5760 1604 5764 1636
rect 5796 1604 5924 1636
rect 5956 1604 5960 1636
rect 5760 1600 5960 1604
rect 6000 1636 6200 1640
rect 6000 1604 6004 1636
rect 6036 1604 6164 1636
rect 6196 1604 6200 1636
rect 6000 1600 6200 1604
rect 4240 1556 4440 1560
rect 4240 1524 4244 1556
rect 4276 1524 4404 1556
rect 4436 1524 4440 1556
rect 4240 1520 4440 1524
rect 4480 1556 4680 1560
rect 4480 1524 4484 1556
rect 4516 1524 4644 1556
rect 4676 1524 4680 1556
rect 4480 1520 4680 1524
rect 4720 1556 5720 1560
rect 4720 1524 4724 1556
rect 4756 1524 4884 1556
rect 4916 1524 5044 1556
rect 5076 1524 5204 1556
rect 5236 1524 5364 1556
rect 5396 1524 5524 1556
rect 5556 1524 5684 1556
rect 5716 1524 5720 1556
rect 4720 1520 5720 1524
rect 5760 1556 5960 1560
rect 5760 1524 5764 1556
rect 5796 1524 5924 1556
rect 5956 1524 5960 1556
rect 5760 1520 5960 1524
rect 6000 1556 6200 1560
rect 6000 1524 6004 1556
rect 6036 1524 6164 1556
rect 6196 1524 6200 1556
rect 6000 1520 6200 1524
rect 4240 1476 4440 1480
rect 4240 1444 4244 1476
rect 4276 1444 4404 1476
rect 4436 1444 4440 1476
rect 4240 1440 4440 1444
rect 4480 1476 4680 1480
rect 4480 1444 4484 1476
rect 4516 1444 4644 1476
rect 4676 1444 4680 1476
rect 4480 1440 4680 1444
rect 4720 1476 5720 1480
rect 4720 1444 4724 1476
rect 4756 1444 4884 1476
rect 4916 1444 5044 1476
rect 5076 1444 5204 1476
rect 5236 1444 5364 1476
rect 5396 1444 5524 1476
rect 5556 1444 5684 1476
rect 5716 1444 5720 1476
rect 4720 1440 5720 1444
rect 5760 1476 5960 1480
rect 5760 1444 5764 1476
rect 5796 1444 5924 1476
rect 5956 1444 5960 1476
rect 5760 1440 5960 1444
rect 6000 1476 6200 1480
rect 6000 1444 6004 1476
rect 6036 1444 6164 1476
rect 6196 1444 6200 1476
rect 6000 1440 6200 1444
rect 4240 1396 4440 1400
rect 4240 1364 4244 1396
rect 4276 1364 4404 1396
rect 4436 1364 4440 1396
rect 4240 1360 4440 1364
rect 4480 1396 4680 1400
rect 4480 1364 4484 1396
rect 4516 1364 4644 1396
rect 4676 1364 4680 1396
rect 4480 1360 4680 1364
rect 4720 1396 5720 1400
rect 4720 1364 4724 1396
rect 4756 1364 4884 1396
rect 4916 1364 5044 1396
rect 5076 1364 5204 1396
rect 5236 1364 5364 1396
rect 5396 1364 5524 1396
rect 5556 1364 5684 1396
rect 5716 1364 5720 1396
rect 4720 1360 5720 1364
rect 5760 1396 5960 1400
rect 5760 1364 5764 1396
rect 5796 1364 5924 1396
rect 5956 1364 5960 1396
rect 5760 1360 5960 1364
rect 6000 1396 6200 1400
rect 6000 1364 6004 1396
rect 6036 1364 6164 1396
rect 6196 1364 6200 1396
rect 6000 1360 6200 1364
rect 4240 1316 4440 1320
rect 4240 1284 4244 1316
rect 4276 1284 4404 1316
rect 4436 1284 4440 1316
rect 4240 1280 4440 1284
rect 4480 1316 4680 1320
rect 4480 1284 4484 1316
rect 4516 1284 4644 1316
rect 4676 1284 4680 1316
rect 4480 1280 4680 1284
rect 4720 1316 5720 1320
rect 4720 1284 4724 1316
rect 4756 1284 4884 1316
rect 4916 1284 5044 1316
rect 5076 1284 5204 1316
rect 5236 1284 5364 1316
rect 5396 1284 5524 1316
rect 5556 1284 5684 1316
rect 5716 1284 5720 1316
rect 4720 1280 5720 1284
rect 5760 1316 5960 1320
rect 5760 1284 5764 1316
rect 5796 1284 5924 1316
rect 5956 1284 5960 1316
rect 5760 1280 5960 1284
rect 6000 1316 6200 1320
rect 6000 1284 6004 1316
rect 6036 1284 6164 1316
rect 6196 1284 6200 1316
rect 6000 1280 6200 1284
rect 4240 1236 4440 1240
rect 4240 1204 4244 1236
rect 4276 1204 4404 1236
rect 4436 1204 4440 1236
rect 4240 1200 4440 1204
rect 4480 1236 4680 1240
rect 4480 1204 4484 1236
rect 4516 1204 4644 1236
rect 4676 1204 4680 1236
rect 4480 1200 4680 1204
rect 4720 1236 5720 1240
rect 4720 1204 4724 1236
rect 4756 1204 4884 1236
rect 4916 1204 5044 1236
rect 5076 1204 5204 1236
rect 5236 1204 5364 1236
rect 5396 1204 5524 1236
rect 5556 1204 5684 1236
rect 5716 1204 5720 1236
rect 4720 1200 5720 1204
rect 5760 1236 5960 1240
rect 5760 1204 5764 1236
rect 5796 1204 5924 1236
rect 5956 1204 5960 1236
rect 5760 1200 5960 1204
rect 6000 1236 6200 1240
rect 6000 1204 6004 1236
rect 6036 1204 6164 1236
rect 6196 1204 6200 1236
rect 6000 1200 6200 1204
rect 4240 1156 4440 1160
rect 4240 1124 4244 1156
rect 4276 1124 4404 1156
rect 4436 1124 4440 1156
rect 4240 1120 4440 1124
rect 4480 1156 4680 1160
rect 4480 1124 4484 1156
rect 4516 1124 4644 1156
rect 4676 1124 4680 1156
rect 4480 1120 4680 1124
rect 4720 1156 5720 1160
rect 4720 1124 4724 1156
rect 4756 1124 4884 1156
rect 4916 1124 5044 1156
rect 5076 1124 5204 1156
rect 5236 1124 5364 1156
rect 5396 1124 5524 1156
rect 5556 1124 5684 1156
rect 5716 1124 5720 1156
rect 4720 1120 5720 1124
rect 5760 1156 5960 1160
rect 5760 1124 5764 1156
rect 5796 1124 5924 1156
rect 5956 1124 5960 1156
rect 5760 1120 5960 1124
rect 6000 1156 6200 1160
rect 6000 1124 6004 1156
rect 6036 1124 6164 1156
rect 6196 1124 6200 1156
rect 6000 1120 6200 1124
rect 4240 1076 4440 1080
rect 4240 1044 4244 1076
rect 4276 1044 4404 1076
rect 4436 1044 4440 1076
rect 4240 1040 4440 1044
rect 4480 1076 4680 1080
rect 4480 1044 4484 1076
rect 4516 1044 4644 1076
rect 4676 1044 4680 1076
rect 4480 1040 4680 1044
rect 4720 1076 5720 1080
rect 4720 1044 4724 1076
rect 4756 1044 4884 1076
rect 4916 1044 5044 1076
rect 5076 1044 5204 1076
rect 5236 1044 5364 1076
rect 5396 1044 5524 1076
rect 5556 1044 5684 1076
rect 5716 1044 5720 1076
rect 4720 1040 5720 1044
rect 5760 1076 5960 1080
rect 5760 1044 5764 1076
rect 5796 1044 5924 1076
rect 5956 1044 5960 1076
rect 5760 1040 5960 1044
rect 6000 1076 6200 1080
rect 6000 1044 6004 1076
rect 6036 1044 6164 1076
rect 6196 1044 6200 1076
rect 6000 1040 6200 1044
rect 4240 996 4440 1000
rect 4240 964 4244 996
rect 4276 964 4404 996
rect 4436 964 4440 996
rect 4240 960 4440 964
rect 4480 996 4680 1000
rect 4480 964 4484 996
rect 4516 964 4644 996
rect 4676 964 4680 996
rect 4480 960 4680 964
rect 4720 996 5720 1000
rect 4720 964 4724 996
rect 4756 964 4884 996
rect 4916 964 5044 996
rect 5076 964 5204 996
rect 5236 964 5364 996
rect 5396 964 5524 996
rect 5556 964 5684 996
rect 5716 964 5720 996
rect 4720 960 5720 964
rect 5760 996 5960 1000
rect 5760 964 5764 996
rect 5796 964 5924 996
rect 5956 964 5960 996
rect 5760 960 5960 964
rect 6000 996 6200 1000
rect 6000 964 6004 996
rect 6036 964 6164 996
rect 6196 964 6200 996
rect 6000 960 6200 964
rect 4240 916 4440 920
rect 4240 884 4244 916
rect 4276 884 4404 916
rect 4436 884 4440 916
rect 4240 880 4440 884
rect 4480 916 4680 920
rect 4480 884 4484 916
rect 4516 884 4644 916
rect 4676 884 4680 916
rect 4480 880 4680 884
rect 4720 916 5720 920
rect 4720 884 4724 916
rect 4756 884 4884 916
rect 4916 884 5044 916
rect 5076 884 5204 916
rect 5236 884 5364 916
rect 5396 884 5524 916
rect 5556 884 5684 916
rect 5716 884 5720 916
rect 4720 880 5720 884
rect 5760 916 5960 920
rect 5760 884 5764 916
rect 5796 884 5924 916
rect 5956 884 5960 916
rect 5760 880 5960 884
rect 6000 916 6200 920
rect 6000 884 6004 916
rect 6036 884 6164 916
rect 6196 884 6200 916
rect 6000 880 6200 884
rect 4240 836 4440 840
rect 4240 804 4244 836
rect 4276 804 4404 836
rect 4436 804 4440 836
rect 4240 800 4440 804
rect 4480 836 4680 840
rect 4480 804 4484 836
rect 4516 804 4644 836
rect 4676 804 4680 836
rect 4480 800 4680 804
rect 4720 836 5720 840
rect 4720 804 4724 836
rect 4756 804 4884 836
rect 4916 804 5044 836
rect 5076 804 5204 836
rect 5236 804 5364 836
rect 5396 804 5524 836
rect 5556 804 5684 836
rect 5716 804 5720 836
rect 4720 800 5720 804
rect 5760 836 5960 840
rect 5760 804 5764 836
rect 5796 804 5924 836
rect 5956 804 5960 836
rect 5760 800 5960 804
rect 6000 836 6200 840
rect 6000 804 6004 836
rect 6036 804 6164 836
rect 6196 804 6200 836
rect 6000 800 6200 804
rect 4240 756 4440 760
rect 4240 724 4244 756
rect 4276 724 4404 756
rect 4436 724 4440 756
rect 4240 720 4440 724
rect 4480 756 4680 760
rect 4480 724 4484 756
rect 4516 724 4644 756
rect 4676 724 4680 756
rect 4480 720 4680 724
rect 4720 756 5720 760
rect 4720 724 4724 756
rect 4756 724 4884 756
rect 4916 724 5044 756
rect 5076 724 5204 756
rect 5236 724 5364 756
rect 5396 724 5524 756
rect 5556 724 5684 756
rect 5716 724 5720 756
rect 4720 720 5720 724
rect 5760 756 5960 760
rect 5760 724 5764 756
rect 5796 724 5924 756
rect 5956 724 5960 756
rect 5760 720 5960 724
rect 6000 756 6200 760
rect 6000 724 6004 756
rect 6036 724 6164 756
rect 6196 724 6200 756
rect 6000 720 6200 724
rect 4240 676 4440 680
rect 4240 644 4244 676
rect 4276 644 4404 676
rect 4436 644 4440 676
rect 4240 640 4440 644
rect 4480 676 4680 680
rect 4480 644 4484 676
rect 4516 644 4644 676
rect 4676 644 4680 676
rect 4480 640 4680 644
rect 4720 676 5720 680
rect 4720 644 4724 676
rect 4756 644 4884 676
rect 4916 644 5044 676
rect 5076 644 5204 676
rect 5236 644 5364 676
rect 5396 644 5524 676
rect 5556 644 5684 676
rect 5716 644 5720 676
rect 4720 640 5720 644
rect 5760 676 5960 680
rect 5760 644 5764 676
rect 5796 644 5924 676
rect 5956 644 5960 676
rect 5760 640 5960 644
rect 6000 676 6200 680
rect 6000 644 6004 676
rect 6036 644 6164 676
rect 6196 644 6200 676
rect 6000 640 6200 644
rect 4240 596 4440 600
rect 4240 564 4244 596
rect 4276 564 4404 596
rect 4436 564 4440 596
rect 4240 560 4440 564
rect 4480 596 4680 600
rect 4480 564 4484 596
rect 4516 564 4644 596
rect 4676 564 4680 596
rect 4480 560 4680 564
rect 4720 596 5720 600
rect 4720 564 4724 596
rect 4756 564 4884 596
rect 4916 564 5044 596
rect 5076 564 5204 596
rect 5236 564 5364 596
rect 5396 564 5524 596
rect 5556 564 5684 596
rect 5716 564 5720 596
rect 4720 560 5720 564
rect 5760 596 5960 600
rect 5760 564 5764 596
rect 5796 564 5924 596
rect 5956 564 5960 596
rect 5760 560 5960 564
rect 6000 596 6200 600
rect 6000 564 6004 596
rect 6036 564 6164 596
rect 6196 564 6200 596
rect 6000 560 6200 564
rect 4240 516 4440 520
rect 4240 484 4244 516
rect 4276 484 4404 516
rect 4436 484 4440 516
rect 4240 480 4440 484
rect 4480 516 4680 520
rect 4480 484 4484 516
rect 4516 484 4644 516
rect 4676 484 4680 516
rect 4480 480 4680 484
rect 4720 516 5720 520
rect 4720 484 4724 516
rect 4756 484 4884 516
rect 4916 484 5044 516
rect 5076 484 5204 516
rect 5236 484 5364 516
rect 5396 484 5524 516
rect 5556 484 5684 516
rect 5716 484 5720 516
rect 4720 480 5720 484
rect 5760 516 5960 520
rect 5760 484 5764 516
rect 5796 484 5924 516
rect 5956 484 5960 516
rect 5760 480 5960 484
rect 6000 516 6200 520
rect 6000 484 6004 516
rect 6036 484 6164 516
rect 6196 484 6200 516
rect 6000 480 6200 484
rect 4240 436 4440 440
rect 4240 404 4244 436
rect 4276 404 4404 436
rect 4436 404 4440 436
rect 4240 400 4440 404
rect 4480 436 4680 440
rect 4480 404 4484 436
rect 4516 404 4644 436
rect 4676 404 4680 436
rect 4480 400 4680 404
rect 4720 436 5720 440
rect 4720 404 4724 436
rect 4756 404 4884 436
rect 4916 404 5044 436
rect 5076 404 5204 436
rect 5236 404 5364 436
rect 5396 404 5524 436
rect 5556 404 5684 436
rect 5716 404 5720 436
rect 4720 400 5720 404
rect 5760 436 5960 440
rect 5760 404 5764 436
rect 5796 404 5924 436
rect 5956 404 5960 436
rect 5760 400 5960 404
rect 6000 436 6200 440
rect 6000 404 6004 436
rect 6036 404 6164 436
rect 6196 404 6200 436
rect 6000 400 6200 404
rect 4240 356 4440 360
rect 4240 324 4244 356
rect 4276 324 4404 356
rect 4436 324 4440 356
rect 4240 320 4440 324
rect 4480 356 4680 360
rect 4480 324 4484 356
rect 4516 324 4644 356
rect 4676 324 4680 356
rect 4480 320 4680 324
rect 4720 356 5720 360
rect 4720 324 4724 356
rect 4756 324 4884 356
rect 4916 324 5044 356
rect 5076 324 5204 356
rect 5236 324 5364 356
rect 5396 324 5524 356
rect 5556 324 5684 356
rect 5716 324 5720 356
rect 4720 320 5720 324
rect 5760 356 5960 360
rect 5760 324 5764 356
rect 5796 324 5924 356
rect 5956 324 5960 356
rect 5760 320 5960 324
rect 6000 356 6200 360
rect 6000 324 6004 356
rect 6036 324 6164 356
rect 6196 324 6200 356
rect 6000 320 6200 324
rect 4240 276 4440 280
rect 4240 244 4244 276
rect 4276 244 4404 276
rect 4436 244 4440 276
rect 4240 240 4440 244
rect 4480 276 4680 280
rect 4480 244 4484 276
rect 4516 244 4644 276
rect 4676 244 4680 276
rect 4480 240 4680 244
rect 4720 276 5720 280
rect 4720 244 4724 276
rect 4756 244 4884 276
rect 4916 244 5044 276
rect 5076 244 5204 276
rect 5236 244 5364 276
rect 5396 244 5524 276
rect 5556 244 5684 276
rect 5716 244 5720 276
rect 4720 240 5720 244
rect 5760 276 5960 280
rect 5760 244 5764 276
rect 5796 244 5924 276
rect 5956 244 5960 276
rect 5760 240 5960 244
rect 6000 276 6200 280
rect 6000 244 6004 276
rect 6036 244 6164 276
rect 6196 244 6200 276
rect 6000 240 6200 244
rect 4240 196 4440 200
rect 4240 164 4244 196
rect 4276 164 4404 196
rect 4436 164 4440 196
rect 4240 160 4440 164
rect 4480 196 4680 200
rect 4480 164 4484 196
rect 4516 164 4644 196
rect 4676 164 4680 196
rect 4480 160 4680 164
rect 4720 196 5720 200
rect 4720 164 4724 196
rect 4756 164 4884 196
rect 4916 164 5044 196
rect 5076 164 5204 196
rect 5236 164 5364 196
rect 5396 164 5524 196
rect 5556 164 5684 196
rect 5716 164 5720 196
rect 4720 160 5720 164
rect 5760 196 5960 200
rect 5760 164 5764 196
rect 5796 164 5924 196
rect 5956 164 5960 196
rect 5760 160 5960 164
rect 6000 196 6200 200
rect 6000 164 6004 196
rect 6036 164 6164 196
rect 6196 164 6200 196
rect 6000 160 6200 164
rect 4240 116 4440 120
rect 4240 84 4244 116
rect 4276 84 4404 116
rect 4436 84 4440 116
rect 4240 80 4440 84
rect 4480 116 4680 120
rect 4480 84 4484 116
rect 4516 84 4644 116
rect 4676 84 4680 116
rect 4480 80 4680 84
rect 4720 116 5720 120
rect 4720 84 4724 116
rect 4756 84 4884 116
rect 4916 84 5044 116
rect 5076 84 5204 116
rect 5236 84 5364 116
rect 5396 84 5524 116
rect 5556 84 5684 116
rect 5716 84 5720 116
rect 4720 80 5720 84
rect 5760 116 5960 120
rect 5760 84 5764 116
rect 5796 84 5924 116
rect 5956 84 5960 116
rect 5760 80 5960 84
rect 6000 116 6200 120
rect 6000 84 6004 116
rect 6036 84 6164 116
rect 6196 84 6200 116
rect 6000 80 6200 84
rect 4240 36 4440 40
rect 4240 4 4244 36
rect 4276 4 4404 36
rect 4436 4 4440 36
rect 4240 0 4440 4
rect 4480 36 4680 40
rect 4480 4 4484 36
rect 4516 4 4644 36
rect 4676 4 4680 36
rect 4480 0 4680 4
rect 4720 36 5720 40
rect 4720 4 4724 36
rect 4756 4 4884 36
rect 4916 4 5044 36
rect 5076 4 5204 36
rect 5236 4 5364 36
rect 5396 4 5524 36
rect 5556 4 5684 36
rect 5716 4 5720 36
rect 4720 0 5720 4
rect 5760 36 5960 40
rect 5760 4 5764 36
rect 5796 4 5924 36
rect 5956 4 5960 36
rect 5760 0 5960 4
rect 6000 36 6200 40
rect 6000 4 6004 36
rect 6036 4 6164 36
rect 6196 4 6200 36
rect 6000 0 6200 4
rect 0 -44 10440 -40
rect 0 -80 5764 -44
rect 0 -200 120 -80
rect 240 -200 3960 -80
rect 4080 -200 5764 -80
rect 0 -236 5764 -200
rect 5796 -236 5924 -44
rect 5956 -80 10440 -44
rect 5956 -200 6360 -80
rect 6480 -200 10200 -80
rect 10320 -200 10440 -80
rect 5956 -236 10440 -200
rect 0 -240 10440 -236
rect 0 -284 10440 -280
rect 0 -320 4484 -284
rect 0 -440 600 -320
rect 720 -440 3480 -320
rect 3600 -440 4484 -320
rect 0 -476 4484 -440
rect 4516 -476 4644 -284
rect 4676 -320 10440 -284
rect 4676 -440 6840 -320
rect 6960 -440 9720 -320
rect 9840 -440 10440 -320
rect 4676 -476 10440 -440
rect 0 -480 10440 -476
rect 0 -524 10440 -520
rect 0 -560 4724 -524
rect 0 -680 1080 -560
rect 1200 -680 2040 -560
rect 2160 -680 3000 -560
rect 3120 -680 4724 -560
rect 0 -716 4724 -680
rect 4756 -716 4884 -524
rect 4916 -716 5044 -524
rect 5076 -716 5204 -524
rect 5236 -716 5364 -524
rect 5396 -716 5524 -524
rect 5556 -716 5684 -524
rect 5716 -716 6004 -524
rect 6036 -716 6164 -524
rect 6196 -560 10440 -524
rect 6196 -680 7320 -560
rect 7440 -680 8280 -560
rect 8400 -680 9240 -560
rect 9360 -680 10440 -560
rect 6196 -716 10440 -680
rect 0 -720 10440 -716
rect 0 -764 10440 -760
rect 0 -800 4244 -764
rect 0 -920 1560 -800
rect 1680 -920 2520 -800
rect 2640 -920 4244 -800
rect 0 -956 4244 -920
rect 4276 -956 4404 -764
rect 4436 -800 10440 -764
rect 4436 -920 7800 -800
rect 7920 -920 8760 -800
rect 8880 -920 10440 -800
rect 4436 -956 10440 -920
rect 0 -960 10440 -956
rect 120 -1004 10320 -1000
rect 120 -1036 124 -1004
rect 156 -1036 4484 -1004
rect 4516 -1036 4644 -1004
rect 4676 -1036 10284 -1004
rect 10316 -1036 10320 -1004
rect 120 -1040 10320 -1036
rect 240 -1084 10280 -1080
rect 240 -1116 244 -1084
rect 276 -1116 1204 -1084
rect 1236 -1116 1364 -1084
rect 1396 -1116 2324 -1084
rect 2356 -1116 2484 -1084
rect 2516 -1116 3444 -1084
rect 3476 -1116 3604 -1084
rect 3636 -1116 4564 -1084
rect 4596 -1116 4724 -1084
rect 4756 -1116 5684 -1084
rect 5716 -1116 5844 -1084
rect 5876 -1116 6804 -1084
rect 6836 -1116 6964 -1084
rect 6996 -1116 7924 -1084
rect 7956 -1116 8084 -1084
rect 8116 -1116 9044 -1084
rect 9076 -1116 9204 -1084
rect 9236 -1116 10164 -1084
rect 10196 -1116 10280 -1084
rect 240 -1120 10280 -1116
rect 240 -1240 1240 -1160
rect 240 -2160 320 -1240
rect 1160 -2160 1240 -1240
rect 240 -2240 1240 -2160
rect 240 -2280 280 -2240
rect 1200 -2280 1240 -2240
rect 1360 -1240 2360 -1160
rect 1360 -2160 1440 -1240
rect 2280 -2160 2360 -1240
rect 1360 -2240 2360 -2160
rect 1360 -2280 1400 -2240
rect 2320 -2280 2360 -2240
rect 2480 -1240 3480 -1160
rect 2480 -2160 2560 -1240
rect 3400 -2160 3480 -1240
rect 2480 -2240 3480 -2160
rect 2480 -2280 2520 -2240
rect 3440 -2280 3480 -2240
rect 3600 -1240 4600 -1160
rect 3600 -2160 3680 -1240
rect 4520 -2160 4600 -1240
rect 3600 -2240 4600 -2160
rect 3600 -2280 3640 -2240
rect 4560 -2280 4600 -2240
rect 4720 -1240 5720 -1160
rect 4720 -2160 4800 -1240
rect 5640 -2160 5720 -1240
rect 4720 -2240 5720 -2160
rect 4720 -2280 4760 -2240
rect 5680 -2280 5720 -2240
rect 5840 -1240 6840 -1160
rect 5840 -2160 5920 -1240
rect 6760 -2160 6840 -1240
rect 5840 -2240 6840 -2160
rect 5840 -2280 5880 -2240
rect 6800 -2280 6840 -2240
rect 6960 -1240 7960 -1160
rect 6960 -2160 7040 -1240
rect 7880 -2160 7960 -1240
rect 6960 -2240 7960 -2160
rect 6960 -2280 7000 -2240
rect 7920 -2280 7960 -2240
rect 8080 -1240 9080 -1160
rect 8080 -2160 8160 -1240
rect 9000 -2160 9080 -1240
rect 8080 -2240 9080 -2160
rect 8080 -2280 8120 -2240
rect 9040 -2280 9080 -2240
rect 9200 -1240 10200 -1160
rect 9200 -2160 9280 -1240
rect 10120 -2160 10200 -1240
rect 9200 -2240 10200 -2160
rect 9200 -2280 9240 -2240
rect 10160 -2280 10200 -2240
rect 120 -2284 10320 -2280
rect 120 -2316 124 -2284
rect 156 -2316 10284 -2284
rect 10316 -2316 10320 -2284
rect 120 -2320 10320 -2316
<< via4 >>
rect 120 -200 240 -80
rect 3960 -200 4080 -80
rect 6360 -200 6480 -80
rect 10200 -200 10320 -80
rect 600 -440 720 -320
rect 3480 -440 3600 -320
rect 6840 -440 6960 -320
rect 9720 -440 9840 -320
rect 1080 -680 1200 -560
rect 2040 -680 2160 -560
rect 3000 -680 3120 -560
rect 7320 -680 7440 -560
rect 8280 -680 8400 -560
rect 9240 -680 9360 -560
rect 1560 -920 1680 -800
rect 2520 -920 2640 -800
rect 7800 -920 7920 -800
rect 8760 -920 8880 -800
<< metal5 >>
rect 80 -80 280 15800
rect 80 -200 120 -80
rect 240 -200 280 -80
rect 80 -960 280 -200
rect 560 -320 760 15800
rect 560 -440 600 -320
rect 720 -440 760 -320
rect 560 -960 760 -440
rect 1040 -560 1240 15800
rect 1040 -680 1080 -560
rect 1200 -680 1240 -560
rect 1040 -960 1240 -680
rect 1520 -800 1720 15800
rect 1520 -920 1560 -800
rect 1680 -920 1720 -800
rect 1520 -960 1720 -920
rect 2000 -560 2200 15800
rect 2000 -680 2040 -560
rect 2160 -680 2200 -560
rect 2000 -960 2200 -680
rect 2480 -800 2680 15800
rect 2480 -920 2520 -800
rect 2640 -920 2680 -800
rect 2480 -960 2680 -920
rect 2960 -560 3160 15800
rect 2960 -680 3000 -560
rect 3120 -680 3160 -560
rect 2960 -960 3160 -680
rect 3440 -320 3640 15800
rect 3440 -440 3480 -320
rect 3600 -440 3640 -320
rect 3440 -960 3640 -440
rect 3920 -80 4120 15800
rect 3920 -200 3960 -80
rect 4080 -200 4120 -80
rect 3920 -960 4120 -200
rect 6320 -80 6520 15800
rect 6320 -200 6360 -80
rect 6480 -200 6520 -80
rect 6320 -960 6520 -200
rect 6800 -320 7000 15800
rect 6800 -440 6840 -320
rect 6960 -440 7000 -320
rect 6800 -960 7000 -440
rect 7280 -560 7480 15800
rect 7280 -680 7320 -560
rect 7440 -680 7480 -560
rect 7280 -960 7480 -680
rect 7760 -800 7960 15800
rect 7760 -920 7800 -800
rect 7920 -920 7960 -800
rect 7760 -960 7960 -920
rect 8240 -560 8440 15800
rect 8240 -680 8280 -560
rect 8400 -680 8440 -560
rect 8240 -960 8440 -680
rect 8720 -800 8920 15800
rect 8720 -920 8760 -800
rect 8880 -920 8920 -800
rect 8720 -960 8920 -920
rect 9200 -560 9400 15800
rect 9200 -680 9240 -560
rect 9360 -680 9400 -560
rect 9200 -960 9400 -680
rect 9680 -320 9880 15800
rect 9680 -440 9720 -320
rect 9840 -440 9880 -320
rect 9680 -960 9880 -440
rect 10160 -80 10360 15800
rect 10160 -200 10200 -80
rect 10320 -200 10360 -80
rect 10160 -960 10360 -200
use inv_bias  biasp ../../inv1v8/mag
timestamp 1638390070
transform 1 0 0 0 1 520
box 0 -520 4200 5040
use inv_bias  biasm
timestamp 1638390070
transform -1 0 10440 0 1 520
box 0 -520 4200 5040
use inv_1_4  bp ../../inv1v8/mag
timestamp 1638390070
transform 1 0 0 0 -1 9640
box 0 0 4200 2000
use inv_1_4  cp
timestamp 1638390070
transform 1 0 0 0 1 9680
box 0 0 4200 2000
use inv_2_2  ap ../../inv1v8/mag
timestamp 1638390070
transform 1 0 0 0 1 5600
box 0 0 4200 2000
use inv_1_4  bm
timestamp 1638390070
transform -1 0 10440 0 -1 9640
box 0 0 4200 2000
use inv_1_4  cm
timestamp 1638390070
transform -1 0 10440 0 1 9680
box 0 0 4200 2000
use inv_2_2  am
timestamp 1638390070
transform -1 0 10440 0 1 5600
box 0 0 4200 2000
use inv_1_4  d
timestamp 1638390070
transform 1 0 0 0 -1 13720
box 0 0 4200 2000
use inv_2_2  fp
timestamp 1638390070
transform 1 0 0 0 1 13760
box 0 0 4200 2000
use inv_1_4  e
timestamp 1638390070
transform -1 0 10440 0 -1 13720
box 0 0 4200 2000
use inv_2_2  fm
timestamp 1638390070
transform -1 0 10440 0 1 13760
box 0 0 4200 2000
<< labels >>
rlabel metal3 5600 0 5640 15760 0 im
port 1 nsew
rlabel metal3 4800 0 4840 15760 0 ip
port 2 nsew
rlabel metal3 5440 0 5480 15760 0 op
port 3 nsew
rlabel metal3 4960 0 5000 15760 0 om
port 4 nsew
rlabel metal3 5120 0 5160 15760 0 x
port 5 nsew
rlabel metal3 5280 0 5320 15760 0 y
port 6 nsew
rlabel metal3 4320 0 4360 15760 0 ib
port 7 nsew
rlabel metal3 6080 0 6120 15760 0 q
port 8 nsew
rlabel metal3 5840 0 5880 15760 0 z
port 9 nsew
rlabel metal3 4560 0 4600 15760 0 bp
port 10 nsew
rlabel metal5 80 -960 280 15760 0 vdda
port 11 nsew
rlabel metal5 560 -960 760 15760 0 vddx
port 12 nsew
rlabel metal5 1040 -960 1240 15760 0 gnda
port 13 nsew
rlabel metal5 1520 -960 1720 15760 0 vssa
port 14 nsew
<< end >>
