magic
tech sky130A
magscale 1 2
timestamp 1634821592
<< error_p >>
rect -317 692 -259 698
rect -317 658 -305 692
rect -317 652 -259 658
<< pwell >>
rect -439 -526 439 526
<< nmos >>
rect -351 -500 -321 500
rect -255 -500 -225 500
rect -159 -500 -129 500
rect -63 -500 -33 500
rect 33 -500 63 500
rect 129 -500 159 500
rect 225 -500 255 500
rect 321 -500 351 500
<< ndiff >>
rect -413 459 -351 500
rect -413 425 -401 459
rect -367 425 -351 459
rect -413 391 -351 425
rect -413 357 -401 391
rect -367 357 -351 391
rect -413 323 -351 357
rect -413 289 -401 323
rect -367 289 -351 323
rect -413 255 -351 289
rect -413 221 -401 255
rect -367 221 -351 255
rect -413 187 -351 221
rect -413 153 -401 187
rect -367 153 -351 187
rect -413 119 -351 153
rect -413 85 -401 119
rect -367 85 -351 119
rect -413 51 -351 85
rect -413 17 -401 51
rect -367 17 -351 51
rect -413 -17 -351 17
rect -413 -51 -401 -17
rect -367 -51 -351 -17
rect -413 -85 -351 -51
rect -413 -119 -401 -85
rect -367 -119 -351 -85
rect -413 -153 -351 -119
rect -413 -187 -401 -153
rect -367 -187 -351 -153
rect -413 -221 -351 -187
rect -413 -255 -401 -221
rect -367 -255 -351 -221
rect -413 -289 -351 -255
rect -413 -323 -401 -289
rect -367 -323 -351 -289
rect -413 -357 -351 -323
rect -413 -391 -401 -357
rect -367 -391 -351 -357
rect -413 -425 -351 -391
rect -413 -459 -401 -425
rect -367 -459 -351 -425
rect -413 -500 -351 -459
rect -321 459 -255 500
rect -321 425 -305 459
rect -271 425 -255 459
rect -321 391 -255 425
rect -321 357 -305 391
rect -271 357 -255 391
rect -321 323 -255 357
rect -321 289 -305 323
rect -271 289 -255 323
rect -321 255 -255 289
rect -321 221 -305 255
rect -271 221 -255 255
rect -321 187 -255 221
rect -321 153 -305 187
rect -271 153 -255 187
rect -321 119 -255 153
rect -321 85 -305 119
rect -271 85 -255 119
rect -321 51 -255 85
rect -321 17 -305 51
rect -271 17 -255 51
rect -321 -17 -255 17
rect -321 -51 -305 -17
rect -271 -51 -255 -17
rect -321 -85 -255 -51
rect -321 -119 -305 -85
rect -271 -119 -255 -85
rect -321 -153 -255 -119
rect -321 -187 -305 -153
rect -271 -187 -255 -153
rect -321 -221 -255 -187
rect -321 -255 -305 -221
rect -271 -255 -255 -221
rect -321 -289 -255 -255
rect -321 -323 -305 -289
rect -271 -323 -255 -289
rect -321 -357 -255 -323
rect -321 -391 -305 -357
rect -271 -391 -255 -357
rect -321 -425 -255 -391
rect -321 -459 -305 -425
rect -271 -459 -255 -425
rect -321 -500 -255 -459
rect -225 459 -159 500
rect -225 425 -209 459
rect -175 425 -159 459
rect -225 391 -159 425
rect -225 357 -209 391
rect -175 357 -159 391
rect -225 323 -159 357
rect -225 289 -209 323
rect -175 289 -159 323
rect -225 255 -159 289
rect -225 221 -209 255
rect -175 221 -159 255
rect -225 187 -159 221
rect -225 153 -209 187
rect -175 153 -159 187
rect -225 119 -159 153
rect -225 85 -209 119
rect -175 85 -159 119
rect -225 51 -159 85
rect -225 17 -209 51
rect -175 17 -159 51
rect -225 -17 -159 17
rect -225 -51 -209 -17
rect -175 -51 -159 -17
rect -225 -85 -159 -51
rect -225 -119 -209 -85
rect -175 -119 -159 -85
rect -225 -153 -159 -119
rect -225 -187 -209 -153
rect -175 -187 -159 -153
rect -225 -221 -159 -187
rect -225 -255 -209 -221
rect -175 -255 -159 -221
rect -225 -289 -159 -255
rect -225 -323 -209 -289
rect -175 -323 -159 -289
rect -225 -357 -159 -323
rect -225 -391 -209 -357
rect -175 -391 -159 -357
rect -225 -425 -159 -391
rect -225 -459 -209 -425
rect -175 -459 -159 -425
rect -225 -500 -159 -459
rect -129 459 -63 500
rect -129 425 -113 459
rect -79 425 -63 459
rect -129 391 -63 425
rect -129 357 -113 391
rect -79 357 -63 391
rect -129 323 -63 357
rect -129 289 -113 323
rect -79 289 -63 323
rect -129 255 -63 289
rect -129 221 -113 255
rect -79 221 -63 255
rect -129 187 -63 221
rect -129 153 -113 187
rect -79 153 -63 187
rect -129 119 -63 153
rect -129 85 -113 119
rect -79 85 -63 119
rect -129 51 -63 85
rect -129 17 -113 51
rect -79 17 -63 51
rect -129 -17 -63 17
rect -129 -51 -113 -17
rect -79 -51 -63 -17
rect -129 -85 -63 -51
rect -129 -119 -113 -85
rect -79 -119 -63 -85
rect -129 -153 -63 -119
rect -129 -187 -113 -153
rect -79 -187 -63 -153
rect -129 -221 -63 -187
rect -129 -255 -113 -221
rect -79 -255 -63 -221
rect -129 -289 -63 -255
rect -129 -323 -113 -289
rect -79 -323 -63 -289
rect -129 -357 -63 -323
rect -129 -391 -113 -357
rect -79 -391 -63 -357
rect -129 -425 -63 -391
rect -129 -459 -113 -425
rect -79 -459 -63 -425
rect -129 -500 -63 -459
rect -33 459 33 500
rect -33 425 -17 459
rect 17 425 33 459
rect -33 391 33 425
rect -33 357 -17 391
rect 17 357 33 391
rect -33 323 33 357
rect -33 289 -17 323
rect 17 289 33 323
rect -33 255 33 289
rect -33 221 -17 255
rect 17 221 33 255
rect -33 187 33 221
rect -33 153 -17 187
rect 17 153 33 187
rect -33 119 33 153
rect -33 85 -17 119
rect 17 85 33 119
rect -33 51 33 85
rect -33 17 -17 51
rect 17 17 33 51
rect -33 -17 33 17
rect -33 -51 -17 -17
rect 17 -51 33 -17
rect -33 -85 33 -51
rect -33 -119 -17 -85
rect 17 -119 33 -85
rect -33 -153 33 -119
rect -33 -187 -17 -153
rect 17 -187 33 -153
rect -33 -221 33 -187
rect -33 -255 -17 -221
rect 17 -255 33 -221
rect -33 -289 33 -255
rect -33 -323 -17 -289
rect 17 -323 33 -289
rect -33 -357 33 -323
rect -33 -391 -17 -357
rect 17 -391 33 -357
rect -33 -425 33 -391
rect -33 -459 -17 -425
rect 17 -459 33 -425
rect -33 -500 33 -459
rect 63 459 129 500
rect 63 425 79 459
rect 113 425 129 459
rect 63 391 129 425
rect 63 357 79 391
rect 113 357 129 391
rect 63 323 129 357
rect 63 289 79 323
rect 113 289 129 323
rect 63 255 129 289
rect 63 221 79 255
rect 113 221 129 255
rect 63 187 129 221
rect 63 153 79 187
rect 113 153 129 187
rect 63 119 129 153
rect 63 85 79 119
rect 113 85 129 119
rect 63 51 129 85
rect 63 17 79 51
rect 113 17 129 51
rect 63 -17 129 17
rect 63 -51 79 -17
rect 113 -51 129 -17
rect 63 -85 129 -51
rect 63 -119 79 -85
rect 113 -119 129 -85
rect 63 -153 129 -119
rect 63 -187 79 -153
rect 113 -187 129 -153
rect 63 -221 129 -187
rect 63 -255 79 -221
rect 113 -255 129 -221
rect 63 -289 129 -255
rect 63 -323 79 -289
rect 113 -323 129 -289
rect 63 -357 129 -323
rect 63 -391 79 -357
rect 113 -391 129 -357
rect 63 -425 129 -391
rect 63 -459 79 -425
rect 113 -459 129 -425
rect 63 -500 129 -459
rect 159 459 225 500
rect 159 425 175 459
rect 209 425 225 459
rect 159 391 225 425
rect 159 357 175 391
rect 209 357 225 391
rect 159 323 225 357
rect 159 289 175 323
rect 209 289 225 323
rect 159 255 225 289
rect 159 221 175 255
rect 209 221 225 255
rect 159 187 225 221
rect 159 153 175 187
rect 209 153 225 187
rect 159 119 225 153
rect 159 85 175 119
rect 209 85 225 119
rect 159 51 225 85
rect 159 17 175 51
rect 209 17 225 51
rect 159 -17 225 17
rect 159 -51 175 -17
rect 209 -51 225 -17
rect 159 -85 225 -51
rect 159 -119 175 -85
rect 209 -119 225 -85
rect 159 -153 225 -119
rect 159 -187 175 -153
rect 209 -187 225 -153
rect 159 -221 225 -187
rect 159 -255 175 -221
rect 209 -255 225 -221
rect 159 -289 225 -255
rect 159 -323 175 -289
rect 209 -323 225 -289
rect 159 -357 225 -323
rect 159 -391 175 -357
rect 209 -391 225 -357
rect 159 -425 225 -391
rect 159 -459 175 -425
rect 209 -459 225 -425
rect 159 -500 225 -459
rect 255 459 321 500
rect 255 425 271 459
rect 305 425 321 459
rect 255 391 321 425
rect 255 357 271 391
rect 305 357 321 391
rect 255 323 321 357
rect 255 289 271 323
rect 305 289 321 323
rect 255 255 321 289
rect 255 221 271 255
rect 305 221 321 255
rect 255 187 321 221
rect 255 153 271 187
rect 305 153 321 187
rect 255 119 321 153
rect 255 85 271 119
rect 305 85 321 119
rect 255 51 321 85
rect 255 17 271 51
rect 305 17 321 51
rect 255 -17 321 17
rect 255 -51 271 -17
rect 305 -51 321 -17
rect 255 -85 321 -51
rect 255 -119 271 -85
rect 305 -119 321 -85
rect 255 -153 321 -119
rect 255 -187 271 -153
rect 305 -187 321 -153
rect 255 -221 321 -187
rect 255 -255 271 -221
rect 305 -255 321 -221
rect 255 -289 321 -255
rect 255 -323 271 -289
rect 305 -323 321 -289
rect 255 -357 321 -323
rect 255 -391 271 -357
rect 305 -391 321 -357
rect 255 -425 321 -391
rect 255 -459 271 -425
rect 305 -459 321 -425
rect 255 -500 321 -459
rect 351 459 413 500
rect 351 425 367 459
rect 401 425 413 459
rect 351 391 413 425
rect 351 357 367 391
rect 401 357 413 391
rect 351 323 413 357
rect 351 289 367 323
rect 401 289 413 323
rect 351 255 413 289
rect 351 221 367 255
rect 401 221 413 255
rect 351 187 413 221
rect 351 153 367 187
rect 401 153 413 187
rect 351 119 413 153
rect 351 85 367 119
rect 401 85 413 119
rect 351 51 413 85
rect 351 17 367 51
rect 401 17 413 51
rect 351 -17 413 17
rect 351 -51 367 -17
rect 401 -51 413 -17
rect 351 -85 413 -51
rect 351 -119 367 -85
rect 401 -119 413 -85
rect 351 -153 413 -119
rect 351 -187 367 -153
rect 401 -187 413 -153
rect 351 -221 413 -187
rect 351 -255 367 -221
rect 401 -255 413 -221
rect 351 -289 413 -255
rect 351 -323 367 -289
rect 401 -323 413 -289
rect 351 -357 413 -323
rect 351 -391 367 -357
rect 401 -391 413 -357
rect 351 -425 413 -391
rect 351 -459 367 -425
rect 401 -459 413 -425
rect 351 -500 413 -459
<< ndiffc >>
rect -401 425 -367 459
rect -401 357 -367 391
rect -401 289 -367 323
rect -401 221 -367 255
rect -401 153 -367 187
rect -401 85 -367 119
rect -401 17 -367 51
rect -401 -51 -367 -17
rect -401 -119 -367 -85
rect -401 -187 -367 -153
rect -401 -255 -367 -221
rect -401 -323 -367 -289
rect -401 -391 -367 -357
rect -401 -459 -367 -425
rect -305 425 -271 459
rect -305 357 -271 391
rect -305 289 -271 323
rect -305 221 -271 255
rect -305 153 -271 187
rect -305 85 -271 119
rect -305 17 -271 51
rect -305 -51 -271 -17
rect -305 -119 -271 -85
rect -305 -187 -271 -153
rect -305 -255 -271 -221
rect -305 -323 -271 -289
rect -305 -391 -271 -357
rect -305 -459 -271 -425
rect -209 425 -175 459
rect -209 357 -175 391
rect -209 289 -175 323
rect -209 221 -175 255
rect -209 153 -175 187
rect -209 85 -175 119
rect -209 17 -175 51
rect -209 -51 -175 -17
rect -209 -119 -175 -85
rect -209 -187 -175 -153
rect -209 -255 -175 -221
rect -209 -323 -175 -289
rect -209 -391 -175 -357
rect -209 -459 -175 -425
rect -113 425 -79 459
rect -113 357 -79 391
rect -113 289 -79 323
rect -113 221 -79 255
rect -113 153 -79 187
rect -113 85 -79 119
rect -113 17 -79 51
rect -113 -51 -79 -17
rect -113 -119 -79 -85
rect -113 -187 -79 -153
rect -113 -255 -79 -221
rect -113 -323 -79 -289
rect -113 -391 -79 -357
rect -113 -459 -79 -425
rect -17 425 17 459
rect -17 357 17 391
rect -17 289 17 323
rect -17 221 17 255
rect -17 153 17 187
rect -17 85 17 119
rect -17 17 17 51
rect -17 -51 17 -17
rect -17 -119 17 -85
rect -17 -187 17 -153
rect -17 -255 17 -221
rect -17 -323 17 -289
rect -17 -391 17 -357
rect -17 -459 17 -425
rect 79 425 113 459
rect 79 357 113 391
rect 79 289 113 323
rect 79 221 113 255
rect 79 153 113 187
rect 79 85 113 119
rect 79 17 113 51
rect 79 -51 113 -17
rect 79 -119 113 -85
rect 79 -187 113 -153
rect 79 -255 113 -221
rect 79 -323 113 -289
rect 79 -391 113 -357
rect 79 -459 113 -425
rect 175 425 209 459
rect 175 357 209 391
rect 175 289 209 323
rect 175 221 209 255
rect 175 153 209 187
rect 175 85 209 119
rect 175 17 209 51
rect 175 -51 209 -17
rect 175 -119 209 -85
rect 175 -187 209 -153
rect 175 -255 209 -221
rect 175 -323 209 -289
rect 175 -391 209 -357
rect 175 -459 209 -425
rect 271 425 305 459
rect 271 357 305 391
rect 271 289 305 323
rect 271 221 305 255
rect 271 153 305 187
rect 271 85 305 119
rect 271 17 305 51
rect 271 -51 305 -17
rect 271 -119 305 -85
rect 271 -187 305 -153
rect 271 -255 305 -221
rect 271 -323 305 -289
rect 271 -391 305 -357
rect 271 -459 305 -425
rect 367 425 401 459
rect 367 357 401 391
rect 367 289 401 323
rect 367 221 401 255
rect 367 153 401 187
rect 367 85 401 119
rect 367 17 401 51
rect 367 -51 401 -17
rect 367 -119 401 -85
rect 367 -187 401 -153
rect 367 -255 401 -221
rect 367 -323 401 -289
rect 367 -391 401 -357
rect 367 -459 401 -425
<< poly >>
rect -321 692 -255 708
rect -321 658 -305 692
rect -271 658 -255 692
rect -321 642 -255 658
rect -305 600 -275 642
rect -351 564 351 600
rect -351 500 -321 564
rect -255 500 -225 564
rect -159 500 -129 564
rect -63 500 -33 564
rect 33 500 63 564
rect 129 500 159 564
rect 225 500 255 564
rect 321 500 351 564
rect -351 -526 -321 -500
rect -255 -526 -225 -500
rect -159 -526 -129 -500
rect -63 -526 -33 -500
rect 33 -526 63 -500
rect 129 -526 159 -500
rect 225 -526 255 -500
rect 321 -526 351 -500
<< polycont >>
rect -305 658 -271 692
<< locali >>
rect -321 658 -305 692
rect -271 658 -255 692
rect -305 554 305 588
rect -401 485 -367 504
rect -401 413 -367 425
rect -401 341 -367 357
rect -401 269 -367 289
rect -401 197 -367 221
rect -401 125 -367 153
rect -401 53 -367 85
rect -401 -17 -367 17
rect -401 -85 -367 -53
rect -401 -153 -367 -125
rect -401 -221 -367 -197
rect -401 -289 -367 -269
rect -401 -357 -367 -341
rect -401 -425 -367 -413
rect -401 -564 -367 -485
rect -305 485 -271 554
rect -305 413 -271 425
rect -305 341 -271 357
rect -305 269 -271 289
rect -305 197 -271 221
rect -305 125 -271 153
rect -305 53 -271 85
rect -305 -17 -271 17
rect -305 -85 -271 -53
rect -305 -153 -271 -125
rect -305 -221 -271 -197
rect -305 -289 -271 -269
rect -305 -357 -271 -341
rect -305 -425 -271 -413
rect -305 -504 -271 -485
rect -209 485 -175 504
rect -209 413 -175 425
rect -209 341 -175 357
rect -209 269 -175 289
rect -209 197 -175 221
rect -209 125 -175 153
rect -209 53 -175 85
rect -209 -17 -175 17
rect -209 -85 -175 -53
rect -209 -153 -175 -125
rect -209 -221 -175 -197
rect -209 -289 -175 -269
rect -209 -357 -175 -341
rect -209 -425 -175 -413
rect -209 -564 -175 -485
rect -113 485 -79 554
rect -113 413 -79 425
rect -113 341 -79 357
rect -113 269 -79 289
rect -113 197 -79 221
rect -113 125 -79 153
rect -113 53 -79 85
rect -113 -17 -79 17
rect -113 -85 -79 -53
rect -113 -153 -79 -125
rect -113 -221 -79 -197
rect -113 -289 -79 -269
rect -113 -357 -79 -341
rect -113 -425 -79 -413
rect -113 -504 -79 -485
rect -17 485 17 504
rect -17 413 17 425
rect -17 341 17 357
rect -17 269 17 289
rect -17 197 17 221
rect -17 125 17 153
rect -17 53 17 85
rect -17 -17 17 17
rect -17 -85 17 -53
rect -17 -153 17 -125
rect -17 -221 17 -197
rect -17 -289 17 -269
rect -17 -357 17 -341
rect -17 -425 17 -413
rect -17 -564 17 -485
rect 79 485 113 554
rect 79 413 113 425
rect 79 341 113 357
rect 79 269 113 289
rect 79 197 113 221
rect 79 125 113 153
rect 79 53 113 85
rect 79 -17 113 17
rect 79 -85 113 -53
rect 79 -153 113 -125
rect 79 -221 113 -197
rect 79 -289 113 -269
rect 79 -357 113 -341
rect 79 -425 113 -413
rect 79 -504 113 -485
rect 175 485 209 504
rect 175 413 209 425
rect 175 341 209 357
rect 175 269 209 289
rect 175 197 209 221
rect 175 125 209 153
rect 175 53 209 85
rect 175 -17 209 17
rect 175 -85 209 -53
rect 175 -153 209 -125
rect 175 -221 209 -197
rect 175 -289 209 -269
rect 175 -357 209 -341
rect 175 -425 209 -413
rect 175 -564 209 -485
rect 271 485 305 554
rect 271 413 305 425
rect 271 341 305 357
rect 271 269 305 289
rect 271 197 305 221
rect 271 125 305 153
rect 271 53 305 85
rect 271 -17 305 17
rect 271 -85 305 -53
rect 271 -153 305 -125
rect 271 -221 305 -197
rect 271 -289 305 -269
rect 271 -357 305 -341
rect 271 -425 305 -413
rect 271 -504 305 -485
rect 367 485 401 504
rect 367 413 401 425
rect 367 341 401 357
rect 367 269 401 289
rect 367 197 401 221
rect 367 125 401 153
rect 367 53 401 85
rect 367 -17 401 17
rect 367 -85 401 -53
rect 367 -153 401 -125
rect 367 -221 401 -197
rect 367 -289 401 -269
rect 367 -357 401 -341
rect 367 -425 401 -413
rect 367 -564 401 -485
rect -401 -598 401 -564
<< viali >>
rect -305 658 -271 692
rect -401 459 -367 485
rect -401 451 -367 459
rect -401 391 -367 413
rect -401 379 -367 391
rect -401 323 -367 341
rect -401 307 -367 323
rect -401 255 -367 269
rect -401 235 -367 255
rect -401 187 -367 197
rect -401 163 -367 187
rect -401 119 -367 125
rect -401 91 -367 119
rect -401 51 -367 53
rect -401 19 -367 51
rect -401 -51 -367 -19
rect -401 -53 -367 -51
rect -401 -119 -367 -91
rect -401 -125 -367 -119
rect -401 -187 -367 -163
rect -401 -197 -367 -187
rect -401 -255 -367 -235
rect -401 -269 -367 -255
rect -401 -323 -367 -307
rect -401 -341 -367 -323
rect -401 -391 -367 -379
rect -401 -413 -367 -391
rect -401 -459 -367 -451
rect -401 -485 -367 -459
rect -305 459 -271 485
rect -305 451 -271 459
rect -305 391 -271 413
rect -305 379 -271 391
rect -305 323 -271 341
rect -305 307 -271 323
rect -305 255 -271 269
rect -305 235 -271 255
rect -305 187 -271 197
rect -305 163 -271 187
rect -305 119 -271 125
rect -305 91 -271 119
rect -305 51 -271 53
rect -305 19 -271 51
rect -305 -51 -271 -19
rect -305 -53 -271 -51
rect -305 -119 -271 -91
rect -305 -125 -271 -119
rect -305 -187 -271 -163
rect -305 -197 -271 -187
rect -305 -255 -271 -235
rect -305 -269 -271 -255
rect -305 -323 -271 -307
rect -305 -341 -271 -323
rect -305 -391 -271 -379
rect -305 -413 -271 -391
rect -305 -459 -271 -451
rect -305 -485 -271 -459
rect -209 459 -175 485
rect -209 451 -175 459
rect -209 391 -175 413
rect -209 379 -175 391
rect -209 323 -175 341
rect -209 307 -175 323
rect -209 255 -175 269
rect -209 235 -175 255
rect -209 187 -175 197
rect -209 163 -175 187
rect -209 119 -175 125
rect -209 91 -175 119
rect -209 51 -175 53
rect -209 19 -175 51
rect -209 -51 -175 -19
rect -209 -53 -175 -51
rect -209 -119 -175 -91
rect -209 -125 -175 -119
rect -209 -187 -175 -163
rect -209 -197 -175 -187
rect -209 -255 -175 -235
rect -209 -269 -175 -255
rect -209 -323 -175 -307
rect -209 -341 -175 -323
rect -209 -391 -175 -379
rect -209 -413 -175 -391
rect -209 -459 -175 -451
rect -209 -485 -175 -459
rect -113 459 -79 485
rect -113 451 -79 459
rect -113 391 -79 413
rect -113 379 -79 391
rect -113 323 -79 341
rect -113 307 -79 323
rect -113 255 -79 269
rect -113 235 -79 255
rect -113 187 -79 197
rect -113 163 -79 187
rect -113 119 -79 125
rect -113 91 -79 119
rect -113 51 -79 53
rect -113 19 -79 51
rect -113 -51 -79 -19
rect -113 -53 -79 -51
rect -113 -119 -79 -91
rect -113 -125 -79 -119
rect -113 -187 -79 -163
rect -113 -197 -79 -187
rect -113 -255 -79 -235
rect -113 -269 -79 -255
rect -113 -323 -79 -307
rect -113 -341 -79 -323
rect -113 -391 -79 -379
rect -113 -413 -79 -391
rect -113 -459 -79 -451
rect -113 -485 -79 -459
rect -17 459 17 485
rect -17 451 17 459
rect -17 391 17 413
rect -17 379 17 391
rect -17 323 17 341
rect -17 307 17 323
rect -17 255 17 269
rect -17 235 17 255
rect -17 187 17 197
rect -17 163 17 187
rect -17 119 17 125
rect -17 91 17 119
rect -17 51 17 53
rect -17 19 17 51
rect -17 -51 17 -19
rect -17 -53 17 -51
rect -17 -119 17 -91
rect -17 -125 17 -119
rect -17 -187 17 -163
rect -17 -197 17 -187
rect -17 -255 17 -235
rect -17 -269 17 -255
rect -17 -323 17 -307
rect -17 -341 17 -323
rect -17 -391 17 -379
rect -17 -413 17 -391
rect -17 -459 17 -451
rect -17 -485 17 -459
rect 79 459 113 485
rect 79 451 113 459
rect 79 391 113 413
rect 79 379 113 391
rect 79 323 113 341
rect 79 307 113 323
rect 79 255 113 269
rect 79 235 113 255
rect 79 187 113 197
rect 79 163 113 187
rect 79 119 113 125
rect 79 91 113 119
rect 79 51 113 53
rect 79 19 113 51
rect 79 -51 113 -19
rect 79 -53 113 -51
rect 79 -119 113 -91
rect 79 -125 113 -119
rect 79 -187 113 -163
rect 79 -197 113 -187
rect 79 -255 113 -235
rect 79 -269 113 -255
rect 79 -323 113 -307
rect 79 -341 113 -323
rect 79 -391 113 -379
rect 79 -413 113 -391
rect 79 -459 113 -451
rect 79 -485 113 -459
rect 175 459 209 485
rect 175 451 209 459
rect 175 391 209 413
rect 175 379 209 391
rect 175 323 209 341
rect 175 307 209 323
rect 175 255 209 269
rect 175 235 209 255
rect 175 187 209 197
rect 175 163 209 187
rect 175 119 209 125
rect 175 91 209 119
rect 175 51 209 53
rect 175 19 209 51
rect 175 -51 209 -19
rect 175 -53 209 -51
rect 175 -119 209 -91
rect 175 -125 209 -119
rect 175 -187 209 -163
rect 175 -197 209 -187
rect 175 -255 209 -235
rect 175 -269 209 -255
rect 175 -323 209 -307
rect 175 -341 209 -323
rect 175 -391 209 -379
rect 175 -413 209 -391
rect 175 -459 209 -451
rect 175 -485 209 -459
rect 271 459 305 485
rect 271 451 305 459
rect 271 391 305 413
rect 271 379 305 391
rect 271 323 305 341
rect 271 307 305 323
rect 271 255 305 269
rect 271 235 305 255
rect 271 187 305 197
rect 271 163 305 187
rect 271 119 305 125
rect 271 91 305 119
rect 271 51 305 53
rect 271 19 305 51
rect 271 -51 305 -19
rect 271 -53 305 -51
rect 271 -119 305 -91
rect 271 -125 305 -119
rect 271 -187 305 -163
rect 271 -197 305 -187
rect 271 -255 305 -235
rect 271 -269 305 -255
rect 271 -323 305 -307
rect 271 -341 305 -323
rect 271 -391 305 -379
rect 271 -413 305 -391
rect 271 -459 305 -451
rect 271 -485 305 -459
rect 367 459 401 485
rect 367 451 401 459
rect 367 391 401 413
rect 367 379 401 391
rect 367 323 401 341
rect 367 307 401 323
rect 367 255 401 269
rect 367 235 401 255
rect 367 187 401 197
rect 367 163 401 187
rect 367 119 401 125
rect 367 91 401 119
rect 367 51 401 53
rect 367 19 401 51
rect 367 -51 401 -19
rect 367 -53 401 -51
rect 367 -119 401 -91
rect 367 -125 401 -119
rect 367 -187 401 -163
rect 367 -197 401 -187
rect 367 -255 401 -235
rect 367 -269 401 -255
rect 367 -323 401 -307
rect 367 -341 401 -323
rect 367 -391 401 -379
rect 367 -413 401 -391
rect 367 -459 401 -451
rect 367 -485 401 -459
<< metal1 >>
rect -317 692 -259 698
rect -317 658 -305 692
rect -271 658 -259 692
rect -317 652 -259 658
rect -407 485 -361 500
rect -407 451 -401 485
rect -367 451 -361 485
rect -407 413 -361 451
rect -407 379 -401 413
rect -367 379 -361 413
rect -407 341 -361 379
rect -407 307 -401 341
rect -367 307 -361 341
rect -407 269 -361 307
rect -407 235 -401 269
rect -367 235 -361 269
rect -407 197 -361 235
rect -407 163 -401 197
rect -367 163 -361 197
rect -407 125 -361 163
rect -407 91 -401 125
rect -367 91 -361 125
rect -407 53 -361 91
rect -407 19 -401 53
rect -367 19 -361 53
rect -407 -19 -361 19
rect -407 -53 -401 -19
rect -367 -53 -361 -19
rect -407 -91 -361 -53
rect -407 -125 -401 -91
rect -367 -125 -361 -91
rect -407 -163 -361 -125
rect -407 -197 -401 -163
rect -367 -197 -361 -163
rect -407 -235 -361 -197
rect -407 -269 -401 -235
rect -367 -269 -361 -235
rect -407 -307 -361 -269
rect -407 -341 -401 -307
rect -367 -341 -361 -307
rect -407 -379 -361 -341
rect -407 -413 -401 -379
rect -367 -413 -361 -379
rect -407 -451 -361 -413
rect -407 -485 -401 -451
rect -367 -485 -361 -451
rect -407 -500 -361 -485
rect -311 485 -265 500
rect -311 451 -305 485
rect -271 451 -265 485
rect -311 413 -265 451
rect -311 379 -305 413
rect -271 379 -265 413
rect -311 341 -265 379
rect -311 307 -305 341
rect -271 307 -265 341
rect -311 269 -265 307
rect -311 235 -305 269
rect -271 235 -265 269
rect -311 197 -265 235
rect -311 163 -305 197
rect -271 163 -265 197
rect -311 125 -265 163
rect -311 91 -305 125
rect -271 91 -265 125
rect -311 53 -265 91
rect -311 19 -305 53
rect -271 19 -265 53
rect -311 -19 -265 19
rect -311 -53 -305 -19
rect -271 -53 -265 -19
rect -311 -91 -265 -53
rect -311 -125 -305 -91
rect -271 -125 -265 -91
rect -311 -163 -265 -125
rect -311 -197 -305 -163
rect -271 -197 -265 -163
rect -311 -235 -265 -197
rect -311 -269 -305 -235
rect -271 -269 -265 -235
rect -311 -307 -265 -269
rect -311 -341 -305 -307
rect -271 -341 -265 -307
rect -311 -379 -265 -341
rect -311 -413 -305 -379
rect -271 -413 -265 -379
rect -311 -451 -265 -413
rect -311 -485 -305 -451
rect -271 -485 -265 -451
rect -311 -500 -265 -485
rect -215 485 -169 500
rect -215 451 -209 485
rect -175 451 -169 485
rect -215 413 -169 451
rect -215 379 -209 413
rect -175 379 -169 413
rect -215 341 -169 379
rect -215 307 -209 341
rect -175 307 -169 341
rect -215 269 -169 307
rect -215 235 -209 269
rect -175 235 -169 269
rect -215 197 -169 235
rect -215 163 -209 197
rect -175 163 -169 197
rect -215 125 -169 163
rect -215 91 -209 125
rect -175 91 -169 125
rect -215 53 -169 91
rect -215 19 -209 53
rect -175 19 -169 53
rect -215 -19 -169 19
rect -215 -53 -209 -19
rect -175 -53 -169 -19
rect -215 -91 -169 -53
rect -215 -125 -209 -91
rect -175 -125 -169 -91
rect -215 -163 -169 -125
rect -215 -197 -209 -163
rect -175 -197 -169 -163
rect -215 -235 -169 -197
rect -215 -269 -209 -235
rect -175 -269 -169 -235
rect -215 -307 -169 -269
rect -215 -341 -209 -307
rect -175 -341 -169 -307
rect -215 -379 -169 -341
rect -215 -413 -209 -379
rect -175 -413 -169 -379
rect -215 -451 -169 -413
rect -215 -485 -209 -451
rect -175 -485 -169 -451
rect -215 -500 -169 -485
rect -119 485 -73 500
rect -119 451 -113 485
rect -79 451 -73 485
rect -119 413 -73 451
rect -119 379 -113 413
rect -79 379 -73 413
rect -119 341 -73 379
rect -119 307 -113 341
rect -79 307 -73 341
rect -119 269 -73 307
rect -119 235 -113 269
rect -79 235 -73 269
rect -119 197 -73 235
rect -119 163 -113 197
rect -79 163 -73 197
rect -119 125 -73 163
rect -119 91 -113 125
rect -79 91 -73 125
rect -119 53 -73 91
rect -119 19 -113 53
rect -79 19 -73 53
rect -119 -19 -73 19
rect -119 -53 -113 -19
rect -79 -53 -73 -19
rect -119 -91 -73 -53
rect -119 -125 -113 -91
rect -79 -125 -73 -91
rect -119 -163 -73 -125
rect -119 -197 -113 -163
rect -79 -197 -73 -163
rect -119 -235 -73 -197
rect -119 -269 -113 -235
rect -79 -269 -73 -235
rect -119 -307 -73 -269
rect -119 -341 -113 -307
rect -79 -341 -73 -307
rect -119 -379 -73 -341
rect -119 -413 -113 -379
rect -79 -413 -73 -379
rect -119 -451 -73 -413
rect -119 -485 -113 -451
rect -79 -485 -73 -451
rect -119 -500 -73 -485
rect -23 485 23 500
rect -23 451 -17 485
rect 17 451 23 485
rect -23 413 23 451
rect -23 379 -17 413
rect 17 379 23 413
rect -23 341 23 379
rect -23 307 -17 341
rect 17 307 23 341
rect -23 269 23 307
rect -23 235 -17 269
rect 17 235 23 269
rect -23 197 23 235
rect -23 163 -17 197
rect 17 163 23 197
rect -23 125 23 163
rect -23 91 -17 125
rect 17 91 23 125
rect -23 53 23 91
rect -23 19 -17 53
rect 17 19 23 53
rect -23 -19 23 19
rect -23 -53 -17 -19
rect 17 -53 23 -19
rect -23 -91 23 -53
rect -23 -125 -17 -91
rect 17 -125 23 -91
rect -23 -163 23 -125
rect -23 -197 -17 -163
rect 17 -197 23 -163
rect -23 -235 23 -197
rect -23 -269 -17 -235
rect 17 -269 23 -235
rect -23 -307 23 -269
rect -23 -341 -17 -307
rect 17 -341 23 -307
rect -23 -379 23 -341
rect -23 -413 -17 -379
rect 17 -413 23 -379
rect -23 -451 23 -413
rect -23 -485 -17 -451
rect 17 -485 23 -451
rect -23 -500 23 -485
rect 73 485 119 500
rect 73 451 79 485
rect 113 451 119 485
rect 73 413 119 451
rect 73 379 79 413
rect 113 379 119 413
rect 73 341 119 379
rect 73 307 79 341
rect 113 307 119 341
rect 73 269 119 307
rect 73 235 79 269
rect 113 235 119 269
rect 73 197 119 235
rect 73 163 79 197
rect 113 163 119 197
rect 73 125 119 163
rect 73 91 79 125
rect 113 91 119 125
rect 73 53 119 91
rect 73 19 79 53
rect 113 19 119 53
rect 73 -19 119 19
rect 73 -53 79 -19
rect 113 -53 119 -19
rect 73 -91 119 -53
rect 73 -125 79 -91
rect 113 -125 119 -91
rect 73 -163 119 -125
rect 73 -197 79 -163
rect 113 -197 119 -163
rect 73 -235 119 -197
rect 73 -269 79 -235
rect 113 -269 119 -235
rect 73 -307 119 -269
rect 73 -341 79 -307
rect 113 -341 119 -307
rect 73 -379 119 -341
rect 73 -413 79 -379
rect 113 -413 119 -379
rect 73 -451 119 -413
rect 73 -485 79 -451
rect 113 -485 119 -451
rect 73 -500 119 -485
rect 169 485 215 500
rect 169 451 175 485
rect 209 451 215 485
rect 169 413 215 451
rect 169 379 175 413
rect 209 379 215 413
rect 169 341 215 379
rect 169 307 175 341
rect 209 307 215 341
rect 169 269 215 307
rect 169 235 175 269
rect 209 235 215 269
rect 169 197 215 235
rect 169 163 175 197
rect 209 163 215 197
rect 169 125 215 163
rect 169 91 175 125
rect 209 91 215 125
rect 169 53 215 91
rect 169 19 175 53
rect 209 19 215 53
rect 169 -19 215 19
rect 169 -53 175 -19
rect 209 -53 215 -19
rect 169 -91 215 -53
rect 169 -125 175 -91
rect 209 -125 215 -91
rect 169 -163 215 -125
rect 169 -197 175 -163
rect 209 -197 215 -163
rect 169 -235 215 -197
rect 169 -269 175 -235
rect 209 -269 215 -235
rect 169 -307 215 -269
rect 169 -341 175 -307
rect 209 -341 215 -307
rect 169 -379 215 -341
rect 169 -413 175 -379
rect 209 -413 215 -379
rect 169 -451 215 -413
rect 169 -485 175 -451
rect 209 -485 215 -451
rect 169 -500 215 -485
rect 265 485 311 500
rect 265 451 271 485
rect 305 451 311 485
rect 265 413 311 451
rect 265 379 271 413
rect 305 379 311 413
rect 265 341 311 379
rect 265 307 271 341
rect 305 307 311 341
rect 265 269 311 307
rect 265 235 271 269
rect 305 235 311 269
rect 265 197 311 235
rect 265 163 271 197
rect 305 163 311 197
rect 265 125 311 163
rect 265 91 271 125
rect 305 91 311 125
rect 265 53 311 91
rect 265 19 271 53
rect 305 19 311 53
rect 265 -19 311 19
rect 265 -53 271 -19
rect 305 -53 311 -19
rect 265 -91 311 -53
rect 265 -125 271 -91
rect 305 -125 311 -91
rect 265 -163 311 -125
rect 265 -197 271 -163
rect 305 -197 311 -163
rect 265 -235 311 -197
rect 265 -269 271 -235
rect 305 -269 311 -235
rect 265 -307 311 -269
rect 265 -341 271 -307
rect 305 -341 311 -307
rect 265 -379 311 -341
rect 265 -413 271 -379
rect 305 -413 311 -379
rect 265 -451 311 -413
rect 265 -485 271 -451
rect 305 -485 311 -451
rect 265 -500 311 -485
rect 361 485 407 500
rect 361 451 367 485
rect 401 451 407 485
rect 361 413 407 451
rect 361 379 367 413
rect 401 379 407 413
rect 361 341 407 379
rect 361 307 367 341
rect 401 307 407 341
rect 361 269 407 307
rect 361 235 367 269
rect 401 235 407 269
rect 361 197 407 235
rect 361 163 367 197
rect 401 163 407 197
rect 361 125 407 163
rect 361 91 367 125
rect 401 91 407 125
rect 361 53 407 91
rect 361 19 367 53
rect 401 19 407 53
rect 361 -19 407 19
rect 361 -53 367 -19
rect 401 -53 407 -19
rect 361 -91 407 -53
rect 361 -125 367 -91
rect 401 -125 407 -91
rect 361 -163 407 -125
rect 361 -197 367 -163
rect 401 -197 407 -163
rect 361 -235 407 -197
rect 361 -269 367 -235
rect 401 -269 407 -235
rect 361 -307 407 -269
rect 361 -341 367 -307
rect 401 -341 407 -307
rect 361 -379 407 -341
rect 361 -413 367 -379
rect 401 -413 407 -379
rect 361 -451 407 -413
rect 361 -485 367 -451
rect 401 -485 407 -451
rect 361 -500 407 -485
<< end >>
