magic
tech sky130A
magscale 1 2
timestamp 1634765323
<< nwell >>
rect 1420 -510 1850 -320
rect 1530 -550 1610 -510
rect 1500 -640 1740 -550
rect 1530 -700 1610 -640
rect 1480 -960 1610 -700
rect 1660 -1100 1760 -880
<< pwell >>
rect 710 -1000 900 -990
rect 710 -1010 910 -1000
rect 760 -1050 910 -1010
rect 700 -1200 790 -1110
rect 710 -1240 790 -1200
<< metal1 >>
rect 700 520 900 610
rect 480 300 980 520
rect 1930 380 2130 420
rect 480 150 600 300
rect 1540 270 2130 380
rect 780 190 840 250
rect 480 -110 790 150
rect 1540 120 1630 270
rect 1930 220 2130 270
rect 1660 150 1720 210
rect 1530 100 1660 120
rect 1530 40 1560 100
rect 1620 40 1660 100
rect 1530 20 1660 40
rect 1720 -50 2010 50
rect 1650 -170 1740 -110
rect 840 -390 1740 -170
rect 840 -420 1190 -390
rect 710 -650 910 -490
rect 440 -690 910 -650
rect 440 -820 750 -690
rect 880 -820 910 -690
rect 440 -850 910 -820
rect 710 -1060 910 -850
rect 1030 -1110 1190 -420
rect 1230 -510 1410 -490
rect 1230 -530 1740 -510
rect 1230 -620 1260 -530
rect 1370 -600 1740 -530
rect 1370 -620 1410 -600
rect 1230 -650 1410 -620
rect 1500 -640 1740 -600
rect 1480 -740 1610 -700
rect 1480 -930 1510 -740
rect 1590 -930 1610 -740
rect 1920 -880 2010 -50
rect 1480 -960 1610 -930
rect 1660 -1100 2010 -880
rect 440 -1240 790 -1110
rect 440 -1310 720 -1240
rect 830 -1250 1190 -1110
rect 1830 -1188 2010 -1100
rect 640 -1430 720 -1310
rect 1830 -1280 2006 -1188
rect 780 -1390 850 -1330
rect 1610 -1390 1670 -1320
rect 1830 -1430 2126 -1280
rect 640 -1500 1000 -1430
rect 1540 -1480 2126 -1430
<< via1 >>
rect 1560 40 1620 100
rect 750 -820 880 -690
rect 1260 -620 1370 -530
rect 1510 -930 1590 -740
<< metal2 >>
rect 1530 100 1630 120
rect 1530 40 1560 100
rect 1620 40 1630 100
rect 1530 20 1630 40
rect 1230 -530 1410 -490
rect 1230 -620 1260 -530
rect 1370 -620 1410 -530
rect 1230 -650 1410 -620
rect 700 -690 1410 -650
rect 700 -820 750 -690
rect 880 -820 1410 -690
rect 1530 -700 1610 20
rect 700 -850 1410 -820
rect 1480 -740 1610 -700
rect 1480 -930 1510 -740
rect 1590 -930 1610 -740
rect 1480 -960 1610 -930
use sky130_fd_pr__pfet_01v8_4J4M39  XM2
timestamp 1634485485
transform 1 0 811 0 1 -141
box -211 -519 211 519
use sky130_fd_pr__nfet_01v8_V3CPBF  XM1
timestamp 1634512638
transform 1 0 811 0 1 -1200
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_RJZS2S  XM4
timestamp 1634512638
transform 1 0 1638 0 1 -994
box -211 -519 211 519
use sky130_fd_pr__nfet_01v8_ZBX7X9  XM3
timestamp 1634485485
transform -1 0 1691 0 -1 30
box -211 -310 211 310
<< labels >>
flabel metal1 440 -850 640 -650 0 FreeSans 256 0 0 0 ctrl
port 2 nsew
flabel metal1 1930 220 2130 420 0 FreeSans 256 0 0 0 a
port 5 nsew
flabel metal1 440 -1310 640 -1110 0 FreeSans 256 0 0 0 vgnd
port 3 nsew
flabel metal1 700 410 900 610 5 FreeSans 256 0 0 0 vs
port 1 nsew
flabel metal1 1926 -1480 2126 -1280 0 FreeSans 256 0 0 0 b
port 4 nsew
<< end >>
