magic
tech sky130A
magscale 1 2
timestamp 1635533344
<< checkpaint >>
rect 10412 16858 13334 30410
rect -124 10984 4020 13010
rect -124 8880 6300 10984
rect 2128 7440 6300 8880
rect 2128 6300 5240 7440
<< metal1 >>
rect 40 53160 420 53520
rect 80 52660 360 53160
rect 4440 53100 4820 53460
rect 8840 53100 9220 53460
rect 13260 53100 13640 53460
rect 80 52480 140 52660
rect 300 52480 360 52660
rect 80 52380 360 52480
rect 4500 52660 4780 53100
rect 4500 52480 4540 52660
rect 4700 52480 4780 52660
rect 4500 52380 4780 52480
rect 8940 52640 9160 53100
rect 8940 52460 8980 52640
rect 9140 52460 9160 52640
rect 8940 52420 9160 52460
rect 13340 52680 13560 53100
rect 13340 52500 13380 52680
rect 13540 52500 13560 52680
rect 13340 52440 13560 52500
rect -5720 39970 -5340 40010
rect -5720 39830 -2460 39970
rect -5720 39800 -880 39830
rect -5720 39670 -2460 39800
rect -930 39790 -900 39800
rect -5720 39650 -5340 39670
rect -5720 37560 -5340 37580
rect -5720 37520 -960 37560
rect -5720 37260 -1270 37520
rect -1030 37260 -960 37520
rect -5720 37240 -960 37260
rect -5720 37220 -5340 37240
rect 7900 33040 8100 33100
rect 1280 33000 1500 33040
rect -920 32960 -740 33000
rect -920 32800 -880 32960
rect -780 32800 -740 32960
rect -920 32080 -740 32800
rect 1280 32800 1320 33000
rect 1460 32800 1500 33000
rect 5660 32960 5880 33020
rect 1280 32060 1500 32800
rect 3420 32920 3640 32960
rect 3420 32720 3460 32920
rect 3600 32720 3640 32920
rect 5660 32760 5700 32960
rect 3420 32240 3640 32720
rect 5680 32700 5700 32760
rect 5860 32700 5880 32960
rect 3420 31840 3660 32240
rect 5680 31740 5880 32700
rect 7900 32780 7940 33040
rect 8060 32780 8100 33040
rect 7900 31740 8100 32780
rect 10060 33020 10260 33060
rect 10060 32760 10100 33020
rect 10220 32760 10260 33020
rect 10060 31980 10260 32760
rect 12320 33000 12500 33060
rect 12320 32780 12360 33000
rect 12480 32780 12500 33000
rect 12320 31960 12500 32780
rect 14520 32940 14720 33020
rect 14520 32740 14560 32940
rect 14700 32740 14720 32940
rect 14520 31980 14720 32740
rect -5700 14780 -2420 14880
rect -6060 14420 -2420 14780
rect -5700 14360 -2420 14420
rect -5700 12940 -3200 12980
rect -6080 12880 -3200 12940
rect -6080 12620 -3840 12880
rect -3300 12620 -3200 12880
rect -6080 12580 -3200 12620
rect -5700 12560 -3200 12580
rect -1040 11180 -500 13960
rect 5040 12920 5400 13360
rect 10360 13300 10620 13340
rect 8040 13280 10620 13300
rect 5040 12610 5090 12920
rect 5360 12610 5400 12920
rect 5040 12140 5400 12610
rect 6680 13120 10620 13280
rect 6680 12470 6940 13120
rect 8040 13100 10620 13120
rect 17010 12480 17390 12570
rect 6680 12250 7790 12470
rect 8050 12260 17390 12480
rect 6680 12180 6940 12250
rect 17010 12170 17390 12260
rect 16980 11460 17360 11520
rect 7560 11180 17360 11460
rect -6170 9840 -5730 9880
rect -1040 9840 -260 11180
rect 16980 11120 17360 11180
rect 17000 10200 17380 10260
rect 7760 9920 17380 10200
rect 17000 9860 17380 9920
rect -6170 9760 -260 9840
rect -6170 9660 -280 9760
rect -6170 9560 -500 9660
rect -6170 9520 -5730 9560
rect -6160 7620 -5700 7640
rect -6160 7300 -200 7620
rect -6160 7280 -5700 7300
<< via1 >>
rect 140 52480 300 52660
rect 4540 52480 4700 52660
rect 8980 52460 9140 52640
rect 13380 52500 13540 52680
rect -1270 37260 -1030 37520
rect -880 32800 -780 32960
rect 1320 32800 1460 33000
rect 3460 32720 3600 32920
rect 5700 32700 5860 32960
rect 7940 32780 8060 33040
rect 10100 32760 10220 33020
rect 12360 32780 12480 33000
rect 14560 32740 14700 32940
rect -3840 12620 -3300 12880
rect 5090 12610 5360 12920
<< metal2 >>
rect 80 52660 360 52740
rect 80 52480 140 52660
rect 300 52480 360 52660
rect 80 51820 360 52480
rect 4500 52660 4780 52720
rect 4500 52480 4540 52660
rect 4700 52480 4780 52660
rect 4500 51800 4780 52480
rect 8940 52640 9160 52700
rect 8940 52460 8980 52640
rect 9140 52460 9160 52640
rect 8940 51820 9160 52460
rect 13340 52680 13560 52700
rect 13340 52500 13380 52680
rect 13540 52500 13560 52680
rect 13340 51820 13560 52500
rect -1300 37520 -1020 37570
rect -1300 37260 -1270 37520
rect -1030 37260 -1020 37520
rect -1300 37230 -1020 37260
rect 7900 33040 8100 33100
rect 1280 33000 1500 33040
rect -920 32960 -740 33000
rect -920 32800 -880 32960
rect -780 32800 -740 32960
rect -920 32680 -740 32800
rect 1280 32800 1320 33000
rect 1460 32800 1500 33000
rect 5660 32960 5880 33020
rect 1280 32700 1500 32800
rect 3420 32920 3640 32960
rect 3420 32720 3460 32920
rect 3600 32720 3640 32920
rect 3420 32660 3640 32720
rect 5660 32700 5700 32960
rect 5860 32700 5880 32960
rect 7900 32780 7940 33040
rect 8060 32780 8100 33040
rect 7900 32720 8100 32780
rect 10060 33020 10260 33060
rect 10060 32760 10100 33020
rect 10220 32760 10260 33020
rect 10060 32720 10260 32760
rect 12320 33000 12500 33060
rect 12320 32780 12360 33000
rect 12480 32780 12500 33000
rect 12320 32720 12500 32780
rect 14520 32940 14720 33020
rect 14520 32740 14560 32940
rect 14700 32740 14720 32940
rect 5660 32640 5880 32700
rect 14520 32680 14720 32740
rect -3900 12920 5400 12970
rect -3900 12880 5090 12920
rect -3900 12620 -3840 12880
rect -3300 12620 5090 12880
rect -3900 12610 5090 12620
rect 5360 12610 5400 12920
rect -3900 12560 5400 12610
<< via2 >>
rect -1270 37260 -1030 37520
<< metal3 >>
rect -1300 37520 -1020 37570
rect -1300 37260 -1270 37520
rect -1030 37260 -1020 37520
rect -1300 37230 -1020 37260
<< via3 >>
rect -1270 37260 -1030 37520
<< metal4 >>
rect -1300 37520 -1020 37570
rect -1300 37260 -1270 37520
rect -1030 37260 -1020 37520
rect -1300 37230 -1020 37260
<< via4 >>
rect -1270 37260 -1030 37520
<< metal5 >>
rect -1300 37520 -930 37570
rect -1300 37260 -1270 37520
rect -1030 37260 -930 37520
rect -1300 37230 -930 37260
use sky130_fd_pr__res_high_po_0p35_LN2BL5  XRI
timestamp 1634754066
transform 0 -1 7926 1 0 12351
box -201 -696 201 696
use ota  ota_0 VGA/./ota/mag
timestamp 1635533344
transform -1 0 6440 0 1 2580
box -1540 -300 6960 9860
use digpot  digpot_0 VGA/./digpot/mag
timestamp 1635533344
transform 1 0 1172 0 1 -1182
box -4160 14300 15416 33360
use spi_slave  spi_slave_0 ./spi/magic
timestamp 1635533332
transform 1 0 -2046 0 1 32740
box 1066 0 16727 19884
<< labels >>
flabel metal1 -6170 9520 -5730 9880 5 FreeSans 12800 180 0 0 out
port 5 s
flabel metal1 -6140 7280 -5700 7640 5 FreeSans 12800 180 0 0 vs
port 7 s
flabel metal1 16980 11120 17360 11520 3 FreeSans 12800 0 0 0 in2
port 2 s
flabel metal1 17000 9860 17380 10260 5 FreeSans 12800 0 0 0 ib
port 3 s
flabel metal1 8840 53100 9220 53460 5 FreeSans 12800 180 0 0 sdi
port 10 s
flabel metal1 13260 53100 13640 53460 5 FreeSans 12800 180 0 0 reset
port 11 s
flabel metal1 4440 53100 4820 53460 5 FreeSans 12800 180 0 0 sclk
port 9 s
flabel metal1 40 53160 420 53520 5 FreeSans 12800 180 0 0 ss
port 8 s
flabel metal1 17010 12170 17390 12570 5 FreeSans 12800 180 0 0 in
port 1 s
flabel metal1 -6060 14420 -5680 14780 5 FreeSans 12800 180 0 0 gnd2
port 6 s
flabel metal1 -6080 12580 -5700 12940 5 FreeSans 12800 180 0 0 vd2
port 4 s
flabel metal1 -5720 37220 -5340 37580 5 FreeSans 12800 180 0 0 vd1
port 4 s
flabel metal1 -5720 39650 -5340 40010 5 FreeSans 12800 180 0 0 gnd1
port 9 s
<< end >>
