* OpAmp open-loop dc testbench

* Include SkyWater sky130 device models
.lib "/usr/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice" tt
.param mc_mm_switch=0
.include "../mag/opamp_core.spice"

* supply voltages
vdda  vdda 0 dc 1.0 pulse(1.0 1.8 10m 1u 1u 10 1)
vssa  vssa 0 0.0
egnda gnda vssa ib vssa 1

* input signals
vin in gnda dc 0 ac 1

* DUT
x0 out in out ib q vdda bp vddx gnda vssa xn xp x y z opamp_core
ib vdda ib 2n
cl out gnda 10p
il out gnda 0 

cmp out dp 10p
cmn out dn 10p

*.option METHOD="Gear"
.option gmin=1e-12
.control

	op
	print ib i(vdda)

	dc vin -0.5 0.5 1m
	plot in out xp xn z

	dc il -3u 3u 10n
	plot in out bp vddx
	
	tran 10u 20m
	plot in out vddx vdda

.endc

.end
