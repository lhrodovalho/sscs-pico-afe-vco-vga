magic
tech sky130A
magscale 1 2
timestamp 1634881297
<< nwell >>
rect -2366 7582 16048 8168
rect -2366 6926 16044 7582
rect -2366 3712 16042 6926
rect -2366 3680 4918 3712
rect 4928 3680 4990 3712
rect 5000 3680 16042 3712
rect -2366 3582 16042 3680
rect -2366 3580 -230 3582
<< pwell >>
rect -2426 -1250 16034 3502
<< psubdiff >>
rect -2308 833 -1944 884
rect -2308 255 -2279 833
rect -1973 255 -1944 833
rect -2308 204 -1944 255
<< nsubdiff >>
rect -2310 7123 -1942 7156
rect -2310 6477 -2279 7123
rect -1973 6477 -1942 7123
rect -2310 6444 -1942 6477
<< psubdiffcont >>
rect -2279 255 -1973 833
<< nsubdiffcont >>
rect -2279 6477 -1973 7123
<< locali >>
rect -2310 7123 -1942 7148
rect -2310 6477 -2279 7123
rect -1973 6700 -1942 7123
rect -1973 6666 -1902 6700
rect -1868 6666 294 6700
rect -1973 6477 -1942 6666
rect -2310 6452 -1942 6477
rect -1162 6006 -1128 6666
rect 15614 6032 15648 6148
rect 15518 5996 15744 6032
rect 15518 5926 15552 5996
rect 15710 5928 15744 5996
rect 15614 5926 15648 5928
rect -1158 4768 -1124 4860
rect -1158 4734 -1068 4768
rect 15614 3852 15648 3924
rect 2426 2316 2692 2350
rect 5426 2316 5692 2350
rect 8426 2316 8692 2350
rect 11426 2316 11692 2350
rect 14426 2316 14692 2350
rect 2658 2278 2692 2316
rect 5658 2278 5692 2316
rect 8658 2278 8692 2316
rect 11658 2280 11692 2316
rect 5500 2264 5534 2278
rect 8500 2264 8534 2278
rect 11500 2264 11534 2278
rect 14500 2264 14534 2278
rect 14658 2276 14692 2316
rect -1098 2138 -1097 2172
rect -1063 2138 -1062 2172
rect 2658 2074 2692 2076
rect 2500 1912 2534 2074
rect 2102 1878 2534 1912
rect 1664 1522 1698 1534
rect 2102 1522 2136 1878
rect 5500 1788 5534 2074
rect 5658 2070 5692 2076
rect 8500 1802 8534 2076
rect 8658 2070 8692 2074
rect 1664 1488 2136 1522
rect 4974 1754 5534 1788
rect 8002 1768 8534 1802
rect 4974 1490 5008 1754
rect 8002 1496 8036 1768
rect 11500 1690 11534 2074
rect 11658 2068 11692 2076
rect 10966 1656 11534 1690
rect 10966 1498 11000 1656
rect 14500 1638 14534 2076
rect 14658 2070 14692 2078
rect -2308 833 -1944 876
rect -2308 255 -2279 833
rect -1973 255 -1944 833
rect -2308 236 -1944 255
rect -2308 212 -1942 236
rect -1976 -18 -1942 212
rect -1686 -18 -1652 64
rect -1976 -52 -1564 -18
rect -1490 -40 -1456 64
rect -1294 -40 -1260 64
rect -1098 -40 -1064 64
rect -902 -18 -868 64
rect 626 -18 660 208
rect 1664 24 1698 1488
rect 4664 1456 5008 1490
rect 7664 1462 8036 1496
rect 10664 1464 11000 1498
rect 14152 1604 14534 1638
rect 4664 16 4698 1456
rect 7664 18 7698 1462
rect 4656 13 4708 16
rect -998 -52 660 -18
rect 4656 -21 4665 13
rect 4699 -21 4708 13
rect 4656 -24 4708 -21
rect 7656 15 7708 18
rect 7656 -19 7665 15
rect 7699 -19 7708 15
rect 10664 14 10698 1464
rect 14152 1448 14186 1604
rect 13964 1414 14186 1448
rect 7656 -22 7708 -19
rect 10654 11 10706 14
rect 10654 -23 10663 11
rect 10697 -23 10706 11
rect 13964 -12 13998 1414
rect 15510 52 15544 100
rect 15510 16 15544 18
rect 10654 -26 10706 -23
rect 13956 -15 14008 -12
rect 13956 -49 13965 -15
rect 13999 -49 14008 -15
rect 13956 -52 14008 -49
rect 13964 -56 13998 -52
<< viali >>
rect -1902 6666 -1868 6700
rect 15614 6148 15648 6182
rect 15710 3726 15744 3760
rect -1110 3290 -1076 3324
rect 2392 2316 2426 2350
rect 5392 2316 5426 2350
rect 8392 2316 8426 2350
rect 11392 2316 11426 2350
rect 14392 2316 14426 2350
rect -1097 2138 -1063 2172
rect 1664 -10 1698 24
rect 4665 -21 4699 13
rect 7665 -19 7699 15
rect 10663 -23 10697 11
rect 15510 18 15544 52
rect 13965 -49 13999 -15
<< metal1 >>
rect 4678 7064 4750 7122
rect -550 7002 12578 7064
rect -1916 6700 -1854 6722
rect -1916 6666 -1902 6700
rect -1868 6666 -1854 6700
rect -1916 3442 -1854 6666
rect -550 4780 -488 7002
rect 274 6762 336 7002
rect 1758 6947 1834 6950
rect 1758 6895 1770 6947
rect 1822 6895 1834 6947
rect 1758 6892 1834 6895
rect 2758 6809 2960 6814
rect 2758 6757 2893 6809
rect 2945 6757 2960 6809
rect 2758 6752 2960 6757
rect 3230 6742 3292 7002
rect 4668 6927 4760 6934
rect 4668 6875 4688 6927
rect 4740 6875 4760 6927
rect 4668 6868 4760 6875
rect 5908 6803 5990 6806
rect 5908 6800 5923 6803
rect 5706 6751 5923 6800
rect 5975 6751 5990 6803
rect 5706 6748 5990 6751
rect 5706 6742 5950 6748
rect 6260 6744 6322 7002
rect 7662 6934 7766 6952
rect 7662 6882 7688 6934
rect 7740 6882 7766 6934
rect 7662 6864 7766 6882
rect 8740 6799 8972 6804
rect 8740 6747 8905 6799
rect 8957 6747 8972 6799
rect 8740 6742 8972 6747
rect 9348 6742 9410 7002
rect 10730 6922 10838 6940
rect 10730 6870 10758 6922
rect 10810 6870 10838 6922
rect 10730 6852 10838 6870
rect 11814 6801 12122 6806
rect 11814 6749 12055 6801
rect 12107 6749 12122 6801
rect 11814 6744 12122 6749
rect 12504 6718 12566 7002
rect 13922 6899 14036 6920
rect 13922 6847 13953 6899
rect 14005 6847 14036 6899
rect 13922 6826 14036 6847
rect 14844 6769 14978 6774
rect 14844 6717 14855 6769
rect 14907 6717 14978 6769
rect 14844 6712 14978 6717
rect 15582 6345 15676 6356
rect 15582 6293 15603 6345
rect 15655 6293 15676 6345
rect 15582 6282 15676 6293
rect 15592 6182 15666 6282
rect 15592 6148 15614 6182
rect 15648 6148 15666 6182
rect 15592 6126 15666 6148
rect -1082 4718 -488 4780
rect -1082 3580 -1020 4718
rect 11160 3877 11724 3886
rect 11160 3825 11636 3877
rect 11688 3825 11724 3877
rect 11160 3816 11724 3825
rect 1842 3790 2168 3792
rect 1760 3787 2168 3790
rect 1760 3735 2101 3787
rect 2153 3735 2168 3787
rect 11160 3774 11230 3816
rect 15332 3794 15394 3798
rect 1760 3732 2168 3735
rect 1842 3730 2168 3732
rect 4714 3769 5000 3774
rect 4714 3717 4933 3769
rect 4985 3717 5000 3769
rect 4714 3712 5000 3717
rect 5598 3712 7614 3774
rect 7744 3712 8364 3774
rect 10008 3767 10698 3772
rect 10008 3715 10023 3767
rect 10075 3715 10698 3767
rect -1126 3518 -1020 3580
rect -1916 3380 -1546 3442
rect -1126 3324 -1064 3518
rect -1126 3290 -1110 3324
rect -1076 3290 -1064 3324
rect -1126 3276 -1064 3290
rect 3658 3305 3720 3320
rect 3658 3253 3663 3305
rect 3715 3253 3720 3305
rect 3658 3126 3720 3253
rect 5600 3215 5662 3712
rect 7122 3479 7656 3532
rect 7122 3427 7127 3479
rect 7179 3470 7656 3479
rect 7179 3427 7184 3470
rect 7122 3412 7184 3427
rect 7648 3378 7692 3430
rect 8298 3408 8360 3712
rect 10008 3710 10698 3715
rect 10830 3710 11230 3774
rect 13552 3684 13854 3748
rect 13988 3684 14642 3750
rect 15326 3732 15336 3794
rect 15398 3732 15560 3794
rect 15698 3760 15760 3772
rect 8672 3592 8682 3676
rect 8752 3652 8762 3676
rect 8752 3596 10798 3652
rect 8752 3592 8762 3596
rect 10404 3471 10466 3486
rect 10404 3419 10409 3471
rect 10461 3419 10466 3471
rect 10404 3408 10466 3419
rect 8298 3352 8746 3408
rect 8850 3352 10466 3408
rect 8298 3350 10466 3352
rect 13076 3471 13138 3486
rect 13076 3419 13081 3471
rect 13133 3419 13138 3471
rect 8298 3346 10464 3350
rect 5600 3163 5605 3215
rect 5657 3163 5662 3215
rect 13076 3260 13138 3419
rect 13552 3354 13614 3684
rect 13426 3349 13614 3354
rect 13426 3297 13441 3349
rect 13493 3297 13614 3349
rect 13426 3292 13614 3297
rect 13942 3272 14154 3330
rect 5600 3148 5662 3163
rect 7284 3191 7346 3206
rect 13076 3198 13934 3260
rect 7284 3139 7289 3191
rect 7341 3139 7346 3191
rect 1662 3064 4244 3126
rect 1394 3013 1626 3018
rect 1394 2961 1409 3013
rect 1461 2961 1626 3013
rect 1394 2956 1626 2961
rect 2232 2360 2294 3064
rect 4182 3000 4244 3064
rect 4618 3046 7200 3108
rect 4182 2938 4560 3000
rect 2550 2592 2642 2622
rect 2550 2540 2570 2592
rect 2622 2540 2642 2592
rect 2550 2388 2642 2540
rect 5132 2360 5194 3046
rect 7138 3000 7200 3046
rect 7284 3000 7346 3139
rect 7678 3066 10260 3128
rect 7138 2938 7608 3000
rect 5550 2592 5642 2622
rect 5550 2540 5570 2592
rect 5622 2540 5642 2592
rect 5550 2388 5642 2540
rect 8232 2360 8294 3066
rect 10198 2998 10260 3066
rect 10778 3064 13522 3126
rect 13892 3112 14296 3174
rect 10196 2936 10698 2998
rect 8550 2597 8644 2628
rect 8550 2545 8571 2597
rect 8623 2545 8644 2597
rect 8550 2514 8644 2545
rect 8550 2388 8642 2514
rect 11232 2360 11294 3064
rect 13460 2972 13522 3064
rect 13460 2910 13856 2972
rect 11550 2568 11642 2598
rect 11550 2516 11570 2568
rect 11622 2516 11642 2568
rect 11550 2388 11642 2516
rect 14232 2360 14294 3112
rect 14550 2388 14642 3684
rect 2232 2350 2438 2360
rect 2232 2316 2392 2350
rect 2426 2316 2438 2350
rect 2232 2298 2438 2316
rect 5132 2350 5438 2360
rect 5132 2316 5392 2350
rect 5426 2316 5438 2350
rect 5132 2298 5438 2316
rect 8232 2350 8440 2360
rect 8232 2316 8392 2350
rect 8426 2316 8440 2350
rect 8232 2298 8440 2316
rect 11232 2350 11440 2360
rect 11232 2316 11392 2350
rect 11426 2316 11440 2350
rect 11232 2298 11440 2316
rect 14232 2350 14442 2360
rect 14232 2316 14392 2350
rect 14426 2316 14442 2350
rect 14232 2298 14442 2316
rect -1110 2172 -1048 2190
rect -1110 2138 -1097 2172
rect -1063 2138 -1048 2172
rect -1110 1256 -1048 2138
rect 15332 1326 15394 3732
rect 15698 3726 15710 3760
rect 15744 3726 15760 3760
rect 15452 1671 15514 1686
rect 15452 1619 15457 1671
rect 15509 1619 15514 1671
rect 15452 1444 15514 1619
rect -914 1250 -458 1312
rect -522 -130 -458 1250
rect 142 -76 204 144
rect 1698 -10 1864 2
rect 1696 -20 1864 -10
rect 2774 -15 2836 144
rect 1700 -45 1774 -20
rect 142 -130 206 -76
rect 1700 -97 1711 -45
rect 1763 -97 1774 -45
rect 2774 -67 2779 -15
rect 2831 -67 2836 -15
rect 2774 -82 2836 -67
rect 3098 -76 3160 128
rect 4656 13 4708 16
rect 4656 -21 4665 13
rect 4699 -21 4708 13
rect 5730 -11 5792 122
rect 4656 -24 4708 -21
rect 4856 -23 4938 -18
rect 4856 -75 4871 -23
rect 4923 -75 4938 -23
rect 1700 -102 1774 -97
rect 3098 -130 3162 -76
rect 4856 -80 4938 -75
rect 5730 -63 5735 -11
rect 5787 -63 5792 -11
rect 5730 -78 5792 -63
rect 6128 -78 6190 126
rect 7656 15 7708 18
rect 7656 -19 7665 15
rect 7699 -19 7708 15
rect 7656 -22 7708 -19
rect 7822 -13 7904 -8
rect 7822 -65 7837 -13
rect 7889 -65 7904 -13
rect 7822 -70 7904 -65
rect 8760 -25 8822 122
rect 6126 -130 6190 -78
rect 8760 -77 8765 -25
rect 8817 -77 8822 -25
rect 8760 -92 8822 -77
rect 9214 -76 9276 128
rect 10654 11 10706 14
rect 10654 -23 10663 11
rect 10697 -23 10706 11
rect 10654 -26 10706 -23
rect 10930 -34 11012 -24
rect 9214 -130 9278 -76
rect 10930 -86 10945 -34
rect 10997 -86 11012 -34
rect 10930 -96 11012 -86
rect 11848 -25 11910 122
rect 11848 -77 11853 -25
rect 11905 -77 11910 -25
rect 11848 -92 11910 -77
rect 12372 -74 12434 96
rect 13956 -15 14008 -12
rect 13956 -49 13965 -15
rect 13999 -49 14008 -15
rect 13956 -52 14008 -49
rect 14106 -45 14188 -38
rect 12372 -130 12436 -74
rect 14106 -97 14121 -45
rect 14173 -97 14188 -45
rect 14106 -104 14188 -97
rect 15002 -66 15064 98
rect 15322 52 15554 64
rect 15322 18 15510 52
rect 15544 18 15554 52
rect 15322 2 15554 18
rect 15322 -66 15384 2
rect 15002 -128 15384 -66
rect -522 -190 12440 -130
rect 6126 -192 6190 -190
rect 2790 -249 2956 -244
rect 2790 -301 2889 -249
rect 2941 -301 2956 -249
rect 15320 -258 15384 -128
rect 15698 -258 15760 3726
rect 2790 -306 2956 -301
rect 8580 -265 8744 -260
rect 2790 -456 2852 -306
rect 5558 -307 5706 -302
rect 5558 -359 5639 -307
rect 5691 -359 5706 -307
rect 8580 -317 8677 -265
rect 8729 -317 8744 -265
rect 8580 -322 8744 -317
rect 11668 -283 11818 -278
rect 5558 -364 5706 -359
rect 5558 -456 5620 -364
rect 8582 -456 8644 -322
rect 11668 -335 11751 -283
rect 11803 -335 11818 -283
rect 11668 -340 11818 -335
rect 15320 -320 15760 -258
rect 11668 -456 11730 -340
rect 15320 -456 15384 -320
rect 2790 -518 15386 -456
<< via1 >>
rect 1770 6895 1822 6947
rect 2893 6757 2945 6809
rect 4688 6875 4740 6927
rect 5923 6751 5975 6803
rect 7688 6882 7740 6934
rect 8905 6747 8957 6799
rect 10758 6870 10810 6922
rect 12055 6749 12107 6801
rect 13953 6847 14005 6899
rect 14855 6717 14907 6769
rect 15603 6293 15655 6345
rect 11636 3825 11688 3877
rect 2101 3735 2153 3787
rect 4933 3717 4985 3769
rect 10023 3715 10075 3767
rect 3663 3253 3715 3305
rect 7127 3427 7179 3479
rect 15336 3732 15398 3794
rect 8682 3592 8752 3676
rect 10409 3419 10461 3471
rect 8746 3352 8850 3408
rect 13081 3419 13133 3471
rect 5605 3163 5657 3215
rect 13441 3297 13493 3349
rect 7289 3139 7341 3191
rect 1409 2961 1461 3013
rect 2570 2540 2622 2592
rect 5570 2540 5622 2592
rect 8571 2545 8623 2597
rect 11570 2516 11622 2568
rect 15457 1619 15509 1671
rect 1711 -97 1763 -45
rect 2779 -67 2831 -15
rect 4871 -75 4923 -23
rect 5735 -63 5787 -11
rect 7837 -65 7889 -13
rect 8765 -77 8817 -25
rect 10945 -86 10997 -34
rect 11853 -77 11905 -25
rect 14121 -97 14173 -45
rect 2889 -301 2941 -249
rect 5639 -359 5691 -307
rect 8677 -317 8729 -265
rect 11751 -335 11803 -283
<< metal2 >>
rect 15058 7404 15120 7434
rect 2888 7344 15130 7404
rect 1768 7163 1824 7174
rect 1768 6947 1824 7107
rect 1768 6895 1770 6947
rect 1822 6895 1824 6947
rect 1768 6882 1824 6895
rect 2888 6809 2950 7344
rect 4678 7173 4750 7190
rect 4678 7117 4686 7173
rect 4742 7117 4750 7173
rect 4678 6927 4750 7117
rect 4678 6875 4688 6927
rect 4740 6875 4750 6927
rect 4678 6858 4750 6875
rect 2888 6757 2893 6809
rect 2945 6757 2950 6809
rect 2888 6742 2950 6757
rect 5918 6803 5980 7344
rect 7672 7238 7756 7264
rect 7672 7182 7686 7238
rect 7742 7182 7756 7238
rect 7672 6934 7756 7182
rect 7672 6882 7688 6934
rect 7740 6882 7756 6934
rect 7672 6854 7756 6882
rect 5918 6751 5923 6803
rect 5975 6751 5980 6803
rect 5918 6738 5980 6751
rect 8900 6799 8962 7344
rect 10740 7202 10828 7228
rect 10740 7146 10756 7202
rect 10812 7146 10828 7202
rect 10740 6922 10828 7146
rect 10740 6870 10758 6922
rect 10810 6870 10828 6922
rect 10740 6842 10828 6870
rect 8900 6747 8905 6799
rect 8957 6747 8962 6799
rect 8900 6732 8962 6747
rect 12050 6801 12112 7344
rect 13932 7135 14026 7164
rect 13932 7079 13951 7135
rect 14007 7079 14026 7135
rect 13932 6899 14026 7079
rect 13932 6847 13953 6899
rect 14005 6847 14026 6899
rect 13932 6816 14026 6847
rect 12050 6749 12055 6801
rect 12107 6749 12112 6801
rect 12050 6734 12112 6749
rect 14850 6769 14912 7344
rect 14850 6717 14855 6769
rect 14907 6717 14912 6769
rect 14850 6702 14912 6717
rect 11610 3877 11714 3896
rect 11610 3825 11636 3877
rect 11688 3825 11714 3877
rect 2096 3787 2158 3802
rect 2096 3735 2101 3787
rect 2153 3735 2158 3787
rect 2096 3484 2158 3735
rect 4928 3769 4990 3784
rect 4928 3717 4933 3769
rect 4985 3717 4990 3769
rect 4928 3666 4990 3717
rect 10018 3767 10080 3782
rect 10018 3715 10023 3767
rect 10075 3715 10080 3767
rect 8682 3676 8752 3686
rect 4928 3664 5082 3666
rect 5484 3664 8682 3666
rect 4928 3646 8682 3664
rect 4928 3604 5364 3646
rect 5458 3604 8682 3646
rect 8682 3582 8752 3592
rect 5364 3556 5458 3566
rect 2096 3479 7194 3484
rect 2096 3427 7127 3479
rect 7179 3427 7194 3479
rect 2096 3422 7194 3427
rect 2886 3364 2950 3422
rect 2710 3360 2950 3364
rect 2710 3304 2744 3360
rect 2800 3304 2950 3360
rect 8746 3408 8850 3418
rect 8746 3342 8850 3352
rect 10018 3310 10080 3715
rect 11610 3776 11714 3825
rect 11610 3720 11634 3776
rect 11690 3720 11714 3776
rect 11610 3700 11714 3720
rect 10394 3471 13148 3476
rect 10394 3419 10409 3471
rect 10461 3419 13081 3471
rect 13133 3419 13148 3471
rect 10394 3414 13148 3419
rect 2710 3300 2950 3304
rect 3648 3305 10080 3310
rect 3648 3253 3663 3305
rect 3715 3253 10080 3305
rect 3648 3248 10080 3253
rect 13436 3349 13498 3364
rect 13436 3297 13441 3349
rect 13493 3297 13498 3349
rect 1404 3215 5680 3220
rect 1404 3163 5605 3215
rect 5657 3163 5680 3215
rect 13436 3196 13498 3297
rect 1404 3158 5680 3163
rect 7274 3191 13498 3196
rect 1404 3013 1466 3158
rect 7274 3139 7289 3191
rect 7341 3139 13498 3191
rect 7274 3134 13498 3139
rect 1404 2961 1409 3013
rect 1461 2961 1466 3013
rect 1404 2946 1466 2961
rect 2540 2594 2828 2612
rect 2540 2592 2744 2594
rect 2540 2540 2570 2592
rect 2622 2540 2744 2592
rect 2540 2538 2744 2540
rect 2800 2538 2828 2594
rect 2540 2520 2828 2538
rect 5356 2594 5652 2612
rect 5356 2538 5384 2594
rect 5440 2592 5652 2594
rect 5440 2540 5570 2592
rect 5622 2540 5652 2592
rect 5440 2538 5652 2540
rect 5356 2520 5652 2538
rect 8540 2599 8856 2618
rect 8540 2597 8771 2599
rect 8540 2545 8571 2597
rect 8623 2545 8771 2597
rect 8540 2543 8771 2545
rect 8827 2543 8856 2599
rect 8540 2524 8856 2543
rect 11540 2570 11836 2588
rect 11540 2568 11752 2570
rect 11540 2516 11570 2568
rect 11622 2516 11752 2568
rect 11540 2514 11752 2516
rect 11808 2514 11836 2570
rect 11540 2496 11836 2514
rect 15058 1676 15120 7344
rect 15592 6653 15666 6672
rect 15592 6597 15601 6653
rect 15657 6597 15666 6653
rect 15592 6345 15666 6597
rect 15592 6293 15603 6345
rect 15655 6293 15666 6345
rect 15592 6272 15666 6293
rect 15336 3794 15398 3804
rect 15336 3676 15398 3732
rect 15336 3614 15946 3676
rect 15548 1676 15610 1686
rect 15058 1673 15610 1676
rect 15058 1671 15551 1673
rect 15058 1619 15457 1671
rect 15509 1619 15551 1671
rect 15058 1617 15551 1619
rect 15607 1617 15610 1673
rect 15058 1614 15610 1617
rect 15548 1604 15610 1614
rect 2764 -15 2946 -10
rect 1706 -45 1768 -30
rect 1706 -97 1711 -45
rect 1763 -97 1768 -45
rect 2764 -67 2779 -15
rect 2831 -67 2946 -15
rect 2764 -72 2946 -67
rect 1706 -223 1768 -97
rect 1706 -279 1709 -223
rect 1765 -279 1768 -223
rect 1706 -292 1768 -279
rect 2884 -249 2946 -72
rect 2884 -301 2889 -249
rect 2941 -301 2946 -249
rect 2884 -316 2946 -301
rect 4866 -23 4928 -8
rect 4866 -75 4871 -23
rect 4923 -75 4928 -23
rect 4866 -237 4928 -75
rect 4866 -293 4869 -237
rect 4925 -293 4928 -237
rect 4866 -306 4928 -293
rect 5634 -11 5802 -6
rect 5634 -63 5735 -11
rect 5787 -63 5802 -11
rect 5634 -68 5802 -63
rect 7832 -13 7894 2
rect 7832 -65 7837 -13
rect 7889 -65 7894 -13
rect 5634 -307 5696 -68
rect 7832 -225 7894 -65
rect 7832 -281 7835 -225
rect 7891 -281 7894 -225
rect 7832 -294 7894 -281
rect 8672 -25 8832 -20
rect 8672 -77 8765 -25
rect 8817 -77 8832 -25
rect 8672 -82 8832 -77
rect 10940 -34 11002 -14
rect 8672 -265 8734 -82
rect 5634 -359 5639 -307
rect 5691 -359 5696 -307
rect 8672 -317 8677 -265
rect 8729 -317 8734 -265
rect 10940 -86 10945 -34
rect 10997 -86 11002 -34
rect 10940 -238 11002 -86
rect 10940 -294 10943 -238
rect 10999 -294 11002 -238
rect 10940 -312 11002 -294
rect 11746 -25 11920 -20
rect 11746 -77 11853 -25
rect 11905 -77 11920 -25
rect 11746 -82 11920 -77
rect 14116 -45 14178 -28
rect 11746 -283 11808 -82
rect 14116 -97 14121 -45
rect 14173 -97 14178 -45
rect 15882 -60 15946 3614
rect 14116 -177 14178 -97
rect 14116 -233 14119 -177
rect 14175 -233 14178 -177
rect 15576 -116 15946 -60
rect 15576 -184 15626 -116
rect 14116 -248 14178 -233
rect 15572 -194 15630 -184
rect 15572 -250 15573 -194
rect 15629 -250 15630 -194
rect 15572 -260 15630 -250
rect 8672 -332 8734 -317
rect 11746 -335 11751 -283
rect 11803 -335 11808 -283
rect 11746 -350 11808 -335
rect 5634 -374 5696 -359
<< via2 >>
rect 1768 7107 1824 7163
rect 4686 7117 4742 7173
rect 7686 7182 7742 7238
rect 10756 7146 10812 7202
rect 13951 7079 14007 7135
rect 5364 3566 5458 3646
rect 2744 3304 2800 3360
rect 8746 3352 8850 3408
rect 11634 3720 11690 3776
rect 2744 2538 2800 2594
rect 5384 2538 5440 2594
rect 8771 2543 8827 2599
rect 11752 2514 11808 2570
rect 15601 6597 15657 6653
rect 15551 1617 15607 1673
rect 1709 -279 1765 -223
rect 4869 -293 4925 -237
rect 7835 -281 7891 -225
rect 10943 -294 10999 -238
rect 14119 -233 14175 -177
rect 15573 -250 15629 -194
<< metal3 >>
rect 4862 7632 4968 7642
rect 4862 7568 4883 7632
rect 4947 7568 4968 7632
rect 4862 7558 4968 7568
rect 7910 7601 8028 7618
rect 1880 7331 1990 7344
rect 1880 7267 1903 7331
rect 1967 7267 1990 7331
rect 1880 7254 1990 7267
rect 1890 7182 1980 7254
rect 4872 7188 4958 7558
rect 7910 7537 7937 7601
rect 8001 7537 8028 7601
rect 14298 7604 14422 7624
rect 7910 7520 8028 7537
rect 11076 7580 11196 7598
rect 7920 7260 8018 7520
rect 11076 7516 11104 7580
rect 11168 7516 11196 7580
rect 14298 7540 14328 7604
rect 14392 7540 14422 7604
rect 14298 7520 14422 7540
rect 11076 7498 11196 7516
rect 7746 7259 8018 7260
rect 1752 7163 1980 7182
rect 1752 7107 1768 7163
rect 1824 7107 1980 7163
rect 1752 7092 1980 7107
rect 4660 7173 4958 7188
rect 4660 7117 4686 7173
rect 4742 7117 4958 7173
rect 7662 7238 8018 7259
rect 7662 7182 7686 7238
rect 7742 7182 8018 7238
rect 11086 7224 11186 7498
rect 10830 7223 11186 7224
rect 7662 7162 8018 7182
rect 10730 7202 11186 7223
rect 7662 7161 7766 7162
rect 10730 7146 10756 7202
rect 10812 7146 11186 7202
rect 14308 7160 14412 7520
rect 13932 7159 14412 7160
rect 10730 7125 11186 7146
rect 10830 7124 11186 7125
rect 13922 7135 14412 7159
rect 4660 7102 4958 7117
rect 13922 7079 13951 7135
rect 14007 7079 14412 7135
rect 13922 7056 14412 7079
rect 13922 7055 14036 7056
rect 14308 7054 14412 7056
rect 15570 7063 15688 7080
rect 15570 6999 15597 7063
rect 15661 6999 15688 7063
rect 15570 6982 15688 6999
rect 15580 6653 15678 6982
rect 15580 6597 15601 6653
rect 15657 6597 15678 6653
rect 15580 6576 15678 6597
rect 11722 3791 11832 3792
rect 11600 3776 11832 3791
rect 11600 3720 11634 3776
rect 11690 3720 11832 3776
rect 11600 3705 11832 3720
rect 11722 3704 11832 3705
rect 5360 3651 5464 3672
rect 5354 3646 5468 3651
rect 5354 3566 5364 3646
rect 5458 3566 5468 3646
rect 5354 3561 5468 3566
rect 2715 3360 2829 3374
rect 2715 3304 2744 3360
rect 2800 3304 2829 3360
rect 2715 3290 2829 3304
rect 2720 2616 2824 3290
rect 2721 2594 2823 2616
rect 2721 2538 2744 2594
rect 2800 2538 2823 2594
rect 5360 2594 5464 3561
rect 8746 3413 8852 3414
rect 8736 3408 8860 3413
rect 8736 3352 8746 3408
rect 8850 3352 8860 3408
rect 8736 3347 8860 3352
rect 8746 2624 8852 3347
rect 5360 2582 5384 2594
rect 2721 2510 2823 2538
rect 5361 2538 5384 2582
rect 5440 2582 5464 2594
rect 8747 2599 8851 2624
rect 5440 2538 5463 2582
rect 5361 2510 5463 2538
rect 8747 2543 8771 2599
rect 8827 2543 8851 2599
rect 11728 2590 11832 3704
rect 8747 2514 8851 2543
rect 11729 2570 11831 2590
rect 11729 2514 11752 2570
rect 11808 2514 11831 2570
rect 11729 2486 11831 2514
rect 15536 1677 15884 1694
rect 15536 1673 15793 1677
rect 15536 1617 15551 1673
rect 15607 1617 15793 1673
rect 15536 1613 15793 1617
rect 15857 1613 15884 1677
rect 15536 1596 15884 1613
rect 14102 -177 14366 -162
rect 1688 -223 1916 -202
rect 1688 -279 1709 -223
rect 1765 -279 1916 -223
rect 1688 -296 1916 -279
rect 1822 -361 1916 -296
rect 4852 -237 5070 -224
rect 4852 -293 4869 -237
rect 4925 -293 5070 -237
rect 4852 -312 5070 -293
rect 7806 -225 8070 -210
rect 7806 -281 7835 -225
rect 7891 -281 8070 -225
rect 7806 -302 8070 -281
rect 1821 -368 1916 -361
rect 1821 -386 1915 -368
rect 1821 -450 1836 -386
rect 1900 -450 1915 -386
rect 1821 -475 1915 -450
rect 4982 -643 5070 -312
rect 7978 -583 8070 -302
rect 10924 -238 11126 -222
rect 10924 -294 10943 -238
rect 10999 -294 11126 -238
rect 14102 -233 14119 -177
rect 14175 -233 14366 -177
rect 14102 -248 14366 -233
rect 10924 -318 11126 -294
rect 4981 -644 5070 -643
rect 7969 -607 8073 -583
rect 4981 -665 5069 -644
rect 4981 -729 4993 -665
rect 5057 -729 5069 -665
rect 7969 -671 7989 -607
rect 8053 -671 8073 -607
rect 11032 -607 11126 -318
rect 14282 -598 14366 -248
rect 15542 -194 15654 -178
rect 15542 -250 15573 -194
rect 15629 -250 15654 -194
rect 15542 -330 15654 -250
rect 15532 -345 15664 -330
rect 15532 -409 15566 -345
rect 15630 -409 15664 -345
rect 15532 -424 15664 -409
rect 11032 -608 11127 -607
rect 7969 -695 8073 -671
rect 11033 -632 11127 -608
rect 11033 -696 11048 -632
rect 11112 -696 11127 -632
rect 14283 -613 14363 -598
rect 14283 -677 14291 -613
rect 14355 -677 14363 -613
rect 14283 -695 14363 -677
rect 11033 -721 11127 -696
rect 4981 -751 5069 -729
<< via3 >>
rect 4883 7568 4947 7632
rect 1903 7267 1967 7331
rect 7937 7537 8001 7601
rect 11104 7516 11168 7580
rect 14328 7540 14392 7604
rect 15597 6999 15661 7063
rect 15793 1613 15857 1677
rect 1836 -450 1900 -386
rect 4993 -729 5057 -665
rect 7989 -671 8053 -607
rect 15566 -409 15630 -345
rect 11048 -696 11112 -632
rect 14291 -677 14355 -613
<< metal4 >>
rect 908 7790 15998 8014
rect 1884 7331 1984 7790
rect 4864 7632 4964 7790
rect 7916 7706 8020 7790
rect 4864 7568 4883 7632
rect 4947 7568 4964 7632
rect 4864 7552 4964 7568
rect 7918 7601 8020 7706
rect 7918 7537 7937 7601
rect 8001 7537 8020 7601
rect 7918 7518 8020 7537
rect 11084 7580 11188 7790
rect 11084 7516 11104 7580
rect 11168 7516 11188 7580
rect 14306 7604 14414 7790
rect 14306 7540 14328 7604
rect 14392 7540 14414 7604
rect 14306 7518 14414 7540
rect 11084 7496 11188 7516
rect 1884 7267 1903 7331
rect 1967 7267 1984 7331
rect 1884 7252 1984 7267
rect 1884 7250 1982 7252
rect 15578 7063 15680 7790
rect 15578 6999 15597 7063
rect 15661 6999 15680 7063
rect 15578 6980 15680 6999
rect 16036 1764 16284 1770
rect 16036 1696 16042 1764
rect 15774 1677 16042 1696
rect 15774 1613 15793 1677
rect 15857 1613 16042 1677
rect 15774 1596 16042 1613
rect 15775 1595 15875 1596
rect 16036 1528 16042 1596
rect 16278 1528 16284 1764
rect 16036 1522 16284 1528
rect 15541 -345 15655 -329
rect 1812 -386 2086 -366
rect 1812 -450 1836 -386
rect 1900 -450 2086 -386
rect 15541 -409 15566 -345
rect 15630 -409 15655 -345
rect 15541 -425 15655 -409
rect 1812 -470 2086 -450
rect 1982 -826 2086 -470
rect 7968 -607 8232 -592
rect 4976 -665 5228 -648
rect 4976 -729 4993 -665
rect 5057 -729 5228 -665
rect 7968 -671 7989 -607
rect 8053 -671 8232 -607
rect 7968 -686 8232 -671
rect 4976 -748 5228 -729
rect 5128 -826 5228 -748
rect 8126 -826 8232 -686
rect 11028 -632 11290 -612
rect 11028 -696 11048 -632
rect 11112 -696 11290 -632
rect 14280 -613 14520 -602
rect 14280 -677 14291 -613
rect 14355 -677 14520 -613
rect 14280 -688 14520 -677
rect 11028 -714 11290 -696
rect 11196 -826 11290 -714
rect 14436 -826 14520 -688
rect 15542 -826 15654 -425
rect -592 -1040 15686 -826
<< via4 >>
rect 16042 1528 16278 1764
<< metal5 >>
rect 15972 1764 16698 1860
rect 15972 1528 16042 1764
rect 16278 1528 16698 1764
rect 15972 1432 16698 1528
use 5_Stage_MSSRO_PD  5_Stage_MSSRO_PD_0
timestamp 1634821592
transform 1 0 1452 0 1 1758
box -1468 -1778 1646 5200
use sky130_fd_pr__pfet_01v8_DWWSZ5  sky130_fd_pr__pfet_01v8_DWWSZ5_0
timestamp 1634821592
transform 1 0 -1243 0 1 5436
box -511 -720 457 636
use sky130_fd_pr__nfet_01v8_S65HPN  sky130_fd_pr__nfet_01v8_S65HPN_0
timestamp 1634821592
transform 1 0 -1285 0 1 2736
box -439 -598 439 708
use sky130_fd_pr__nfet_01v8_T4KHC3  sky130_fd_pr__nfet_01v8_T4KHC3_0
timestamp 1634821592
transform 1 0 -1277 0 1 566
box -447 -618 447 748
use 5_Stage_MSSRO_PD  5_Stage_MSSRO_PD_1
timestamp 1634821592
transform 1 0 4408 0 1 1742
box -1468 -1778 1646 5200
use sky130_fd_pr__nfet_01v8_U9YZD6  sky130_fd_pr__nfet_01v8_U9YZD6_0
timestamp 1634712416
transform 1 0 2596 0 1 2207
box -134 -157 134 237
use 5_Stage_MSSRO_PD  5_Stage_MSSRO_PD_2
timestamp 1634821592
transform 1 0 7438 0 1 1742
box -1468 -1778 1646 5200
use sky130_fd_pr__nfet_01v8_U9YZD6  sky130_fd_pr__nfet_01v8_U9YZD6_1
timestamp 1634712416
transform 1 0 5596 0 1 2207
box -134 -157 134 237
use 5_Stage_MSSRO_PD  5_Stage_MSSRO_PD_3
timestamp 1634821592
transform 1 0 10526 0 1 1740
box -1468 -1778 1646 5200
use sky130_fd_pr__nfet_01v8_U9YZD6  sky130_fd_pr__nfet_01v8_U9YZD6_2
timestamp 1634712416
transform 1 0 8596 0 1 2207
box -134 -157 134 237
use 5_Stage_MSSRO_PD  5_Stage_MSSRO_PD_4
timestamp 1634821592
transform 1 0 13682 0 1 1714
box -1468 -1778 1646 5200
use sky130_fd_pr__nfet_01v8_U9YZD6  sky130_fd_pr__nfet_01v8_U9YZD6_3
timestamp 1634712416
transform 1 0 11596 0 1 2207
box -134 -157 134 237
use sky130_fd_pr__pfet_01v8_AQ8SEE  sky130_fd_pr__pfet_01v8_AQ8SEE_0
timestamp 1634728397
transform 1 0 15631 0 1 4926
box -259 -1200 263 1100
use sky130_fd_pr__nfet_01v8_NC5H7G  sky130_fd_pr__nfet_01v8_NC5H7G_0
timestamp 1634712416
transform 1 0 15483 0 1 731
box -141 -657 99 777
use sky130_fd_pr__nfet_01v8_U9YZD6  sky130_fd_pr__nfet_01v8_U9YZD6_4
timestamp 1634712416
transform 1 0 14596 0 1 2207
box -134 -157 134 237
<< labels >>
rlabel metal4 7152 7932 7152 7932 1 VP
port 2 n
rlabel metal4 11374 -976 11374 -976 1 VN
port 4 n
rlabel metal5 16574 1566 16574 1566 1 VCT
port 3 n
rlabel metal1 14146 3302 14146 3302 1 OUT
port 1 n
<< end >>
