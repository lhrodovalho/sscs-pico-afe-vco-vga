magic
tech sky130A
timestamp 1638390070
<< psubdiff >>
rect -6440 3880 -6360 3920
rect 7360 3880 7440 3920
rect -6440 3840 -6400 3880
rect -6440 720 -6400 760
rect 7400 3840 7440 3880
rect 7400 720 7440 760
rect -6440 680 -6360 720
rect 7360 680 7440 720
<< psubdiffcont >>
rect -6360 3880 7360 3920
rect -6440 760 -6400 3840
rect 7400 760 7440 3840
rect -6360 680 7360 720
<< locali >>
rect -6440 3880 -6360 3920
rect 7360 3880 7440 3920
rect -6440 3840 -6400 3880
rect -6440 720 -6400 760
rect 7400 3840 7440 3880
rect 7400 720 7440 760
rect -6440 680 -6360 720
rect 7360 680 7440 720
<< metal3 >>
rect -6360 3836 -6160 3840
rect -6360 3804 -6356 3836
rect -6324 3804 -6276 3836
rect -6244 3804 -6196 3836
rect -6164 3804 -6160 3836
rect -6360 3676 -6160 3804
rect 7160 3836 7360 3840
rect 7160 3804 7164 3836
rect 7196 3804 7244 3836
rect 7276 3804 7324 3836
rect 7356 3804 7360 3836
rect -6360 3644 -6356 3676
rect -6324 3644 -6276 3676
rect -6244 3644 -6196 3676
rect -6164 3644 -6160 3676
rect -6360 3516 -6160 3644
rect -5520 3756 -5480 3760
rect -5520 3724 -5516 3756
rect -5484 3724 -5480 3756
rect -6360 3484 -6356 3516
rect -6324 3484 -6276 3516
rect -6244 3484 -6196 3516
rect -6164 3484 -6160 3516
rect -6360 1116 -6160 3484
rect -6120 3516 -6080 3520
rect -6120 3484 -6116 3516
rect -6084 3484 -6080 3516
rect -6120 2360 -6080 3484
rect -5520 3440 -5480 3724
rect -4320 3756 -4280 3760
rect -4320 3724 -4316 3756
rect -4284 3724 -4280 3756
rect -4920 3516 -4880 3520
rect -4920 3484 -4916 3516
rect -4884 3484 -4880 3516
rect -6000 2360 -5000 3440
rect -4920 2360 -4880 3484
rect -4320 3440 -4280 3724
rect -3120 3756 -3080 3760
rect -3120 3724 -3116 3756
rect -3084 3724 -3080 3756
rect -3720 3516 -3680 3520
rect -3720 3484 -3716 3516
rect -3684 3484 -3680 3516
rect -4800 2360 -3800 3440
rect -3720 2360 -3680 3484
rect -3120 3440 -3080 3724
rect -1920 3756 -1880 3760
rect -1920 3724 -1916 3756
rect -1884 3724 -1880 3756
rect -2520 3516 -2480 3520
rect -2520 3484 -2516 3516
rect -2484 3484 -2480 3516
rect -3600 2360 -2600 3440
rect -2520 2360 -2480 3484
rect -1920 3440 -1880 3724
rect -720 3756 -680 3760
rect -720 3724 -716 3756
rect -684 3724 -680 3756
rect -1320 3516 -1280 3520
rect -1320 3484 -1316 3516
rect -1284 3484 -1280 3516
rect -2400 2360 -1400 3440
rect -1320 2360 -1280 3484
rect -720 3440 -680 3724
rect 1680 3756 1720 3760
rect 1680 3724 1684 3756
rect 1716 3724 1720 3756
rect 480 3596 520 3600
rect 480 3564 484 3596
rect 516 3564 520 3596
rect -120 3516 -80 3520
rect -120 3484 -116 3516
rect -84 3484 -80 3516
rect -1200 2360 -200 3440
rect -120 2360 -80 3484
rect 480 3440 520 3564
rect 1080 3516 1120 3520
rect 1080 3484 1084 3516
rect 1116 3484 1120 3516
rect 0 2360 1000 3440
rect 1080 2360 1120 3484
rect 1680 3440 1720 3724
rect 2880 3756 2920 3760
rect 2880 3724 2884 3756
rect 2916 3724 2920 3756
rect 2280 3516 2320 3520
rect 2280 3484 2284 3516
rect 2316 3484 2320 3516
rect 1200 2360 2200 3440
rect 2280 2360 2320 3484
rect 2880 3440 2920 3724
rect 4080 3756 4120 3760
rect 4080 3724 4084 3756
rect 4116 3724 4120 3756
rect 3480 3516 3520 3520
rect 3480 3484 3484 3516
rect 3516 3484 3520 3516
rect 2400 2360 3400 3440
rect 3480 2360 3520 3484
rect 4080 3440 4120 3724
rect 5280 3756 5320 3760
rect 5280 3724 5284 3756
rect 5316 3724 5320 3756
rect 4680 3516 4720 3520
rect 4680 3484 4684 3516
rect 4716 3484 4720 3516
rect 3600 2360 4600 3440
rect 4680 2360 4720 3484
rect 5280 3440 5320 3724
rect 6480 3756 6520 3760
rect 6480 3724 6484 3756
rect 6516 3724 6520 3756
rect 5880 3516 5920 3520
rect 5880 3484 5884 3516
rect 5916 3484 5920 3516
rect 4800 2360 5800 3440
rect 5880 2360 5920 3484
rect 6480 3440 6520 3724
rect 7160 3676 7360 3804
rect 7160 3644 7164 3676
rect 7196 3644 7244 3676
rect 7276 3644 7324 3676
rect 7356 3644 7360 3676
rect 7080 3516 7120 3520
rect 7080 3484 7084 3516
rect 7116 3484 7120 3516
rect 6000 2360 7000 3440
rect 7080 2360 7120 3484
rect 7160 3516 7360 3644
rect 7160 3484 7164 3516
rect 7196 3484 7244 3516
rect 7276 3484 7324 3516
rect 7356 3484 7360 3516
rect -6360 1084 -6356 1116
rect -6324 1084 -6276 1116
rect -6244 1084 -6196 1116
rect -6164 1084 -6160 1116
rect -6360 956 -6160 1084
rect -6120 1116 -6080 2240
rect -6000 1160 -5000 2240
rect -6120 1084 -6116 1116
rect -6084 1084 -6080 1116
rect -6120 1080 -6080 1084
rect -6360 924 -6356 956
rect -6324 924 -6276 956
rect -6244 924 -6196 956
rect -6164 924 -6160 956
rect -6360 796 -6160 924
rect -5520 876 -5480 1160
rect -4920 1116 -4880 2240
rect -4800 1160 -3800 2240
rect -4920 1084 -4916 1116
rect -4884 1084 -4880 1116
rect -4920 1080 -4880 1084
rect -5520 844 -5516 876
rect -5484 844 -5480 876
rect -5520 840 -5480 844
rect -4320 876 -4280 1160
rect -3720 1116 -3680 2240
rect -3600 1160 -2600 2240
rect -3720 1084 -3716 1116
rect -3684 1084 -3680 1116
rect -3720 1080 -3680 1084
rect -4320 844 -4316 876
rect -4284 844 -4280 876
rect -4320 840 -4280 844
rect -3120 876 -3080 1160
rect -2520 1116 -2480 2240
rect -2400 1160 -1400 2240
rect -2520 1084 -2516 1116
rect -2484 1084 -2480 1116
rect -2520 1080 -2480 1084
rect -3120 844 -3116 876
rect -3084 844 -3080 876
rect -3120 840 -3080 844
rect -1920 876 -1880 1160
rect -1320 1116 -1280 2240
rect -1200 1160 -200 2240
rect -1320 1084 -1316 1116
rect -1284 1084 -1280 1116
rect -1320 1080 -1280 1084
rect -1920 844 -1916 876
rect -1884 844 -1880 876
rect -1920 840 -1880 844
rect -720 876 -680 1160
rect -120 1116 -80 2240
rect 0 1160 1000 2240
rect -120 1084 -116 1116
rect -84 1084 -80 1116
rect -120 1080 -80 1084
rect 480 1036 520 1160
rect 1080 1116 1120 2240
rect 1200 1160 2200 2240
rect 1080 1084 1084 1116
rect 1116 1084 1120 1116
rect 1080 1080 1120 1084
rect 480 1004 484 1036
rect 516 1004 520 1036
rect 480 1000 520 1004
rect -720 844 -716 876
rect -684 844 -680 876
rect -720 840 -680 844
rect 1680 876 1720 1160
rect 2280 1116 2320 2240
rect 2400 1160 3400 2240
rect 2280 1084 2284 1116
rect 2316 1084 2320 1116
rect 2280 1080 2320 1084
rect 1680 844 1684 876
rect 1716 844 1720 876
rect 1680 840 1720 844
rect 2880 876 2920 1160
rect 3480 1116 3520 2240
rect 3600 1160 4600 2240
rect 3480 1084 3484 1116
rect 3516 1084 3520 1116
rect 3480 1080 3520 1084
rect 2880 844 2884 876
rect 2916 844 2920 876
rect 2880 840 2920 844
rect 4080 876 4120 1160
rect 4680 1116 4720 2240
rect 4800 1160 5800 2240
rect 4680 1084 4684 1116
rect 4716 1084 4720 1116
rect 4680 1080 4720 1084
rect 4080 844 4084 876
rect 4116 844 4120 876
rect 4080 840 4120 844
rect 5280 876 5320 1160
rect 5880 1116 5920 2240
rect 6000 1160 7000 2240
rect 5880 1084 5884 1116
rect 5916 1084 5920 1116
rect 5880 1080 5920 1084
rect 5280 844 5284 876
rect 5316 844 5320 876
rect 5280 840 5320 844
rect 6480 876 6520 1160
rect 7080 1116 7120 2240
rect 7080 1084 7084 1116
rect 7116 1084 7120 1116
rect 7080 1080 7120 1084
rect 7160 1116 7360 3484
rect 7160 1084 7164 1116
rect 7196 1084 7244 1116
rect 7276 1084 7324 1116
rect 7356 1084 7360 1116
rect 6480 844 6484 876
rect 6516 844 6520 876
rect 6480 840 6520 844
rect 7160 956 7360 1084
rect 7160 924 7164 956
rect 7196 924 7244 956
rect 7276 924 7324 956
rect 7356 924 7360 956
rect -6360 764 -6356 796
rect -6324 764 -6276 796
rect -6244 764 -6196 796
rect -6164 764 -6160 796
rect -6360 760 -6160 764
rect 7160 796 7360 924
rect 7160 764 7164 796
rect 7196 764 7244 796
rect 7276 764 7324 796
rect 7356 764 7360 796
rect 7160 760 7360 764
<< via3 >>
rect -6356 3804 -6324 3836
rect -6276 3804 -6244 3836
rect -6196 3804 -6164 3836
rect 7164 3804 7196 3836
rect 7244 3804 7276 3836
rect 7324 3804 7356 3836
rect -6356 3644 -6324 3676
rect -6276 3644 -6244 3676
rect -6196 3644 -6164 3676
rect -5516 3724 -5484 3756
rect -6356 3484 -6324 3516
rect -6276 3484 -6244 3516
rect -6196 3484 -6164 3516
rect -6116 3484 -6084 3516
rect -4316 3724 -4284 3756
rect -4916 3484 -4884 3516
rect -3116 3724 -3084 3756
rect -3716 3484 -3684 3516
rect -1916 3724 -1884 3756
rect -2516 3484 -2484 3516
rect -716 3724 -684 3756
rect -1316 3484 -1284 3516
rect 1684 3724 1716 3756
rect 484 3564 516 3596
rect -116 3484 -84 3516
rect 1084 3484 1116 3516
rect 2884 3724 2916 3756
rect 2284 3484 2316 3516
rect 4084 3724 4116 3756
rect 3484 3484 3516 3516
rect 5284 3724 5316 3756
rect 4684 3484 4716 3516
rect 6484 3724 6516 3756
rect 5884 3484 5916 3516
rect 7164 3644 7196 3676
rect 7244 3644 7276 3676
rect 7324 3644 7356 3676
rect 7084 3484 7116 3516
rect 7164 3484 7196 3516
rect 7244 3484 7276 3516
rect 7324 3484 7356 3516
rect -6356 1084 -6324 1116
rect -6276 1084 -6244 1116
rect -6196 1084 -6164 1116
rect -6116 1084 -6084 1116
rect -6356 924 -6324 956
rect -6276 924 -6244 956
rect -6196 924 -6164 956
rect -4916 1084 -4884 1116
rect -5516 844 -5484 876
rect -3716 1084 -3684 1116
rect -4316 844 -4284 876
rect -2516 1084 -2484 1116
rect -3116 844 -3084 876
rect -1316 1084 -1284 1116
rect -1916 844 -1884 876
rect -116 1084 -84 1116
rect 1084 1084 1116 1116
rect 484 1004 516 1036
rect -716 844 -684 876
rect 2284 1084 2316 1116
rect 1684 844 1716 876
rect 3484 1084 3516 1116
rect 2884 844 2916 876
rect 4684 1084 4716 1116
rect 4084 844 4116 876
rect 5884 1084 5916 1116
rect 5284 844 5316 876
rect 7084 1084 7116 1116
rect 7164 1084 7196 1116
rect 7244 1084 7276 1116
rect 7324 1084 7356 1116
rect 6484 844 6516 876
rect 7164 924 7196 956
rect 7244 924 7276 956
rect 7324 924 7356 956
rect -6356 764 -6324 796
rect -6276 764 -6244 796
rect -6196 764 -6164 796
rect 7164 764 7196 796
rect 7244 764 7276 796
rect 7324 764 7356 796
<< mimcap >>
rect -6320 3360 -6200 3400
rect -6320 2440 -6280 3360
rect -6240 2440 -6200 3360
rect -6320 2400 -6200 2440
rect -5960 3360 -5040 3400
rect -5960 2440 -5920 3360
rect -5080 2440 -5040 3360
rect -5960 2400 -5040 2440
rect -4760 3360 -3840 3400
rect -4760 2440 -4720 3360
rect -3880 2440 -3840 3360
rect -4760 2400 -3840 2440
rect -3560 3360 -2640 3400
rect -3560 2440 -3520 3360
rect -2680 2440 -2640 3360
rect -3560 2400 -2640 2440
rect -2360 3360 -1440 3400
rect -2360 2440 -2320 3360
rect -1480 2440 -1440 3360
rect -2360 2400 -1440 2440
rect -1160 3360 -240 3400
rect -1160 2440 -1120 3360
rect -280 2440 -240 3360
rect -1160 2400 -240 2440
rect 40 3360 960 3400
rect 40 2440 80 3360
rect 920 2440 960 3360
rect 40 2400 960 2440
rect 1240 3360 2160 3400
rect 1240 2440 1280 3360
rect 2120 2440 2160 3360
rect 1240 2400 2160 2440
rect 2440 3360 3360 3400
rect 2440 2440 2480 3360
rect 3320 2440 3360 3360
rect 2440 2400 3360 2440
rect 3640 3360 4560 3400
rect 3640 2440 3680 3360
rect 4520 2440 4560 3360
rect 3640 2400 4560 2440
rect 4840 3360 5760 3400
rect 4840 2440 4880 3360
rect 5720 2440 5760 3360
rect 4840 2400 5760 2440
rect 6040 3360 6960 3400
rect 6040 2440 6080 3360
rect 6920 2440 6960 3360
rect 6040 2400 6960 2440
rect 7200 3360 7320 3400
rect 7200 2440 7240 3360
rect 7280 2440 7320 3360
rect 7200 2400 7320 2440
rect -6320 2160 -6200 2200
rect -6320 1240 -6280 2160
rect -6240 1240 -6200 2160
rect -6320 1200 -6200 1240
rect -5960 2160 -5040 2200
rect -5960 1240 -5920 2160
rect -5080 1240 -5040 2160
rect -5960 1200 -5040 1240
rect -4760 2160 -3840 2200
rect -4760 1240 -4720 2160
rect -3880 1240 -3840 2160
rect -4760 1200 -3840 1240
rect -3560 2160 -2640 2200
rect -3560 1240 -3520 2160
rect -2680 1240 -2640 2160
rect -3560 1200 -2640 1240
rect -2360 2160 -1440 2200
rect -2360 1240 -2320 2160
rect -1480 1240 -1440 2160
rect -2360 1200 -1440 1240
rect -1160 2160 -240 2200
rect -1160 1240 -1120 2160
rect -280 1240 -240 2160
rect -1160 1200 -240 1240
rect 40 2160 960 2200
rect 40 1240 80 2160
rect 920 1240 960 2160
rect 40 1200 960 1240
rect 1240 2160 2160 2200
rect 1240 1240 1280 2160
rect 2120 1240 2160 2160
rect 1240 1200 2160 1240
rect 2440 2160 3360 2200
rect 2440 1240 2480 2160
rect 3320 1240 3360 2160
rect 2440 1200 3360 1240
rect 3640 2160 4560 2200
rect 3640 1240 3680 2160
rect 4520 1240 4560 2160
rect 3640 1200 4560 1240
rect 4840 2160 5760 2200
rect 4840 1240 4880 2160
rect 5720 1240 5760 2160
rect 4840 1200 5760 1240
rect 6040 2160 6960 2200
rect 6040 1240 6080 2160
rect 6920 1240 6960 2160
rect 6040 1200 6960 1240
rect 7200 2160 7320 2200
rect 7200 1240 7240 2160
rect 7280 1240 7320 2160
rect 7200 1200 7320 1240
<< mimcapcontact >>
rect -6280 2440 -6240 3360
rect -5920 2440 -5080 3360
rect -4720 2440 -3880 3360
rect -3520 2440 -2680 3360
rect -2320 2440 -1480 3360
rect -1120 2440 -280 3360
rect 80 2440 920 3360
rect 1280 2440 2120 3360
rect 2480 2440 3320 3360
rect 3680 2440 4520 3360
rect 4880 2440 5720 3360
rect 6080 2440 6920 3360
rect 7240 2440 7280 3360
rect -6280 1240 -6240 2160
rect -5920 1240 -5080 2160
rect -4720 1240 -3880 2160
rect -3520 1240 -2680 2160
rect -2320 1240 -1480 2160
rect -1120 1240 -280 2160
rect 80 1240 920 2160
rect 1280 1240 2120 2160
rect 2480 1240 3320 2160
rect 3680 1240 4520 2160
rect 4880 1240 5720 2160
rect 6080 1240 6920 2160
rect 7240 1240 7280 2160
<< metal4 >>
rect -6360 3836 7440 3840
rect -6360 3804 -6356 3836
rect -6324 3804 -6276 3836
rect -6244 3804 -6196 3836
rect -6164 3804 7164 3836
rect 7196 3804 7244 3836
rect 7276 3804 7324 3836
rect 7356 3804 7440 3836
rect -6360 3800 7440 3804
rect -6360 3756 7440 3760
rect -6360 3724 -5516 3756
rect -5484 3724 -4316 3756
rect -4284 3724 -3116 3756
rect -3084 3724 -1916 3756
rect -1884 3724 -716 3756
rect -684 3724 1684 3756
rect 1716 3724 2884 3756
rect 2916 3724 4084 3756
rect 4116 3724 5284 3756
rect 5316 3724 6484 3756
rect 6516 3724 7440 3756
rect -6360 3720 7440 3724
rect -6360 3676 7440 3680
rect -6360 3644 -6356 3676
rect -6324 3644 -6276 3676
rect -6244 3644 -6196 3676
rect -6164 3644 7164 3676
rect 7196 3644 7244 3676
rect 7276 3644 7324 3676
rect 7356 3644 7440 3676
rect -6360 3640 7440 3644
rect -6360 3596 7440 3600
rect -6360 3564 484 3596
rect 516 3564 7440 3596
rect -6360 3560 7440 3564
rect -6360 3516 7440 3520
rect -6360 3484 -6356 3516
rect -6324 3484 -6276 3516
rect -6244 3484 -6196 3516
rect -6164 3484 -6116 3516
rect -6084 3484 -4916 3516
rect -4884 3484 -3716 3516
rect -3684 3484 -2516 3516
rect -2484 3484 -1316 3516
rect -1284 3484 -116 3516
rect -84 3484 1084 3516
rect 1116 3484 2284 3516
rect 2316 3484 3484 3516
rect 3516 3484 4684 3516
rect 4716 3484 5884 3516
rect 5916 3484 7084 3516
rect 7116 3484 7164 3516
rect 7196 3484 7244 3516
rect 7276 3484 7324 3516
rect 7356 3484 7440 3516
rect -6360 3480 7440 3484
rect -6360 3440 -6320 3480
rect -6280 3440 -6240 3480
rect -6200 3440 -6160 3480
rect -6360 3360 -6160 3440
rect -6360 2440 -6280 3360
rect -6240 2440 -6160 3360
rect -6360 2360 -6160 2440
rect -6120 2360 -6080 3480
rect -6000 3360 -5000 3440
rect -6000 2440 -5920 3360
rect -5080 2440 -5000 3360
rect -6000 2360 -5000 2440
rect -4920 2360 -4880 3480
rect -4800 3360 -3800 3440
rect -4800 2440 -4720 3360
rect -3880 2440 -3800 3360
rect -4800 2360 -3800 2440
rect -3720 2360 -3680 3480
rect -3600 3360 -2600 3440
rect -3600 2440 -3520 3360
rect -2680 2440 -2600 3360
rect -3600 2360 -2600 2440
rect -2520 2360 -2480 3480
rect -2400 3360 -1400 3440
rect -2400 2440 -2320 3360
rect -1480 2440 -1400 3360
rect -2400 2360 -1400 2440
rect -1320 2360 -1280 3480
rect -1200 3360 -200 3440
rect -1200 2440 -1120 3360
rect -280 2440 -200 3360
rect -1200 2360 -200 2440
rect -120 2360 -80 3480
rect 0 3360 1000 3440
rect 0 2440 80 3360
rect 920 2440 1000 3360
rect 0 2360 1000 2440
rect 1080 2360 1120 3480
rect 1200 3360 2200 3440
rect 1200 2440 1280 3360
rect 2120 2440 2200 3360
rect 1200 2360 2200 2440
rect 2280 2360 2320 3480
rect 2400 3360 3400 3440
rect 2400 2440 2480 3360
rect 3320 2440 3400 3360
rect 2400 2360 3400 2440
rect 3480 2360 3520 3480
rect 3600 3360 4600 3440
rect 3600 2440 3680 3360
rect 4520 2440 4600 3360
rect 3600 2360 4600 2440
rect 4680 2360 4720 3480
rect 4800 3360 5800 3440
rect 4800 2440 4880 3360
rect 5720 2440 5800 3360
rect 4800 2360 5800 2440
rect 5880 2360 5920 3480
rect 6000 3360 7000 3440
rect 6000 2440 6080 3360
rect 6920 2440 7000 3360
rect 6000 2360 7000 2440
rect 7080 2360 7120 3480
rect 7160 3440 7200 3480
rect 7240 3440 7280 3480
rect 7320 3440 7360 3480
rect 7160 3360 7360 3440
rect 7160 2440 7240 3360
rect 7280 2440 7360 3360
rect 7160 2360 7360 2440
rect -6000 2320 -5960 2360
rect -5920 2320 -5840 2360
rect -5800 2320 -5760 2360
rect -5720 2320 -5680 2360
rect -5640 2320 -5600 2360
rect -5560 2320 -5520 2360
rect -5480 2320 -5440 2360
rect -5400 2320 -5360 2360
rect -5320 2320 -5280 2360
rect -5240 2320 -5200 2360
rect -5160 2320 -5080 2360
rect -5040 2320 -5000 2360
rect -4800 2320 -4760 2360
rect -4720 2320 -4640 2360
rect -4600 2320 -4560 2360
rect -4520 2320 -4480 2360
rect -4440 2320 -4400 2360
rect -4360 2320 -4320 2360
rect -4280 2320 -4240 2360
rect -4200 2320 -4160 2360
rect -4120 2320 -4080 2360
rect -4040 2320 -4000 2360
rect -3960 2320 -3880 2360
rect -3840 2320 -3800 2360
rect -3600 2320 -3560 2360
rect -3520 2320 -3440 2360
rect -3400 2320 -3360 2360
rect -3320 2320 -3280 2360
rect -3240 2320 -3200 2360
rect -3160 2320 -3120 2360
rect -3080 2320 -3040 2360
rect -3000 2320 -2960 2360
rect -2920 2320 -2880 2360
rect -2840 2320 -2800 2360
rect -2760 2320 -2680 2360
rect -2640 2320 -2600 2360
rect -2400 2320 -2360 2360
rect -2320 2320 -2240 2360
rect -2200 2320 -2160 2360
rect -2120 2320 -2080 2360
rect -2040 2320 -2000 2360
rect -1960 2320 -1920 2360
rect -1880 2320 -1840 2360
rect -1800 2320 -1760 2360
rect -1720 2320 -1680 2360
rect -1640 2320 -1600 2360
rect -1560 2320 -1480 2360
rect -1440 2320 -1400 2360
rect -1200 2320 -1160 2360
rect -1120 2320 -1040 2360
rect -1000 2320 -960 2360
rect -920 2320 -880 2360
rect -840 2320 -800 2360
rect -760 2320 -720 2360
rect -680 2320 -640 2360
rect -600 2320 -560 2360
rect -520 2320 -480 2360
rect -440 2320 -400 2360
rect -360 2320 -280 2360
rect -240 2320 -200 2360
rect 0 2320 40 2360
rect 80 2320 160 2360
rect 200 2320 240 2360
rect 280 2320 320 2360
rect 360 2320 400 2360
rect 440 2320 480 2360
rect 520 2320 560 2360
rect 600 2320 640 2360
rect 680 2320 720 2360
rect 760 2320 800 2360
rect 840 2320 920 2360
rect 960 2320 1000 2360
rect 1200 2320 1240 2360
rect 1280 2320 1360 2360
rect 1400 2320 1440 2360
rect 1480 2320 1520 2360
rect 1560 2320 1600 2360
rect 1640 2320 1680 2360
rect 1720 2320 1760 2360
rect 1800 2320 1840 2360
rect 1880 2320 1920 2360
rect 1960 2320 2000 2360
rect 2040 2320 2120 2360
rect 2160 2320 2200 2360
rect 2400 2320 2440 2360
rect 2480 2320 2560 2360
rect 2600 2320 2640 2360
rect 2680 2320 2720 2360
rect 2760 2320 2800 2360
rect 2840 2320 2880 2360
rect 2920 2320 2960 2360
rect 3000 2320 3040 2360
rect 3080 2320 3120 2360
rect 3160 2320 3200 2360
rect 3240 2320 3320 2360
rect 3360 2320 3400 2360
rect 3600 2320 3640 2360
rect 3680 2320 3760 2360
rect 3800 2320 3840 2360
rect 3880 2320 3920 2360
rect 3960 2320 4000 2360
rect 4040 2320 4080 2360
rect 4120 2320 4160 2360
rect 4200 2320 4240 2360
rect 4280 2320 4320 2360
rect 4360 2320 4400 2360
rect 4440 2320 4520 2360
rect 4560 2320 4600 2360
rect 4800 2320 4840 2360
rect 4880 2320 4960 2360
rect 5000 2320 5040 2360
rect 5080 2320 5120 2360
rect 5160 2320 5200 2360
rect 5240 2320 5280 2360
rect 5320 2320 5360 2360
rect 5400 2320 5440 2360
rect 5480 2320 5520 2360
rect 5560 2320 5600 2360
rect 5640 2320 5720 2360
rect 5760 2320 5800 2360
rect 6000 2320 6040 2360
rect 6080 2320 6160 2360
rect 6200 2320 6240 2360
rect 6280 2320 6320 2360
rect 6360 2320 6400 2360
rect 6440 2320 6480 2360
rect 6520 2320 6560 2360
rect 6600 2320 6640 2360
rect 6680 2320 6720 2360
rect 6760 2320 6800 2360
rect 6840 2320 6920 2360
rect 6960 2320 7000 2360
rect -6400 2280 7440 2320
rect -6000 2240 -5960 2280
rect -5920 2240 -5840 2280
rect -5800 2240 -5760 2280
rect -5720 2240 -5680 2280
rect -5640 2240 -5600 2280
rect -5560 2240 -5520 2280
rect -5480 2240 -5440 2280
rect -5400 2240 -5360 2280
rect -5320 2240 -5280 2280
rect -5240 2240 -5200 2280
rect -5160 2240 -5080 2280
rect -5040 2240 -5000 2280
rect -4800 2240 -4760 2280
rect -4720 2240 -4640 2280
rect -4600 2240 -4560 2280
rect -4520 2240 -4480 2280
rect -4440 2240 -4400 2280
rect -4360 2240 -4320 2280
rect -4280 2240 -4240 2280
rect -4200 2240 -4160 2280
rect -4120 2240 -4080 2280
rect -4040 2240 -4000 2280
rect -3960 2240 -3880 2280
rect -3840 2240 -3800 2280
rect -3600 2240 -3560 2280
rect -3520 2240 -3440 2280
rect -3400 2240 -3360 2280
rect -3320 2240 -3280 2280
rect -3240 2240 -3200 2280
rect -3160 2240 -3120 2280
rect -3080 2240 -3040 2280
rect -3000 2240 -2960 2280
rect -2920 2240 -2880 2280
rect -2840 2240 -2800 2280
rect -2760 2240 -2680 2280
rect -2640 2240 -2600 2280
rect -2400 2240 -2360 2280
rect -2320 2240 -2240 2280
rect -2200 2240 -2160 2280
rect -2120 2240 -2080 2280
rect -2040 2240 -2000 2280
rect -1960 2240 -1920 2280
rect -1880 2240 -1840 2280
rect -1800 2240 -1760 2280
rect -1720 2240 -1680 2280
rect -1640 2240 -1600 2280
rect -1560 2240 -1480 2280
rect -1440 2240 -1400 2280
rect -1200 2240 -1160 2280
rect -1120 2240 -1040 2280
rect -1000 2240 -960 2280
rect -920 2240 -880 2280
rect -840 2240 -800 2280
rect -760 2240 -720 2280
rect -680 2240 -640 2280
rect -600 2240 -560 2280
rect -520 2240 -480 2280
rect -440 2240 -400 2280
rect -360 2240 -280 2280
rect -240 2240 -200 2280
rect 0 2240 40 2280
rect 80 2240 160 2280
rect 200 2240 240 2280
rect 280 2240 320 2280
rect 360 2240 400 2280
rect 440 2240 480 2280
rect 520 2240 560 2280
rect 600 2240 640 2280
rect 680 2240 720 2280
rect 760 2240 800 2280
rect 840 2240 920 2280
rect 960 2240 1000 2280
rect 1200 2240 1240 2280
rect 1280 2240 1360 2280
rect 1400 2240 1440 2280
rect 1480 2240 1520 2280
rect 1560 2240 1600 2280
rect 1640 2240 1680 2280
rect 1720 2240 1760 2280
rect 1800 2240 1840 2280
rect 1880 2240 1920 2280
rect 1960 2240 2000 2280
rect 2040 2240 2120 2280
rect 2160 2240 2200 2280
rect 2400 2240 2440 2280
rect 2480 2240 2560 2280
rect 2600 2240 2640 2280
rect 2680 2240 2720 2280
rect 2760 2240 2800 2280
rect 2840 2240 2880 2280
rect 2920 2240 2960 2280
rect 3000 2240 3040 2280
rect 3080 2240 3120 2280
rect 3160 2240 3200 2280
rect 3240 2240 3320 2280
rect 3360 2240 3400 2280
rect 3600 2240 3640 2280
rect 3680 2240 3760 2280
rect 3800 2240 3840 2280
rect 3880 2240 3920 2280
rect 3960 2240 4000 2280
rect 4040 2240 4080 2280
rect 4120 2240 4160 2280
rect 4200 2240 4240 2280
rect 4280 2240 4320 2280
rect 4360 2240 4400 2280
rect 4440 2240 4520 2280
rect 4560 2240 4600 2280
rect 4800 2240 4840 2280
rect 4880 2240 4960 2280
rect 5000 2240 5040 2280
rect 5080 2240 5120 2280
rect 5160 2240 5200 2280
rect 5240 2240 5280 2280
rect 5320 2240 5360 2280
rect 5400 2240 5440 2280
rect 5480 2240 5520 2280
rect 5560 2240 5600 2280
rect 5640 2240 5720 2280
rect 5760 2240 5800 2280
rect 6000 2240 6040 2280
rect 6080 2240 6160 2280
rect 6200 2240 6240 2280
rect 6280 2240 6320 2280
rect 6360 2240 6400 2280
rect 6440 2240 6480 2280
rect 6520 2240 6560 2280
rect 6600 2240 6640 2280
rect 6680 2240 6720 2280
rect 6760 2240 6800 2280
rect 6840 2240 6920 2280
rect 6960 2240 7000 2280
rect -6360 2160 -6160 2240
rect -6360 1240 -6280 2160
rect -6240 1240 -6160 2160
rect -6360 1160 -6160 1240
rect -6360 1120 -6320 1160
rect -6280 1120 -6240 1160
rect -6200 1120 -6160 1160
rect -6120 1120 -6080 2240
rect -6000 2160 -5000 2240
rect -6000 1240 -5920 2160
rect -5080 1240 -5000 2160
rect -6000 1160 -5000 1240
rect -4920 1120 -4880 2240
rect -4800 2160 -3800 2240
rect -4800 1240 -4720 2160
rect -3880 1240 -3800 2160
rect -4800 1160 -3800 1240
rect -3720 1120 -3680 2240
rect -3600 2160 -2600 2240
rect -3600 1240 -3520 2160
rect -2680 1240 -2600 2160
rect -3600 1160 -2600 1240
rect -2520 1120 -2480 2240
rect -2400 2160 -1400 2240
rect -2400 1240 -2320 2160
rect -1480 1240 -1400 2160
rect -2400 1160 -1400 1240
rect -1320 1120 -1280 2240
rect -1200 2160 -200 2240
rect -1200 1240 -1120 2160
rect -280 1240 -200 2160
rect -1200 1160 -200 1240
rect -120 1120 -80 2240
rect 0 2160 1000 2240
rect 0 1240 80 2160
rect 920 1240 1000 2160
rect 0 1160 1000 1240
rect 1080 1120 1120 2240
rect 1200 2160 2200 2240
rect 1200 1240 1280 2160
rect 2120 1240 2200 2160
rect 1200 1160 2200 1240
rect 2280 1120 2320 2240
rect 2400 2160 3400 2240
rect 2400 1240 2480 2160
rect 3320 1240 3400 2160
rect 2400 1160 3400 1240
rect 3480 1120 3520 2240
rect 3600 2160 4600 2240
rect 3600 1240 3680 2160
rect 4520 1240 4600 2160
rect 3600 1160 4600 1240
rect 4680 1120 4720 2240
rect 4800 2160 5800 2240
rect 4800 1240 4880 2160
rect 5720 1240 5800 2160
rect 4800 1160 5800 1240
rect 5880 1120 5920 2240
rect 6000 2160 7000 2240
rect 6000 1240 6080 2160
rect 6920 1240 7000 2160
rect 6000 1160 7000 1240
rect 7080 1120 7120 2240
rect 7160 2160 7360 2240
rect 7160 1240 7240 2160
rect 7280 1240 7360 2160
rect 7160 1160 7360 1240
rect 7160 1120 7200 1160
rect 7240 1120 7280 1160
rect 7320 1120 7360 1160
rect -6400 1116 7440 1120
rect -6400 1084 -6356 1116
rect -6324 1084 -6276 1116
rect -6244 1084 -6196 1116
rect -6164 1084 -6116 1116
rect -6084 1084 -4916 1116
rect -4884 1084 -3716 1116
rect -3684 1084 -2516 1116
rect -2484 1084 -1316 1116
rect -1284 1084 -116 1116
rect -84 1084 1084 1116
rect 1116 1084 2284 1116
rect 2316 1084 3484 1116
rect 3516 1084 4684 1116
rect 4716 1084 5884 1116
rect 5916 1084 7084 1116
rect 7116 1084 7164 1116
rect 7196 1084 7244 1116
rect 7276 1084 7324 1116
rect 7356 1084 7440 1116
rect -6400 1080 7440 1084
rect -6400 1036 7440 1040
rect -6400 1004 484 1036
rect 516 1004 7440 1036
rect -6400 1000 7440 1004
rect -6400 956 7440 960
rect -6400 924 -6356 956
rect -6324 924 -6276 956
rect -6244 924 -6196 956
rect -6164 924 7164 956
rect 7196 924 7244 956
rect 7276 924 7324 956
rect 7356 924 7440 956
rect -6400 920 7440 924
rect -6400 876 7440 880
rect -6400 844 -5516 876
rect -5484 844 -4316 876
rect -4284 844 -3116 876
rect -3084 844 -1916 876
rect -1884 844 -716 876
rect -684 844 1684 876
rect 1716 844 2884 876
rect 2916 844 4084 876
rect 4116 844 5284 876
rect 5316 844 6484 876
rect 6516 844 7440 876
rect -6400 840 7440 844
rect -6400 796 7440 800
rect -6400 764 -6356 796
rect -6324 764 -6276 796
rect -6244 764 -6196 796
rect -6164 764 7164 796
rect 7196 764 7244 796
rect 7276 764 7324 796
rect 7356 764 7440 796
rect -6400 760 7440 764
<< labels >>
rlabel locali 7400 680 7440 720 0 vssa
port 6 nsew
rlabel metal4 7400 3560 7440 3600 0 b1
port 1 nsew
rlabel metal4 7400 3720 7440 3760 0 c1
port 3 nsew
rlabel metal4 7400 1000 7440 1040 0 b2
port 2 nsew
rlabel metal4 7400 840 7440 880 0 c2
port 4 nsew
rlabel metal4 7400 3640 7440 3680 0 gnda
port 5 nsew
rlabel metal4 7400 2280 7440 2320 0 a
port 0 nsew
<< end >>
