magic
tech sky130A
magscale 1 2
timestamp 1634821592
<< error_p >>
rect 305 -638 363 -632
rect 305 -672 317 -638
rect 305 -678 363 -672
<< pwell >>
rect -583 -526 583 526
<< nmos >>
rect -495 -500 -465 500
rect -399 -500 -369 500
rect -303 -500 -273 500
rect -207 -500 -177 500
rect -111 -500 -81 500
rect -15 -500 15 500
rect 81 -500 111 500
rect 177 -500 207 500
rect 273 -500 303 500
rect 369 -500 399 500
rect 465 -500 495 500
<< ndiff >>
rect -557 459 -495 500
rect -557 425 -545 459
rect -511 425 -495 459
rect -557 391 -495 425
rect -557 357 -545 391
rect -511 357 -495 391
rect -557 323 -495 357
rect -557 289 -545 323
rect -511 289 -495 323
rect -557 255 -495 289
rect -557 221 -545 255
rect -511 221 -495 255
rect -557 187 -495 221
rect -557 153 -545 187
rect -511 153 -495 187
rect -557 119 -495 153
rect -557 85 -545 119
rect -511 85 -495 119
rect -557 51 -495 85
rect -557 17 -545 51
rect -511 17 -495 51
rect -557 -17 -495 17
rect -557 -51 -545 -17
rect -511 -51 -495 -17
rect -557 -85 -495 -51
rect -557 -119 -545 -85
rect -511 -119 -495 -85
rect -557 -153 -495 -119
rect -557 -187 -545 -153
rect -511 -187 -495 -153
rect -557 -221 -495 -187
rect -557 -255 -545 -221
rect -511 -255 -495 -221
rect -557 -289 -495 -255
rect -557 -323 -545 -289
rect -511 -323 -495 -289
rect -557 -357 -495 -323
rect -557 -391 -545 -357
rect -511 -391 -495 -357
rect -557 -425 -495 -391
rect -557 -459 -545 -425
rect -511 -459 -495 -425
rect -557 -500 -495 -459
rect -465 459 -399 500
rect -465 425 -449 459
rect -415 425 -399 459
rect -465 391 -399 425
rect -465 357 -449 391
rect -415 357 -399 391
rect -465 323 -399 357
rect -465 289 -449 323
rect -415 289 -399 323
rect -465 255 -399 289
rect -465 221 -449 255
rect -415 221 -399 255
rect -465 187 -399 221
rect -465 153 -449 187
rect -415 153 -399 187
rect -465 119 -399 153
rect -465 85 -449 119
rect -415 85 -399 119
rect -465 51 -399 85
rect -465 17 -449 51
rect -415 17 -399 51
rect -465 -17 -399 17
rect -465 -51 -449 -17
rect -415 -51 -399 -17
rect -465 -85 -399 -51
rect -465 -119 -449 -85
rect -415 -119 -399 -85
rect -465 -153 -399 -119
rect -465 -187 -449 -153
rect -415 -187 -399 -153
rect -465 -221 -399 -187
rect -465 -255 -449 -221
rect -415 -255 -399 -221
rect -465 -289 -399 -255
rect -465 -323 -449 -289
rect -415 -323 -399 -289
rect -465 -357 -399 -323
rect -465 -391 -449 -357
rect -415 -391 -399 -357
rect -465 -425 -399 -391
rect -465 -459 -449 -425
rect -415 -459 -399 -425
rect -465 -500 -399 -459
rect -369 459 -303 500
rect -369 425 -353 459
rect -319 425 -303 459
rect -369 391 -303 425
rect -369 357 -353 391
rect -319 357 -303 391
rect -369 323 -303 357
rect -369 289 -353 323
rect -319 289 -303 323
rect -369 255 -303 289
rect -369 221 -353 255
rect -319 221 -303 255
rect -369 187 -303 221
rect -369 153 -353 187
rect -319 153 -303 187
rect -369 119 -303 153
rect -369 85 -353 119
rect -319 85 -303 119
rect -369 51 -303 85
rect -369 17 -353 51
rect -319 17 -303 51
rect -369 -17 -303 17
rect -369 -51 -353 -17
rect -319 -51 -303 -17
rect -369 -85 -303 -51
rect -369 -119 -353 -85
rect -319 -119 -303 -85
rect -369 -153 -303 -119
rect -369 -187 -353 -153
rect -319 -187 -303 -153
rect -369 -221 -303 -187
rect -369 -255 -353 -221
rect -319 -255 -303 -221
rect -369 -289 -303 -255
rect -369 -323 -353 -289
rect -319 -323 -303 -289
rect -369 -357 -303 -323
rect -369 -391 -353 -357
rect -319 -391 -303 -357
rect -369 -425 -303 -391
rect -369 -459 -353 -425
rect -319 -459 -303 -425
rect -369 -500 -303 -459
rect -273 459 -207 500
rect -273 425 -257 459
rect -223 425 -207 459
rect -273 391 -207 425
rect -273 357 -257 391
rect -223 357 -207 391
rect -273 323 -207 357
rect -273 289 -257 323
rect -223 289 -207 323
rect -273 255 -207 289
rect -273 221 -257 255
rect -223 221 -207 255
rect -273 187 -207 221
rect -273 153 -257 187
rect -223 153 -207 187
rect -273 119 -207 153
rect -273 85 -257 119
rect -223 85 -207 119
rect -273 51 -207 85
rect -273 17 -257 51
rect -223 17 -207 51
rect -273 -17 -207 17
rect -273 -51 -257 -17
rect -223 -51 -207 -17
rect -273 -85 -207 -51
rect -273 -119 -257 -85
rect -223 -119 -207 -85
rect -273 -153 -207 -119
rect -273 -187 -257 -153
rect -223 -187 -207 -153
rect -273 -221 -207 -187
rect -273 -255 -257 -221
rect -223 -255 -207 -221
rect -273 -289 -207 -255
rect -273 -323 -257 -289
rect -223 -323 -207 -289
rect -273 -357 -207 -323
rect -273 -391 -257 -357
rect -223 -391 -207 -357
rect -273 -425 -207 -391
rect -273 -459 -257 -425
rect -223 -459 -207 -425
rect -273 -500 -207 -459
rect -177 459 -111 500
rect -177 425 -161 459
rect -127 425 -111 459
rect -177 391 -111 425
rect -177 357 -161 391
rect -127 357 -111 391
rect -177 323 -111 357
rect -177 289 -161 323
rect -127 289 -111 323
rect -177 255 -111 289
rect -177 221 -161 255
rect -127 221 -111 255
rect -177 187 -111 221
rect -177 153 -161 187
rect -127 153 -111 187
rect -177 119 -111 153
rect -177 85 -161 119
rect -127 85 -111 119
rect -177 51 -111 85
rect -177 17 -161 51
rect -127 17 -111 51
rect -177 -17 -111 17
rect -177 -51 -161 -17
rect -127 -51 -111 -17
rect -177 -85 -111 -51
rect -177 -119 -161 -85
rect -127 -119 -111 -85
rect -177 -153 -111 -119
rect -177 -187 -161 -153
rect -127 -187 -111 -153
rect -177 -221 -111 -187
rect -177 -255 -161 -221
rect -127 -255 -111 -221
rect -177 -289 -111 -255
rect -177 -323 -161 -289
rect -127 -323 -111 -289
rect -177 -357 -111 -323
rect -177 -391 -161 -357
rect -127 -391 -111 -357
rect -177 -425 -111 -391
rect -177 -459 -161 -425
rect -127 -459 -111 -425
rect -177 -500 -111 -459
rect -81 459 -15 500
rect -81 425 -65 459
rect -31 425 -15 459
rect -81 391 -15 425
rect -81 357 -65 391
rect -31 357 -15 391
rect -81 323 -15 357
rect -81 289 -65 323
rect -31 289 -15 323
rect -81 255 -15 289
rect -81 221 -65 255
rect -31 221 -15 255
rect -81 187 -15 221
rect -81 153 -65 187
rect -31 153 -15 187
rect -81 119 -15 153
rect -81 85 -65 119
rect -31 85 -15 119
rect -81 51 -15 85
rect -81 17 -65 51
rect -31 17 -15 51
rect -81 -17 -15 17
rect -81 -51 -65 -17
rect -31 -51 -15 -17
rect -81 -85 -15 -51
rect -81 -119 -65 -85
rect -31 -119 -15 -85
rect -81 -153 -15 -119
rect -81 -187 -65 -153
rect -31 -187 -15 -153
rect -81 -221 -15 -187
rect -81 -255 -65 -221
rect -31 -255 -15 -221
rect -81 -289 -15 -255
rect -81 -323 -65 -289
rect -31 -323 -15 -289
rect -81 -357 -15 -323
rect -81 -391 -65 -357
rect -31 -391 -15 -357
rect -81 -425 -15 -391
rect -81 -459 -65 -425
rect -31 -459 -15 -425
rect -81 -500 -15 -459
rect 15 459 81 500
rect 15 425 31 459
rect 65 425 81 459
rect 15 391 81 425
rect 15 357 31 391
rect 65 357 81 391
rect 15 323 81 357
rect 15 289 31 323
rect 65 289 81 323
rect 15 255 81 289
rect 15 221 31 255
rect 65 221 81 255
rect 15 187 81 221
rect 15 153 31 187
rect 65 153 81 187
rect 15 119 81 153
rect 15 85 31 119
rect 65 85 81 119
rect 15 51 81 85
rect 15 17 31 51
rect 65 17 81 51
rect 15 -17 81 17
rect 15 -51 31 -17
rect 65 -51 81 -17
rect 15 -85 81 -51
rect 15 -119 31 -85
rect 65 -119 81 -85
rect 15 -153 81 -119
rect 15 -187 31 -153
rect 65 -187 81 -153
rect 15 -221 81 -187
rect 15 -255 31 -221
rect 65 -255 81 -221
rect 15 -289 81 -255
rect 15 -323 31 -289
rect 65 -323 81 -289
rect 15 -357 81 -323
rect 15 -391 31 -357
rect 65 -391 81 -357
rect 15 -425 81 -391
rect 15 -459 31 -425
rect 65 -459 81 -425
rect 15 -500 81 -459
rect 111 459 177 500
rect 111 425 127 459
rect 161 425 177 459
rect 111 391 177 425
rect 111 357 127 391
rect 161 357 177 391
rect 111 323 177 357
rect 111 289 127 323
rect 161 289 177 323
rect 111 255 177 289
rect 111 221 127 255
rect 161 221 177 255
rect 111 187 177 221
rect 111 153 127 187
rect 161 153 177 187
rect 111 119 177 153
rect 111 85 127 119
rect 161 85 177 119
rect 111 51 177 85
rect 111 17 127 51
rect 161 17 177 51
rect 111 -17 177 17
rect 111 -51 127 -17
rect 161 -51 177 -17
rect 111 -85 177 -51
rect 111 -119 127 -85
rect 161 -119 177 -85
rect 111 -153 177 -119
rect 111 -187 127 -153
rect 161 -187 177 -153
rect 111 -221 177 -187
rect 111 -255 127 -221
rect 161 -255 177 -221
rect 111 -289 177 -255
rect 111 -323 127 -289
rect 161 -323 177 -289
rect 111 -357 177 -323
rect 111 -391 127 -357
rect 161 -391 177 -357
rect 111 -425 177 -391
rect 111 -459 127 -425
rect 161 -459 177 -425
rect 111 -500 177 -459
rect 207 459 273 500
rect 207 425 223 459
rect 257 425 273 459
rect 207 391 273 425
rect 207 357 223 391
rect 257 357 273 391
rect 207 323 273 357
rect 207 289 223 323
rect 257 289 273 323
rect 207 255 273 289
rect 207 221 223 255
rect 257 221 273 255
rect 207 187 273 221
rect 207 153 223 187
rect 257 153 273 187
rect 207 119 273 153
rect 207 85 223 119
rect 257 85 273 119
rect 207 51 273 85
rect 207 17 223 51
rect 257 17 273 51
rect 207 -17 273 17
rect 207 -51 223 -17
rect 257 -51 273 -17
rect 207 -85 273 -51
rect 207 -119 223 -85
rect 257 -119 273 -85
rect 207 -153 273 -119
rect 207 -187 223 -153
rect 257 -187 273 -153
rect 207 -221 273 -187
rect 207 -255 223 -221
rect 257 -255 273 -221
rect 207 -289 273 -255
rect 207 -323 223 -289
rect 257 -323 273 -289
rect 207 -357 273 -323
rect 207 -391 223 -357
rect 257 -391 273 -357
rect 207 -425 273 -391
rect 207 -459 223 -425
rect 257 -459 273 -425
rect 207 -500 273 -459
rect 303 459 369 500
rect 303 425 319 459
rect 353 425 369 459
rect 303 391 369 425
rect 303 357 319 391
rect 353 357 369 391
rect 303 323 369 357
rect 303 289 319 323
rect 353 289 369 323
rect 303 255 369 289
rect 303 221 319 255
rect 353 221 369 255
rect 303 187 369 221
rect 303 153 319 187
rect 353 153 369 187
rect 303 119 369 153
rect 303 85 319 119
rect 353 85 369 119
rect 303 51 369 85
rect 303 17 319 51
rect 353 17 369 51
rect 303 -17 369 17
rect 303 -51 319 -17
rect 353 -51 369 -17
rect 303 -85 369 -51
rect 303 -119 319 -85
rect 353 -119 369 -85
rect 303 -153 369 -119
rect 303 -187 319 -153
rect 353 -187 369 -153
rect 303 -221 369 -187
rect 303 -255 319 -221
rect 353 -255 369 -221
rect 303 -289 369 -255
rect 303 -323 319 -289
rect 353 -323 369 -289
rect 303 -357 369 -323
rect 303 -391 319 -357
rect 353 -391 369 -357
rect 303 -425 369 -391
rect 303 -459 319 -425
rect 353 -459 369 -425
rect 303 -500 369 -459
rect 399 459 465 500
rect 399 425 415 459
rect 449 425 465 459
rect 399 391 465 425
rect 399 357 415 391
rect 449 357 465 391
rect 399 323 465 357
rect 399 289 415 323
rect 449 289 465 323
rect 399 255 465 289
rect 399 221 415 255
rect 449 221 465 255
rect 399 187 465 221
rect 399 153 415 187
rect 449 153 465 187
rect 399 119 465 153
rect 399 85 415 119
rect 449 85 465 119
rect 399 51 465 85
rect 399 17 415 51
rect 449 17 465 51
rect 399 -17 465 17
rect 399 -51 415 -17
rect 449 -51 465 -17
rect 399 -85 465 -51
rect 399 -119 415 -85
rect 449 -119 465 -85
rect 399 -153 465 -119
rect 399 -187 415 -153
rect 449 -187 465 -153
rect 399 -221 465 -187
rect 399 -255 415 -221
rect 449 -255 465 -221
rect 399 -289 465 -255
rect 399 -323 415 -289
rect 449 -323 465 -289
rect 399 -357 465 -323
rect 399 -391 415 -357
rect 449 -391 465 -357
rect 399 -425 465 -391
rect 399 -459 415 -425
rect 449 -459 465 -425
rect 399 -500 465 -459
rect 495 459 557 500
rect 495 425 511 459
rect 545 425 557 459
rect 495 391 557 425
rect 495 357 511 391
rect 545 357 557 391
rect 495 323 557 357
rect 495 289 511 323
rect 545 289 557 323
rect 495 255 557 289
rect 495 221 511 255
rect 545 221 557 255
rect 495 187 557 221
rect 495 153 511 187
rect 545 153 557 187
rect 495 119 557 153
rect 495 85 511 119
rect 545 85 557 119
rect 495 51 557 85
rect 495 17 511 51
rect 545 17 557 51
rect 495 -17 557 17
rect 495 -51 511 -17
rect 545 -51 557 -17
rect 495 -85 557 -51
rect 495 -119 511 -85
rect 545 -119 557 -85
rect 495 -153 557 -119
rect 495 -187 511 -153
rect 545 -187 557 -153
rect 495 -221 557 -187
rect 495 -255 511 -221
rect 545 -255 557 -221
rect 495 -289 557 -255
rect 495 -323 511 -289
rect 545 -323 557 -289
rect 495 -357 557 -323
rect 495 -391 511 -357
rect 545 -391 557 -357
rect 495 -425 557 -391
rect 495 -459 511 -425
rect 545 -459 557 -425
rect 495 -500 557 -459
<< ndiffc >>
rect -545 425 -511 459
rect -545 357 -511 391
rect -545 289 -511 323
rect -545 221 -511 255
rect -545 153 -511 187
rect -545 85 -511 119
rect -545 17 -511 51
rect -545 -51 -511 -17
rect -545 -119 -511 -85
rect -545 -187 -511 -153
rect -545 -255 -511 -221
rect -545 -323 -511 -289
rect -545 -391 -511 -357
rect -545 -459 -511 -425
rect -449 425 -415 459
rect -449 357 -415 391
rect -449 289 -415 323
rect -449 221 -415 255
rect -449 153 -415 187
rect -449 85 -415 119
rect -449 17 -415 51
rect -449 -51 -415 -17
rect -449 -119 -415 -85
rect -449 -187 -415 -153
rect -449 -255 -415 -221
rect -449 -323 -415 -289
rect -449 -391 -415 -357
rect -449 -459 -415 -425
rect -353 425 -319 459
rect -353 357 -319 391
rect -353 289 -319 323
rect -353 221 -319 255
rect -353 153 -319 187
rect -353 85 -319 119
rect -353 17 -319 51
rect -353 -51 -319 -17
rect -353 -119 -319 -85
rect -353 -187 -319 -153
rect -353 -255 -319 -221
rect -353 -323 -319 -289
rect -353 -391 -319 -357
rect -353 -459 -319 -425
rect -257 425 -223 459
rect -257 357 -223 391
rect -257 289 -223 323
rect -257 221 -223 255
rect -257 153 -223 187
rect -257 85 -223 119
rect -257 17 -223 51
rect -257 -51 -223 -17
rect -257 -119 -223 -85
rect -257 -187 -223 -153
rect -257 -255 -223 -221
rect -257 -323 -223 -289
rect -257 -391 -223 -357
rect -257 -459 -223 -425
rect -161 425 -127 459
rect -161 357 -127 391
rect -161 289 -127 323
rect -161 221 -127 255
rect -161 153 -127 187
rect -161 85 -127 119
rect -161 17 -127 51
rect -161 -51 -127 -17
rect -161 -119 -127 -85
rect -161 -187 -127 -153
rect -161 -255 -127 -221
rect -161 -323 -127 -289
rect -161 -391 -127 -357
rect -161 -459 -127 -425
rect -65 425 -31 459
rect -65 357 -31 391
rect -65 289 -31 323
rect -65 221 -31 255
rect -65 153 -31 187
rect -65 85 -31 119
rect -65 17 -31 51
rect -65 -51 -31 -17
rect -65 -119 -31 -85
rect -65 -187 -31 -153
rect -65 -255 -31 -221
rect -65 -323 -31 -289
rect -65 -391 -31 -357
rect -65 -459 -31 -425
rect 31 425 65 459
rect 31 357 65 391
rect 31 289 65 323
rect 31 221 65 255
rect 31 153 65 187
rect 31 85 65 119
rect 31 17 65 51
rect 31 -51 65 -17
rect 31 -119 65 -85
rect 31 -187 65 -153
rect 31 -255 65 -221
rect 31 -323 65 -289
rect 31 -391 65 -357
rect 31 -459 65 -425
rect 127 425 161 459
rect 127 357 161 391
rect 127 289 161 323
rect 127 221 161 255
rect 127 153 161 187
rect 127 85 161 119
rect 127 17 161 51
rect 127 -51 161 -17
rect 127 -119 161 -85
rect 127 -187 161 -153
rect 127 -255 161 -221
rect 127 -323 161 -289
rect 127 -391 161 -357
rect 127 -459 161 -425
rect 223 425 257 459
rect 223 357 257 391
rect 223 289 257 323
rect 223 221 257 255
rect 223 153 257 187
rect 223 85 257 119
rect 223 17 257 51
rect 223 -51 257 -17
rect 223 -119 257 -85
rect 223 -187 257 -153
rect 223 -255 257 -221
rect 223 -323 257 -289
rect 223 -391 257 -357
rect 223 -459 257 -425
rect 319 425 353 459
rect 319 357 353 391
rect 319 289 353 323
rect 319 221 353 255
rect 319 153 353 187
rect 319 85 353 119
rect 319 17 353 51
rect 319 -51 353 -17
rect 319 -119 353 -85
rect 319 -187 353 -153
rect 319 -255 353 -221
rect 319 -323 353 -289
rect 319 -391 353 -357
rect 319 -459 353 -425
rect 415 425 449 459
rect 415 357 449 391
rect 415 289 449 323
rect 415 221 449 255
rect 415 153 449 187
rect 415 85 449 119
rect 415 17 449 51
rect 415 -51 449 -17
rect 415 -119 449 -85
rect 415 -187 449 -153
rect 415 -255 449 -221
rect 415 -323 449 -289
rect 415 -391 449 -357
rect 415 -459 449 -425
rect 511 425 545 459
rect 511 357 545 391
rect 511 289 545 323
rect 511 221 545 255
rect 511 153 545 187
rect 511 85 545 119
rect 511 17 545 51
rect 511 -51 545 -17
rect 511 -119 545 -85
rect 511 -187 545 -153
rect 511 -255 545 -221
rect 511 -323 545 -289
rect 511 -391 545 -357
rect 511 -459 545 -425
<< poly >>
rect -495 542 495 572
rect -495 500 -465 542
rect -399 500 -369 542
rect -303 500 -273 542
rect -207 500 -177 542
rect -111 500 -81 542
rect -15 500 15 542
rect 81 500 111 542
rect 177 500 207 542
rect 273 500 303 542
rect 369 500 399 542
rect 465 500 495 542
rect -495 -526 -465 -500
rect -399 -526 -369 -500
rect -303 -526 -273 -500
rect -207 -526 -177 -500
rect -111 -526 -81 -500
rect -15 -526 15 -500
rect 81 -526 111 -500
rect 177 -526 207 -500
rect 273 -560 303 -500
rect 369 -526 399 -500
rect 465 -526 495 -500
rect 273 -590 331 -560
rect 301 -622 331 -590
rect 301 -638 367 -622
rect 301 -672 317 -638
rect 351 -672 367 -638
rect 301 -688 367 -672
<< polycont >>
rect 317 -672 351 -638
<< locali >>
rect -449 566 545 600
rect -545 485 -511 504
rect -545 413 -511 425
rect -545 341 -511 357
rect -545 269 -511 289
rect -545 197 -511 221
rect -545 125 -511 153
rect -545 53 -511 85
rect -545 -17 -511 17
rect -545 -85 -511 -53
rect -545 -153 -511 -125
rect -545 -221 -511 -197
rect -545 -289 -511 -269
rect -545 -357 -511 -341
rect -545 -425 -511 -413
rect -545 -552 -511 -485
rect -449 485 -415 566
rect -449 413 -415 425
rect -449 341 -415 357
rect -449 269 -415 289
rect -449 197 -415 221
rect -449 125 -415 153
rect -449 53 -415 85
rect -449 -17 -415 17
rect -449 -85 -415 -53
rect -449 -153 -415 -125
rect -449 -221 -415 -197
rect -449 -289 -415 -269
rect -449 -357 -415 -341
rect -449 -425 -415 -413
rect -449 -504 -415 -485
rect -353 485 -319 504
rect -353 413 -319 425
rect -353 341 -319 357
rect -353 269 -319 289
rect -353 197 -319 221
rect -353 125 -319 153
rect -353 53 -319 85
rect -353 -17 -319 17
rect -353 -85 -319 -53
rect -353 -153 -319 -125
rect -353 -221 -319 -197
rect -353 -289 -319 -269
rect -353 -357 -319 -341
rect -353 -425 -319 -413
rect -353 -552 -319 -485
rect -257 485 -223 566
rect -257 413 -223 425
rect -257 341 -223 357
rect -257 269 -223 289
rect -257 197 -223 221
rect -257 125 -223 153
rect -257 53 -223 85
rect -257 -17 -223 17
rect -257 -85 -223 -53
rect -257 -153 -223 -125
rect -257 -221 -223 -197
rect -257 -289 -223 -269
rect -257 -357 -223 -341
rect -257 -425 -223 -413
rect -257 -504 -223 -485
rect -161 485 -127 504
rect -161 413 -127 425
rect -161 341 -127 357
rect -161 269 -127 289
rect -161 197 -127 221
rect -161 125 -127 153
rect -161 53 -127 85
rect -161 -17 -127 17
rect -161 -85 -127 -53
rect -161 -153 -127 -125
rect -161 -221 -127 -197
rect -161 -289 -127 -269
rect -161 -357 -127 -341
rect -161 -425 -127 -413
rect -161 -552 -127 -485
rect -65 485 -31 566
rect -65 413 -31 425
rect -65 341 -31 357
rect -65 269 -31 289
rect -65 197 -31 221
rect -65 125 -31 153
rect -65 53 -31 85
rect -65 -17 -31 17
rect -65 -85 -31 -53
rect -65 -153 -31 -125
rect -65 -221 -31 -197
rect -65 -289 -31 -269
rect -65 -357 -31 -341
rect -65 -425 -31 -413
rect -65 -504 -31 -485
rect 31 485 65 504
rect 31 413 65 425
rect 31 341 65 357
rect 31 269 65 289
rect 31 197 65 221
rect 31 125 65 153
rect 31 53 65 85
rect 31 -17 65 17
rect 31 -85 65 -53
rect 31 -153 65 -125
rect 31 -221 65 -197
rect 31 -289 65 -269
rect 31 -357 65 -341
rect 31 -425 65 -413
rect 31 -552 65 -485
rect 127 485 161 566
rect 127 413 161 425
rect 127 341 161 357
rect 127 269 161 289
rect 127 197 161 221
rect 127 125 161 153
rect 127 53 161 85
rect 127 -17 161 17
rect 127 -85 161 -53
rect 127 -153 161 -125
rect 127 -221 161 -197
rect 127 -289 161 -269
rect 127 -357 161 -341
rect 127 -425 161 -413
rect 127 -502 161 -485
rect 223 485 257 504
rect 223 413 257 425
rect 223 341 257 357
rect 223 269 257 289
rect 223 197 257 221
rect 223 125 257 153
rect 223 53 257 85
rect 223 -17 257 17
rect 223 -85 257 -53
rect 223 -153 257 -125
rect 223 -221 257 -197
rect 223 -289 257 -269
rect 223 -357 257 -341
rect 223 -425 257 -413
rect 223 -552 257 -485
rect 319 485 353 566
rect 319 413 353 425
rect 319 341 353 357
rect 319 269 353 289
rect 319 197 353 221
rect 319 125 353 153
rect 319 53 353 85
rect 319 -17 353 17
rect 319 -85 353 -53
rect 319 -153 353 -125
rect 319 -221 353 -197
rect 319 -289 353 -269
rect 319 -357 353 -341
rect 319 -425 353 -413
rect 319 -502 353 -485
rect 415 485 449 504
rect 415 413 449 425
rect 415 341 449 357
rect 415 269 449 289
rect 415 197 449 221
rect 415 125 449 153
rect 415 53 449 85
rect 415 -17 449 17
rect 415 -85 449 -53
rect 415 -153 449 -125
rect 415 -221 449 -197
rect 415 -289 449 -269
rect 415 -357 449 -341
rect 415 -425 449 -413
rect 415 -552 449 -485
rect 511 485 545 566
rect 511 413 545 425
rect 511 341 545 357
rect 511 269 545 289
rect 511 197 545 221
rect 511 125 545 153
rect 511 53 545 85
rect 511 -17 545 17
rect 511 -85 545 -53
rect 511 -153 545 -125
rect 511 -221 545 -197
rect 511 -289 545 -269
rect 511 -357 545 -341
rect 511 -425 545 -413
rect 511 -502 545 -485
rect -545 -586 449 -552
rect 301 -672 317 -638
rect 351 -672 367 -638
<< viali >>
rect -545 459 -511 485
rect -545 451 -511 459
rect -545 391 -511 413
rect -545 379 -511 391
rect -545 323 -511 341
rect -545 307 -511 323
rect -545 255 -511 269
rect -545 235 -511 255
rect -545 187 -511 197
rect -545 163 -511 187
rect -545 119 -511 125
rect -545 91 -511 119
rect -545 51 -511 53
rect -545 19 -511 51
rect -545 -51 -511 -19
rect -545 -53 -511 -51
rect -545 -119 -511 -91
rect -545 -125 -511 -119
rect -545 -187 -511 -163
rect -545 -197 -511 -187
rect -545 -255 -511 -235
rect -545 -269 -511 -255
rect -545 -323 -511 -307
rect -545 -341 -511 -323
rect -545 -391 -511 -379
rect -545 -413 -511 -391
rect -545 -459 -511 -451
rect -545 -485 -511 -459
rect -449 459 -415 485
rect -449 451 -415 459
rect -449 391 -415 413
rect -449 379 -415 391
rect -449 323 -415 341
rect -449 307 -415 323
rect -449 255 -415 269
rect -449 235 -415 255
rect -449 187 -415 197
rect -449 163 -415 187
rect -449 119 -415 125
rect -449 91 -415 119
rect -449 51 -415 53
rect -449 19 -415 51
rect -449 -51 -415 -19
rect -449 -53 -415 -51
rect -449 -119 -415 -91
rect -449 -125 -415 -119
rect -449 -187 -415 -163
rect -449 -197 -415 -187
rect -449 -255 -415 -235
rect -449 -269 -415 -255
rect -449 -323 -415 -307
rect -449 -341 -415 -323
rect -449 -391 -415 -379
rect -449 -413 -415 -391
rect -449 -459 -415 -451
rect -449 -485 -415 -459
rect -353 459 -319 485
rect -353 451 -319 459
rect -353 391 -319 413
rect -353 379 -319 391
rect -353 323 -319 341
rect -353 307 -319 323
rect -353 255 -319 269
rect -353 235 -319 255
rect -353 187 -319 197
rect -353 163 -319 187
rect -353 119 -319 125
rect -353 91 -319 119
rect -353 51 -319 53
rect -353 19 -319 51
rect -353 -51 -319 -19
rect -353 -53 -319 -51
rect -353 -119 -319 -91
rect -353 -125 -319 -119
rect -353 -187 -319 -163
rect -353 -197 -319 -187
rect -353 -255 -319 -235
rect -353 -269 -319 -255
rect -353 -323 -319 -307
rect -353 -341 -319 -323
rect -353 -391 -319 -379
rect -353 -413 -319 -391
rect -353 -459 -319 -451
rect -353 -485 -319 -459
rect -257 459 -223 485
rect -257 451 -223 459
rect -257 391 -223 413
rect -257 379 -223 391
rect -257 323 -223 341
rect -257 307 -223 323
rect -257 255 -223 269
rect -257 235 -223 255
rect -257 187 -223 197
rect -257 163 -223 187
rect -257 119 -223 125
rect -257 91 -223 119
rect -257 51 -223 53
rect -257 19 -223 51
rect -257 -51 -223 -19
rect -257 -53 -223 -51
rect -257 -119 -223 -91
rect -257 -125 -223 -119
rect -257 -187 -223 -163
rect -257 -197 -223 -187
rect -257 -255 -223 -235
rect -257 -269 -223 -255
rect -257 -323 -223 -307
rect -257 -341 -223 -323
rect -257 -391 -223 -379
rect -257 -413 -223 -391
rect -257 -459 -223 -451
rect -257 -485 -223 -459
rect -161 459 -127 485
rect -161 451 -127 459
rect -161 391 -127 413
rect -161 379 -127 391
rect -161 323 -127 341
rect -161 307 -127 323
rect -161 255 -127 269
rect -161 235 -127 255
rect -161 187 -127 197
rect -161 163 -127 187
rect -161 119 -127 125
rect -161 91 -127 119
rect -161 51 -127 53
rect -161 19 -127 51
rect -161 -51 -127 -19
rect -161 -53 -127 -51
rect -161 -119 -127 -91
rect -161 -125 -127 -119
rect -161 -187 -127 -163
rect -161 -197 -127 -187
rect -161 -255 -127 -235
rect -161 -269 -127 -255
rect -161 -323 -127 -307
rect -161 -341 -127 -323
rect -161 -391 -127 -379
rect -161 -413 -127 -391
rect -161 -459 -127 -451
rect -161 -485 -127 -459
rect -65 459 -31 485
rect -65 451 -31 459
rect -65 391 -31 413
rect -65 379 -31 391
rect -65 323 -31 341
rect -65 307 -31 323
rect -65 255 -31 269
rect -65 235 -31 255
rect -65 187 -31 197
rect -65 163 -31 187
rect -65 119 -31 125
rect -65 91 -31 119
rect -65 51 -31 53
rect -65 19 -31 51
rect -65 -51 -31 -19
rect -65 -53 -31 -51
rect -65 -119 -31 -91
rect -65 -125 -31 -119
rect -65 -187 -31 -163
rect -65 -197 -31 -187
rect -65 -255 -31 -235
rect -65 -269 -31 -255
rect -65 -323 -31 -307
rect -65 -341 -31 -323
rect -65 -391 -31 -379
rect -65 -413 -31 -391
rect -65 -459 -31 -451
rect -65 -485 -31 -459
rect 31 459 65 485
rect 31 451 65 459
rect 31 391 65 413
rect 31 379 65 391
rect 31 323 65 341
rect 31 307 65 323
rect 31 255 65 269
rect 31 235 65 255
rect 31 187 65 197
rect 31 163 65 187
rect 31 119 65 125
rect 31 91 65 119
rect 31 51 65 53
rect 31 19 65 51
rect 31 -51 65 -19
rect 31 -53 65 -51
rect 31 -119 65 -91
rect 31 -125 65 -119
rect 31 -187 65 -163
rect 31 -197 65 -187
rect 31 -255 65 -235
rect 31 -269 65 -255
rect 31 -323 65 -307
rect 31 -341 65 -323
rect 31 -391 65 -379
rect 31 -413 65 -391
rect 31 -459 65 -451
rect 31 -485 65 -459
rect 127 459 161 485
rect 127 451 161 459
rect 127 391 161 413
rect 127 379 161 391
rect 127 323 161 341
rect 127 307 161 323
rect 127 255 161 269
rect 127 235 161 255
rect 127 187 161 197
rect 127 163 161 187
rect 127 119 161 125
rect 127 91 161 119
rect 127 51 161 53
rect 127 19 161 51
rect 127 -51 161 -19
rect 127 -53 161 -51
rect 127 -119 161 -91
rect 127 -125 161 -119
rect 127 -187 161 -163
rect 127 -197 161 -187
rect 127 -255 161 -235
rect 127 -269 161 -255
rect 127 -323 161 -307
rect 127 -341 161 -323
rect 127 -391 161 -379
rect 127 -413 161 -391
rect 127 -459 161 -451
rect 127 -485 161 -459
rect 223 459 257 485
rect 223 451 257 459
rect 223 391 257 413
rect 223 379 257 391
rect 223 323 257 341
rect 223 307 257 323
rect 223 255 257 269
rect 223 235 257 255
rect 223 187 257 197
rect 223 163 257 187
rect 223 119 257 125
rect 223 91 257 119
rect 223 51 257 53
rect 223 19 257 51
rect 223 -51 257 -19
rect 223 -53 257 -51
rect 223 -119 257 -91
rect 223 -125 257 -119
rect 223 -187 257 -163
rect 223 -197 257 -187
rect 223 -255 257 -235
rect 223 -269 257 -255
rect 223 -323 257 -307
rect 223 -341 257 -323
rect 223 -391 257 -379
rect 223 -413 257 -391
rect 223 -459 257 -451
rect 223 -485 257 -459
rect 319 459 353 485
rect 319 451 353 459
rect 319 391 353 413
rect 319 379 353 391
rect 319 323 353 341
rect 319 307 353 323
rect 319 255 353 269
rect 319 235 353 255
rect 319 187 353 197
rect 319 163 353 187
rect 319 119 353 125
rect 319 91 353 119
rect 319 51 353 53
rect 319 19 353 51
rect 319 -51 353 -19
rect 319 -53 353 -51
rect 319 -119 353 -91
rect 319 -125 353 -119
rect 319 -187 353 -163
rect 319 -197 353 -187
rect 319 -255 353 -235
rect 319 -269 353 -255
rect 319 -323 353 -307
rect 319 -341 353 -323
rect 319 -391 353 -379
rect 319 -413 353 -391
rect 319 -459 353 -451
rect 319 -485 353 -459
rect 415 459 449 485
rect 415 451 449 459
rect 415 391 449 413
rect 415 379 449 391
rect 415 323 449 341
rect 415 307 449 323
rect 415 255 449 269
rect 415 235 449 255
rect 415 187 449 197
rect 415 163 449 187
rect 415 119 449 125
rect 415 91 449 119
rect 415 51 449 53
rect 415 19 449 51
rect 415 -51 449 -19
rect 415 -53 449 -51
rect 415 -119 449 -91
rect 415 -125 449 -119
rect 415 -187 449 -163
rect 415 -197 449 -187
rect 415 -255 449 -235
rect 415 -269 449 -255
rect 415 -323 449 -307
rect 415 -341 449 -323
rect 415 -391 449 -379
rect 415 -413 449 -391
rect 415 -459 449 -451
rect 415 -485 449 -459
rect 511 459 545 485
rect 511 451 545 459
rect 511 391 545 413
rect 511 379 545 391
rect 511 323 545 341
rect 511 307 545 323
rect 511 255 545 269
rect 511 235 545 255
rect 511 187 545 197
rect 511 163 545 187
rect 511 119 545 125
rect 511 91 545 119
rect 511 51 545 53
rect 511 19 545 51
rect 511 -51 545 -19
rect 511 -53 545 -51
rect 511 -119 545 -91
rect 511 -125 545 -119
rect 511 -187 545 -163
rect 511 -197 545 -187
rect 511 -255 545 -235
rect 511 -269 545 -255
rect 511 -323 545 -307
rect 511 -341 545 -323
rect 511 -391 545 -379
rect 511 -413 545 -391
rect 511 -459 545 -451
rect 511 -485 545 -459
rect 317 -672 351 -638
<< metal1 >>
rect -551 485 -505 500
rect -551 451 -545 485
rect -511 451 -505 485
rect -551 413 -505 451
rect -551 379 -545 413
rect -511 379 -505 413
rect -551 341 -505 379
rect -551 307 -545 341
rect -511 307 -505 341
rect -551 269 -505 307
rect -551 235 -545 269
rect -511 235 -505 269
rect -551 197 -505 235
rect -551 163 -545 197
rect -511 163 -505 197
rect -551 125 -505 163
rect -551 91 -545 125
rect -511 91 -505 125
rect -551 53 -505 91
rect -551 19 -545 53
rect -511 19 -505 53
rect -551 -19 -505 19
rect -551 -53 -545 -19
rect -511 -53 -505 -19
rect -551 -91 -505 -53
rect -551 -125 -545 -91
rect -511 -125 -505 -91
rect -551 -163 -505 -125
rect -551 -197 -545 -163
rect -511 -197 -505 -163
rect -551 -235 -505 -197
rect -551 -269 -545 -235
rect -511 -269 -505 -235
rect -551 -307 -505 -269
rect -551 -341 -545 -307
rect -511 -341 -505 -307
rect -551 -379 -505 -341
rect -551 -413 -545 -379
rect -511 -413 -505 -379
rect -551 -451 -505 -413
rect -551 -485 -545 -451
rect -511 -485 -505 -451
rect -551 -500 -505 -485
rect -455 485 -409 500
rect -455 451 -449 485
rect -415 451 -409 485
rect -455 413 -409 451
rect -455 379 -449 413
rect -415 379 -409 413
rect -455 341 -409 379
rect -455 307 -449 341
rect -415 307 -409 341
rect -455 269 -409 307
rect -455 235 -449 269
rect -415 235 -409 269
rect -455 197 -409 235
rect -455 163 -449 197
rect -415 163 -409 197
rect -455 125 -409 163
rect -455 91 -449 125
rect -415 91 -409 125
rect -455 53 -409 91
rect -455 19 -449 53
rect -415 19 -409 53
rect -455 -19 -409 19
rect -455 -53 -449 -19
rect -415 -53 -409 -19
rect -455 -91 -409 -53
rect -455 -125 -449 -91
rect -415 -125 -409 -91
rect -455 -163 -409 -125
rect -455 -197 -449 -163
rect -415 -197 -409 -163
rect -455 -235 -409 -197
rect -455 -269 -449 -235
rect -415 -269 -409 -235
rect -455 -307 -409 -269
rect -455 -341 -449 -307
rect -415 -341 -409 -307
rect -455 -379 -409 -341
rect -455 -413 -449 -379
rect -415 -413 -409 -379
rect -455 -451 -409 -413
rect -455 -485 -449 -451
rect -415 -485 -409 -451
rect -455 -500 -409 -485
rect -359 485 -313 500
rect -359 451 -353 485
rect -319 451 -313 485
rect -359 413 -313 451
rect -359 379 -353 413
rect -319 379 -313 413
rect -359 341 -313 379
rect -359 307 -353 341
rect -319 307 -313 341
rect -359 269 -313 307
rect -359 235 -353 269
rect -319 235 -313 269
rect -359 197 -313 235
rect -359 163 -353 197
rect -319 163 -313 197
rect -359 125 -313 163
rect -359 91 -353 125
rect -319 91 -313 125
rect -359 53 -313 91
rect -359 19 -353 53
rect -319 19 -313 53
rect -359 -19 -313 19
rect -359 -53 -353 -19
rect -319 -53 -313 -19
rect -359 -91 -313 -53
rect -359 -125 -353 -91
rect -319 -125 -313 -91
rect -359 -163 -313 -125
rect -359 -197 -353 -163
rect -319 -197 -313 -163
rect -359 -235 -313 -197
rect -359 -269 -353 -235
rect -319 -269 -313 -235
rect -359 -307 -313 -269
rect -359 -341 -353 -307
rect -319 -341 -313 -307
rect -359 -379 -313 -341
rect -359 -413 -353 -379
rect -319 -413 -313 -379
rect -359 -451 -313 -413
rect -359 -485 -353 -451
rect -319 -485 -313 -451
rect -359 -500 -313 -485
rect -263 485 -217 500
rect -263 451 -257 485
rect -223 451 -217 485
rect -263 413 -217 451
rect -263 379 -257 413
rect -223 379 -217 413
rect -263 341 -217 379
rect -263 307 -257 341
rect -223 307 -217 341
rect -263 269 -217 307
rect -263 235 -257 269
rect -223 235 -217 269
rect -263 197 -217 235
rect -263 163 -257 197
rect -223 163 -217 197
rect -263 125 -217 163
rect -263 91 -257 125
rect -223 91 -217 125
rect -263 53 -217 91
rect -263 19 -257 53
rect -223 19 -217 53
rect -263 -19 -217 19
rect -263 -53 -257 -19
rect -223 -53 -217 -19
rect -263 -91 -217 -53
rect -263 -125 -257 -91
rect -223 -125 -217 -91
rect -263 -163 -217 -125
rect -263 -197 -257 -163
rect -223 -197 -217 -163
rect -263 -235 -217 -197
rect -263 -269 -257 -235
rect -223 -269 -217 -235
rect -263 -307 -217 -269
rect -263 -341 -257 -307
rect -223 -341 -217 -307
rect -263 -379 -217 -341
rect -263 -413 -257 -379
rect -223 -413 -217 -379
rect -263 -451 -217 -413
rect -263 -485 -257 -451
rect -223 -485 -217 -451
rect -263 -500 -217 -485
rect -167 485 -121 500
rect -167 451 -161 485
rect -127 451 -121 485
rect -167 413 -121 451
rect -167 379 -161 413
rect -127 379 -121 413
rect -167 341 -121 379
rect -167 307 -161 341
rect -127 307 -121 341
rect -167 269 -121 307
rect -167 235 -161 269
rect -127 235 -121 269
rect -167 197 -121 235
rect -167 163 -161 197
rect -127 163 -121 197
rect -167 125 -121 163
rect -167 91 -161 125
rect -127 91 -121 125
rect -167 53 -121 91
rect -167 19 -161 53
rect -127 19 -121 53
rect -167 -19 -121 19
rect -167 -53 -161 -19
rect -127 -53 -121 -19
rect -167 -91 -121 -53
rect -167 -125 -161 -91
rect -127 -125 -121 -91
rect -167 -163 -121 -125
rect -167 -197 -161 -163
rect -127 -197 -121 -163
rect -167 -235 -121 -197
rect -167 -269 -161 -235
rect -127 -269 -121 -235
rect -167 -307 -121 -269
rect -167 -341 -161 -307
rect -127 -341 -121 -307
rect -167 -379 -121 -341
rect -167 -413 -161 -379
rect -127 -413 -121 -379
rect -167 -451 -121 -413
rect -167 -485 -161 -451
rect -127 -485 -121 -451
rect -167 -500 -121 -485
rect -71 485 -25 500
rect -71 451 -65 485
rect -31 451 -25 485
rect -71 413 -25 451
rect -71 379 -65 413
rect -31 379 -25 413
rect -71 341 -25 379
rect -71 307 -65 341
rect -31 307 -25 341
rect -71 269 -25 307
rect -71 235 -65 269
rect -31 235 -25 269
rect -71 197 -25 235
rect -71 163 -65 197
rect -31 163 -25 197
rect -71 125 -25 163
rect -71 91 -65 125
rect -31 91 -25 125
rect -71 53 -25 91
rect -71 19 -65 53
rect -31 19 -25 53
rect -71 -19 -25 19
rect -71 -53 -65 -19
rect -31 -53 -25 -19
rect -71 -91 -25 -53
rect -71 -125 -65 -91
rect -31 -125 -25 -91
rect -71 -163 -25 -125
rect -71 -197 -65 -163
rect -31 -197 -25 -163
rect -71 -235 -25 -197
rect -71 -269 -65 -235
rect -31 -269 -25 -235
rect -71 -307 -25 -269
rect -71 -341 -65 -307
rect -31 -341 -25 -307
rect -71 -379 -25 -341
rect -71 -413 -65 -379
rect -31 -413 -25 -379
rect -71 -451 -25 -413
rect -71 -485 -65 -451
rect -31 -485 -25 -451
rect -71 -500 -25 -485
rect 25 485 71 500
rect 25 451 31 485
rect 65 451 71 485
rect 25 413 71 451
rect 25 379 31 413
rect 65 379 71 413
rect 25 341 71 379
rect 25 307 31 341
rect 65 307 71 341
rect 25 269 71 307
rect 25 235 31 269
rect 65 235 71 269
rect 25 197 71 235
rect 25 163 31 197
rect 65 163 71 197
rect 25 125 71 163
rect 25 91 31 125
rect 65 91 71 125
rect 25 53 71 91
rect 25 19 31 53
rect 65 19 71 53
rect 25 -19 71 19
rect 25 -53 31 -19
rect 65 -53 71 -19
rect 25 -91 71 -53
rect 25 -125 31 -91
rect 65 -125 71 -91
rect 25 -163 71 -125
rect 25 -197 31 -163
rect 65 -197 71 -163
rect 25 -235 71 -197
rect 25 -269 31 -235
rect 65 -269 71 -235
rect 25 -307 71 -269
rect 25 -341 31 -307
rect 65 -341 71 -307
rect 25 -379 71 -341
rect 25 -413 31 -379
rect 65 -413 71 -379
rect 25 -451 71 -413
rect 25 -485 31 -451
rect 65 -485 71 -451
rect 25 -500 71 -485
rect 121 485 167 500
rect 121 451 127 485
rect 161 451 167 485
rect 121 413 167 451
rect 121 379 127 413
rect 161 379 167 413
rect 121 341 167 379
rect 121 307 127 341
rect 161 307 167 341
rect 121 269 167 307
rect 121 235 127 269
rect 161 235 167 269
rect 121 197 167 235
rect 121 163 127 197
rect 161 163 167 197
rect 121 125 167 163
rect 121 91 127 125
rect 161 91 167 125
rect 121 53 167 91
rect 121 19 127 53
rect 161 19 167 53
rect 121 -19 167 19
rect 121 -53 127 -19
rect 161 -53 167 -19
rect 121 -91 167 -53
rect 121 -125 127 -91
rect 161 -125 167 -91
rect 121 -163 167 -125
rect 121 -197 127 -163
rect 161 -197 167 -163
rect 121 -235 167 -197
rect 121 -269 127 -235
rect 161 -269 167 -235
rect 121 -307 167 -269
rect 121 -341 127 -307
rect 161 -341 167 -307
rect 121 -379 167 -341
rect 121 -413 127 -379
rect 161 -413 167 -379
rect 121 -451 167 -413
rect 121 -485 127 -451
rect 161 -485 167 -451
rect 121 -500 167 -485
rect 217 485 263 500
rect 217 451 223 485
rect 257 451 263 485
rect 217 413 263 451
rect 217 379 223 413
rect 257 379 263 413
rect 217 341 263 379
rect 217 307 223 341
rect 257 307 263 341
rect 217 269 263 307
rect 217 235 223 269
rect 257 235 263 269
rect 217 197 263 235
rect 217 163 223 197
rect 257 163 263 197
rect 217 125 263 163
rect 217 91 223 125
rect 257 91 263 125
rect 217 53 263 91
rect 217 19 223 53
rect 257 19 263 53
rect 217 -19 263 19
rect 217 -53 223 -19
rect 257 -53 263 -19
rect 217 -91 263 -53
rect 217 -125 223 -91
rect 257 -125 263 -91
rect 217 -163 263 -125
rect 217 -197 223 -163
rect 257 -197 263 -163
rect 217 -235 263 -197
rect 217 -269 223 -235
rect 257 -269 263 -235
rect 217 -307 263 -269
rect 217 -341 223 -307
rect 257 -341 263 -307
rect 217 -379 263 -341
rect 217 -413 223 -379
rect 257 -413 263 -379
rect 217 -451 263 -413
rect 217 -485 223 -451
rect 257 -485 263 -451
rect 217 -500 263 -485
rect 313 485 359 500
rect 313 451 319 485
rect 353 451 359 485
rect 313 413 359 451
rect 313 379 319 413
rect 353 379 359 413
rect 313 341 359 379
rect 313 307 319 341
rect 353 307 359 341
rect 313 269 359 307
rect 313 235 319 269
rect 353 235 359 269
rect 313 197 359 235
rect 313 163 319 197
rect 353 163 359 197
rect 313 125 359 163
rect 313 91 319 125
rect 353 91 359 125
rect 313 53 359 91
rect 313 19 319 53
rect 353 19 359 53
rect 313 -19 359 19
rect 313 -53 319 -19
rect 353 -53 359 -19
rect 313 -91 359 -53
rect 313 -125 319 -91
rect 353 -125 359 -91
rect 313 -163 359 -125
rect 313 -197 319 -163
rect 353 -197 359 -163
rect 313 -235 359 -197
rect 313 -269 319 -235
rect 353 -269 359 -235
rect 313 -307 359 -269
rect 313 -341 319 -307
rect 353 -341 359 -307
rect 313 -379 359 -341
rect 313 -413 319 -379
rect 353 -413 359 -379
rect 313 -451 359 -413
rect 313 -485 319 -451
rect 353 -485 359 -451
rect 313 -500 359 -485
rect 409 485 455 500
rect 409 451 415 485
rect 449 451 455 485
rect 409 413 455 451
rect 409 379 415 413
rect 449 379 455 413
rect 409 341 455 379
rect 409 307 415 341
rect 449 307 455 341
rect 409 269 455 307
rect 409 235 415 269
rect 449 235 455 269
rect 409 197 455 235
rect 409 163 415 197
rect 449 163 455 197
rect 409 125 455 163
rect 409 91 415 125
rect 449 91 455 125
rect 409 53 455 91
rect 409 19 415 53
rect 449 19 455 53
rect 409 -19 455 19
rect 409 -53 415 -19
rect 449 -53 455 -19
rect 409 -91 455 -53
rect 409 -125 415 -91
rect 449 -125 455 -91
rect 409 -163 455 -125
rect 409 -197 415 -163
rect 449 -197 455 -163
rect 409 -235 455 -197
rect 409 -269 415 -235
rect 449 -269 455 -235
rect 409 -307 455 -269
rect 409 -341 415 -307
rect 449 -341 455 -307
rect 409 -379 455 -341
rect 409 -413 415 -379
rect 449 -413 455 -379
rect 409 -451 455 -413
rect 409 -485 415 -451
rect 449 -485 455 -451
rect 409 -500 455 -485
rect 505 485 551 500
rect 505 451 511 485
rect 545 451 551 485
rect 505 413 551 451
rect 505 379 511 413
rect 545 379 551 413
rect 505 341 551 379
rect 505 307 511 341
rect 545 307 551 341
rect 505 269 551 307
rect 505 235 511 269
rect 545 235 551 269
rect 505 197 551 235
rect 505 163 511 197
rect 545 163 551 197
rect 505 125 551 163
rect 505 91 511 125
rect 545 91 551 125
rect 505 53 551 91
rect 505 19 511 53
rect 545 19 551 53
rect 505 -19 551 19
rect 505 -53 511 -19
rect 545 -53 551 -19
rect 505 -91 551 -53
rect 505 -125 511 -91
rect 545 -125 551 -91
rect 505 -163 551 -125
rect 505 -197 511 -163
rect 545 -197 551 -163
rect 505 -235 551 -197
rect 505 -269 511 -235
rect 545 -269 551 -235
rect 505 -307 551 -269
rect 505 -341 511 -307
rect 545 -341 551 -307
rect 505 -379 551 -341
rect 505 -413 511 -379
rect 545 -413 551 -379
rect 505 -451 551 -413
rect 505 -485 511 -451
rect 545 -485 551 -451
rect 505 -500 551 -485
rect 305 -638 363 -632
rect 305 -672 317 -638
rect 351 -672 363 -638
rect 305 -678 363 -672
<< end >>
