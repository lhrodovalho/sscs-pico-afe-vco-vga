magic
tech sky130A
timestamp 1638390070
<< nwell >>
rect 60 1380 4140 1940
rect 60 660 4140 1220
<< nmos >>
rect 260 80 1060 180
rect 1220 80 2020 180
rect 2180 80 2980 180
rect 3140 80 3940 180
<< pmoslvt >>
rect 260 1540 1060 1840
rect 1220 1540 2020 1840
rect 2180 1540 2980 1840
rect 3140 1540 3940 1840
rect 260 820 1060 1120
rect 1220 820 2020 1120
rect 2180 820 2980 1120
rect 3140 820 3940 1120
<< ndiff >>
rect 160 170 260 180
rect 160 90 165 170
rect 195 90 260 170
rect 160 80 260 90
rect 1060 170 1220 180
rect 1060 90 1125 170
rect 1155 90 1220 170
rect 1060 80 1220 90
rect 2020 170 2180 180
rect 2020 90 2085 170
rect 2115 90 2180 170
rect 2020 80 2180 90
rect 2980 170 3140 180
rect 2980 90 3045 170
rect 3075 90 3140 170
rect 2980 80 3140 90
rect 3940 170 4040 180
rect 3940 90 4005 170
rect 4035 90 4040 170
rect 3940 80 4040 90
<< pdiff >>
rect 160 1830 260 1840
rect 160 1550 165 1830
rect 195 1550 260 1830
rect 160 1540 260 1550
rect 1060 1830 1220 1840
rect 1060 1550 1125 1830
rect 1155 1550 1220 1830
rect 1060 1540 1220 1550
rect 2020 1830 2180 1840
rect 2020 1550 2085 1830
rect 2115 1550 2180 1830
rect 2020 1540 2180 1550
rect 2980 1830 3140 1840
rect 2980 1550 3045 1830
rect 3075 1550 3140 1830
rect 2980 1540 3140 1550
rect 3940 1830 4040 1840
rect 3940 1550 4005 1830
rect 4035 1550 4040 1830
rect 3940 1540 4040 1550
rect 160 1110 260 1120
rect 160 830 165 1110
rect 195 830 260 1110
rect 160 820 260 830
rect 1060 1110 1220 1120
rect 1060 830 1125 1110
rect 1155 830 1220 1110
rect 1060 820 1220 830
rect 2020 1110 2180 1120
rect 2020 830 2085 1110
rect 2115 830 2180 1110
rect 2020 820 2180 830
rect 2980 1110 3140 1120
rect 2980 830 3045 1110
rect 3075 830 3140 1110
rect 2980 820 3140 830
rect 3940 1110 4040 1120
rect 3940 830 4005 1110
rect 4035 830 4040 1110
rect 3940 820 4040 830
<< ndiffc >>
rect 165 90 195 170
rect 1125 90 1155 170
rect 2085 90 2115 170
rect 3045 90 3075 170
rect 4005 90 4035 170
<< pdiffc >>
rect 165 1550 195 1830
rect 1125 1550 1155 1830
rect 2085 1550 2115 1830
rect 3045 1550 3075 1830
rect 4005 1550 4035 1830
rect 165 830 195 1110
rect 1125 830 1155 1110
rect 2085 830 2115 1110
rect 3045 830 3075 1110
rect 4005 830 4035 1110
<< psubdiff >>
rect 0 1960 60 2000
rect 4140 1960 4200 2000
rect 0 1940 40 1960
rect 4160 1940 4200 1960
rect 0 1360 40 1380
rect 4160 1360 4200 1380
rect 0 1320 60 1360
rect 4120 1320 4200 1360
rect 0 1240 60 1280
rect 4120 1240 4200 1280
rect 0 1220 40 1240
rect 4160 1220 4200 1240
rect 0 640 40 660
rect 4160 640 4200 660
rect 0 600 60 640
rect 4140 600 4200 640
rect 0 280 60 320
rect 4140 280 4200 320
rect 0 260 40 280
rect 4160 260 4200 280
rect 0 40 40 60
rect 4160 40 4200 60
rect 0 0 60 40
rect 4140 0 4200 40
<< nsubdiff >>
rect 80 1880 140 1920
rect 4060 1880 4120 1920
rect 80 1860 120 1880
rect 4080 1860 4120 1880
rect 80 1440 120 1460
rect 4080 1440 4120 1460
rect 80 1400 140 1440
rect 4060 1400 4120 1440
rect 80 1160 140 1200
rect 4060 1160 4120 1200
rect 80 1140 120 1160
rect 4080 1140 4120 1160
rect 80 720 120 740
rect 4080 720 4120 740
rect 80 680 140 720
rect 4060 680 4120 720
<< psubdiffcont >>
rect 60 1960 4140 2000
rect 0 1380 40 1940
rect 4160 1380 4200 1940
rect 60 1320 4120 1360
rect 60 1240 4120 1280
rect 0 660 40 1220
rect 4160 660 4200 1220
rect 60 600 4140 640
rect 60 280 4140 320
rect 0 60 40 260
rect 4160 60 4200 260
rect 60 0 4140 40
<< nsubdiffcont >>
rect 140 1880 4060 1920
rect 80 1460 120 1860
rect 4080 1460 4120 1860
rect 140 1400 4060 1440
rect 140 1160 4060 1200
rect 80 740 120 1140
rect 4080 740 4120 1140
rect 140 680 4060 720
<< poly >>
rect 260 1840 1060 1860
rect 1220 1840 2020 1860
rect 2180 1840 2980 1860
rect 3140 1840 3940 1860
rect 260 1515 1060 1540
rect 260 1485 270 1515
rect 1050 1485 1060 1515
rect 260 1480 1060 1485
rect 1220 1515 2020 1540
rect 1220 1485 1230 1515
rect 2010 1485 2020 1515
rect 1220 1480 2020 1485
rect 2180 1515 2980 1540
rect 2180 1485 2190 1515
rect 2970 1485 2980 1515
rect 2180 1480 2980 1485
rect 3140 1515 3940 1540
rect 3140 1485 3150 1515
rect 3930 1485 3940 1515
rect 3140 1480 3940 1485
rect 260 1120 1060 1140
rect 1220 1120 2020 1140
rect 2180 1120 2980 1140
rect 3140 1120 3940 1140
rect 260 795 1060 820
rect 260 765 270 795
rect 1050 765 1060 795
rect 260 760 1060 765
rect 1220 795 2020 820
rect 1220 765 1230 795
rect 2010 765 2020 795
rect 1220 760 2020 765
rect 2180 795 2980 820
rect 2180 765 2190 795
rect 2970 765 2980 795
rect 2180 760 2980 765
rect 3140 795 3940 820
rect 3140 765 3150 795
rect 3930 765 3940 795
rect 3140 760 3940 765
rect 260 235 1060 240
rect 260 205 270 235
rect 1050 205 1060 235
rect 260 180 1060 205
rect 1220 235 2020 240
rect 1220 205 1230 235
rect 2010 205 2020 235
rect 1220 180 2020 205
rect 2180 235 2980 240
rect 2180 205 2190 235
rect 2970 205 2980 235
rect 2180 180 2980 205
rect 3140 235 3940 240
rect 3140 205 3150 235
rect 3930 205 3940 235
rect 3140 180 3940 205
rect 260 60 1060 80
rect 1220 60 2020 80
rect 2180 60 2980 80
rect 3140 60 3940 80
<< polycont >>
rect 270 1485 1050 1515
rect 1230 1485 2010 1515
rect 2190 1485 2970 1515
rect 3150 1485 3930 1515
rect 270 765 1050 795
rect 1230 765 2010 795
rect 2190 765 2970 795
rect 3150 765 3930 795
rect 270 205 1050 235
rect 1230 205 2010 235
rect 2190 205 2970 235
rect 3150 205 3930 235
<< locali >>
rect 0 1960 60 2000
rect 4140 1960 4200 2000
rect 0 1940 40 1960
rect 4160 1940 4200 1960
rect 80 1880 140 1920
rect 4060 1880 4120 1920
rect 80 1860 120 1880
rect 160 1830 200 1840
rect 160 1550 165 1830
rect 195 1550 200 1830
rect 160 1540 200 1550
rect 1120 1830 1160 1840
rect 1120 1550 1125 1830
rect 1155 1550 1160 1830
rect 1120 1540 1160 1550
rect 2080 1830 2120 1880
rect 4080 1860 4120 1880
rect 2080 1550 2085 1830
rect 2115 1550 2120 1830
rect 2080 1540 2120 1550
rect 3040 1830 3080 1840
rect 3040 1550 3045 1830
rect 3075 1550 3080 1830
rect 3040 1540 3080 1550
rect 4000 1830 4040 1840
rect 4000 1550 4005 1830
rect 4035 1550 4040 1830
rect 4000 1540 4040 1550
rect 260 1515 1060 1520
rect 260 1485 270 1515
rect 1050 1485 1060 1515
rect 260 1480 1060 1485
rect 1220 1515 2020 1520
rect 1220 1485 1230 1515
rect 2010 1485 2020 1515
rect 1220 1480 2020 1485
rect 2180 1515 2980 1520
rect 2180 1485 2190 1515
rect 2970 1485 2980 1515
rect 2180 1480 2980 1485
rect 3140 1515 3940 1520
rect 3140 1485 3150 1515
rect 3930 1485 3940 1515
rect 3140 1480 3940 1485
rect 80 1440 120 1460
rect 4080 1440 4120 1460
rect 80 1400 140 1440
rect 4060 1400 4120 1440
rect 0 1360 40 1380
rect 4160 1360 4200 1380
rect 0 1320 60 1360
rect 4120 1320 4200 1360
rect 0 1280 40 1320
rect 4160 1280 4200 1320
rect 0 1240 60 1280
rect 4120 1240 4200 1280
rect 0 1220 40 1240
rect 4160 1220 4200 1240
rect 80 1160 140 1200
rect 4060 1160 4120 1200
rect 80 1140 120 1160
rect 160 1110 200 1160
rect 160 830 165 1110
rect 195 830 200 1110
rect 160 820 200 830
rect 1120 1110 1160 1120
rect 1120 830 1125 1110
rect 1155 830 1160 1110
rect 1120 820 1160 830
rect 2080 1110 2120 1120
rect 2080 830 2085 1110
rect 2115 830 2120 1110
rect 2080 820 2120 830
rect 3040 1110 3080 1120
rect 3040 830 3045 1110
rect 3075 830 3080 1110
rect 3040 820 3080 830
rect 4000 1110 4040 1160
rect 4000 830 4005 1110
rect 4035 830 4040 1110
rect 4000 820 4040 830
rect 4080 1140 4120 1160
rect 260 795 1060 800
rect 260 765 270 795
rect 1050 765 1060 795
rect 260 760 1060 765
rect 1220 795 2020 800
rect 1220 765 1230 795
rect 2010 765 2020 795
rect 1220 760 2020 765
rect 2180 795 2980 800
rect 2180 765 2190 795
rect 2970 765 2980 795
rect 2180 760 2980 765
rect 3140 795 3940 800
rect 3140 765 3150 795
rect 3930 765 3940 795
rect 3140 760 3940 765
rect 80 720 120 740
rect 4080 720 4120 740
rect 80 680 140 720
rect 4060 680 4120 720
rect 0 640 40 660
rect 4160 640 4200 660
rect 0 600 60 640
rect 4140 600 4200 640
rect 0 320 40 600
rect 80 470 4120 560
rect 80 450 90 470
rect 110 450 170 470
rect 190 450 250 470
rect 270 450 330 470
rect 350 450 410 470
rect 430 450 490 470
rect 510 450 570 470
rect 590 450 730 470
rect 750 450 810 470
rect 830 450 890 470
rect 910 450 970 470
rect 990 450 1050 470
rect 1070 450 1130 470
rect 1150 450 1210 470
rect 1230 450 1290 470
rect 1310 450 1370 470
rect 1390 450 1450 470
rect 1470 450 1530 470
rect 1550 450 1690 470
rect 1710 450 1770 470
rect 1790 450 1850 470
rect 1870 450 1930 470
rect 1950 450 2010 470
rect 2030 450 2170 470
rect 2190 450 2250 470
rect 2270 450 2330 470
rect 2350 450 2410 470
rect 2430 450 2490 470
rect 2510 450 2650 470
rect 2670 450 2730 470
rect 2750 450 2810 470
rect 2830 450 2890 470
rect 2910 450 2970 470
rect 2990 450 3050 470
rect 3070 450 3130 470
rect 3150 450 3210 470
rect 3230 450 3290 470
rect 3310 450 3370 470
rect 3390 450 3450 470
rect 3470 450 3610 470
rect 3630 450 3690 470
rect 3710 450 3770 470
rect 3790 450 3850 470
rect 3870 450 3930 470
rect 3950 450 4010 470
rect 4030 450 4090 470
rect 4110 450 4120 470
rect 80 360 4120 450
rect 4160 320 4200 600
rect 0 280 60 320
rect 4140 280 4200 320
rect 0 260 40 280
rect 4160 260 4200 280
rect 260 235 1060 240
rect 260 205 270 235
rect 1050 205 1060 235
rect 260 200 1060 205
rect 1220 235 2020 240
rect 1220 205 1230 235
rect 2010 205 2020 235
rect 1220 200 2020 205
rect 2180 235 2980 240
rect 2180 205 2190 235
rect 2970 205 2980 235
rect 2180 200 2980 205
rect 3140 235 3940 240
rect 3140 205 3150 235
rect 3930 205 3940 235
rect 3140 200 3940 205
rect 0 40 40 60
rect 160 170 200 180
rect 160 90 165 170
rect 195 90 200 170
rect 160 40 200 90
rect 1120 170 1160 180
rect 1120 90 1125 170
rect 1155 90 1160 170
rect 1120 80 1160 90
rect 2080 170 2120 180
rect 2080 90 2085 170
rect 2115 90 2120 170
rect 2080 80 2120 90
rect 3040 170 3080 180
rect 3040 90 3045 170
rect 3075 90 3080 170
rect 3040 80 3080 90
rect 4000 170 4040 180
rect 4000 90 4005 170
rect 4035 90 4040 170
rect 4000 40 4040 90
rect 4160 40 4200 60
rect 0 0 60 40
rect 4140 0 4200 40
<< viali >>
rect 165 1550 195 1830
rect 1125 1550 1155 1830
rect 2085 1550 2115 1830
rect 3045 1550 3075 1830
rect 4005 1550 4035 1830
rect 270 1485 1050 1515
rect 1230 1485 2010 1515
rect 2190 1485 2970 1515
rect 3150 1485 3930 1515
rect 165 830 195 1110
rect 1125 830 1155 1110
rect 2085 830 2115 1110
rect 3045 830 3075 1110
rect 4005 830 4035 1110
rect 270 765 1050 795
rect 1230 765 2010 795
rect 2190 765 2970 795
rect 3150 765 3930 795
rect 90 450 110 470
rect 170 450 190 470
rect 250 450 270 470
rect 330 450 350 470
rect 410 450 430 470
rect 490 450 510 470
rect 570 450 590 470
rect 730 450 750 470
rect 810 450 830 470
rect 890 450 910 470
rect 970 450 990 470
rect 1050 450 1070 470
rect 1130 450 1150 470
rect 1210 450 1230 470
rect 1290 450 1310 470
rect 1370 450 1390 470
rect 1450 450 1470 470
rect 1530 450 1550 470
rect 1690 450 1710 470
rect 1770 450 1790 470
rect 1850 450 1870 470
rect 1930 450 1950 470
rect 2010 450 2030 470
rect 2170 450 2190 470
rect 2250 450 2270 470
rect 2330 450 2350 470
rect 2410 450 2430 470
rect 2490 450 2510 470
rect 2650 450 2670 470
rect 2730 450 2750 470
rect 2810 450 2830 470
rect 2890 450 2910 470
rect 2970 450 2990 470
rect 3050 450 3070 470
rect 3130 450 3150 470
rect 3210 450 3230 470
rect 3290 450 3310 470
rect 3370 450 3390 470
rect 3450 450 3470 470
rect 3610 450 3630 470
rect 3690 450 3710 470
rect 3770 450 3790 470
rect 3850 450 3870 470
rect 3930 450 3950 470
rect 4010 450 4030 470
rect 4090 450 4110 470
rect 270 205 1050 235
rect 1230 205 2010 235
rect 2190 205 2970 235
rect 3150 205 3930 235
rect 165 90 195 170
rect 1125 90 1155 170
rect 2085 90 2115 170
rect 3045 90 3075 170
rect 4005 90 4035 170
<< metal1 >>
rect 160 1830 200 1840
rect 160 1550 165 1830
rect 195 1550 200 1830
rect 0 1395 40 1400
rect 0 1365 5 1395
rect 35 1365 40 1395
rect 0 1235 40 1365
rect 0 1205 5 1235
rect 35 1205 40 1235
rect 0 1200 40 1205
rect 80 1395 120 1400
rect 80 1365 85 1395
rect 115 1365 120 1395
rect 80 1235 120 1365
rect 80 1205 85 1235
rect 115 1205 120 1235
rect 80 1200 120 1205
rect 160 1395 200 1550
rect 1120 1830 1160 1840
rect 1120 1550 1125 1830
rect 1155 1550 1160 1830
rect 1120 1540 1160 1550
rect 2080 1830 2120 1840
rect 2080 1550 2085 1830
rect 2115 1550 2120 1830
rect 2080 1540 2120 1550
rect 3040 1830 3080 1840
rect 3040 1550 3045 1830
rect 3075 1550 3080 1830
rect 3040 1540 3080 1550
rect 4000 1830 4040 1840
rect 4000 1550 4005 1830
rect 4035 1550 4040 1830
rect 260 1515 1060 1520
rect 260 1485 270 1515
rect 1050 1485 1060 1515
rect 260 1480 1060 1485
rect 1220 1515 2020 1520
rect 1220 1485 1230 1515
rect 2010 1485 2020 1515
rect 1220 1480 2020 1485
rect 2180 1515 2980 1520
rect 2180 1485 2190 1515
rect 2970 1485 2980 1515
rect 2180 1480 2980 1485
rect 3140 1515 3940 1520
rect 3140 1485 3150 1515
rect 3930 1485 3940 1515
rect 3140 1480 3940 1485
rect 160 1365 165 1395
rect 195 1365 200 1395
rect 160 1235 200 1365
rect 160 1205 165 1235
rect 195 1205 200 1235
rect 160 1110 200 1205
rect 240 1395 280 1400
rect 240 1365 245 1395
rect 275 1365 280 1395
rect 240 1235 280 1365
rect 240 1205 245 1235
rect 275 1205 280 1235
rect 240 1200 280 1205
rect 320 1395 360 1400
rect 320 1365 325 1395
rect 355 1365 360 1395
rect 320 1235 360 1365
rect 320 1205 325 1235
rect 355 1205 360 1235
rect 320 1200 360 1205
rect 400 1395 440 1400
rect 400 1365 405 1395
rect 435 1365 440 1395
rect 400 1235 440 1365
rect 400 1205 405 1235
rect 435 1205 440 1235
rect 400 1200 440 1205
rect 480 1395 520 1400
rect 480 1365 485 1395
rect 515 1365 520 1395
rect 480 1235 520 1365
rect 480 1205 485 1235
rect 515 1205 520 1235
rect 480 1200 520 1205
rect 560 1395 600 1400
rect 560 1365 565 1395
rect 595 1365 600 1395
rect 560 1235 600 1365
rect 640 1315 680 1480
rect 640 1285 645 1315
rect 675 1285 680 1315
rect 640 1280 680 1285
rect 720 1395 760 1400
rect 720 1365 725 1395
rect 755 1365 760 1395
rect 560 1205 565 1235
rect 595 1205 600 1235
rect 560 1200 600 1205
rect 720 1235 760 1365
rect 720 1205 725 1235
rect 755 1205 760 1235
rect 720 1200 760 1205
rect 800 1395 840 1400
rect 800 1365 805 1395
rect 835 1365 840 1395
rect 800 1235 840 1365
rect 800 1205 805 1235
rect 835 1205 840 1235
rect 800 1200 840 1205
rect 880 1395 920 1400
rect 880 1365 885 1395
rect 915 1365 920 1395
rect 880 1235 920 1365
rect 880 1205 885 1235
rect 915 1205 920 1235
rect 880 1200 920 1205
rect 960 1395 1000 1400
rect 960 1365 965 1395
rect 995 1365 1000 1395
rect 960 1235 1000 1365
rect 960 1205 965 1235
rect 995 1205 1000 1235
rect 960 1200 1000 1205
rect 1040 1395 1080 1400
rect 1040 1365 1045 1395
rect 1075 1365 1080 1395
rect 1040 1235 1080 1365
rect 1040 1205 1045 1235
rect 1075 1205 1080 1235
rect 1040 1200 1080 1205
rect 1120 1395 1160 1400
rect 1120 1365 1125 1395
rect 1155 1365 1160 1395
rect 1120 1235 1160 1365
rect 1120 1205 1125 1235
rect 1155 1205 1160 1235
rect 1120 1200 1160 1205
rect 1200 1395 1240 1400
rect 1200 1365 1205 1395
rect 1235 1365 1240 1395
rect 1200 1235 1240 1365
rect 1200 1205 1205 1235
rect 1235 1205 1240 1235
rect 1200 1200 1240 1205
rect 1280 1395 1320 1400
rect 1280 1365 1285 1395
rect 1315 1365 1320 1395
rect 1280 1235 1320 1365
rect 1280 1205 1285 1235
rect 1315 1205 1320 1235
rect 1280 1200 1320 1205
rect 1360 1395 1400 1400
rect 1360 1365 1365 1395
rect 1395 1365 1400 1395
rect 1360 1235 1400 1365
rect 1360 1205 1365 1235
rect 1395 1205 1400 1235
rect 1360 1200 1400 1205
rect 1440 1395 1480 1400
rect 1440 1365 1445 1395
rect 1475 1365 1480 1395
rect 1440 1235 1480 1365
rect 1440 1205 1445 1235
rect 1475 1205 1480 1235
rect 1440 1200 1480 1205
rect 1520 1395 1560 1400
rect 1520 1365 1525 1395
rect 1555 1365 1560 1395
rect 1520 1235 1560 1365
rect 1600 1315 1640 1480
rect 1600 1285 1605 1315
rect 1635 1285 1640 1315
rect 1600 1280 1640 1285
rect 1680 1395 1720 1400
rect 1680 1365 1685 1395
rect 1715 1365 1720 1395
rect 1520 1205 1525 1235
rect 1555 1205 1560 1235
rect 1520 1200 1560 1205
rect 1680 1235 1720 1365
rect 1680 1205 1685 1235
rect 1715 1205 1720 1235
rect 1680 1200 1720 1205
rect 1760 1395 1800 1400
rect 1760 1365 1765 1395
rect 1795 1365 1800 1395
rect 1760 1235 1800 1365
rect 1760 1205 1765 1235
rect 1795 1205 1800 1235
rect 1760 1200 1800 1205
rect 1840 1395 1880 1400
rect 1840 1365 1845 1395
rect 1875 1365 1880 1395
rect 1840 1235 1880 1365
rect 1840 1205 1845 1235
rect 1875 1205 1880 1235
rect 1840 1200 1880 1205
rect 1920 1395 1960 1400
rect 1920 1365 1925 1395
rect 1955 1365 1960 1395
rect 1920 1235 1960 1365
rect 1920 1205 1925 1235
rect 1955 1205 1960 1235
rect 1920 1200 1960 1205
rect 2000 1395 2040 1400
rect 2000 1365 2005 1395
rect 2035 1365 2040 1395
rect 2000 1235 2040 1365
rect 2000 1205 2005 1235
rect 2035 1205 2040 1235
rect 2000 1200 2040 1205
rect 2080 1395 2120 1400
rect 2080 1365 2085 1395
rect 2115 1365 2120 1395
rect 2080 1235 2120 1365
rect 2080 1205 2085 1235
rect 2115 1205 2120 1235
rect 2080 1200 2120 1205
rect 2160 1395 2200 1400
rect 2160 1365 2165 1395
rect 2195 1365 2200 1395
rect 2160 1235 2200 1365
rect 2160 1205 2165 1235
rect 2195 1205 2200 1235
rect 2160 1200 2200 1205
rect 2240 1395 2280 1400
rect 2240 1365 2245 1395
rect 2275 1365 2280 1395
rect 2240 1235 2280 1365
rect 2240 1205 2245 1235
rect 2275 1205 2280 1235
rect 2240 1200 2280 1205
rect 2320 1395 2360 1400
rect 2320 1365 2325 1395
rect 2355 1365 2360 1395
rect 2320 1235 2360 1365
rect 2320 1205 2325 1235
rect 2355 1205 2360 1235
rect 2320 1200 2360 1205
rect 2400 1395 2440 1400
rect 2400 1365 2405 1395
rect 2435 1365 2440 1395
rect 2400 1235 2440 1365
rect 2400 1205 2405 1235
rect 2435 1205 2440 1235
rect 2400 1200 2440 1205
rect 2480 1395 2520 1400
rect 2480 1365 2485 1395
rect 2515 1365 2520 1395
rect 2480 1235 2520 1365
rect 2560 1315 2600 1480
rect 2560 1285 2565 1315
rect 2595 1285 2600 1315
rect 2560 1280 2600 1285
rect 2640 1395 2680 1400
rect 2640 1365 2645 1395
rect 2675 1365 2680 1395
rect 2480 1205 2485 1235
rect 2515 1205 2520 1235
rect 2480 1200 2520 1205
rect 2640 1235 2680 1365
rect 2640 1205 2645 1235
rect 2675 1205 2680 1235
rect 2640 1200 2680 1205
rect 2720 1395 2760 1400
rect 2720 1365 2725 1395
rect 2755 1365 2760 1395
rect 2720 1235 2760 1365
rect 2720 1205 2725 1235
rect 2755 1205 2760 1235
rect 2720 1200 2760 1205
rect 2800 1395 2840 1400
rect 2800 1365 2805 1395
rect 2835 1365 2840 1395
rect 2800 1235 2840 1365
rect 2800 1205 2805 1235
rect 2835 1205 2840 1235
rect 2800 1200 2840 1205
rect 2880 1395 2920 1400
rect 2880 1365 2885 1395
rect 2915 1365 2920 1395
rect 2880 1235 2920 1365
rect 2880 1205 2885 1235
rect 2915 1205 2920 1235
rect 2880 1200 2920 1205
rect 2960 1395 3000 1400
rect 2960 1365 2965 1395
rect 2995 1365 3000 1395
rect 2960 1235 3000 1365
rect 2960 1205 2965 1235
rect 2995 1205 3000 1235
rect 2960 1200 3000 1205
rect 3040 1395 3080 1400
rect 3040 1365 3045 1395
rect 3075 1365 3080 1395
rect 3040 1235 3080 1365
rect 3040 1205 3045 1235
rect 3075 1205 3080 1235
rect 3040 1200 3080 1205
rect 3120 1395 3160 1400
rect 3120 1365 3125 1395
rect 3155 1365 3160 1395
rect 3120 1235 3160 1365
rect 3120 1205 3125 1235
rect 3155 1205 3160 1235
rect 3120 1200 3160 1205
rect 3200 1395 3240 1400
rect 3200 1365 3205 1395
rect 3235 1365 3240 1395
rect 3200 1235 3240 1365
rect 3200 1205 3205 1235
rect 3235 1205 3240 1235
rect 3200 1200 3240 1205
rect 3280 1395 3320 1400
rect 3280 1365 3285 1395
rect 3315 1365 3320 1395
rect 3280 1235 3320 1365
rect 3280 1205 3285 1235
rect 3315 1205 3320 1235
rect 3280 1200 3320 1205
rect 3360 1395 3400 1400
rect 3360 1365 3365 1395
rect 3395 1365 3400 1395
rect 3360 1235 3400 1365
rect 3360 1205 3365 1235
rect 3395 1205 3400 1235
rect 3360 1200 3400 1205
rect 3440 1395 3480 1400
rect 3440 1365 3445 1395
rect 3475 1365 3480 1395
rect 3440 1235 3480 1365
rect 3520 1315 3560 1480
rect 3520 1285 3525 1315
rect 3555 1285 3560 1315
rect 3520 1280 3560 1285
rect 3600 1395 3640 1400
rect 3600 1365 3605 1395
rect 3635 1365 3640 1395
rect 3440 1205 3445 1235
rect 3475 1205 3480 1235
rect 3440 1200 3480 1205
rect 3600 1235 3640 1365
rect 3600 1205 3605 1235
rect 3635 1205 3640 1235
rect 3600 1200 3640 1205
rect 3680 1395 3720 1400
rect 3680 1365 3685 1395
rect 3715 1365 3720 1395
rect 3680 1235 3720 1365
rect 3680 1205 3685 1235
rect 3715 1205 3720 1235
rect 3680 1200 3720 1205
rect 3760 1395 3800 1400
rect 3760 1365 3765 1395
rect 3795 1365 3800 1395
rect 3760 1235 3800 1365
rect 3760 1205 3765 1235
rect 3795 1205 3800 1235
rect 3760 1200 3800 1205
rect 3840 1395 3880 1400
rect 3840 1365 3845 1395
rect 3875 1365 3880 1395
rect 3840 1235 3880 1365
rect 3840 1205 3845 1235
rect 3875 1205 3880 1235
rect 3840 1200 3880 1205
rect 3920 1395 3960 1400
rect 3920 1365 3925 1395
rect 3955 1365 3960 1395
rect 3920 1235 3960 1365
rect 3920 1205 3925 1235
rect 3955 1205 3960 1235
rect 3920 1200 3960 1205
rect 4000 1395 4040 1550
rect 4000 1365 4005 1395
rect 4035 1365 4040 1395
rect 4000 1235 4040 1365
rect 4000 1205 4005 1235
rect 4035 1205 4040 1235
rect 160 830 165 1110
rect 195 830 200 1110
rect 160 820 200 830
rect 1120 1110 1160 1120
rect 1120 830 1125 1110
rect 1155 830 1160 1110
rect 1120 820 1160 830
rect 2080 1110 2120 1120
rect 2080 830 2085 1110
rect 2115 830 2120 1110
rect 260 795 1060 800
rect 260 765 270 795
rect 1050 765 1060 795
rect 260 760 1060 765
rect 1220 795 2020 800
rect 1220 765 1230 795
rect 2010 765 2020 795
rect 1220 760 2020 765
rect 640 555 680 760
rect 640 525 645 555
rect 675 525 680 555
rect 80 475 120 480
rect 80 445 85 475
rect 115 445 120 475
rect 80 440 120 445
rect 160 470 200 480
rect 160 450 170 470
rect 190 450 200 470
rect 160 440 200 450
rect 240 470 280 480
rect 240 450 250 470
rect 270 450 280 470
rect 240 440 280 450
rect 320 470 360 480
rect 320 450 330 470
rect 350 450 360 470
rect 320 440 360 450
rect 400 470 440 480
rect 400 450 410 470
rect 430 450 440 470
rect 400 440 440 450
rect 480 470 520 480
rect 480 450 490 470
rect 510 450 520 470
rect 480 440 520 450
rect 560 470 600 480
rect 560 450 570 470
rect 590 450 600 470
rect 560 440 600 450
rect 640 240 680 525
rect 1600 555 1640 760
rect 1600 525 1605 555
rect 1635 525 1640 555
rect 720 470 760 480
rect 720 450 730 470
rect 750 450 760 470
rect 720 440 760 450
rect 800 470 840 480
rect 800 450 810 470
rect 830 450 840 470
rect 800 440 840 450
rect 880 470 920 480
rect 880 450 890 470
rect 910 450 920 470
rect 880 440 920 450
rect 960 470 1000 480
rect 960 450 970 470
rect 990 450 1000 470
rect 960 440 1000 450
rect 1040 470 1080 480
rect 1040 450 1050 470
rect 1070 450 1080 470
rect 1040 440 1080 450
rect 1120 470 1160 480
rect 1120 450 1130 470
rect 1150 450 1160 470
rect 1120 440 1160 450
rect 1200 470 1240 480
rect 1200 450 1210 470
rect 1230 450 1240 470
rect 1200 440 1240 450
rect 1280 470 1320 480
rect 1280 450 1290 470
rect 1310 450 1320 470
rect 1280 440 1320 450
rect 1360 470 1400 480
rect 1360 450 1370 470
rect 1390 450 1400 470
rect 1360 440 1400 450
rect 1440 470 1480 480
rect 1440 450 1450 470
rect 1470 450 1480 470
rect 1440 440 1480 450
rect 1520 470 1560 480
rect 1520 450 1530 470
rect 1550 450 1560 470
rect 1520 440 1560 450
rect 1600 240 1640 525
rect 1680 470 1720 480
rect 1680 450 1690 470
rect 1710 450 1720 470
rect 1680 440 1720 450
rect 1760 470 1800 480
rect 1760 450 1770 470
rect 1790 450 1800 470
rect 1760 440 1800 450
rect 1840 470 1880 480
rect 1840 450 1850 470
rect 1870 450 1880 470
rect 1840 440 1880 450
rect 1920 470 1960 480
rect 1920 450 1930 470
rect 1950 450 1960 470
rect 1920 440 1960 450
rect 2000 470 2040 480
rect 2000 450 2010 470
rect 2030 450 2040 470
rect 2000 440 2040 450
rect 2080 395 2120 830
rect 3040 1110 3080 1120
rect 3040 830 3045 1110
rect 3075 830 3080 1110
rect 3040 820 3080 830
rect 4000 1110 4040 1205
rect 4080 1395 4120 1400
rect 4080 1365 4085 1395
rect 4115 1365 4120 1395
rect 4080 1235 4120 1365
rect 4080 1205 4085 1235
rect 4115 1205 4120 1235
rect 4080 1200 4120 1205
rect 4160 1395 4200 1400
rect 4160 1365 4165 1395
rect 4195 1365 4200 1395
rect 4160 1235 4200 1365
rect 4160 1205 4165 1235
rect 4195 1205 4200 1235
rect 4160 1200 4200 1205
rect 4000 830 4005 1110
rect 4035 830 4040 1110
rect 4000 820 4040 830
rect 2180 795 2980 800
rect 2180 765 2190 795
rect 2970 765 2980 795
rect 2180 760 2980 765
rect 3140 795 3940 800
rect 3140 765 3150 795
rect 3930 765 3940 795
rect 3140 760 3940 765
rect 2560 555 2600 760
rect 2560 525 2565 555
rect 2595 525 2600 555
rect 2160 470 2200 480
rect 2160 450 2170 470
rect 2190 450 2200 470
rect 2160 440 2200 450
rect 2240 470 2280 480
rect 2240 450 2250 470
rect 2270 450 2280 470
rect 2240 440 2280 450
rect 2320 470 2360 480
rect 2320 450 2330 470
rect 2350 450 2360 470
rect 2320 440 2360 450
rect 2400 470 2440 480
rect 2400 450 2410 470
rect 2430 450 2440 470
rect 2400 440 2440 450
rect 2480 470 2520 480
rect 2480 450 2490 470
rect 2510 450 2520 470
rect 2480 440 2520 450
rect 2080 365 2085 395
rect 2115 365 2120 395
rect 260 235 1060 240
rect 260 205 270 235
rect 1050 205 1060 235
rect 260 200 1060 205
rect 1220 235 2020 240
rect 1220 205 1230 235
rect 2010 205 2020 235
rect 1220 200 2020 205
rect 160 170 200 180
rect 160 90 165 170
rect 195 90 200 170
rect 160 80 200 90
rect 1120 170 1160 180
rect 1120 90 1125 170
rect 1155 90 1160 170
rect 1120 80 1160 90
rect 2080 170 2120 365
rect 2560 240 2600 525
rect 3520 555 3560 760
rect 3520 525 3525 555
rect 3555 525 3560 555
rect 2640 470 2680 480
rect 2640 450 2650 470
rect 2670 450 2680 470
rect 2640 440 2680 450
rect 2720 470 2760 480
rect 2720 450 2730 470
rect 2750 450 2760 470
rect 2720 440 2760 450
rect 2800 470 2840 480
rect 2800 450 2810 470
rect 2830 450 2840 470
rect 2800 440 2840 450
rect 2880 470 2920 480
rect 2880 450 2890 470
rect 2910 450 2920 470
rect 2880 440 2920 450
rect 2960 470 3000 480
rect 2960 450 2970 470
rect 2990 450 3000 470
rect 2960 440 3000 450
rect 3040 470 3080 480
rect 3040 450 3050 470
rect 3070 450 3080 470
rect 3040 440 3080 450
rect 3120 470 3160 480
rect 3120 450 3130 470
rect 3150 450 3160 470
rect 3120 440 3160 450
rect 3200 470 3240 480
rect 3200 450 3210 470
rect 3230 450 3240 470
rect 3200 440 3240 450
rect 3280 470 3320 480
rect 3280 450 3290 470
rect 3310 450 3320 470
rect 3280 440 3320 450
rect 3360 470 3400 480
rect 3360 450 3370 470
rect 3390 450 3400 470
rect 3360 440 3400 450
rect 3440 470 3480 480
rect 3440 450 3450 470
rect 3470 450 3480 470
rect 3440 440 3480 450
rect 3520 240 3560 525
rect 3600 470 3640 480
rect 3600 450 3610 470
rect 3630 450 3640 470
rect 3600 440 3640 450
rect 3680 470 3720 480
rect 3680 450 3690 470
rect 3710 450 3720 470
rect 3680 440 3720 450
rect 3760 470 3800 480
rect 3760 450 3770 470
rect 3790 450 3800 470
rect 3760 440 3800 450
rect 3840 470 3880 480
rect 3840 450 3850 470
rect 3870 450 3880 470
rect 3840 440 3880 450
rect 3920 470 3960 480
rect 3920 450 3930 470
rect 3950 450 3960 470
rect 3920 440 3960 450
rect 4000 470 4040 480
rect 4000 450 4010 470
rect 4030 450 4040 470
rect 4000 440 4040 450
rect 4080 470 4120 480
rect 4080 450 4090 470
rect 4110 450 4120 470
rect 4080 440 4120 450
rect 2180 235 2980 240
rect 2180 205 2190 235
rect 2970 205 2980 235
rect 2180 200 2980 205
rect 3140 235 3940 240
rect 3140 205 3150 235
rect 3930 205 3940 235
rect 3140 200 3940 205
rect 2080 90 2085 170
rect 2115 90 2120 170
rect 2080 80 2120 90
rect 3040 170 3080 180
rect 3040 90 3045 170
rect 3075 90 3080 170
rect 3040 80 3080 90
rect 4000 170 4040 180
rect 4000 90 4005 170
rect 4035 90 4040 170
rect 4000 80 4040 90
<< via1 >>
rect 5 1365 35 1395
rect 5 1205 35 1235
rect 85 1365 115 1395
rect 85 1205 115 1235
rect 2085 1650 2115 1830
rect 165 1365 195 1395
rect 165 1205 195 1235
rect 245 1365 275 1395
rect 245 1205 275 1235
rect 325 1365 355 1395
rect 325 1205 355 1235
rect 405 1365 435 1395
rect 405 1205 435 1235
rect 485 1365 515 1395
rect 485 1205 515 1235
rect 565 1365 595 1395
rect 645 1285 675 1315
rect 725 1365 755 1395
rect 565 1205 595 1235
rect 725 1205 755 1235
rect 805 1365 835 1395
rect 805 1205 835 1235
rect 885 1365 915 1395
rect 885 1205 915 1235
rect 965 1365 995 1395
rect 965 1205 995 1235
rect 1045 1365 1075 1395
rect 1045 1205 1075 1235
rect 1125 1365 1155 1395
rect 1125 1205 1155 1235
rect 1205 1365 1235 1395
rect 1205 1205 1235 1235
rect 1285 1365 1315 1395
rect 1285 1205 1315 1235
rect 1365 1365 1395 1395
rect 1365 1205 1395 1235
rect 1445 1365 1475 1395
rect 1445 1205 1475 1235
rect 1525 1365 1555 1395
rect 1605 1285 1635 1315
rect 1685 1365 1715 1395
rect 1525 1205 1555 1235
rect 1685 1205 1715 1235
rect 1765 1365 1795 1395
rect 1765 1205 1795 1235
rect 1845 1365 1875 1395
rect 1845 1205 1875 1235
rect 1925 1365 1955 1395
rect 1925 1205 1955 1235
rect 2005 1365 2035 1395
rect 2005 1205 2035 1235
rect 2085 1365 2115 1395
rect 2085 1205 2115 1235
rect 2165 1365 2195 1395
rect 2165 1205 2195 1235
rect 2245 1365 2275 1395
rect 2245 1205 2275 1235
rect 2325 1365 2355 1395
rect 2325 1205 2355 1235
rect 2405 1365 2435 1395
rect 2405 1205 2435 1235
rect 2485 1365 2515 1395
rect 2565 1285 2595 1315
rect 2645 1365 2675 1395
rect 2485 1205 2515 1235
rect 2645 1205 2675 1235
rect 2725 1365 2755 1395
rect 2725 1205 2755 1235
rect 2805 1365 2835 1395
rect 2805 1205 2835 1235
rect 2885 1365 2915 1395
rect 2885 1205 2915 1235
rect 2965 1365 2995 1395
rect 2965 1205 2995 1235
rect 3045 1365 3075 1395
rect 3045 1205 3075 1235
rect 3125 1365 3155 1395
rect 3125 1205 3155 1235
rect 3205 1365 3235 1395
rect 3205 1205 3235 1235
rect 3285 1365 3315 1395
rect 3285 1205 3315 1235
rect 3365 1365 3395 1395
rect 3365 1205 3395 1235
rect 3445 1365 3475 1395
rect 3525 1285 3555 1315
rect 3605 1365 3635 1395
rect 3445 1205 3475 1235
rect 3605 1205 3635 1235
rect 3685 1365 3715 1395
rect 3685 1205 3715 1235
rect 3765 1365 3795 1395
rect 3765 1205 3795 1235
rect 3845 1365 3875 1395
rect 3845 1205 3875 1235
rect 3925 1365 3955 1395
rect 3925 1205 3955 1235
rect 4005 1365 4035 1395
rect 4005 1205 4035 1235
rect 645 525 675 555
rect 85 470 115 475
rect 85 450 90 470
rect 90 450 110 470
rect 110 450 115 470
rect 85 445 115 450
rect 1605 525 1635 555
rect 4085 1365 4115 1395
rect 4085 1205 4115 1235
rect 4165 1365 4195 1395
rect 4165 1205 4195 1235
rect 2565 525 2595 555
rect 2085 365 2115 395
rect 165 90 195 170
rect 3525 525 3555 555
rect 4005 90 4035 170
<< metal2 >>
rect 2080 1830 2120 1840
rect 2080 1650 2085 1830
rect 2115 1650 2120 1830
rect 2080 1640 2120 1650
rect 0 1395 4200 1400
rect 0 1365 5 1395
rect 35 1365 85 1395
rect 115 1365 165 1395
rect 195 1365 245 1395
rect 275 1365 325 1395
rect 355 1365 405 1395
rect 435 1365 485 1395
rect 515 1365 565 1395
rect 595 1365 725 1395
rect 755 1365 805 1395
rect 835 1365 885 1395
rect 915 1365 965 1395
rect 995 1365 1045 1395
rect 1075 1365 1125 1395
rect 1155 1365 1205 1395
rect 1235 1365 1285 1395
rect 1315 1365 1365 1395
rect 1395 1365 1445 1395
rect 1475 1365 1525 1395
rect 1555 1365 1685 1395
rect 1715 1365 1765 1395
rect 1795 1365 1845 1395
rect 1875 1365 1925 1395
rect 1955 1365 2005 1395
rect 2035 1365 2085 1395
rect 2115 1365 2165 1395
rect 2195 1365 2245 1395
rect 2275 1365 2325 1395
rect 2355 1365 2405 1395
rect 2435 1365 2485 1395
rect 2515 1365 2645 1395
rect 2675 1365 2725 1395
rect 2755 1365 2805 1395
rect 2835 1365 2885 1395
rect 2915 1365 2965 1395
rect 2995 1365 3045 1395
rect 3075 1365 3125 1395
rect 3155 1365 3205 1395
rect 3235 1365 3285 1395
rect 3315 1365 3365 1395
rect 3395 1365 3445 1395
rect 3475 1365 3605 1395
rect 3635 1365 3685 1395
rect 3715 1365 3765 1395
rect 3795 1365 3845 1395
rect 3875 1365 3925 1395
rect 3955 1365 4005 1395
rect 4035 1365 4085 1395
rect 4115 1365 4165 1395
rect 4195 1365 4200 1395
rect 0 1360 4200 1365
rect 0 1315 4200 1320
rect 0 1285 645 1315
rect 675 1285 1605 1315
rect 1635 1285 2565 1315
rect 2595 1285 3525 1315
rect 3555 1285 4200 1315
rect 0 1280 4200 1285
rect 0 1235 4200 1240
rect 0 1205 5 1235
rect 35 1205 85 1235
rect 115 1205 165 1235
rect 195 1205 245 1235
rect 275 1205 325 1235
rect 355 1205 405 1235
rect 435 1205 485 1235
rect 515 1205 565 1235
rect 595 1205 725 1235
rect 755 1205 805 1235
rect 835 1205 885 1235
rect 915 1205 965 1235
rect 995 1205 1045 1235
rect 1075 1205 1125 1235
rect 1155 1205 1205 1235
rect 1235 1205 1285 1235
rect 1315 1205 1365 1235
rect 1395 1205 1445 1235
rect 1475 1205 1525 1235
rect 1555 1205 1685 1235
rect 1715 1205 1765 1235
rect 1795 1205 1845 1235
rect 1875 1205 1925 1235
rect 1955 1205 2005 1235
rect 2035 1205 2085 1235
rect 2115 1205 2165 1235
rect 2195 1205 2245 1235
rect 2275 1205 2325 1235
rect 2355 1205 2405 1235
rect 2435 1205 2485 1235
rect 2515 1205 2645 1235
rect 2675 1205 2725 1235
rect 2755 1205 2805 1235
rect 2835 1205 2885 1235
rect 2915 1205 2965 1235
rect 2995 1205 3045 1235
rect 3075 1205 3125 1235
rect 3155 1205 3205 1235
rect 3235 1205 3285 1235
rect 3315 1205 3365 1235
rect 3395 1205 3445 1235
rect 3475 1205 3605 1235
rect 3635 1205 3685 1235
rect 3715 1205 3765 1235
rect 3795 1205 3845 1235
rect 3875 1205 3925 1235
rect 3955 1205 4005 1235
rect 4035 1205 4085 1235
rect 4115 1205 4165 1235
rect 4195 1205 4200 1235
rect 0 1200 4200 1205
rect 0 635 4200 640
rect 0 605 85 635
rect 115 605 165 635
rect 195 605 245 635
rect 275 605 325 635
rect 355 605 405 635
rect 435 605 485 635
rect 515 605 565 635
rect 595 605 725 635
rect 755 605 805 635
rect 835 605 885 635
rect 915 605 965 635
rect 995 605 1045 635
rect 1075 605 1125 635
rect 1155 605 1205 635
rect 1235 605 1285 635
rect 1315 605 1365 635
rect 1395 605 1445 635
rect 1475 605 1525 635
rect 1555 605 1685 635
rect 1715 605 1765 635
rect 1795 605 1845 635
rect 1875 605 1925 635
rect 1955 605 2005 635
rect 2035 605 2165 635
rect 2195 605 2245 635
rect 2275 605 2325 635
rect 2355 605 2405 635
rect 2435 605 2485 635
rect 2515 605 2645 635
rect 2675 605 2725 635
rect 2755 605 2805 635
rect 2835 605 2885 635
rect 2915 605 2965 635
rect 2995 605 3045 635
rect 3075 605 3125 635
rect 3155 605 3205 635
rect 3235 605 3285 635
rect 3315 605 3365 635
rect 3395 605 3445 635
rect 3475 605 3605 635
rect 3635 605 3685 635
rect 3715 605 3765 635
rect 3795 605 3845 635
rect 3875 605 3925 635
rect 3955 605 4005 635
rect 4035 605 4085 635
rect 4115 605 4200 635
rect 0 600 4200 605
rect 0 555 4200 560
rect 0 525 645 555
rect 675 525 1605 555
rect 1635 525 2565 555
rect 2595 525 3525 555
rect 3555 525 4200 555
rect 0 520 4200 525
rect 0 475 4200 480
rect 0 445 85 475
rect 115 445 165 475
rect 195 445 245 475
rect 275 445 325 475
rect 355 445 405 475
rect 435 445 485 475
rect 515 445 565 475
rect 595 445 725 475
rect 755 445 805 475
rect 835 445 885 475
rect 915 445 965 475
rect 995 445 1045 475
rect 1075 445 1125 475
rect 1155 445 1205 475
rect 1235 445 1285 475
rect 1315 445 1365 475
rect 1395 445 1445 475
rect 1475 445 1525 475
rect 1555 445 1685 475
rect 1715 445 1765 475
rect 1795 445 1845 475
rect 1875 445 1925 475
rect 1955 445 2005 475
rect 2035 445 2165 475
rect 2195 445 2245 475
rect 2275 445 2325 475
rect 2355 445 2405 475
rect 2435 445 2485 475
rect 2515 445 2645 475
rect 2675 445 2725 475
rect 2755 445 2805 475
rect 2835 445 2885 475
rect 2915 445 2965 475
rect 2995 445 3045 475
rect 3075 445 3125 475
rect 3155 445 3205 475
rect 3235 445 3285 475
rect 3315 445 3365 475
rect 3395 445 3445 475
rect 3475 445 3605 475
rect 3635 445 3685 475
rect 3715 445 3765 475
rect 3795 445 3845 475
rect 3875 445 3925 475
rect 3955 445 4005 475
rect 4035 445 4085 475
rect 4115 445 4200 475
rect 0 440 4200 445
rect 0 395 4200 400
rect 0 365 2085 395
rect 2115 365 4200 395
rect 0 360 4200 365
rect 0 315 4200 320
rect 0 285 85 315
rect 115 285 165 315
rect 195 285 245 315
rect 275 285 325 315
rect 355 285 405 315
rect 435 285 485 315
rect 515 285 565 315
rect 595 285 725 315
rect 755 285 805 315
rect 835 285 885 315
rect 915 285 965 315
rect 995 285 1045 315
rect 1075 285 1125 315
rect 1155 285 1205 315
rect 1235 285 1285 315
rect 1315 285 1365 315
rect 1395 285 1445 315
rect 1475 285 1525 315
rect 1555 285 1685 315
rect 1715 285 1765 315
rect 1795 285 1845 315
rect 1875 285 1925 315
rect 1955 285 2005 315
rect 2035 285 2165 315
rect 2195 285 2245 315
rect 2275 285 2325 315
rect 2355 285 2405 315
rect 2435 285 2485 315
rect 2515 285 2645 315
rect 2675 285 2725 315
rect 2755 285 2805 315
rect 2835 285 2885 315
rect 2915 285 2965 315
rect 2995 285 3045 315
rect 3075 285 3125 315
rect 3155 285 3205 315
rect 3235 285 3285 315
rect 3315 285 3365 315
rect 3395 285 3445 315
rect 3475 285 3605 315
rect 3635 285 3685 315
rect 3715 285 3765 315
rect 3795 285 3845 315
rect 3875 285 3925 315
rect 3955 285 4005 315
rect 4035 285 4085 315
rect 4115 285 4200 315
rect 0 280 4200 285
rect 160 170 200 180
rect 160 90 165 170
rect 195 90 200 170
rect 160 80 200 90
rect 4000 170 4040 180
rect 4000 90 4005 170
rect 4035 90 4040 170
rect 4000 80 4040 90
<< via2 >>
rect 2085 1650 2115 1830
rect 5 1365 35 1395
rect 85 1365 115 1395
rect 165 1365 195 1395
rect 245 1365 275 1395
rect 325 1365 355 1395
rect 405 1365 435 1395
rect 485 1365 515 1395
rect 565 1365 595 1395
rect 725 1365 755 1395
rect 805 1365 835 1395
rect 885 1365 915 1395
rect 965 1365 995 1395
rect 1045 1365 1075 1395
rect 1125 1365 1155 1395
rect 1205 1365 1235 1395
rect 1285 1365 1315 1395
rect 1365 1365 1395 1395
rect 1445 1365 1475 1395
rect 1525 1365 1555 1395
rect 1685 1365 1715 1395
rect 1765 1365 1795 1395
rect 1845 1365 1875 1395
rect 1925 1365 1955 1395
rect 2005 1365 2035 1395
rect 2085 1365 2115 1395
rect 2165 1365 2195 1395
rect 2245 1365 2275 1395
rect 2325 1365 2355 1395
rect 2405 1365 2435 1395
rect 2485 1365 2515 1395
rect 2645 1365 2675 1395
rect 2725 1365 2755 1395
rect 2805 1365 2835 1395
rect 2885 1365 2915 1395
rect 2965 1365 2995 1395
rect 3045 1365 3075 1395
rect 3125 1365 3155 1395
rect 3205 1365 3235 1395
rect 3285 1365 3315 1395
rect 3365 1365 3395 1395
rect 3445 1365 3475 1395
rect 3605 1365 3635 1395
rect 3685 1365 3715 1395
rect 3765 1365 3795 1395
rect 3845 1365 3875 1395
rect 3925 1365 3955 1395
rect 4005 1365 4035 1395
rect 4085 1365 4115 1395
rect 4165 1365 4195 1395
rect 5 1205 35 1235
rect 85 1205 115 1235
rect 165 1205 195 1235
rect 245 1205 275 1235
rect 325 1205 355 1235
rect 405 1205 435 1235
rect 485 1205 515 1235
rect 565 1205 595 1235
rect 725 1205 755 1235
rect 805 1205 835 1235
rect 885 1205 915 1235
rect 965 1205 995 1235
rect 1045 1205 1075 1235
rect 1125 1205 1155 1235
rect 1205 1205 1235 1235
rect 1285 1205 1315 1235
rect 1365 1205 1395 1235
rect 1445 1205 1475 1235
rect 1525 1205 1555 1235
rect 1685 1205 1715 1235
rect 1765 1205 1795 1235
rect 1845 1205 1875 1235
rect 1925 1205 1955 1235
rect 2005 1205 2035 1235
rect 2085 1205 2115 1235
rect 2165 1205 2195 1235
rect 2245 1205 2275 1235
rect 2325 1205 2355 1235
rect 2405 1205 2435 1235
rect 2485 1205 2515 1235
rect 2645 1205 2675 1235
rect 2725 1205 2755 1235
rect 2805 1205 2835 1235
rect 2885 1205 2915 1235
rect 2965 1205 2995 1235
rect 3045 1205 3075 1235
rect 3125 1205 3155 1235
rect 3205 1205 3235 1235
rect 3285 1205 3315 1235
rect 3365 1205 3395 1235
rect 3445 1205 3475 1235
rect 3605 1205 3635 1235
rect 3685 1205 3715 1235
rect 3765 1205 3795 1235
rect 3845 1205 3875 1235
rect 3925 1205 3955 1235
rect 4005 1205 4035 1235
rect 4085 1205 4115 1235
rect 4165 1205 4195 1235
rect 85 605 115 635
rect 165 605 195 635
rect 245 605 275 635
rect 325 605 355 635
rect 405 605 435 635
rect 485 605 515 635
rect 565 605 595 635
rect 725 605 755 635
rect 805 605 835 635
rect 885 605 915 635
rect 965 605 995 635
rect 1045 605 1075 635
rect 1125 605 1155 635
rect 1205 605 1235 635
rect 1285 605 1315 635
rect 1365 605 1395 635
rect 1445 605 1475 635
rect 1525 605 1555 635
rect 1685 605 1715 635
rect 1765 605 1795 635
rect 1845 605 1875 635
rect 1925 605 1955 635
rect 2005 605 2035 635
rect 2165 605 2195 635
rect 2245 605 2275 635
rect 2325 605 2355 635
rect 2405 605 2435 635
rect 2485 605 2515 635
rect 2645 605 2675 635
rect 2725 605 2755 635
rect 2805 605 2835 635
rect 2885 605 2915 635
rect 2965 605 2995 635
rect 3045 605 3075 635
rect 3125 605 3155 635
rect 3205 605 3235 635
rect 3285 605 3315 635
rect 3365 605 3395 635
rect 3445 605 3475 635
rect 3605 605 3635 635
rect 3685 605 3715 635
rect 3765 605 3795 635
rect 3845 605 3875 635
rect 3925 605 3955 635
rect 4005 605 4035 635
rect 4085 605 4115 635
rect 85 445 115 475
rect 165 445 195 475
rect 245 445 275 475
rect 325 445 355 475
rect 405 445 435 475
rect 485 445 515 475
rect 565 445 595 475
rect 725 445 755 475
rect 805 445 835 475
rect 885 445 915 475
rect 965 445 995 475
rect 1045 445 1075 475
rect 1125 445 1155 475
rect 1205 445 1235 475
rect 1285 445 1315 475
rect 1365 445 1395 475
rect 1445 445 1475 475
rect 1525 445 1555 475
rect 1685 445 1715 475
rect 1765 445 1795 475
rect 1845 445 1875 475
rect 1925 445 1955 475
rect 2005 445 2035 475
rect 2165 445 2195 475
rect 2245 445 2275 475
rect 2325 445 2355 475
rect 2405 445 2435 475
rect 2485 445 2515 475
rect 2645 445 2675 475
rect 2725 445 2755 475
rect 2805 445 2835 475
rect 2885 445 2915 475
rect 2965 445 2995 475
rect 3045 445 3075 475
rect 3125 445 3155 475
rect 3205 445 3235 475
rect 3285 445 3315 475
rect 3365 445 3395 475
rect 3445 445 3475 475
rect 3605 445 3635 475
rect 3685 445 3715 475
rect 3765 445 3795 475
rect 3845 445 3875 475
rect 3925 445 3955 475
rect 4005 445 4035 475
rect 4085 445 4115 475
rect 85 285 115 315
rect 165 285 195 315
rect 245 285 275 315
rect 325 285 355 315
rect 405 285 435 315
rect 485 285 515 315
rect 565 285 595 315
rect 725 285 755 315
rect 805 285 835 315
rect 885 285 915 315
rect 965 285 995 315
rect 1045 285 1075 315
rect 1125 285 1155 315
rect 1205 285 1235 315
rect 1285 285 1315 315
rect 1365 285 1395 315
rect 1445 285 1475 315
rect 1525 285 1555 315
rect 1685 285 1715 315
rect 1765 285 1795 315
rect 1845 285 1875 315
rect 1925 285 1955 315
rect 2005 285 2035 315
rect 2165 285 2195 315
rect 2245 285 2275 315
rect 2325 285 2355 315
rect 2405 285 2435 315
rect 2485 285 2515 315
rect 2645 285 2675 315
rect 2725 285 2755 315
rect 2805 285 2835 315
rect 2885 285 2915 315
rect 2965 285 2995 315
rect 3045 285 3075 315
rect 3125 285 3155 315
rect 3205 285 3235 315
rect 3285 285 3315 315
rect 3365 285 3395 315
rect 3445 285 3475 315
rect 3605 285 3635 315
rect 3685 285 3715 315
rect 3765 285 3795 315
rect 3845 285 3875 315
rect 3925 285 3955 315
rect 4005 285 4035 315
rect 4085 285 4115 315
rect 165 90 195 170
rect 4005 90 4035 170
<< metal3 >>
rect 2080 1831 2120 1840
rect 2080 1649 2084 1831
rect 2116 1649 2120 1831
rect 2080 1640 2120 1649
rect 0 1396 40 1400
rect 0 1364 4 1396
rect 36 1364 40 1396
rect 0 1236 40 1364
rect 0 1204 4 1236
rect 36 1204 40 1236
rect 0 1200 40 1204
rect 80 1396 120 1400
rect 80 1364 84 1396
rect 116 1364 120 1396
rect 80 1236 120 1364
rect 80 1204 84 1236
rect 116 1204 120 1236
rect 80 1200 120 1204
rect 160 1396 200 1400
rect 160 1364 164 1396
rect 196 1364 200 1396
rect 160 1236 200 1364
rect 160 1204 164 1236
rect 196 1204 200 1236
rect 160 1200 200 1204
rect 240 1396 280 1400
rect 240 1364 244 1396
rect 276 1364 280 1396
rect 240 1236 280 1364
rect 240 1204 244 1236
rect 276 1204 280 1236
rect 240 1200 280 1204
rect 320 1396 360 1400
rect 320 1364 324 1396
rect 356 1364 360 1396
rect 320 1236 360 1364
rect 320 1204 324 1236
rect 356 1204 360 1236
rect 320 1200 360 1204
rect 400 1396 440 1400
rect 400 1364 404 1396
rect 436 1364 440 1396
rect 400 1236 440 1364
rect 400 1204 404 1236
rect 436 1204 440 1236
rect 400 1200 440 1204
rect 480 1396 520 1400
rect 480 1364 484 1396
rect 516 1364 520 1396
rect 480 1236 520 1364
rect 480 1204 484 1236
rect 516 1204 520 1236
rect 480 1200 520 1204
rect 560 1396 600 1400
rect 560 1364 564 1396
rect 596 1364 600 1396
rect 560 1236 600 1364
rect 560 1204 564 1236
rect 596 1204 600 1236
rect 560 1200 600 1204
rect 720 1396 760 1400
rect 720 1364 724 1396
rect 756 1364 760 1396
rect 720 1236 760 1364
rect 720 1204 724 1236
rect 756 1204 760 1236
rect 720 1200 760 1204
rect 800 1396 840 1400
rect 800 1364 804 1396
rect 836 1364 840 1396
rect 800 1236 840 1364
rect 800 1204 804 1236
rect 836 1204 840 1236
rect 800 1200 840 1204
rect 880 1396 920 1400
rect 880 1364 884 1396
rect 916 1364 920 1396
rect 880 1236 920 1364
rect 880 1204 884 1236
rect 916 1204 920 1236
rect 880 1200 920 1204
rect 960 1396 1000 1400
rect 960 1364 964 1396
rect 996 1364 1000 1396
rect 960 1236 1000 1364
rect 960 1204 964 1236
rect 996 1204 1000 1236
rect 960 1200 1000 1204
rect 1040 1396 1080 1400
rect 1040 1364 1044 1396
rect 1076 1364 1080 1396
rect 1040 1236 1080 1364
rect 1040 1204 1044 1236
rect 1076 1204 1080 1236
rect 1040 1200 1080 1204
rect 1120 1396 1160 1400
rect 1120 1364 1124 1396
rect 1156 1364 1160 1396
rect 1120 1236 1160 1364
rect 1120 1204 1124 1236
rect 1156 1204 1160 1236
rect 1120 1200 1160 1204
rect 1200 1396 1240 1400
rect 1200 1364 1204 1396
rect 1236 1364 1240 1396
rect 1200 1236 1240 1364
rect 1200 1204 1204 1236
rect 1236 1204 1240 1236
rect 1200 1200 1240 1204
rect 1280 1396 1320 1400
rect 1280 1364 1284 1396
rect 1316 1364 1320 1396
rect 1280 1236 1320 1364
rect 1280 1204 1284 1236
rect 1316 1204 1320 1236
rect 1280 1200 1320 1204
rect 1360 1396 1400 1400
rect 1360 1364 1364 1396
rect 1396 1364 1400 1396
rect 1360 1236 1400 1364
rect 1360 1204 1364 1236
rect 1396 1204 1400 1236
rect 1360 1200 1400 1204
rect 1440 1396 1480 1400
rect 1440 1364 1444 1396
rect 1476 1364 1480 1396
rect 1440 1236 1480 1364
rect 1440 1204 1444 1236
rect 1476 1204 1480 1236
rect 1440 1200 1480 1204
rect 1520 1396 1560 1400
rect 1520 1364 1524 1396
rect 1556 1364 1560 1396
rect 1520 1236 1560 1364
rect 1520 1204 1524 1236
rect 1556 1204 1560 1236
rect 1520 1200 1560 1204
rect 1680 1396 1720 1400
rect 1680 1364 1684 1396
rect 1716 1364 1720 1396
rect 1680 1236 1720 1364
rect 1680 1204 1684 1236
rect 1716 1204 1720 1236
rect 1680 1200 1720 1204
rect 1760 1396 1800 1400
rect 1760 1364 1764 1396
rect 1796 1364 1800 1396
rect 1760 1236 1800 1364
rect 1760 1204 1764 1236
rect 1796 1204 1800 1236
rect 1760 1200 1800 1204
rect 1840 1396 1880 1400
rect 1840 1364 1844 1396
rect 1876 1364 1880 1396
rect 1840 1236 1880 1364
rect 1840 1204 1844 1236
rect 1876 1204 1880 1236
rect 1840 1200 1880 1204
rect 1920 1396 1960 1400
rect 1920 1364 1924 1396
rect 1956 1364 1960 1396
rect 1920 1236 1960 1364
rect 1920 1204 1924 1236
rect 1956 1204 1960 1236
rect 1920 1200 1960 1204
rect 2000 1396 2040 1400
rect 2000 1364 2004 1396
rect 2036 1364 2040 1396
rect 2000 1236 2040 1364
rect 2000 1204 2004 1236
rect 2036 1204 2040 1236
rect 2000 1200 2040 1204
rect 2080 1396 2120 1400
rect 2080 1364 2084 1396
rect 2116 1364 2120 1396
rect 2080 1236 2120 1364
rect 2080 1204 2084 1236
rect 2116 1204 2120 1236
rect 2080 1200 2120 1204
rect 2160 1396 2200 1400
rect 2160 1364 2164 1396
rect 2196 1364 2200 1396
rect 2160 1236 2200 1364
rect 2160 1204 2164 1236
rect 2196 1204 2200 1236
rect 2160 1200 2200 1204
rect 2240 1396 2280 1400
rect 2240 1364 2244 1396
rect 2276 1364 2280 1396
rect 2240 1236 2280 1364
rect 2240 1204 2244 1236
rect 2276 1204 2280 1236
rect 2240 1200 2280 1204
rect 2320 1396 2360 1400
rect 2320 1364 2324 1396
rect 2356 1364 2360 1396
rect 2320 1236 2360 1364
rect 2320 1204 2324 1236
rect 2356 1204 2360 1236
rect 2320 1200 2360 1204
rect 2400 1396 2440 1400
rect 2400 1364 2404 1396
rect 2436 1364 2440 1396
rect 2400 1236 2440 1364
rect 2400 1204 2404 1236
rect 2436 1204 2440 1236
rect 2400 1200 2440 1204
rect 2480 1396 2520 1400
rect 2480 1364 2484 1396
rect 2516 1364 2520 1396
rect 2480 1236 2520 1364
rect 2480 1204 2484 1236
rect 2516 1204 2520 1236
rect 2480 1200 2520 1204
rect 2640 1396 2680 1400
rect 2640 1364 2644 1396
rect 2676 1364 2680 1396
rect 2640 1236 2680 1364
rect 2640 1204 2644 1236
rect 2676 1204 2680 1236
rect 2640 1200 2680 1204
rect 2720 1396 2760 1400
rect 2720 1364 2724 1396
rect 2756 1364 2760 1396
rect 2720 1236 2760 1364
rect 2720 1204 2724 1236
rect 2756 1204 2760 1236
rect 2720 1200 2760 1204
rect 2800 1396 2840 1400
rect 2800 1364 2804 1396
rect 2836 1364 2840 1396
rect 2800 1236 2840 1364
rect 2800 1204 2804 1236
rect 2836 1204 2840 1236
rect 2800 1200 2840 1204
rect 2880 1396 2920 1400
rect 2880 1364 2884 1396
rect 2916 1364 2920 1396
rect 2880 1236 2920 1364
rect 2880 1204 2884 1236
rect 2916 1204 2920 1236
rect 2880 1200 2920 1204
rect 2960 1396 3000 1400
rect 2960 1364 2964 1396
rect 2996 1364 3000 1396
rect 2960 1236 3000 1364
rect 2960 1204 2964 1236
rect 2996 1204 3000 1236
rect 2960 1200 3000 1204
rect 3040 1396 3080 1400
rect 3040 1364 3044 1396
rect 3076 1364 3080 1396
rect 3040 1236 3080 1364
rect 3040 1204 3044 1236
rect 3076 1204 3080 1236
rect 3040 1200 3080 1204
rect 3120 1396 3160 1400
rect 3120 1364 3124 1396
rect 3156 1364 3160 1396
rect 3120 1236 3160 1364
rect 3120 1204 3124 1236
rect 3156 1204 3160 1236
rect 3120 1200 3160 1204
rect 3200 1396 3240 1400
rect 3200 1364 3204 1396
rect 3236 1364 3240 1396
rect 3200 1236 3240 1364
rect 3200 1204 3204 1236
rect 3236 1204 3240 1236
rect 3200 1200 3240 1204
rect 3280 1396 3320 1400
rect 3280 1364 3284 1396
rect 3316 1364 3320 1396
rect 3280 1236 3320 1364
rect 3280 1204 3284 1236
rect 3316 1204 3320 1236
rect 3280 1200 3320 1204
rect 3360 1396 3400 1400
rect 3360 1364 3364 1396
rect 3396 1364 3400 1396
rect 3360 1236 3400 1364
rect 3360 1204 3364 1236
rect 3396 1204 3400 1236
rect 3360 1200 3400 1204
rect 3440 1396 3480 1400
rect 3440 1364 3444 1396
rect 3476 1364 3480 1396
rect 3440 1236 3480 1364
rect 3440 1204 3444 1236
rect 3476 1204 3480 1236
rect 3440 1200 3480 1204
rect 3600 1396 3640 1400
rect 3600 1364 3604 1396
rect 3636 1364 3640 1396
rect 3600 1236 3640 1364
rect 3600 1204 3604 1236
rect 3636 1204 3640 1236
rect 3600 1200 3640 1204
rect 3680 1396 3720 1400
rect 3680 1364 3684 1396
rect 3716 1364 3720 1396
rect 3680 1236 3720 1364
rect 3680 1204 3684 1236
rect 3716 1204 3720 1236
rect 3680 1200 3720 1204
rect 3760 1396 3800 1400
rect 3760 1364 3764 1396
rect 3796 1364 3800 1396
rect 3760 1236 3800 1364
rect 3760 1204 3764 1236
rect 3796 1204 3800 1236
rect 3760 1200 3800 1204
rect 3840 1396 3880 1400
rect 3840 1364 3844 1396
rect 3876 1364 3880 1396
rect 3840 1236 3880 1364
rect 3840 1204 3844 1236
rect 3876 1204 3880 1236
rect 3840 1200 3880 1204
rect 3920 1396 3960 1400
rect 3920 1364 3924 1396
rect 3956 1364 3960 1396
rect 3920 1236 3960 1364
rect 3920 1204 3924 1236
rect 3956 1204 3960 1236
rect 3920 1200 3960 1204
rect 4000 1396 4040 1400
rect 4000 1364 4004 1396
rect 4036 1364 4040 1396
rect 4000 1236 4040 1364
rect 4000 1204 4004 1236
rect 4036 1204 4040 1236
rect 4000 1200 4040 1204
rect 4080 1396 4120 1400
rect 4080 1364 4084 1396
rect 4116 1364 4120 1396
rect 4080 1236 4120 1364
rect 4080 1204 4084 1236
rect 4116 1204 4120 1236
rect 4080 1200 4120 1204
rect 4160 1396 4200 1400
rect 4160 1364 4164 1396
rect 4196 1364 4200 1396
rect 4160 1236 4200 1364
rect 4160 1204 4164 1236
rect 4196 1204 4200 1236
rect 4160 1200 4200 1204
rect 80 635 120 640
rect 80 605 85 635
rect 115 605 120 635
rect 80 556 120 605
rect 80 524 84 556
rect 116 524 120 556
rect 80 476 120 524
rect 80 444 84 476
rect 116 444 120 476
rect 80 396 120 444
rect 80 364 84 396
rect 116 364 120 396
rect 80 315 120 364
rect 80 285 85 315
rect 115 285 120 315
rect 80 280 120 285
rect 160 635 200 640
rect 160 605 165 635
rect 195 605 200 635
rect 160 556 200 605
rect 160 524 164 556
rect 196 524 200 556
rect 160 476 200 524
rect 160 444 164 476
rect 196 444 200 476
rect 160 396 200 444
rect 160 364 164 396
rect 196 364 200 396
rect 160 315 200 364
rect 160 285 165 315
rect 195 285 200 315
rect 160 280 200 285
rect 240 635 280 640
rect 240 605 245 635
rect 275 605 280 635
rect 240 556 280 605
rect 240 524 244 556
rect 276 524 280 556
rect 240 476 280 524
rect 240 444 244 476
rect 276 444 280 476
rect 240 396 280 444
rect 240 364 244 396
rect 276 364 280 396
rect 240 315 280 364
rect 240 285 245 315
rect 275 285 280 315
rect 240 280 280 285
rect 320 635 360 640
rect 320 605 325 635
rect 355 605 360 635
rect 320 556 360 605
rect 320 524 324 556
rect 356 524 360 556
rect 320 476 360 524
rect 320 444 324 476
rect 356 444 360 476
rect 320 396 360 444
rect 320 364 324 396
rect 356 364 360 396
rect 320 315 360 364
rect 320 285 325 315
rect 355 285 360 315
rect 320 280 360 285
rect 400 635 440 640
rect 400 605 405 635
rect 435 605 440 635
rect 400 556 440 605
rect 400 524 404 556
rect 436 524 440 556
rect 400 476 440 524
rect 400 444 404 476
rect 436 444 440 476
rect 400 396 440 444
rect 400 364 404 396
rect 436 364 440 396
rect 400 315 440 364
rect 400 285 405 315
rect 435 285 440 315
rect 400 280 440 285
rect 480 635 520 640
rect 480 605 485 635
rect 515 605 520 635
rect 480 556 520 605
rect 480 524 484 556
rect 516 524 520 556
rect 480 476 520 524
rect 480 444 484 476
rect 516 444 520 476
rect 480 396 520 444
rect 480 364 484 396
rect 516 364 520 396
rect 480 315 520 364
rect 480 285 485 315
rect 515 285 520 315
rect 480 280 520 285
rect 560 635 600 640
rect 560 605 565 635
rect 595 605 600 635
rect 560 556 600 605
rect 560 524 564 556
rect 596 524 600 556
rect 560 476 600 524
rect 560 444 564 476
rect 596 444 600 476
rect 560 396 600 444
rect 560 364 564 396
rect 596 364 600 396
rect 560 315 600 364
rect 560 285 565 315
rect 595 285 600 315
rect 560 280 600 285
rect 720 635 760 640
rect 720 605 725 635
rect 755 605 760 635
rect 720 556 760 605
rect 720 524 724 556
rect 756 524 760 556
rect 720 476 760 524
rect 720 444 724 476
rect 756 444 760 476
rect 720 396 760 444
rect 720 364 724 396
rect 756 364 760 396
rect 720 315 760 364
rect 720 285 725 315
rect 755 285 760 315
rect 720 280 760 285
rect 800 635 840 640
rect 800 605 805 635
rect 835 605 840 635
rect 800 556 840 605
rect 800 524 804 556
rect 836 524 840 556
rect 800 476 840 524
rect 800 444 804 476
rect 836 444 840 476
rect 800 396 840 444
rect 800 364 804 396
rect 836 364 840 396
rect 800 315 840 364
rect 800 285 805 315
rect 835 285 840 315
rect 800 280 840 285
rect 880 635 920 640
rect 880 605 885 635
rect 915 605 920 635
rect 880 556 920 605
rect 880 524 884 556
rect 916 524 920 556
rect 880 476 920 524
rect 880 444 884 476
rect 916 444 920 476
rect 880 396 920 444
rect 880 364 884 396
rect 916 364 920 396
rect 880 315 920 364
rect 880 285 885 315
rect 915 285 920 315
rect 880 280 920 285
rect 960 635 1000 640
rect 960 605 965 635
rect 995 605 1000 635
rect 960 556 1000 605
rect 960 524 964 556
rect 996 524 1000 556
rect 960 476 1000 524
rect 960 444 964 476
rect 996 444 1000 476
rect 960 396 1000 444
rect 960 364 964 396
rect 996 364 1000 396
rect 960 315 1000 364
rect 960 285 965 315
rect 995 285 1000 315
rect 960 280 1000 285
rect 1040 635 1080 640
rect 1040 605 1045 635
rect 1075 605 1080 635
rect 1040 556 1080 605
rect 1040 524 1044 556
rect 1076 524 1080 556
rect 1040 476 1080 524
rect 1040 444 1044 476
rect 1076 444 1080 476
rect 1040 396 1080 444
rect 1040 364 1044 396
rect 1076 364 1080 396
rect 1040 315 1080 364
rect 1040 285 1045 315
rect 1075 285 1080 315
rect 1040 280 1080 285
rect 1120 635 1160 640
rect 1120 605 1125 635
rect 1155 605 1160 635
rect 1120 556 1160 605
rect 1120 524 1124 556
rect 1156 524 1160 556
rect 1120 476 1160 524
rect 1120 444 1124 476
rect 1156 444 1160 476
rect 1120 396 1160 444
rect 1120 364 1124 396
rect 1156 364 1160 396
rect 1120 315 1160 364
rect 1120 285 1125 315
rect 1155 285 1160 315
rect 1120 280 1160 285
rect 1200 635 1240 640
rect 1200 605 1205 635
rect 1235 605 1240 635
rect 1200 556 1240 605
rect 1200 524 1204 556
rect 1236 524 1240 556
rect 1200 476 1240 524
rect 1200 444 1204 476
rect 1236 444 1240 476
rect 1200 396 1240 444
rect 1200 364 1204 396
rect 1236 364 1240 396
rect 1200 315 1240 364
rect 1200 285 1205 315
rect 1235 285 1240 315
rect 1200 280 1240 285
rect 1280 635 1320 640
rect 1280 605 1285 635
rect 1315 605 1320 635
rect 1280 556 1320 605
rect 1280 524 1284 556
rect 1316 524 1320 556
rect 1280 476 1320 524
rect 1280 444 1284 476
rect 1316 444 1320 476
rect 1280 396 1320 444
rect 1280 364 1284 396
rect 1316 364 1320 396
rect 1280 315 1320 364
rect 1280 285 1285 315
rect 1315 285 1320 315
rect 1280 280 1320 285
rect 1360 635 1400 640
rect 1360 605 1365 635
rect 1395 605 1400 635
rect 1360 556 1400 605
rect 1360 524 1364 556
rect 1396 524 1400 556
rect 1360 476 1400 524
rect 1360 444 1364 476
rect 1396 444 1400 476
rect 1360 396 1400 444
rect 1360 364 1364 396
rect 1396 364 1400 396
rect 1360 315 1400 364
rect 1360 285 1365 315
rect 1395 285 1400 315
rect 1360 280 1400 285
rect 1440 635 1480 640
rect 1440 605 1445 635
rect 1475 605 1480 635
rect 1440 556 1480 605
rect 1440 524 1444 556
rect 1476 524 1480 556
rect 1440 476 1480 524
rect 1440 444 1444 476
rect 1476 444 1480 476
rect 1440 396 1480 444
rect 1440 364 1444 396
rect 1476 364 1480 396
rect 1440 315 1480 364
rect 1440 285 1445 315
rect 1475 285 1480 315
rect 1440 280 1480 285
rect 1520 635 1560 640
rect 1520 605 1525 635
rect 1555 605 1560 635
rect 1520 556 1560 605
rect 1520 524 1524 556
rect 1556 524 1560 556
rect 1520 476 1560 524
rect 1520 444 1524 476
rect 1556 444 1560 476
rect 1520 396 1560 444
rect 1520 364 1524 396
rect 1556 364 1560 396
rect 1520 315 1560 364
rect 1520 285 1525 315
rect 1555 285 1560 315
rect 1520 280 1560 285
rect 1680 635 1720 640
rect 1680 605 1685 635
rect 1715 605 1720 635
rect 1680 556 1720 605
rect 1680 524 1684 556
rect 1716 524 1720 556
rect 1680 476 1720 524
rect 1680 444 1684 476
rect 1716 444 1720 476
rect 1680 396 1720 444
rect 1680 364 1684 396
rect 1716 364 1720 396
rect 1680 315 1720 364
rect 1680 285 1685 315
rect 1715 285 1720 315
rect 1680 280 1720 285
rect 1760 635 1800 640
rect 1760 605 1765 635
rect 1795 605 1800 635
rect 1760 556 1800 605
rect 1760 524 1764 556
rect 1796 524 1800 556
rect 1760 476 1800 524
rect 1760 444 1764 476
rect 1796 444 1800 476
rect 1760 396 1800 444
rect 1760 364 1764 396
rect 1796 364 1800 396
rect 1760 315 1800 364
rect 1760 285 1765 315
rect 1795 285 1800 315
rect 1760 280 1800 285
rect 1840 635 1880 640
rect 1840 605 1845 635
rect 1875 605 1880 635
rect 1840 556 1880 605
rect 1840 524 1844 556
rect 1876 524 1880 556
rect 1840 476 1880 524
rect 1840 444 1844 476
rect 1876 444 1880 476
rect 1840 396 1880 444
rect 1840 364 1844 396
rect 1876 364 1880 396
rect 1840 315 1880 364
rect 1840 285 1845 315
rect 1875 285 1880 315
rect 1840 280 1880 285
rect 1920 635 1960 640
rect 1920 605 1925 635
rect 1955 605 1960 635
rect 1920 556 1960 605
rect 1920 524 1924 556
rect 1956 524 1960 556
rect 1920 476 1960 524
rect 1920 444 1924 476
rect 1956 444 1960 476
rect 1920 396 1960 444
rect 1920 364 1924 396
rect 1956 364 1960 396
rect 1920 315 1960 364
rect 1920 285 1925 315
rect 1955 285 1960 315
rect 1920 280 1960 285
rect 2000 635 2040 640
rect 2000 605 2005 635
rect 2035 605 2040 635
rect 2000 556 2040 605
rect 2000 524 2004 556
rect 2036 524 2040 556
rect 2000 476 2040 524
rect 2000 444 2004 476
rect 2036 444 2040 476
rect 2000 396 2040 444
rect 2000 364 2004 396
rect 2036 364 2040 396
rect 2000 315 2040 364
rect 2000 285 2005 315
rect 2035 285 2040 315
rect 2000 280 2040 285
rect 2160 635 2200 640
rect 2160 605 2165 635
rect 2195 605 2200 635
rect 2160 556 2200 605
rect 2160 524 2164 556
rect 2196 524 2200 556
rect 2160 476 2200 524
rect 2160 444 2164 476
rect 2196 444 2200 476
rect 2160 396 2200 444
rect 2160 364 2164 396
rect 2196 364 2200 396
rect 2160 315 2200 364
rect 2160 285 2165 315
rect 2195 285 2200 315
rect 2160 280 2200 285
rect 2240 635 2280 640
rect 2240 605 2245 635
rect 2275 605 2280 635
rect 2240 556 2280 605
rect 2240 524 2244 556
rect 2276 524 2280 556
rect 2240 476 2280 524
rect 2240 444 2244 476
rect 2276 444 2280 476
rect 2240 396 2280 444
rect 2240 364 2244 396
rect 2276 364 2280 396
rect 2240 315 2280 364
rect 2240 285 2245 315
rect 2275 285 2280 315
rect 2240 280 2280 285
rect 2320 635 2360 640
rect 2320 605 2325 635
rect 2355 605 2360 635
rect 2320 556 2360 605
rect 2320 524 2324 556
rect 2356 524 2360 556
rect 2320 476 2360 524
rect 2320 444 2324 476
rect 2356 444 2360 476
rect 2320 396 2360 444
rect 2320 364 2324 396
rect 2356 364 2360 396
rect 2320 315 2360 364
rect 2320 285 2325 315
rect 2355 285 2360 315
rect 2320 280 2360 285
rect 2400 635 2440 640
rect 2400 605 2405 635
rect 2435 605 2440 635
rect 2400 556 2440 605
rect 2400 524 2404 556
rect 2436 524 2440 556
rect 2400 476 2440 524
rect 2400 444 2404 476
rect 2436 444 2440 476
rect 2400 396 2440 444
rect 2400 364 2404 396
rect 2436 364 2440 396
rect 2400 315 2440 364
rect 2400 285 2405 315
rect 2435 285 2440 315
rect 2400 280 2440 285
rect 2480 635 2520 640
rect 2480 605 2485 635
rect 2515 605 2520 635
rect 2480 556 2520 605
rect 2480 524 2484 556
rect 2516 524 2520 556
rect 2480 476 2520 524
rect 2480 444 2484 476
rect 2516 444 2520 476
rect 2480 396 2520 444
rect 2480 364 2484 396
rect 2516 364 2520 396
rect 2480 315 2520 364
rect 2480 285 2485 315
rect 2515 285 2520 315
rect 2480 280 2520 285
rect 2640 635 2680 640
rect 2640 605 2645 635
rect 2675 605 2680 635
rect 2640 556 2680 605
rect 2640 524 2644 556
rect 2676 524 2680 556
rect 2640 476 2680 524
rect 2640 444 2644 476
rect 2676 444 2680 476
rect 2640 396 2680 444
rect 2640 364 2644 396
rect 2676 364 2680 396
rect 2640 315 2680 364
rect 2640 285 2645 315
rect 2675 285 2680 315
rect 2640 280 2680 285
rect 2720 635 2760 640
rect 2720 605 2725 635
rect 2755 605 2760 635
rect 2720 556 2760 605
rect 2720 524 2724 556
rect 2756 524 2760 556
rect 2720 476 2760 524
rect 2720 444 2724 476
rect 2756 444 2760 476
rect 2720 396 2760 444
rect 2720 364 2724 396
rect 2756 364 2760 396
rect 2720 315 2760 364
rect 2720 285 2725 315
rect 2755 285 2760 315
rect 2720 280 2760 285
rect 2800 635 2840 640
rect 2800 605 2805 635
rect 2835 605 2840 635
rect 2800 556 2840 605
rect 2800 524 2804 556
rect 2836 524 2840 556
rect 2800 476 2840 524
rect 2800 444 2804 476
rect 2836 444 2840 476
rect 2800 396 2840 444
rect 2800 364 2804 396
rect 2836 364 2840 396
rect 2800 315 2840 364
rect 2800 285 2805 315
rect 2835 285 2840 315
rect 2800 280 2840 285
rect 2880 635 2920 640
rect 2880 605 2885 635
rect 2915 605 2920 635
rect 2880 556 2920 605
rect 2880 524 2884 556
rect 2916 524 2920 556
rect 2880 476 2920 524
rect 2880 444 2884 476
rect 2916 444 2920 476
rect 2880 396 2920 444
rect 2880 364 2884 396
rect 2916 364 2920 396
rect 2880 315 2920 364
rect 2880 285 2885 315
rect 2915 285 2920 315
rect 2880 280 2920 285
rect 2960 635 3000 640
rect 2960 605 2965 635
rect 2995 605 3000 635
rect 2960 556 3000 605
rect 2960 524 2964 556
rect 2996 524 3000 556
rect 2960 476 3000 524
rect 2960 444 2964 476
rect 2996 444 3000 476
rect 2960 396 3000 444
rect 2960 364 2964 396
rect 2996 364 3000 396
rect 2960 315 3000 364
rect 2960 285 2965 315
rect 2995 285 3000 315
rect 2960 280 3000 285
rect 3040 635 3080 640
rect 3040 605 3045 635
rect 3075 605 3080 635
rect 3040 556 3080 605
rect 3040 524 3044 556
rect 3076 524 3080 556
rect 3040 476 3080 524
rect 3040 444 3044 476
rect 3076 444 3080 476
rect 3040 396 3080 444
rect 3040 364 3044 396
rect 3076 364 3080 396
rect 3040 315 3080 364
rect 3040 285 3045 315
rect 3075 285 3080 315
rect 3040 280 3080 285
rect 3120 635 3160 640
rect 3120 605 3125 635
rect 3155 605 3160 635
rect 3120 556 3160 605
rect 3120 524 3124 556
rect 3156 524 3160 556
rect 3120 476 3160 524
rect 3120 444 3124 476
rect 3156 444 3160 476
rect 3120 396 3160 444
rect 3120 364 3124 396
rect 3156 364 3160 396
rect 3120 315 3160 364
rect 3120 285 3125 315
rect 3155 285 3160 315
rect 3120 280 3160 285
rect 3200 635 3240 640
rect 3200 605 3205 635
rect 3235 605 3240 635
rect 3200 556 3240 605
rect 3200 524 3204 556
rect 3236 524 3240 556
rect 3200 476 3240 524
rect 3200 444 3204 476
rect 3236 444 3240 476
rect 3200 396 3240 444
rect 3200 364 3204 396
rect 3236 364 3240 396
rect 3200 315 3240 364
rect 3200 285 3205 315
rect 3235 285 3240 315
rect 3200 280 3240 285
rect 3280 635 3320 640
rect 3280 605 3285 635
rect 3315 605 3320 635
rect 3280 556 3320 605
rect 3280 524 3284 556
rect 3316 524 3320 556
rect 3280 476 3320 524
rect 3280 444 3284 476
rect 3316 444 3320 476
rect 3280 396 3320 444
rect 3280 364 3284 396
rect 3316 364 3320 396
rect 3280 315 3320 364
rect 3280 285 3285 315
rect 3315 285 3320 315
rect 3280 280 3320 285
rect 3360 635 3400 640
rect 3360 605 3365 635
rect 3395 605 3400 635
rect 3360 556 3400 605
rect 3360 524 3364 556
rect 3396 524 3400 556
rect 3360 476 3400 524
rect 3360 444 3364 476
rect 3396 444 3400 476
rect 3360 396 3400 444
rect 3360 364 3364 396
rect 3396 364 3400 396
rect 3360 315 3400 364
rect 3360 285 3365 315
rect 3395 285 3400 315
rect 3360 280 3400 285
rect 3440 635 3480 640
rect 3440 605 3445 635
rect 3475 605 3480 635
rect 3440 556 3480 605
rect 3440 524 3444 556
rect 3476 524 3480 556
rect 3440 476 3480 524
rect 3440 444 3444 476
rect 3476 444 3480 476
rect 3440 396 3480 444
rect 3440 364 3444 396
rect 3476 364 3480 396
rect 3440 315 3480 364
rect 3440 285 3445 315
rect 3475 285 3480 315
rect 3440 280 3480 285
rect 3600 635 3640 640
rect 3600 605 3605 635
rect 3635 605 3640 635
rect 3600 556 3640 605
rect 3600 524 3604 556
rect 3636 524 3640 556
rect 3600 476 3640 524
rect 3600 444 3604 476
rect 3636 444 3640 476
rect 3600 396 3640 444
rect 3600 364 3604 396
rect 3636 364 3640 396
rect 3600 315 3640 364
rect 3600 285 3605 315
rect 3635 285 3640 315
rect 3600 280 3640 285
rect 3680 635 3720 640
rect 3680 605 3685 635
rect 3715 605 3720 635
rect 3680 556 3720 605
rect 3680 524 3684 556
rect 3716 524 3720 556
rect 3680 476 3720 524
rect 3680 444 3684 476
rect 3716 444 3720 476
rect 3680 396 3720 444
rect 3680 364 3684 396
rect 3716 364 3720 396
rect 3680 315 3720 364
rect 3680 285 3685 315
rect 3715 285 3720 315
rect 3680 280 3720 285
rect 3760 635 3800 640
rect 3760 605 3765 635
rect 3795 605 3800 635
rect 3760 556 3800 605
rect 3760 524 3764 556
rect 3796 524 3800 556
rect 3760 476 3800 524
rect 3760 444 3764 476
rect 3796 444 3800 476
rect 3760 396 3800 444
rect 3760 364 3764 396
rect 3796 364 3800 396
rect 3760 315 3800 364
rect 3760 285 3765 315
rect 3795 285 3800 315
rect 3760 280 3800 285
rect 3840 635 3880 640
rect 3840 605 3845 635
rect 3875 605 3880 635
rect 3840 556 3880 605
rect 3840 524 3844 556
rect 3876 524 3880 556
rect 3840 476 3880 524
rect 3840 444 3844 476
rect 3876 444 3880 476
rect 3840 396 3880 444
rect 3840 364 3844 396
rect 3876 364 3880 396
rect 3840 315 3880 364
rect 3840 285 3845 315
rect 3875 285 3880 315
rect 3840 280 3880 285
rect 3920 635 3960 640
rect 3920 605 3925 635
rect 3955 605 3960 635
rect 3920 556 3960 605
rect 3920 524 3924 556
rect 3956 524 3960 556
rect 3920 476 3960 524
rect 3920 444 3924 476
rect 3956 444 3960 476
rect 3920 396 3960 444
rect 3920 364 3924 396
rect 3956 364 3960 396
rect 3920 315 3960 364
rect 3920 285 3925 315
rect 3955 285 3960 315
rect 3920 280 3960 285
rect 4000 635 4040 640
rect 4000 605 4005 635
rect 4035 605 4040 635
rect 4000 556 4040 605
rect 4000 524 4004 556
rect 4036 524 4040 556
rect 4000 476 4040 524
rect 4000 444 4004 476
rect 4036 444 4040 476
rect 4000 396 4040 444
rect 4000 364 4004 396
rect 4036 364 4040 396
rect 4000 315 4040 364
rect 4000 285 4005 315
rect 4035 285 4040 315
rect 4000 280 4040 285
rect 4080 635 4120 640
rect 4080 605 4085 635
rect 4115 605 4120 635
rect 4080 556 4120 605
rect 4080 524 4084 556
rect 4116 524 4120 556
rect 4080 476 4120 524
rect 4080 444 4084 476
rect 4116 444 4120 476
rect 4080 396 4120 444
rect 4080 364 4084 396
rect 4116 364 4120 396
rect 4080 315 4120 364
rect 4080 285 4085 315
rect 4115 285 4120 315
rect 4080 280 4120 285
rect 160 171 200 180
rect 160 89 164 171
rect 196 89 200 171
rect 160 80 200 89
rect 4000 171 4040 180
rect 4000 89 4004 171
rect 4036 89 4040 171
rect 4000 80 4040 89
<< via3 >>
rect 2084 1830 2116 1831
rect 2084 1650 2085 1830
rect 2085 1650 2115 1830
rect 2115 1650 2116 1830
rect 2084 1649 2116 1650
rect 4 1395 36 1396
rect 4 1365 5 1395
rect 5 1365 35 1395
rect 35 1365 36 1395
rect 4 1364 36 1365
rect 4 1235 36 1236
rect 4 1205 5 1235
rect 5 1205 35 1235
rect 35 1205 36 1235
rect 4 1204 36 1205
rect 84 1395 116 1396
rect 84 1365 85 1395
rect 85 1365 115 1395
rect 115 1365 116 1395
rect 84 1364 116 1365
rect 84 1235 116 1236
rect 84 1205 85 1235
rect 85 1205 115 1235
rect 115 1205 116 1235
rect 84 1204 116 1205
rect 164 1395 196 1396
rect 164 1365 165 1395
rect 165 1365 195 1395
rect 195 1365 196 1395
rect 164 1364 196 1365
rect 164 1235 196 1236
rect 164 1205 165 1235
rect 165 1205 195 1235
rect 195 1205 196 1235
rect 164 1204 196 1205
rect 244 1395 276 1396
rect 244 1365 245 1395
rect 245 1365 275 1395
rect 275 1365 276 1395
rect 244 1364 276 1365
rect 244 1235 276 1236
rect 244 1205 245 1235
rect 245 1205 275 1235
rect 275 1205 276 1235
rect 244 1204 276 1205
rect 324 1395 356 1396
rect 324 1365 325 1395
rect 325 1365 355 1395
rect 355 1365 356 1395
rect 324 1364 356 1365
rect 324 1235 356 1236
rect 324 1205 325 1235
rect 325 1205 355 1235
rect 355 1205 356 1235
rect 324 1204 356 1205
rect 404 1395 436 1396
rect 404 1365 405 1395
rect 405 1365 435 1395
rect 435 1365 436 1395
rect 404 1364 436 1365
rect 404 1235 436 1236
rect 404 1205 405 1235
rect 405 1205 435 1235
rect 435 1205 436 1235
rect 404 1204 436 1205
rect 484 1395 516 1396
rect 484 1365 485 1395
rect 485 1365 515 1395
rect 515 1365 516 1395
rect 484 1364 516 1365
rect 484 1235 516 1236
rect 484 1205 485 1235
rect 485 1205 515 1235
rect 515 1205 516 1235
rect 484 1204 516 1205
rect 564 1395 596 1396
rect 564 1365 565 1395
rect 565 1365 595 1395
rect 595 1365 596 1395
rect 564 1364 596 1365
rect 564 1235 596 1236
rect 564 1205 565 1235
rect 565 1205 595 1235
rect 595 1205 596 1235
rect 564 1204 596 1205
rect 724 1395 756 1396
rect 724 1365 725 1395
rect 725 1365 755 1395
rect 755 1365 756 1395
rect 724 1364 756 1365
rect 724 1235 756 1236
rect 724 1205 725 1235
rect 725 1205 755 1235
rect 755 1205 756 1235
rect 724 1204 756 1205
rect 804 1395 836 1396
rect 804 1365 805 1395
rect 805 1365 835 1395
rect 835 1365 836 1395
rect 804 1364 836 1365
rect 804 1235 836 1236
rect 804 1205 805 1235
rect 805 1205 835 1235
rect 835 1205 836 1235
rect 804 1204 836 1205
rect 884 1395 916 1396
rect 884 1365 885 1395
rect 885 1365 915 1395
rect 915 1365 916 1395
rect 884 1364 916 1365
rect 884 1235 916 1236
rect 884 1205 885 1235
rect 885 1205 915 1235
rect 915 1205 916 1235
rect 884 1204 916 1205
rect 964 1395 996 1396
rect 964 1365 965 1395
rect 965 1365 995 1395
rect 995 1365 996 1395
rect 964 1364 996 1365
rect 964 1235 996 1236
rect 964 1205 965 1235
rect 965 1205 995 1235
rect 995 1205 996 1235
rect 964 1204 996 1205
rect 1044 1395 1076 1396
rect 1044 1365 1045 1395
rect 1045 1365 1075 1395
rect 1075 1365 1076 1395
rect 1044 1364 1076 1365
rect 1044 1235 1076 1236
rect 1044 1205 1045 1235
rect 1045 1205 1075 1235
rect 1075 1205 1076 1235
rect 1044 1204 1076 1205
rect 1124 1395 1156 1396
rect 1124 1365 1125 1395
rect 1125 1365 1155 1395
rect 1155 1365 1156 1395
rect 1124 1364 1156 1365
rect 1124 1235 1156 1236
rect 1124 1205 1125 1235
rect 1125 1205 1155 1235
rect 1155 1205 1156 1235
rect 1124 1204 1156 1205
rect 1204 1395 1236 1396
rect 1204 1365 1205 1395
rect 1205 1365 1235 1395
rect 1235 1365 1236 1395
rect 1204 1364 1236 1365
rect 1204 1235 1236 1236
rect 1204 1205 1205 1235
rect 1205 1205 1235 1235
rect 1235 1205 1236 1235
rect 1204 1204 1236 1205
rect 1284 1395 1316 1396
rect 1284 1365 1285 1395
rect 1285 1365 1315 1395
rect 1315 1365 1316 1395
rect 1284 1364 1316 1365
rect 1284 1235 1316 1236
rect 1284 1205 1285 1235
rect 1285 1205 1315 1235
rect 1315 1205 1316 1235
rect 1284 1204 1316 1205
rect 1364 1395 1396 1396
rect 1364 1365 1365 1395
rect 1365 1365 1395 1395
rect 1395 1365 1396 1395
rect 1364 1364 1396 1365
rect 1364 1235 1396 1236
rect 1364 1205 1365 1235
rect 1365 1205 1395 1235
rect 1395 1205 1396 1235
rect 1364 1204 1396 1205
rect 1444 1395 1476 1396
rect 1444 1365 1445 1395
rect 1445 1365 1475 1395
rect 1475 1365 1476 1395
rect 1444 1364 1476 1365
rect 1444 1235 1476 1236
rect 1444 1205 1445 1235
rect 1445 1205 1475 1235
rect 1475 1205 1476 1235
rect 1444 1204 1476 1205
rect 1524 1395 1556 1396
rect 1524 1365 1525 1395
rect 1525 1365 1555 1395
rect 1555 1365 1556 1395
rect 1524 1364 1556 1365
rect 1524 1235 1556 1236
rect 1524 1205 1525 1235
rect 1525 1205 1555 1235
rect 1555 1205 1556 1235
rect 1524 1204 1556 1205
rect 1684 1395 1716 1396
rect 1684 1365 1685 1395
rect 1685 1365 1715 1395
rect 1715 1365 1716 1395
rect 1684 1364 1716 1365
rect 1684 1235 1716 1236
rect 1684 1205 1685 1235
rect 1685 1205 1715 1235
rect 1715 1205 1716 1235
rect 1684 1204 1716 1205
rect 1764 1395 1796 1396
rect 1764 1365 1765 1395
rect 1765 1365 1795 1395
rect 1795 1365 1796 1395
rect 1764 1364 1796 1365
rect 1764 1235 1796 1236
rect 1764 1205 1765 1235
rect 1765 1205 1795 1235
rect 1795 1205 1796 1235
rect 1764 1204 1796 1205
rect 1844 1395 1876 1396
rect 1844 1365 1845 1395
rect 1845 1365 1875 1395
rect 1875 1365 1876 1395
rect 1844 1364 1876 1365
rect 1844 1235 1876 1236
rect 1844 1205 1845 1235
rect 1845 1205 1875 1235
rect 1875 1205 1876 1235
rect 1844 1204 1876 1205
rect 1924 1395 1956 1396
rect 1924 1365 1925 1395
rect 1925 1365 1955 1395
rect 1955 1365 1956 1395
rect 1924 1364 1956 1365
rect 1924 1235 1956 1236
rect 1924 1205 1925 1235
rect 1925 1205 1955 1235
rect 1955 1205 1956 1235
rect 1924 1204 1956 1205
rect 2004 1395 2036 1396
rect 2004 1365 2005 1395
rect 2005 1365 2035 1395
rect 2035 1365 2036 1395
rect 2004 1364 2036 1365
rect 2004 1235 2036 1236
rect 2004 1205 2005 1235
rect 2005 1205 2035 1235
rect 2035 1205 2036 1235
rect 2004 1204 2036 1205
rect 2084 1395 2116 1396
rect 2084 1365 2085 1395
rect 2085 1365 2115 1395
rect 2115 1365 2116 1395
rect 2084 1364 2116 1365
rect 2084 1235 2116 1236
rect 2084 1205 2085 1235
rect 2085 1205 2115 1235
rect 2115 1205 2116 1235
rect 2084 1204 2116 1205
rect 2164 1395 2196 1396
rect 2164 1365 2165 1395
rect 2165 1365 2195 1395
rect 2195 1365 2196 1395
rect 2164 1364 2196 1365
rect 2164 1235 2196 1236
rect 2164 1205 2165 1235
rect 2165 1205 2195 1235
rect 2195 1205 2196 1235
rect 2164 1204 2196 1205
rect 2244 1395 2276 1396
rect 2244 1365 2245 1395
rect 2245 1365 2275 1395
rect 2275 1365 2276 1395
rect 2244 1364 2276 1365
rect 2244 1235 2276 1236
rect 2244 1205 2245 1235
rect 2245 1205 2275 1235
rect 2275 1205 2276 1235
rect 2244 1204 2276 1205
rect 2324 1395 2356 1396
rect 2324 1365 2325 1395
rect 2325 1365 2355 1395
rect 2355 1365 2356 1395
rect 2324 1364 2356 1365
rect 2324 1235 2356 1236
rect 2324 1205 2325 1235
rect 2325 1205 2355 1235
rect 2355 1205 2356 1235
rect 2324 1204 2356 1205
rect 2404 1395 2436 1396
rect 2404 1365 2405 1395
rect 2405 1365 2435 1395
rect 2435 1365 2436 1395
rect 2404 1364 2436 1365
rect 2404 1235 2436 1236
rect 2404 1205 2405 1235
rect 2405 1205 2435 1235
rect 2435 1205 2436 1235
rect 2404 1204 2436 1205
rect 2484 1395 2516 1396
rect 2484 1365 2485 1395
rect 2485 1365 2515 1395
rect 2515 1365 2516 1395
rect 2484 1364 2516 1365
rect 2484 1235 2516 1236
rect 2484 1205 2485 1235
rect 2485 1205 2515 1235
rect 2515 1205 2516 1235
rect 2484 1204 2516 1205
rect 2644 1395 2676 1396
rect 2644 1365 2645 1395
rect 2645 1365 2675 1395
rect 2675 1365 2676 1395
rect 2644 1364 2676 1365
rect 2644 1235 2676 1236
rect 2644 1205 2645 1235
rect 2645 1205 2675 1235
rect 2675 1205 2676 1235
rect 2644 1204 2676 1205
rect 2724 1395 2756 1396
rect 2724 1365 2725 1395
rect 2725 1365 2755 1395
rect 2755 1365 2756 1395
rect 2724 1364 2756 1365
rect 2724 1235 2756 1236
rect 2724 1205 2725 1235
rect 2725 1205 2755 1235
rect 2755 1205 2756 1235
rect 2724 1204 2756 1205
rect 2804 1395 2836 1396
rect 2804 1365 2805 1395
rect 2805 1365 2835 1395
rect 2835 1365 2836 1395
rect 2804 1364 2836 1365
rect 2804 1235 2836 1236
rect 2804 1205 2805 1235
rect 2805 1205 2835 1235
rect 2835 1205 2836 1235
rect 2804 1204 2836 1205
rect 2884 1395 2916 1396
rect 2884 1365 2885 1395
rect 2885 1365 2915 1395
rect 2915 1365 2916 1395
rect 2884 1364 2916 1365
rect 2884 1235 2916 1236
rect 2884 1205 2885 1235
rect 2885 1205 2915 1235
rect 2915 1205 2916 1235
rect 2884 1204 2916 1205
rect 2964 1395 2996 1396
rect 2964 1365 2965 1395
rect 2965 1365 2995 1395
rect 2995 1365 2996 1395
rect 2964 1364 2996 1365
rect 2964 1235 2996 1236
rect 2964 1205 2965 1235
rect 2965 1205 2995 1235
rect 2995 1205 2996 1235
rect 2964 1204 2996 1205
rect 3044 1395 3076 1396
rect 3044 1365 3045 1395
rect 3045 1365 3075 1395
rect 3075 1365 3076 1395
rect 3044 1364 3076 1365
rect 3044 1235 3076 1236
rect 3044 1205 3045 1235
rect 3045 1205 3075 1235
rect 3075 1205 3076 1235
rect 3044 1204 3076 1205
rect 3124 1395 3156 1396
rect 3124 1365 3125 1395
rect 3125 1365 3155 1395
rect 3155 1365 3156 1395
rect 3124 1364 3156 1365
rect 3124 1235 3156 1236
rect 3124 1205 3125 1235
rect 3125 1205 3155 1235
rect 3155 1205 3156 1235
rect 3124 1204 3156 1205
rect 3204 1395 3236 1396
rect 3204 1365 3205 1395
rect 3205 1365 3235 1395
rect 3235 1365 3236 1395
rect 3204 1364 3236 1365
rect 3204 1235 3236 1236
rect 3204 1205 3205 1235
rect 3205 1205 3235 1235
rect 3235 1205 3236 1235
rect 3204 1204 3236 1205
rect 3284 1395 3316 1396
rect 3284 1365 3285 1395
rect 3285 1365 3315 1395
rect 3315 1365 3316 1395
rect 3284 1364 3316 1365
rect 3284 1235 3316 1236
rect 3284 1205 3285 1235
rect 3285 1205 3315 1235
rect 3315 1205 3316 1235
rect 3284 1204 3316 1205
rect 3364 1395 3396 1396
rect 3364 1365 3365 1395
rect 3365 1365 3395 1395
rect 3395 1365 3396 1395
rect 3364 1364 3396 1365
rect 3364 1235 3396 1236
rect 3364 1205 3365 1235
rect 3365 1205 3395 1235
rect 3395 1205 3396 1235
rect 3364 1204 3396 1205
rect 3444 1395 3476 1396
rect 3444 1365 3445 1395
rect 3445 1365 3475 1395
rect 3475 1365 3476 1395
rect 3444 1364 3476 1365
rect 3444 1235 3476 1236
rect 3444 1205 3445 1235
rect 3445 1205 3475 1235
rect 3475 1205 3476 1235
rect 3444 1204 3476 1205
rect 3604 1395 3636 1396
rect 3604 1365 3605 1395
rect 3605 1365 3635 1395
rect 3635 1365 3636 1395
rect 3604 1364 3636 1365
rect 3604 1235 3636 1236
rect 3604 1205 3605 1235
rect 3605 1205 3635 1235
rect 3635 1205 3636 1235
rect 3604 1204 3636 1205
rect 3684 1395 3716 1396
rect 3684 1365 3685 1395
rect 3685 1365 3715 1395
rect 3715 1365 3716 1395
rect 3684 1364 3716 1365
rect 3684 1235 3716 1236
rect 3684 1205 3685 1235
rect 3685 1205 3715 1235
rect 3715 1205 3716 1235
rect 3684 1204 3716 1205
rect 3764 1395 3796 1396
rect 3764 1365 3765 1395
rect 3765 1365 3795 1395
rect 3795 1365 3796 1395
rect 3764 1364 3796 1365
rect 3764 1235 3796 1236
rect 3764 1205 3765 1235
rect 3765 1205 3795 1235
rect 3795 1205 3796 1235
rect 3764 1204 3796 1205
rect 3844 1395 3876 1396
rect 3844 1365 3845 1395
rect 3845 1365 3875 1395
rect 3875 1365 3876 1395
rect 3844 1364 3876 1365
rect 3844 1235 3876 1236
rect 3844 1205 3845 1235
rect 3845 1205 3875 1235
rect 3875 1205 3876 1235
rect 3844 1204 3876 1205
rect 3924 1395 3956 1396
rect 3924 1365 3925 1395
rect 3925 1365 3955 1395
rect 3955 1365 3956 1395
rect 3924 1364 3956 1365
rect 3924 1235 3956 1236
rect 3924 1205 3925 1235
rect 3925 1205 3955 1235
rect 3955 1205 3956 1235
rect 3924 1204 3956 1205
rect 4004 1395 4036 1396
rect 4004 1365 4005 1395
rect 4005 1365 4035 1395
rect 4035 1365 4036 1395
rect 4004 1364 4036 1365
rect 4004 1235 4036 1236
rect 4004 1205 4005 1235
rect 4005 1205 4035 1235
rect 4035 1205 4036 1235
rect 4004 1204 4036 1205
rect 4084 1395 4116 1396
rect 4084 1365 4085 1395
rect 4085 1365 4115 1395
rect 4115 1365 4116 1395
rect 4084 1364 4116 1365
rect 4084 1235 4116 1236
rect 4084 1205 4085 1235
rect 4085 1205 4115 1235
rect 4115 1205 4116 1235
rect 4084 1204 4116 1205
rect 4164 1395 4196 1396
rect 4164 1365 4165 1395
rect 4165 1365 4195 1395
rect 4195 1365 4196 1395
rect 4164 1364 4196 1365
rect 4164 1235 4196 1236
rect 4164 1205 4165 1235
rect 4165 1205 4195 1235
rect 4195 1205 4196 1235
rect 4164 1204 4196 1205
rect 84 524 116 556
rect 84 475 116 476
rect 84 445 85 475
rect 85 445 115 475
rect 115 445 116 475
rect 84 444 116 445
rect 84 364 116 396
rect 164 524 196 556
rect 164 475 196 476
rect 164 445 165 475
rect 165 445 195 475
rect 195 445 196 475
rect 164 444 196 445
rect 164 364 196 396
rect 244 524 276 556
rect 244 475 276 476
rect 244 445 245 475
rect 245 445 275 475
rect 275 445 276 475
rect 244 444 276 445
rect 244 364 276 396
rect 324 524 356 556
rect 324 475 356 476
rect 324 445 325 475
rect 325 445 355 475
rect 355 445 356 475
rect 324 444 356 445
rect 324 364 356 396
rect 404 524 436 556
rect 404 475 436 476
rect 404 445 405 475
rect 405 445 435 475
rect 435 445 436 475
rect 404 444 436 445
rect 404 364 436 396
rect 484 524 516 556
rect 484 475 516 476
rect 484 445 485 475
rect 485 445 515 475
rect 515 445 516 475
rect 484 444 516 445
rect 484 364 516 396
rect 564 524 596 556
rect 564 475 596 476
rect 564 445 565 475
rect 565 445 595 475
rect 595 445 596 475
rect 564 444 596 445
rect 564 364 596 396
rect 724 524 756 556
rect 724 475 756 476
rect 724 445 725 475
rect 725 445 755 475
rect 755 445 756 475
rect 724 444 756 445
rect 724 364 756 396
rect 804 524 836 556
rect 804 475 836 476
rect 804 445 805 475
rect 805 445 835 475
rect 835 445 836 475
rect 804 444 836 445
rect 804 364 836 396
rect 884 524 916 556
rect 884 475 916 476
rect 884 445 885 475
rect 885 445 915 475
rect 915 445 916 475
rect 884 444 916 445
rect 884 364 916 396
rect 964 524 996 556
rect 964 475 996 476
rect 964 445 965 475
rect 965 445 995 475
rect 995 445 996 475
rect 964 444 996 445
rect 964 364 996 396
rect 1044 524 1076 556
rect 1044 475 1076 476
rect 1044 445 1045 475
rect 1045 445 1075 475
rect 1075 445 1076 475
rect 1044 444 1076 445
rect 1044 364 1076 396
rect 1124 524 1156 556
rect 1124 475 1156 476
rect 1124 445 1125 475
rect 1125 445 1155 475
rect 1155 445 1156 475
rect 1124 444 1156 445
rect 1124 364 1156 396
rect 1204 524 1236 556
rect 1204 475 1236 476
rect 1204 445 1205 475
rect 1205 445 1235 475
rect 1235 445 1236 475
rect 1204 444 1236 445
rect 1204 364 1236 396
rect 1284 524 1316 556
rect 1284 475 1316 476
rect 1284 445 1285 475
rect 1285 445 1315 475
rect 1315 445 1316 475
rect 1284 444 1316 445
rect 1284 364 1316 396
rect 1364 524 1396 556
rect 1364 475 1396 476
rect 1364 445 1365 475
rect 1365 445 1395 475
rect 1395 445 1396 475
rect 1364 444 1396 445
rect 1364 364 1396 396
rect 1444 524 1476 556
rect 1444 475 1476 476
rect 1444 445 1445 475
rect 1445 445 1475 475
rect 1475 445 1476 475
rect 1444 444 1476 445
rect 1444 364 1476 396
rect 1524 524 1556 556
rect 1524 475 1556 476
rect 1524 445 1525 475
rect 1525 445 1555 475
rect 1555 445 1556 475
rect 1524 444 1556 445
rect 1524 364 1556 396
rect 1684 524 1716 556
rect 1684 475 1716 476
rect 1684 445 1685 475
rect 1685 445 1715 475
rect 1715 445 1716 475
rect 1684 444 1716 445
rect 1684 364 1716 396
rect 1764 524 1796 556
rect 1764 475 1796 476
rect 1764 445 1765 475
rect 1765 445 1795 475
rect 1795 445 1796 475
rect 1764 444 1796 445
rect 1764 364 1796 396
rect 1844 524 1876 556
rect 1844 475 1876 476
rect 1844 445 1845 475
rect 1845 445 1875 475
rect 1875 445 1876 475
rect 1844 444 1876 445
rect 1844 364 1876 396
rect 1924 524 1956 556
rect 1924 475 1956 476
rect 1924 445 1925 475
rect 1925 445 1955 475
rect 1955 445 1956 475
rect 1924 444 1956 445
rect 1924 364 1956 396
rect 2004 524 2036 556
rect 2004 475 2036 476
rect 2004 445 2005 475
rect 2005 445 2035 475
rect 2035 445 2036 475
rect 2004 444 2036 445
rect 2004 364 2036 396
rect 2164 524 2196 556
rect 2164 475 2196 476
rect 2164 445 2165 475
rect 2165 445 2195 475
rect 2195 445 2196 475
rect 2164 444 2196 445
rect 2164 364 2196 396
rect 2244 524 2276 556
rect 2244 475 2276 476
rect 2244 445 2245 475
rect 2245 445 2275 475
rect 2275 445 2276 475
rect 2244 444 2276 445
rect 2244 364 2276 396
rect 2324 524 2356 556
rect 2324 475 2356 476
rect 2324 445 2325 475
rect 2325 445 2355 475
rect 2355 445 2356 475
rect 2324 444 2356 445
rect 2324 364 2356 396
rect 2404 524 2436 556
rect 2404 475 2436 476
rect 2404 445 2405 475
rect 2405 445 2435 475
rect 2435 445 2436 475
rect 2404 444 2436 445
rect 2404 364 2436 396
rect 2484 524 2516 556
rect 2484 475 2516 476
rect 2484 445 2485 475
rect 2485 445 2515 475
rect 2515 445 2516 475
rect 2484 444 2516 445
rect 2484 364 2516 396
rect 2644 524 2676 556
rect 2644 475 2676 476
rect 2644 445 2645 475
rect 2645 445 2675 475
rect 2675 445 2676 475
rect 2644 444 2676 445
rect 2644 364 2676 396
rect 2724 524 2756 556
rect 2724 475 2756 476
rect 2724 445 2725 475
rect 2725 445 2755 475
rect 2755 445 2756 475
rect 2724 444 2756 445
rect 2724 364 2756 396
rect 2804 524 2836 556
rect 2804 475 2836 476
rect 2804 445 2805 475
rect 2805 445 2835 475
rect 2835 445 2836 475
rect 2804 444 2836 445
rect 2804 364 2836 396
rect 2884 524 2916 556
rect 2884 475 2916 476
rect 2884 445 2885 475
rect 2885 445 2915 475
rect 2915 445 2916 475
rect 2884 444 2916 445
rect 2884 364 2916 396
rect 2964 524 2996 556
rect 2964 475 2996 476
rect 2964 445 2965 475
rect 2965 445 2995 475
rect 2995 445 2996 475
rect 2964 444 2996 445
rect 2964 364 2996 396
rect 3044 524 3076 556
rect 3044 475 3076 476
rect 3044 445 3045 475
rect 3045 445 3075 475
rect 3075 445 3076 475
rect 3044 444 3076 445
rect 3044 364 3076 396
rect 3124 524 3156 556
rect 3124 475 3156 476
rect 3124 445 3125 475
rect 3125 445 3155 475
rect 3155 445 3156 475
rect 3124 444 3156 445
rect 3124 364 3156 396
rect 3204 524 3236 556
rect 3204 475 3236 476
rect 3204 445 3205 475
rect 3205 445 3235 475
rect 3235 445 3236 475
rect 3204 444 3236 445
rect 3204 364 3236 396
rect 3284 524 3316 556
rect 3284 475 3316 476
rect 3284 445 3285 475
rect 3285 445 3315 475
rect 3315 445 3316 475
rect 3284 444 3316 445
rect 3284 364 3316 396
rect 3364 524 3396 556
rect 3364 475 3396 476
rect 3364 445 3365 475
rect 3365 445 3395 475
rect 3395 445 3396 475
rect 3364 444 3396 445
rect 3364 364 3396 396
rect 3444 524 3476 556
rect 3444 475 3476 476
rect 3444 445 3445 475
rect 3445 445 3475 475
rect 3475 445 3476 475
rect 3444 444 3476 445
rect 3444 364 3476 396
rect 3604 524 3636 556
rect 3604 475 3636 476
rect 3604 445 3605 475
rect 3605 445 3635 475
rect 3635 445 3636 475
rect 3604 444 3636 445
rect 3604 364 3636 396
rect 3684 524 3716 556
rect 3684 475 3716 476
rect 3684 445 3685 475
rect 3685 445 3715 475
rect 3715 445 3716 475
rect 3684 444 3716 445
rect 3684 364 3716 396
rect 3764 524 3796 556
rect 3764 475 3796 476
rect 3764 445 3765 475
rect 3765 445 3795 475
rect 3795 445 3796 475
rect 3764 444 3796 445
rect 3764 364 3796 396
rect 3844 524 3876 556
rect 3844 475 3876 476
rect 3844 445 3845 475
rect 3845 445 3875 475
rect 3875 445 3876 475
rect 3844 444 3876 445
rect 3844 364 3876 396
rect 3924 524 3956 556
rect 3924 475 3956 476
rect 3924 445 3925 475
rect 3925 445 3955 475
rect 3955 445 3956 475
rect 3924 444 3956 445
rect 3924 364 3956 396
rect 4004 524 4036 556
rect 4004 475 4036 476
rect 4004 445 4005 475
rect 4005 445 4035 475
rect 4035 445 4036 475
rect 4004 444 4036 445
rect 4004 364 4036 396
rect 4084 524 4116 556
rect 4084 475 4116 476
rect 4084 445 4085 475
rect 4085 445 4115 475
rect 4115 445 4116 475
rect 4084 444 4116 445
rect 4084 364 4116 396
rect 164 170 196 171
rect 164 90 165 170
rect 165 90 195 170
rect 195 90 196 170
rect 164 89 196 90
rect 4004 170 4036 171
rect 4004 90 4005 170
rect 4005 90 4035 170
rect 4035 90 4036 170
rect 4004 89 4036 90
<< metal4 >>
rect 0 1831 4200 1840
rect 0 1800 2084 1831
rect 0 1680 120 1800
rect 240 1680 2084 1800
rect 0 1649 2084 1680
rect 2116 1800 4200 1831
rect 2116 1680 3960 1800
rect 4080 1680 4200 1800
rect 2116 1649 4200 1680
rect 0 1640 4200 1649
rect 0 1396 4200 1400
rect 0 1364 4 1396
rect 36 1364 84 1396
rect 116 1364 164 1396
rect 196 1364 244 1396
rect 276 1364 324 1396
rect 356 1364 404 1396
rect 436 1364 484 1396
rect 516 1364 564 1396
rect 596 1364 724 1396
rect 756 1364 804 1396
rect 836 1364 884 1396
rect 916 1364 964 1396
rect 996 1364 1044 1396
rect 1076 1364 1124 1396
rect 1156 1364 1204 1396
rect 1236 1364 1284 1396
rect 1316 1364 1364 1396
rect 1396 1364 1444 1396
rect 1476 1364 1524 1396
rect 1556 1364 1684 1396
rect 1716 1364 1764 1396
rect 1796 1364 1844 1396
rect 1876 1364 1924 1396
rect 1956 1364 2004 1396
rect 2036 1364 2084 1396
rect 2116 1364 2164 1396
rect 2196 1364 2244 1396
rect 2276 1364 2324 1396
rect 2356 1364 2404 1396
rect 2436 1364 2484 1396
rect 2516 1364 2644 1396
rect 2676 1364 2724 1396
rect 2756 1364 2804 1396
rect 2836 1364 2884 1396
rect 2916 1364 2964 1396
rect 2996 1364 3044 1396
rect 3076 1364 3124 1396
rect 3156 1364 3204 1396
rect 3236 1364 3284 1396
rect 3316 1364 3364 1396
rect 3396 1364 3444 1396
rect 3476 1364 3604 1396
rect 3636 1364 3684 1396
rect 3716 1364 3764 1396
rect 3796 1364 3844 1396
rect 3876 1364 3924 1396
rect 3956 1364 4004 1396
rect 4036 1364 4084 1396
rect 4116 1364 4164 1396
rect 4196 1364 4200 1396
rect 0 1360 4200 1364
rect 0 1240 600 1360
rect 720 1240 3480 1360
rect 3600 1240 4200 1360
rect 0 1236 4200 1240
rect 0 1204 4 1236
rect 36 1204 84 1236
rect 116 1204 164 1236
rect 196 1204 244 1236
rect 276 1204 324 1236
rect 356 1204 404 1236
rect 436 1204 484 1236
rect 516 1204 564 1236
rect 596 1204 724 1236
rect 756 1204 804 1236
rect 836 1204 884 1236
rect 916 1204 964 1236
rect 996 1204 1044 1236
rect 1076 1204 1124 1236
rect 1156 1204 1204 1236
rect 1236 1204 1284 1236
rect 1316 1204 1364 1236
rect 1396 1204 1444 1236
rect 1476 1204 1524 1236
rect 1556 1204 1684 1236
rect 1716 1204 1764 1236
rect 1796 1204 1844 1236
rect 1876 1204 1924 1236
rect 1956 1204 2004 1236
rect 2036 1204 2084 1236
rect 2116 1204 2164 1236
rect 2196 1204 2244 1236
rect 2276 1204 2324 1236
rect 2356 1204 2404 1236
rect 2436 1204 2484 1236
rect 2516 1204 2644 1236
rect 2676 1204 2724 1236
rect 2756 1204 2804 1236
rect 2836 1204 2884 1236
rect 2916 1204 2964 1236
rect 2996 1204 3044 1236
rect 3076 1204 3124 1236
rect 3156 1204 3204 1236
rect 3236 1204 3284 1236
rect 3316 1204 3364 1236
rect 3396 1204 3444 1236
rect 3476 1204 3604 1236
rect 3636 1204 3684 1236
rect 3716 1204 3764 1236
rect 3796 1204 3844 1236
rect 3876 1204 3924 1236
rect 3956 1204 4004 1236
rect 4036 1204 4084 1236
rect 4116 1204 4164 1236
rect 4196 1204 4200 1236
rect 0 1200 4200 1204
rect 0 556 4200 560
rect 0 524 84 556
rect 116 524 164 556
rect 196 524 244 556
rect 276 524 324 556
rect 356 524 404 556
rect 436 524 484 556
rect 516 524 564 556
rect 596 524 724 556
rect 756 524 804 556
rect 836 524 884 556
rect 916 524 964 556
rect 996 524 1044 556
rect 1076 524 1124 556
rect 1156 524 1204 556
rect 1236 524 1284 556
rect 1316 524 1364 556
rect 1396 524 1444 556
rect 1476 524 1524 556
rect 1556 524 1684 556
rect 1716 524 1764 556
rect 1796 524 1844 556
rect 1876 524 1924 556
rect 1956 524 2004 556
rect 2036 524 2164 556
rect 2196 524 2244 556
rect 2276 524 2324 556
rect 2356 524 2404 556
rect 2436 524 2484 556
rect 2516 524 2644 556
rect 2676 524 2724 556
rect 2756 524 2804 556
rect 2836 524 2884 556
rect 2916 524 2964 556
rect 2996 524 3044 556
rect 3076 524 3124 556
rect 3156 524 3204 556
rect 3236 524 3284 556
rect 3316 524 3364 556
rect 3396 524 3444 556
rect 3476 524 3604 556
rect 3636 524 3684 556
rect 3716 524 3764 556
rect 3796 524 3844 556
rect 3876 524 3924 556
rect 3956 524 4004 556
rect 4036 524 4084 556
rect 4116 524 4200 556
rect 0 520 4200 524
rect 0 476 1080 520
rect 1200 476 2040 520
rect 0 444 84 476
rect 116 444 164 476
rect 196 444 244 476
rect 276 444 324 476
rect 356 444 404 476
rect 436 444 484 476
rect 516 444 564 476
rect 596 444 724 476
rect 756 444 804 476
rect 836 444 884 476
rect 916 444 964 476
rect 996 444 1044 476
rect 1076 444 1080 476
rect 1200 444 1204 476
rect 1236 444 1284 476
rect 1316 444 1364 476
rect 1396 444 1444 476
rect 1476 444 1524 476
rect 1556 444 1684 476
rect 1716 444 1764 476
rect 1796 444 1844 476
rect 1876 444 1924 476
rect 1956 444 2004 476
rect 2036 444 2040 476
rect 0 400 1080 444
rect 1200 400 2040 444
rect 2160 476 3000 520
rect 3120 476 4200 520
rect 2160 444 2164 476
rect 2196 444 2244 476
rect 2276 444 2324 476
rect 2356 444 2404 476
rect 2436 444 2484 476
rect 2516 444 2644 476
rect 2676 444 2724 476
rect 2756 444 2804 476
rect 2836 444 2884 476
rect 2916 444 2964 476
rect 2996 444 3000 476
rect 3120 444 3124 476
rect 3156 444 3204 476
rect 3236 444 3284 476
rect 3316 444 3364 476
rect 3396 444 3444 476
rect 3476 444 3604 476
rect 3636 444 3684 476
rect 3716 444 3764 476
rect 3796 444 3844 476
rect 3876 444 3924 476
rect 3956 444 4004 476
rect 4036 444 4084 476
rect 4116 444 4200 476
rect 2160 400 3000 444
rect 3120 400 4200 444
rect 0 396 4200 400
rect 0 364 84 396
rect 116 364 164 396
rect 196 364 244 396
rect 276 364 324 396
rect 356 364 404 396
rect 436 364 484 396
rect 516 364 564 396
rect 596 364 724 396
rect 756 364 804 396
rect 836 364 884 396
rect 916 364 964 396
rect 996 364 1044 396
rect 1076 364 1124 396
rect 1156 364 1204 396
rect 1236 364 1284 396
rect 1316 364 1364 396
rect 1396 364 1444 396
rect 1476 364 1524 396
rect 1556 364 1684 396
rect 1716 364 1764 396
rect 1796 364 1844 396
rect 1876 364 1924 396
rect 1956 364 2004 396
rect 2036 364 2164 396
rect 2196 364 2244 396
rect 2276 364 2324 396
rect 2356 364 2404 396
rect 2436 364 2484 396
rect 2516 364 2644 396
rect 2676 364 2724 396
rect 2756 364 2804 396
rect 2836 364 2884 396
rect 2916 364 2964 396
rect 2996 364 3044 396
rect 3076 364 3124 396
rect 3156 364 3204 396
rect 3236 364 3284 396
rect 3316 364 3364 396
rect 3396 364 3444 396
rect 3476 364 3604 396
rect 3636 364 3684 396
rect 3716 364 3764 396
rect 3796 364 3844 396
rect 3876 364 3924 396
rect 3956 364 4004 396
rect 4036 364 4084 396
rect 4116 364 4200 396
rect 0 360 4200 364
rect 0 171 4200 200
rect 0 89 164 171
rect 196 160 4004 171
rect 196 89 1560 160
rect 0 40 1560 89
rect 1680 40 2520 160
rect 2640 89 4004 160
rect 4036 89 4200 171
rect 2640 40 4200 89
rect 0 0 4200 40
<< via4 >>
rect 120 1680 240 1800
rect 3960 1680 4080 1800
rect 600 1240 720 1360
rect 3480 1240 3600 1360
rect 1080 476 1200 520
rect 1080 444 1124 476
rect 1124 444 1156 476
rect 1156 444 1200 476
rect 1080 400 1200 444
rect 2040 400 2160 520
rect 3000 476 3120 520
rect 3000 444 3044 476
rect 3044 444 3076 476
rect 3076 444 3120 476
rect 3000 400 3120 444
rect 1560 40 1680 160
rect 2520 40 2640 160
<< metal5 >>
rect 80 1800 280 2000
rect 80 1680 120 1800
rect 240 1680 280 1800
rect 80 0 280 1680
rect 560 1360 760 2000
rect 560 1240 600 1360
rect 720 1240 760 1360
rect 560 0 760 1240
rect 1040 520 1240 2000
rect 1040 400 1080 520
rect 1200 400 1240 520
rect 1040 0 1240 400
rect 1520 160 1720 2000
rect 1520 40 1560 160
rect 1680 40 1720 160
rect 1520 0 1720 40
rect 2000 520 2200 2000
rect 2000 400 2040 520
rect 2160 400 2200 520
rect 2000 0 2200 400
rect 2480 160 2680 2000
rect 2480 40 2520 160
rect 2640 40 2680 160
rect 2480 0 2680 40
rect 2960 520 3160 2000
rect 2960 400 3000 520
rect 3120 400 3160 520
rect 2960 0 3160 400
rect 3440 1360 3640 2000
rect 3440 1240 3480 1360
rect 3600 1240 3640 1360
rect 3440 0 3640 1240
rect 3920 1800 4120 2000
rect 3920 1680 3960 1800
rect 4080 1680 4120 1800
rect 3920 0 4120 1680
<< labels >>
rlabel metal2 0 520 4200 560 0 in
port 1 nsew
rlabel metal2 0 360 4200 400 0 out
port 2 nsew
rlabel metal5 80 0 280 2000 0 vdda
port 3 nsew
rlabel metal2 0 1280 4200 1320 0 bp
port 4 nsew
rlabel metal5 560 0 760 2000 0 vddx
port 5 nsew
rlabel metal5 1040 0 1240 2000 0 gnda
port 6 nsew
rlabel metal5 1520 0 1720 2000 0 vssa
port 7 nsew
rlabel metal1 1120 1540 1160 1840 0 pa1
rlabel metal1 1120 820 1160 1120 0 pb1
rlabel metal1 3040 820 3080 1120 0 pb2
rlabel metal1 1120 80 1160 180 0 n1
rlabel metal1 3040 80 3080 180 0 n2
rlabel metal1 3040 1540 3080 1840 0 pa2
<< end >>
