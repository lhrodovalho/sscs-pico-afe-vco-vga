magic
tech sky130A
timestamp 1638409393
<< locali >>
rect -480 20950 -440 20960
rect -480 20930 -470 20950
rect -450 20930 -440 20950
rect -480 20790 -440 20930
rect -480 20770 -470 20790
rect -450 20770 -440 20790
rect -480 20760 -440 20770
rect -400 20950 -360 20960
rect -400 20930 -390 20950
rect -370 20930 -360 20950
rect -400 20790 -360 20930
rect -400 20770 -390 20790
rect -370 20770 -360 20790
rect -400 20760 -360 20770
rect -320 20950 -280 20960
rect -320 20930 -310 20950
rect -290 20930 -280 20950
rect -320 20790 -280 20930
rect -320 20770 -310 20790
rect -290 20770 -280 20790
rect -320 20760 -280 20770
rect -240 20950 -200 20960
rect -240 20930 -230 20950
rect -210 20930 -200 20950
rect -240 20790 -200 20930
rect -240 20770 -230 20790
rect -210 20770 -200 20790
rect -240 20760 -200 20770
rect -160 20950 -120 20960
rect -160 20930 -150 20950
rect -130 20930 -120 20950
rect -160 20790 -120 20930
rect -160 20770 -150 20790
rect -130 20770 -120 20790
rect -160 20760 -120 20770
rect -80 20950 -40 20960
rect -80 20930 -70 20950
rect -50 20930 -40 20950
rect -80 20790 -40 20930
rect -80 20770 -70 20790
rect -50 20770 -40 20790
rect -80 20760 -40 20770
rect 0 20950 40 20960
rect 0 20930 10 20950
rect 30 20930 40 20950
rect 0 20790 40 20930
rect 0 20770 10 20790
rect 30 20770 40 20790
rect 0 20760 40 20770
rect 38360 20310 38400 20320
rect 38360 20290 38370 20310
rect 38390 20290 38400 20310
rect 38360 20150 38400 20290
rect 38360 20130 38370 20150
rect 38390 20130 38400 20150
rect 38360 20120 38400 20130
rect 38440 20310 38480 20320
rect 38440 20290 38450 20310
rect 38470 20290 38480 20310
rect 38440 20150 38480 20290
rect 38440 20130 38450 20150
rect 38470 20130 38480 20150
rect 38440 20120 38480 20130
rect -3520 19150 -3480 19160
rect -3520 19130 -3510 19150
rect -3490 19130 -3480 19150
rect -3520 18990 -3480 19130
rect -3520 18970 -3510 18990
rect -3490 18970 -3480 18990
rect -3520 18830 -3480 18970
rect -3520 18810 -3510 18830
rect -3490 18810 -3480 18830
rect -3520 18800 -3480 18810
rect -3440 19150 -3400 19160
rect -3440 19130 -3430 19150
rect -3410 19130 -3400 19150
rect -3440 18990 -3400 19130
rect -3440 18970 -3430 18990
rect -3410 18970 -3400 18990
rect -3440 18830 -3400 18970
rect -3440 18810 -3430 18830
rect -3410 18810 -3400 18830
rect -3440 18800 -3400 18810
rect -3360 19150 -3320 19160
rect -3360 19130 -3350 19150
rect -3330 19130 -3320 19150
rect -3360 18990 -3320 19130
rect -3360 18970 -3350 18990
rect -3330 18970 -3320 18990
rect -3360 18830 -3320 18970
rect -3360 18810 -3350 18830
rect -3330 18810 -3320 18830
rect -3360 18800 -3320 18810
rect -3280 19150 -3240 19160
rect -3280 19130 -3270 19150
rect -3250 19130 -3240 19150
rect -3280 18990 -3240 19130
rect -3280 18970 -3270 18990
rect -3250 18970 -3240 18990
rect -3280 18830 -3240 18970
rect -3280 18810 -3270 18830
rect -3250 18810 -3240 18830
rect -3280 18800 -3240 18810
rect -3200 19150 -3160 19160
rect -3200 19130 -3190 19150
rect -3170 19130 -3160 19150
rect -3200 18990 -3160 19130
rect -3200 18970 -3190 18990
rect -3170 18970 -3160 18990
rect -3200 18830 -3160 18970
rect -3200 18810 -3190 18830
rect -3170 18810 -3160 18830
rect -3200 18800 -3160 18810
rect -3120 19150 -3080 19160
rect -3120 19130 -3110 19150
rect -3090 19130 -3080 19150
rect -3120 18990 -3080 19130
rect -3120 18970 -3110 18990
rect -3090 18970 -3080 18990
rect -3120 18830 -3080 18970
rect -3120 18810 -3110 18830
rect -3090 18810 -3080 18830
rect -3120 18800 -3080 18810
rect -3040 19150 -3000 19160
rect -3040 19130 -3030 19150
rect -3010 19130 -3000 19150
rect -3040 18990 -3000 19130
rect -3040 18970 -3030 18990
rect -3010 18970 -3000 18990
rect -3040 18830 -3000 18970
rect -3040 18810 -3030 18830
rect -3010 18810 -3000 18830
rect -3040 18800 -3000 18810
rect -2960 19150 -2920 19160
rect -2960 19130 -2950 19150
rect -2930 19130 -2920 19150
rect -2960 18990 -2920 19130
rect -2960 18970 -2950 18990
rect -2930 18970 -2920 18990
rect -2960 18830 -2920 18970
rect -2960 18810 -2950 18830
rect -2930 18810 -2920 18830
rect -2960 18800 -2920 18810
rect -2880 19150 -2840 19160
rect -2880 19130 -2870 19150
rect -2850 19130 -2840 19150
rect -2880 18990 -2840 19130
rect -2880 18970 -2870 18990
rect -2850 18970 -2840 18990
rect -2880 18830 -2840 18970
rect -2880 18810 -2870 18830
rect -2850 18810 -2840 18830
rect -2880 18800 -2840 18810
rect -2800 19150 -2760 19160
rect -2800 19130 -2790 19150
rect -2770 19130 -2760 19150
rect -2800 18990 -2760 19130
rect -2800 18970 -2790 18990
rect -2770 18970 -2760 18990
rect -2800 18830 -2760 18970
rect -2800 18810 -2790 18830
rect -2770 18810 -2760 18830
rect -2800 18800 -2760 18810
rect -2720 19150 -2680 19160
rect -2720 19130 -2710 19150
rect -2690 19130 -2680 19150
rect -2720 18990 -2680 19130
rect -2720 18970 -2710 18990
rect -2690 18970 -2680 18990
rect -2720 18830 -2680 18970
rect -2720 18810 -2710 18830
rect -2690 18810 -2680 18830
rect -2720 18800 -2680 18810
rect -2640 19150 -2600 19160
rect -2640 19130 -2630 19150
rect -2610 19130 -2600 19150
rect -2640 18990 -2600 19130
rect -2640 18970 -2630 18990
rect -2610 18970 -2600 18990
rect -2640 18830 -2600 18970
rect -2640 18810 -2630 18830
rect -2610 18810 -2600 18830
rect -2640 18800 -2600 18810
rect -2560 19150 -2520 19160
rect -2560 19130 -2550 19150
rect -2530 19130 -2520 19150
rect -2560 18990 -2520 19130
rect -2560 18970 -2550 18990
rect -2530 18970 -2520 18990
rect -2560 18830 -2520 18970
rect -2560 18810 -2550 18830
rect -2530 18810 -2520 18830
rect -2560 18800 -2520 18810
rect -2480 19150 -2440 19160
rect -2480 19130 -2470 19150
rect -2450 19130 -2440 19150
rect -2480 18990 -2440 19130
rect -2480 18970 -2470 18990
rect -2450 18970 -2440 18990
rect -2480 18830 -2440 18970
rect -2480 18810 -2470 18830
rect -2450 18810 -2440 18830
rect -2480 18800 -2440 18810
rect -2400 19150 -2360 19160
rect -2400 19130 -2390 19150
rect -2370 19130 -2360 19150
rect -2400 18990 -2360 19130
rect -2400 18970 -2390 18990
rect -2370 18970 -2360 18990
rect -2400 18830 -2360 18970
rect -2400 18810 -2390 18830
rect -2370 18810 -2360 18830
rect -2400 18800 -2360 18810
rect -2320 19150 -2280 19160
rect -2320 19130 -2310 19150
rect -2290 19130 -2280 19150
rect -2320 18990 -2280 19130
rect -2320 18970 -2310 18990
rect -2290 18970 -2280 18990
rect -2320 18830 -2280 18970
rect -2320 18810 -2310 18830
rect -2290 18810 -2280 18830
rect -2320 18800 -2280 18810
rect -2240 19150 -2200 19160
rect -2240 19130 -2230 19150
rect -2210 19130 -2200 19150
rect -2240 18990 -2200 19130
rect -2240 18970 -2230 18990
rect -2210 18970 -2200 18990
rect -2240 18830 -2200 18970
rect -2240 18810 -2230 18830
rect -2210 18810 -2200 18830
rect -2240 18800 -2200 18810
rect -2160 19150 -2120 19160
rect -2160 19130 -2150 19150
rect -2130 19130 -2120 19150
rect -2160 18990 -2120 19130
rect -2160 18970 -2150 18990
rect -2130 18970 -2120 18990
rect -2160 18830 -2120 18970
rect -2160 18810 -2150 18830
rect -2130 18810 -2120 18830
rect -2160 18800 -2120 18810
rect -2080 19150 -2040 19160
rect -2080 19130 -2070 19150
rect -2050 19130 -2040 19150
rect -2080 18990 -2040 19130
rect -2080 18970 -2070 18990
rect -2050 18970 -2040 18990
rect -2080 18830 -2040 18970
rect -2080 18810 -2070 18830
rect -2050 18810 -2040 18830
rect -2080 18800 -2040 18810
rect -2000 19150 -1960 19160
rect -2000 19130 -1990 19150
rect -1970 19130 -1960 19150
rect -2000 18990 -1960 19130
rect -2000 18970 -1990 18990
rect -1970 18970 -1960 18990
rect -2000 18830 -1960 18970
rect -2000 18810 -1990 18830
rect -1970 18810 -1960 18830
rect -2000 18800 -1960 18810
rect -1920 19150 -1880 19160
rect -1920 19130 -1910 19150
rect -1890 19130 -1880 19150
rect -1920 18990 -1880 19130
rect -1920 18970 -1910 18990
rect -1890 18970 -1880 18990
rect -1920 18830 -1880 18970
rect -1920 18810 -1910 18830
rect -1890 18810 -1880 18830
rect -1920 18800 -1880 18810
rect -1840 19150 -1800 19160
rect -1840 19130 -1830 19150
rect -1810 19130 -1800 19150
rect -1840 18990 -1800 19130
rect -1840 18970 -1830 18990
rect -1810 18970 -1800 18990
rect -1840 18830 -1800 18970
rect -1840 18810 -1830 18830
rect -1810 18810 -1800 18830
rect -1840 18800 -1800 18810
rect -1760 19150 -1720 19160
rect -1760 19130 -1750 19150
rect -1730 19130 -1720 19150
rect -1760 18990 -1720 19130
rect -1760 18970 -1750 18990
rect -1730 18970 -1720 18990
rect -1760 18830 -1720 18970
rect -1760 18810 -1750 18830
rect -1730 18810 -1720 18830
rect -1760 18800 -1720 18810
rect -1680 19150 -1640 19160
rect -1680 19130 -1670 19150
rect -1650 19130 -1640 19150
rect -1680 18990 -1640 19130
rect -1680 18970 -1670 18990
rect -1650 18970 -1640 18990
rect -1680 18830 -1640 18970
rect -1680 18810 -1670 18830
rect -1650 18810 -1640 18830
rect -1680 18800 -1640 18810
rect -1600 19150 -1560 19160
rect -1600 19130 -1590 19150
rect -1570 19130 -1560 19150
rect -1600 18990 -1560 19130
rect -1600 18970 -1590 18990
rect -1570 18970 -1560 18990
rect -1600 18830 -1560 18970
rect -1600 18810 -1590 18830
rect -1570 18810 -1560 18830
rect -1600 18800 -1560 18810
rect -1520 19150 -1480 19160
rect -1520 19130 -1510 19150
rect -1490 19130 -1480 19150
rect -1520 18990 -1480 19130
rect -1520 18970 -1510 18990
rect -1490 18970 -1480 18990
rect -1520 18830 -1480 18970
rect -1520 18810 -1510 18830
rect -1490 18810 -1480 18830
rect -1520 18800 -1480 18810
rect -1440 19150 -1400 19160
rect -1440 19130 -1430 19150
rect -1410 19130 -1400 19150
rect -1440 18990 -1400 19130
rect -1440 18970 -1430 18990
rect -1410 18970 -1400 18990
rect -1440 18830 -1400 18970
rect -1440 18810 -1430 18830
rect -1410 18810 -1400 18830
rect -1440 18800 -1400 18810
rect -1360 19150 -1320 19160
rect -1360 19130 -1350 19150
rect -1330 19130 -1320 19150
rect -1360 18990 -1320 19130
rect -1360 18970 -1350 18990
rect -1330 18970 -1320 18990
rect -1360 18830 -1320 18970
rect -1360 18810 -1350 18830
rect -1330 18810 -1320 18830
rect -1360 18800 -1320 18810
rect -1280 19150 -1240 19160
rect -1280 19130 -1270 19150
rect -1250 19130 -1240 19150
rect -1280 18990 -1240 19130
rect -1280 18970 -1270 18990
rect -1250 18970 -1240 18990
rect -1280 18830 -1240 18970
rect -1280 18810 -1270 18830
rect -1250 18810 -1240 18830
rect -1280 18800 -1240 18810
rect -1200 19150 -1160 19160
rect -1200 19130 -1190 19150
rect -1170 19130 -1160 19150
rect -1200 18990 -1160 19130
rect -1200 18970 -1190 18990
rect -1170 18970 -1160 18990
rect -1200 18830 -1160 18970
rect -1200 18810 -1190 18830
rect -1170 18810 -1160 18830
rect -1200 18800 -1160 18810
rect -1120 19150 -1080 19160
rect -1120 19130 -1110 19150
rect -1090 19130 -1080 19150
rect -1120 18990 -1080 19130
rect -1120 18970 -1110 18990
rect -1090 18970 -1080 18990
rect -1120 18830 -1080 18970
rect -1120 18810 -1110 18830
rect -1090 18810 -1080 18830
rect -1120 18800 -1080 18810
rect -1040 19150 -1000 19160
rect -1040 19130 -1030 19150
rect -1010 19130 -1000 19150
rect -1040 18990 -1000 19130
rect -1040 18970 -1030 18990
rect -1010 18970 -1000 18990
rect -1040 18830 -1000 18970
rect -1040 18810 -1030 18830
rect -1010 18810 -1000 18830
rect -1040 18800 -1000 18810
rect -960 19150 -920 19160
rect -960 19130 -950 19150
rect -930 19130 -920 19150
rect -960 18990 -920 19130
rect -960 18970 -950 18990
rect -930 18970 -920 18990
rect -960 18830 -920 18970
rect -960 18810 -950 18830
rect -930 18810 -920 18830
rect -960 18800 -920 18810
rect -880 19150 -840 19160
rect -880 19130 -870 19150
rect -850 19130 -840 19150
rect -880 18990 -840 19130
rect -880 18970 -870 18990
rect -850 18970 -840 18990
rect -880 18830 -840 18970
rect -880 18810 -870 18830
rect -850 18810 -840 18830
rect -880 18800 -840 18810
rect -800 19150 -760 19160
rect -800 19130 -790 19150
rect -770 19130 -760 19150
rect -800 18990 -760 19130
rect -800 18970 -790 18990
rect -770 18970 -760 18990
rect -800 18830 -760 18970
rect -800 18810 -790 18830
rect -770 18810 -760 18830
rect -800 18800 -760 18810
rect -720 19150 -680 19160
rect -720 19130 -710 19150
rect -690 19130 -680 19150
rect -720 18990 -680 19130
rect -720 18970 -710 18990
rect -690 18970 -680 18990
rect -720 18830 -680 18970
rect -720 18810 -710 18830
rect -690 18810 -680 18830
rect -720 18800 -680 18810
rect -640 19150 -600 19160
rect -640 19130 -630 19150
rect -610 19130 -600 19150
rect -640 18990 -600 19130
rect -640 18970 -630 18990
rect -610 18970 -600 18990
rect -640 18830 -600 18970
rect -640 18810 -630 18830
rect -610 18810 -600 18830
rect -640 18800 -600 18810
rect -560 19150 -520 19160
rect -560 19130 -550 19150
rect -530 19130 -520 19150
rect -560 18990 -520 19130
rect -560 18970 -550 18990
rect -530 18970 -520 18990
rect -560 18830 -520 18970
rect -560 18810 -550 18830
rect -530 18810 -520 18830
rect -560 18800 -520 18810
rect -480 19150 -440 19160
rect -480 19130 -470 19150
rect -450 19130 -440 19150
rect -480 18990 -440 19130
rect -480 18970 -470 18990
rect -450 18970 -440 18990
rect -480 18830 -440 18970
rect -480 18810 -470 18830
rect -450 18810 -440 18830
rect -480 18800 -440 18810
rect -400 19150 -360 19160
rect -400 19130 -390 19150
rect -370 19130 -360 19150
rect -400 18990 -360 19130
rect -400 18970 -390 18990
rect -370 18970 -360 18990
rect -400 18830 -360 18970
rect -400 18810 -390 18830
rect -370 18810 -360 18830
rect -400 18800 -360 18810
rect -320 19150 -280 19160
rect -320 19130 -310 19150
rect -290 19130 -280 19150
rect -320 18990 -280 19130
rect -320 18970 -310 18990
rect -290 18970 -280 18990
rect -320 18830 -280 18970
rect -320 18810 -310 18830
rect -290 18810 -280 18830
rect -320 18800 -280 18810
rect -240 19150 -200 19160
rect -240 19130 -230 19150
rect -210 19130 -200 19150
rect -240 18990 -200 19130
rect -240 18970 -230 18990
rect -210 18970 -200 18990
rect -240 18830 -200 18970
rect -240 18810 -230 18830
rect -210 18810 -200 18830
rect -240 18800 -200 18810
rect -160 19150 -120 19160
rect -160 19130 -150 19150
rect -130 19130 -120 19150
rect -160 18990 -120 19130
rect -160 18970 -150 18990
rect -130 18970 -120 18990
rect -160 18830 -120 18970
rect -160 18810 -150 18830
rect -130 18810 -120 18830
rect -160 18800 -120 18810
rect -80 19150 -40 19160
rect -80 19130 -70 19150
rect -50 19130 -40 19150
rect -80 18990 -40 19130
rect -80 18970 -70 18990
rect -50 18970 -40 18990
rect -80 18830 -40 18970
rect -80 18810 -70 18830
rect -50 18810 -40 18830
rect -80 18800 -40 18810
rect 0 19150 40 19160
rect 0 19130 10 19150
rect 30 19130 40 19150
rect 0 18990 40 19130
rect 0 18970 10 18990
rect 30 18970 40 18990
rect 0 18830 40 18970
rect 0 18810 10 18830
rect 30 18810 40 18830
rect 0 18800 40 18810
rect 38360 18310 38400 18320
rect 38360 18290 38370 18310
rect 38390 18290 38400 18310
rect 38360 18150 38400 18290
rect 38360 18130 38370 18150
rect 38390 18130 38400 18150
rect 38360 18120 38400 18130
rect 38440 18310 38480 18320
rect 38440 18290 38450 18310
rect 38470 18290 38480 18310
rect 38440 18150 38480 18290
rect 38440 18130 38450 18150
rect 38470 18130 38480 18150
rect 38440 18120 38480 18130
rect -1280 17630 -1240 17640
rect -1280 17610 -1270 17630
rect -1250 17610 -1240 17630
rect -1280 17470 -1240 17610
rect -1280 17450 -1270 17470
rect -1250 17450 -1240 17470
rect -1280 17440 -1240 17450
rect -1200 17630 -1160 17640
rect -1200 17610 -1190 17630
rect -1170 17610 -1160 17630
rect -1200 17470 -1160 17610
rect -1200 17450 -1190 17470
rect -1170 17450 -1160 17470
rect -1200 17440 -1160 17450
rect -1120 17630 -1080 17640
rect -1120 17610 -1110 17630
rect -1090 17610 -1080 17630
rect -1120 17470 -1080 17610
rect -1120 17450 -1110 17470
rect -1090 17450 -1080 17470
rect -1120 17440 -1080 17450
rect -1040 17630 -1000 17640
rect -1040 17610 -1030 17630
rect -1010 17610 -1000 17630
rect -1040 17470 -1000 17610
rect -1040 17450 -1030 17470
rect -1010 17450 -1000 17470
rect -1040 17440 -1000 17450
rect -960 17630 -920 17640
rect -960 17610 -950 17630
rect -930 17610 -920 17630
rect -960 17470 -920 17610
rect -960 17450 -950 17470
rect -930 17450 -920 17470
rect -960 17440 -920 17450
rect -880 17630 -840 17640
rect -880 17610 -870 17630
rect -850 17610 -840 17630
rect -880 17470 -840 17610
rect -880 17450 -870 17470
rect -850 17450 -840 17470
rect -880 17440 -840 17450
rect -800 17630 -760 17640
rect -800 17610 -790 17630
rect -770 17610 -760 17630
rect -800 17470 -760 17610
rect -800 17450 -790 17470
rect -770 17450 -760 17470
rect -800 17440 -760 17450
rect -720 17630 -680 17640
rect -720 17610 -710 17630
rect -690 17610 -680 17630
rect -720 17470 -680 17610
rect -720 17450 -710 17470
rect -690 17450 -680 17470
rect -720 17440 -680 17450
rect -640 17630 -600 17640
rect -640 17610 -630 17630
rect -610 17610 -600 17630
rect -640 17470 -600 17610
rect -640 17450 -630 17470
rect -610 17450 -600 17470
rect -640 17440 -600 17450
rect -560 17630 -520 17640
rect -560 17610 -550 17630
rect -530 17610 -520 17630
rect -560 17470 -520 17610
rect -560 17450 -550 17470
rect -530 17450 -520 17470
rect -560 17440 -520 17450
rect -480 17630 -440 17640
rect -480 17610 -470 17630
rect -450 17610 -440 17630
rect -480 17470 -440 17610
rect -480 17450 -470 17470
rect -450 17450 -440 17470
rect -480 17440 -440 17450
rect -400 17630 -360 17640
rect -400 17610 -390 17630
rect -370 17610 -360 17630
rect -400 17470 -360 17610
rect -400 17450 -390 17470
rect -370 17450 -360 17470
rect -400 17440 -360 17450
rect -320 17630 -280 17640
rect -320 17610 -310 17630
rect -290 17610 -280 17630
rect -320 17470 -280 17610
rect -320 17450 -310 17470
rect -290 17450 -280 17470
rect -320 17440 -280 17450
rect -240 17630 -200 17640
rect -240 17610 -230 17630
rect -210 17610 -200 17630
rect -240 17470 -200 17610
rect -240 17450 -230 17470
rect -210 17450 -200 17470
rect -240 17440 -200 17450
rect -160 17630 -120 17640
rect -160 17610 -150 17630
rect -130 17610 -120 17630
rect -160 17470 -120 17610
rect -160 17450 -150 17470
rect -130 17450 -120 17470
rect -160 17440 -120 17450
rect -80 17630 -40 17640
rect -80 17610 -70 17630
rect -50 17610 -40 17630
rect -80 17470 -40 17610
rect -80 17450 -70 17470
rect -50 17450 -40 17470
rect -80 17440 -40 17450
rect 0 17630 40 17640
rect 0 17610 10 17630
rect 30 17610 40 17630
rect 0 17470 40 17610
rect 0 17450 10 17470
rect 30 17450 40 17470
rect 0 17440 40 17450
<< viali >>
rect -470 20930 -450 20950
rect -470 20770 -450 20790
rect -390 20930 -370 20950
rect -390 20770 -370 20790
rect -310 20930 -290 20950
rect -310 20770 -290 20790
rect -230 20930 -210 20950
rect -230 20770 -210 20790
rect -150 20930 -130 20950
rect -150 20770 -130 20790
rect -70 20930 -50 20950
rect -70 20770 -50 20790
rect 10 20930 30 20950
rect 10 20770 30 20790
rect 38370 20290 38390 20310
rect 38370 20130 38390 20150
rect 38450 20290 38470 20310
rect 38450 20130 38470 20150
rect -3510 19130 -3490 19150
rect -3510 18970 -3490 18990
rect -3510 18810 -3490 18830
rect -3430 19130 -3410 19150
rect -3430 18970 -3410 18990
rect -3430 18810 -3410 18830
rect -3350 19130 -3330 19150
rect -3350 18970 -3330 18990
rect -3350 18810 -3330 18830
rect -3270 19130 -3250 19150
rect -3270 18970 -3250 18990
rect -3270 18810 -3250 18830
rect -3190 19130 -3170 19150
rect -3190 18970 -3170 18990
rect -3190 18810 -3170 18830
rect -3110 19130 -3090 19150
rect -3110 18970 -3090 18990
rect -3110 18810 -3090 18830
rect -3030 19130 -3010 19150
rect -3030 18970 -3010 18990
rect -3030 18810 -3010 18830
rect -2950 19130 -2930 19150
rect -2950 18970 -2930 18990
rect -2950 18810 -2930 18830
rect -2870 19130 -2850 19150
rect -2870 18970 -2850 18990
rect -2870 18810 -2850 18830
rect -2790 19130 -2770 19150
rect -2790 18970 -2770 18990
rect -2790 18810 -2770 18830
rect -2710 19130 -2690 19150
rect -2710 18970 -2690 18990
rect -2710 18810 -2690 18830
rect -2630 19130 -2610 19150
rect -2630 18970 -2610 18990
rect -2630 18810 -2610 18830
rect -2550 19130 -2530 19150
rect -2550 18970 -2530 18990
rect -2550 18810 -2530 18830
rect -2470 19130 -2450 19150
rect -2470 18970 -2450 18990
rect -2470 18810 -2450 18830
rect -2390 19130 -2370 19150
rect -2390 18970 -2370 18990
rect -2390 18810 -2370 18830
rect -2310 19130 -2290 19150
rect -2310 18970 -2290 18990
rect -2310 18810 -2290 18830
rect -2230 19130 -2210 19150
rect -2230 18970 -2210 18990
rect -2230 18810 -2210 18830
rect -2150 19130 -2130 19150
rect -2150 18970 -2130 18990
rect -2150 18810 -2130 18830
rect -2070 19130 -2050 19150
rect -2070 18970 -2050 18990
rect -2070 18810 -2050 18830
rect -1990 19130 -1970 19150
rect -1990 18970 -1970 18990
rect -1990 18810 -1970 18830
rect -1910 19130 -1890 19150
rect -1910 18970 -1890 18990
rect -1910 18810 -1890 18830
rect -1830 19130 -1810 19150
rect -1830 18970 -1810 18990
rect -1830 18810 -1810 18830
rect -1750 19130 -1730 19150
rect -1750 18970 -1730 18990
rect -1750 18810 -1730 18830
rect -1670 19130 -1650 19150
rect -1670 18970 -1650 18990
rect -1670 18810 -1650 18830
rect -1590 19130 -1570 19150
rect -1590 18970 -1570 18990
rect -1590 18810 -1570 18830
rect -1510 19130 -1490 19150
rect -1510 18970 -1490 18990
rect -1510 18810 -1490 18830
rect -1430 19130 -1410 19150
rect -1430 18970 -1410 18990
rect -1430 18810 -1410 18830
rect -1350 19130 -1330 19150
rect -1350 18970 -1330 18990
rect -1350 18810 -1330 18830
rect -1270 19130 -1250 19150
rect -1270 18970 -1250 18990
rect -1270 18810 -1250 18830
rect -1190 19130 -1170 19150
rect -1190 18970 -1170 18990
rect -1190 18810 -1170 18830
rect -1110 19130 -1090 19150
rect -1110 18970 -1090 18990
rect -1110 18810 -1090 18830
rect -1030 19130 -1010 19150
rect -1030 18970 -1010 18990
rect -1030 18810 -1010 18830
rect -950 19130 -930 19150
rect -950 18970 -930 18990
rect -950 18810 -930 18830
rect -870 19130 -850 19150
rect -870 18970 -850 18990
rect -870 18810 -850 18830
rect -790 19130 -770 19150
rect -790 18970 -770 18990
rect -790 18810 -770 18830
rect -710 19130 -690 19150
rect -710 18970 -690 18990
rect -710 18810 -690 18830
rect -630 19130 -610 19150
rect -630 18970 -610 18990
rect -630 18810 -610 18830
rect -550 19130 -530 19150
rect -550 18970 -530 18990
rect -550 18810 -530 18830
rect -470 19130 -450 19150
rect -470 18970 -450 18990
rect -470 18810 -450 18830
rect -390 19130 -370 19150
rect -390 18970 -370 18990
rect -390 18810 -370 18830
rect -310 19130 -290 19150
rect -310 18970 -290 18990
rect -310 18810 -290 18830
rect -230 19130 -210 19150
rect -230 18970 -210 18990
rect -230 18810 -210 18830
rect -150 19130 -130 19150
rect -150 18970 -130 18990
rect -150 18810 -130 18830
rect -70 19130 -50 19150
rect -70 18970 -50 18990
rect -70 18810 -50 18830
rect 10 19130 30 19150
rect 10 18970 30 18990
rect 10 18810 30 18830
rect 38370 18290 38390 18310
rect 38370 18130 38390 18150
rect 38450 18290 38470 18310
rect 38450 18130 38470 18150
rect -1270 17610 -1250 17630
rect -1270 17450 -1250 17470
rect -1190 17610 -1170 17630
rect -1190 17450 -1170 17470
rect -1110 17610 -1090 17630
rect -1110 17450 -1090 17470
rect -1030 17610 -1010 17630
rect -1030 17450 -1010 17470
rect -950 17610 -930 17630
rect -950 17450 -930 17470
rect -870 17610 -850 17630
rect -870 17450 -850 17470
rect -790 17610 -770 17630
rect -790 17450 -770 17470
rect -710 17610 -690 17630
rect -710 17450 -690 17470
rect -630 17610 -610 17630
rect -630 17450 -610 17470
rect -550 17610 -530 17630
rect -550 17450 -530 17470
rect -470 17610 -450 17630
rect -470 17450 -450 17470
rect -390 17610 -370 17630
rect -390 17450 -370 17470
rect -310 17610 -290 17630
rect -310 17450 -290 17470
rect -230 17610 -210 17630
rect -230 17450 -210 17470
rect -150 17610 -130 17630
rect -150 17450 -130 17470
rect -70 17610 -50 17630
rect -70 17450 -50 17470
rect 10 17610 30 17630
rect 10 17450 30 17470
<< metal1 >>
rect -480 20955 -440 20960
rect -480 20925 -475 20955
rect -445 20925 -440 20955
rect -480 20920 -440 20925
rect -400 20955 -360 20960
rect -400 20925 -395 20955
rect -365 20925 -360 20955
rect -400 20920 -360 20925
rect -320 20955 -280 20960
rect -320 20925 -315 20955
rect -285 20925 -280 20955
rect -320 20920 -280 20925
rect -240 20955 -200 20960
rect -240 20925 -235 20955
rect -205 20925 -200 20955
rect -240 20920 -200 20925
rect -160 20955 -120 20960
rect -160 20925 -155 20955
rect -125 20925 -120 20955
rect -160 20920 -120 20925
rect -80 20955 -40 20960
rect -80 20925 -75 20955
rect -45 20925 -40 20955
rect -80 20920 -40 20925
rect 0 20955 40 20960
rect 0 20925 5 20955
rect 35 20925 40 20955
rect 0 20920 40 20925
rect -480 20795 -440 20800
rect -480 20765 -475 20795
rect -445 20765 -440 20795
rect -480 20760 -440 20765
rect -400 20795 -360 20800
rect -400 20765 -395 20795
rect -365 20765 -360 20795
rect -400 20760 -360 20765
rect -320 20795 -280 20800
rect -320 20765 -315 20795
rect -285 20765 -280 20795
rect -320 20760 -280 20765
rect -240 20795 -200 20800
rect -240 20765 -235 20795
rect -205 20765 -200 20795
rect -240 20760 -200 20765
rect -160 20795 -120 20800
rect -160 20765 -155 20795
rect -125 20765 -120 20795
rect -160 20760 -120 20765
rect -80 20795 -40 20800
rect -80 20765 -75 20795
rect -45 20765 -40 20795
rect -80 20760 -40 20765
rect 0 20795 40 20800
rect 0 20765 5 20795
rect 35 20765 40 20795
rect 0 20760 40 20765
rect 38360 20315 38400 20320
rect 38360 20285 38365 20315
rect 38395 20285 38400 20315
rect 38360 20280 38400 20285
rect 38440 20315 38480 20320
rect 38440 20285 38445 20315
rect 38475 20285 38480 20315
rect 38440 20280 38480 20285
rect 38360 20155 38400 20160
rect 38360 20125 38365 20155
rect 38395 20125 38400 20155
rect 38360 20120 38400 20125
rect 38440 20155 38480 20160
rect 38440 20125 38445 20155
rect 38475 20125 38480 20155
rect 38440 20120 38480 20125
rect -3520 19155 -3480 19160
rect -3520 19125 -3515 19155
rect -3485 19125 -3480 19155
rect -3520 19120 -3480 19125
rect -3440 19155 -3400 19160
rect -3440 19125 -3435 19155
rect -3405 19125 -3400 19155
rect -3440 19120 -3400 19125
rect -3360 19155 -3320 19160
rect -3360 19125 -3355 19155
rect -3325 19125 -3320 19155
rect -3360 19120 -3320 19125
rect -3280 19155 -3240 19160
rect -3280 19125 -3275 19155
rect -3245 19125 -3240 19155
rect -3280 19120 -3240 19125
rect -3200 19155 -3160 19160
rect -3200 19125 -3195 19155
rect -3165 19125 -3160 19155
rect -3200 19120 -3160 19125
rect -3120 19155 -3080 19160
rect -3120 19125 -3115 19155
rect -3085 19125 -3080 19155
rect -3120 19120 -3080 19125
rect -3040 19155 -3000 19160
rect -3040 19125 -3035 19155
rect -3005 19125 -3000 19155
rect -3040 19120 -3000 19125
rect -2960 19155 -2920 19160
rect -2960 19125 -2955 19155
rect -2925 19125 -2920 19155
rect -2960 19120 -2920 19125
rect -2880 19155 -2840 19160
rect -2880 19125 -2875 19155
rect -2845 19125 -2840 19155
rect -2880 19120 -2840 19125
rect -2800 19155 -2760 19160
rect -2800 19125 -2795 19155
rect -2765 19125 -2760 19155
rect -2800 19120 -2760 19125
rect -2720 19155 -2680 19160
rect -2720 19125 -2715 19155
rect -2685 19125 -2680 19155
rect -2720 19120 -2680 19125
rect -2640 19155 -2600 19160
rect -2640 19125 -2635 19155
rect -2605 19125 -2600 19155
rect -2640 19120 -2600 19125
rect -2560 19155 -2520 19160
rect -2560 19125 -2555 19155
rect -2525 19125 -2520 19155
rect -2560 19120 -2520 19125
rect -2480 19155 -2440 19160
rect -2480 19125 -2475 19155
rect -2445 19125 -2440 19155
rect -2480 19120 -2440 19125
rect -2400 19155 -2360 19160
rect -2400 19125 -2395 19155
rect -2365 19125 -2360 19155
rect -2400 19120 -2360 19125
rect -2320 19155 -2280 19160
rect -2320 19125 -2315 19155
rect -2285 19125 -2280 19155
rect -2320 19120 -2280 19125
rect -2240 19155 -2200 19160
rect -2240 19125 -2235 19155
rect -2205 19125 -2200 19155
rect -2240 19120 -2200 19125
rect -2160 19155 -2120 19160
rect -2160 19125 -2155 19155
rect -2125 19125 -2120 19155
rect -2160 19120 -2120 19125
rect -2080 19155 -2040 19160
rect -2080 19125 -2075 19155
rect -2045 19125 -2040 19155
rect -2080 19120 -2040 19125
rect -2000 19155 -1960 19160
rect -2000 19125 -1995 19155
rect -1965 19125 -1960 19155
rect -2000 19120 -1960 19125
rect -1920 19155 -1880 19160
rect -1920 19125 -1915 19155
rect -1885 19125 -1880 19155
rect -1920 19120 -1880 19125
rect -1840 19155 -1800 19160
rect -1840 19125 -1835 19155
rect -1805 19125 -1800 19155
rect -1840 19120 -1800 19125
rect -1760 19155 -1720 19160
rect -1760 19125 -1755 19155
rect -1725 19125 -1720 19155
rect -1760 19120 -1720 19125
rect -1680 19155 -1640 19160
rect -1680 19125 -1675 19155
rect -1645 19125 -1640 19155
rect -1680 19120 -1640 19125
rect -1600 19155 -1560 19160
rect -1600 19125 -1595 19155
rect -1565 19125 -1560 19155
rect -1600 19120 -1560 19125
rect -1520 19155 -1480 19160
rect -1520 19125 -1515 19155
rect -1485 19125 -1480 19155
rect -1520 19120 -1480 19125
rect -1440 19155 -1400 19160
rect -1440 19125 -1435 19155
rect -1405 19125 -1400 19155
rect -1440 19120 -1400 19125
rect -1360 19155 -1320 19160
rect -1360 19125 -1355 19155
rect -1325 19125 -1320 19155
rect -1360 19120 -1320 19125
rect -1280 19155 -1240 19160
rect -1280 19125 -1275 19155
rect -1245 19125 -1240 19155
rect -1280 19120 -1240 19125
rect -1200 19155 -1160 19160
rect -1200 19125 -1195 19155
rect -1165 19125 -1160 19155
rect -1200 19120 -1160 19125
rect -1120 19155 -1080 19160
rect -1120 19125 -1115 19155
rect -1085 19125 -1080 19155
rect -1120 19120 -1080 19125
rect -1040 19155 -1000 19160
rect -1040 19125 -1035 19155
rect -1005 19125 -1000 19155
rect -1040 19120 -1000 19125
rect -960 19155 -920 19160
rect -960 19125 -955 19155
rect -925 19125 -920 19155
rect -960 19120 -920 19125
rect -880 19155 -840 19160
rect -880 19125 -875 19155
rect -845 19125 -840 19155
rect -880 19120 -840 19125
rect -800 19155 -760 19160
rect -800 19125 -795 19155
rect -765 19125 -760 19155
rect -800 19120 -760 19125
rect -720 19155 -680 19160
rect -720 19125 -715 19155
rect -685 19125 -680 19155
rect -720 19120 -680 19125
rect -640 19155 -600 19160
rect -640 19125 -635 19155
rect -605 19125 -600 19155
rect -640 19120 -600 19125
rect -560 19155 -520 19160
rect -560 19125 -555 19155
rect -525 19125 -520 19155
rect -560 19120 -520 19125
rect -480 19155 -440 19160
rect -480 19125 -475 19155
rect -445 19125 -440 19155
rect -480 19120 -440 19125
rect -400 19155 -360 19160
rect -400 19125 -395 19155
rect -365 19125 -360 19155
rect -400 19120 -360 19125
rect -320 19155 -280 19160
rect -320 19125 -315 19155
rect -285 19125 -280 19155
rect -320 19120 -280 19125
rect -240 19155 -200 19160
rect -240 19125 -235 19155
rect -205 19125 -200 19155
rect -240 19120 -200 19125
rect -160 19155 -120 19160
rect -160 19125 -155 19155
rect -125 19125 -120 19155
rect -160 19120 -120 19125
rect -80 19155 -40 19160
rect -80 19125 -75 19155
rect -45 19125 -40 19155
rect -80 19120 -40 19125
rect 0 19155 40 19160
rect 0 19125 5 19155
rect 35 19125 40 19155
rect 0 19120 40 19125
rect -3520 18995 -3480 19000
rect -3520 18965 -3515 18995
rect -3485 18965 -3480 18995
rect -3520 18960 -3480 18965
rect -3440 18995 -3400 19000
rect -3440 18965 -3435 18995
rect -3405 18965 -3400 18995
rect -3440 18960 -3400 18965
rect -3360 18995 -3320 19000
rect -3360 18965 -3355 18995
rect -3325 18965 -3320 18995
rect -3360 18960 -3320 18965
rect -3280 18995 -3240 19000
rect -3280 18965 -3275 18995
rect -3245 18965 -3240 18995
rect -3280 18960 -3240 18965
rect -3200 18995 -3160 19000
rect -3200 18965 -3195 18995
rect -3165 18965 -3160 18995
rect -3200 18960 -3160 18965
rect -3120 18995 -3080 19000
rect -3120 18965 -3115 18995
rect -3085 18965 -3080 18995
rect -3120 18960 -3080 18965
rect -3040 18995 -3000 19000
rect -3040 18965 -3035 18995
rect -3005 18965 -3000 18995
rect -3040 18960 -3000 18965
rect -2960 18995 -2920 19000
rect -2960 18965 -2955 18995
rect -2925 18965 -2920 18995
rect -2960 18960 -2920 18965
rect -2880 18995 -2840 19000
rect -2880 18965 -2875 18995
rect -2845 18965 -2840 18995
rect -2880 18960 -2840 18965
rect -2800 18995 -2760 19000
rect -2800 18965 -2795 18995
rect -2765 18965 -2760 18995
rect -2800 18960 -2760 18965
rect -2720 18995 -2680 19000
rect -2720 18965 -2715 18995
rect -2685 18965 -2680 18995
rect -2720 18960 -2680 18965
rect -2640 18995 -2600 19000
rect -2640 18965 -2635 18995
rect -2605 18965 -2600 18995
rect -2640 18960 -2600 18965
rect -2560 18995 -2520 19000
rect -2560 18965 -2555 18995
rect -2525 18965 -2520 18995
rect -2560 18960 -2520 18965
rect -2480 18995 -2440 19000
rect -2480 18965 -2475 18995
rect -2445 18965 -2440 18995
rect -2480 18960 -2440 18965
rect -2400 18995 -2360 19000
rect -2400 18965 -2395 18995
rect -2365 18965 -2360 18995
rect -2400 18960 -2360 18965
rect -2320 18995 -2280 19000
rect -2320 18965 -2315 18995
rect -2285 18965 -2280 18995
rect -2320 18960 -2280 18965
rect -2240 18995 -2200 19000
rect -2240 18965 -2235 18995
rect -2205 18965 -2200 18995
rect -2240 18960 -2200 18965
rect -2160 18995 -2120 19000
rect -2160 18965 -2155 18995
rect -2125 18965 -2120 18995
rect -2160 18960 -2120 18965
rect -2080 18995 -2040 19000
rect -2080 18965 -2075 18995
rect -2045 18965 -2040 18995
rect -2080 18960 -2040 18965
rect -2000 18995 -1960 19000
rect -2000 18965 -1995 18995
rect -1965 18965 -1960 18995
rect -2000 18960 -1960 18965
rect -1920 18995 -1880 19000
rect -1920 18965 -1915 18995
rect -1885 18965 -1880 18995
rect -1920 18960 -1880 18965
rect -1840 18995 -1800 19000
rect -1840 18965 -1835 18995
rect -1805 18965 -1800 18995
rect -1840 18960 -1800 18965
rect -1760 18995 -1720 19000
rect -1760 18965 -1755 18995
rect -1725 18965 -1720 18995
rect -1760 18960 -1720 18965
rect -1680 18995 -1640 19000
rect -1680 18965 -1675 18995
rect -1645 18965 -1640 18995
rect -1680 18960 -1640 18965
rect -1600 18995 -1560 19000
rect -1600 18965 -1595 18995
rect -1565 18965 -1560 18995
rect -1600 18960 -1560 18965
rect -1520 18995 -1480 19000
rect -1520 18965 -1515 18995
rect -1485 18965 -1480 18995
rect -1520 18960 -1480 18965
rect -1440 18995 -1400 19000
rect -1440 18965 -1435 18995
rect -1405 18965 -1400 18995
rect -1440 18960 -1400 18965
rect -1360 18995 -1320 19000
rect -1360 18965 -1355 18995
rect -1325 18965 -1320 18995
rect -1360 18960 -1320 18965
rect -1280 18995 -1240 19000
rect -1280 18965 -1275 18995
rect -1245 18965 -1240 18995
rect -1280 18960 -1240 18965
rect -1200 18995 -1160 19000
rect -1200 18965 -1195 18995
rect -1165 18965 -1160 18995
rect -1200 18960 -1160 18965
rect -1120 18995 -1080 19000
rect -1120 18965 -1115 18995
rect -1085 18965 -1080 18995
rect -1120 18960 -1080 18965
rect -1040 18995 -1000 19000
rect -1040 18965 -1035 18995
rect -1005 18965 -1000 18995
rect -1040 18960 -1000 18965
rect -960 18995 -920 19000
rect -960 18965 -955 18995
rect -925 18965 -920 18995
rect -960 18960 -920 18965
rect -880 18995 -840 19000
rect -880 18965 -875 18995
rect -845 18965 -840 18995
rect -880 18960 -840 18965
rect -800 18995 -760 19000
rect -800 18965 -795 18995
rect -765 18965 -760 18995
rect -800 18960 -760 18965
rect -720 18995 -680 19000
rect -720 18965 -715 18995
rect -685 18965 -680 18995
rect -720 18960 -680 18965
rect -640 18995 -600 19000
rect -640 18965 -635 18995
rect -605 18965 -600 18995
rect -640 18960 -600 18965
rect -560 18995 -520 19000
rect -560 18965 -555 18995
rect -525 18965 -520 18995
rect -560 18960 -520 18965
rect -480 18995 -440 19000
rect -480 18965 -475 18995
rect -445 18965 -440 18995
rect -480 18960 -440 18965
rect -400 18995 -360 19000
rect -400 18965 -395 18995
rect -365 18965 -360 18995
rect -400 18960 -360 18965
rect -320 18995 -280 19000
rect -320 18965 -315 18995
rect -285 18965 -280 18995
rect -320 18960 -280 18965
rect -240 18995 -200 19000
rect -240 18965 -235 18995
rect -205 18965 -200 18995
rect -240 18960 -200 18965
rect -160 18995 -120 19000
rect -160 18965 -155 18995
rect -125 18965 -120 18995
rect -160 18960 -120 18965
rect -80 18995 -40 19000
rect -80 18965 -75 18995
rect -45 18965 -40 18995
rect -80 18960 -40 18965
rect 0 18995 40 19000
rect 0 18965 5 18995
rect 35 18965 40 18995
rect 0 18960 40 18965
rect -3520 18835 -3480 18840
rect -3520 18805 -3515 18835
rect -3485 18805 -3480 18835
rect -3520 18800 -3480 18805
rect -3440 18835 -3400 18840
rect -3440 18805 -3435 18835
rect -3405 18805 -3400 18835
rect -3440 18800 -3400 18805
rect -3360 18835 -3320 18840
rect -3360 18805 -3355 18835
rect -3325 18805 -3320 18835
rect -3360 18800 -3320 18805
rect -3280 18835 -3240 18840
rect -3280 18805 -3275 18835
rect -3245 18805 -3240 18835
rect -3280 18800 -3240 18805
rect -3200 18835 -3160 18840
rect -3200 18805 -3195 18835
rect -3165 18805 -3160 18835
rect -3200 18800 -3160 18805
rect -3120 18835 -3080 18840
rect -3120 18805 -3115 18835
rect -3085 18805 -3080 18835
rect -3120 18800 -3080 18805
rect -3040 18835 -3000 18840
rect -3040 18805 -3035 18835
rect -3005 18805 -3000 18835
rect -3040 18800 -3000 18805
rect -2960 18835 -2920 18840
rect -2960 18805 -2955 18835
rect -2925 18805 -2920 18835
rect -2960 18800 -2920 18805
rect -2880 18835 -2840 18840
rect -2880 18805 -2875 18835
rect -2845 18805 -2840 18835
rect -2880 18800 -2840 18805
rect -2800 18835 -2760 18840
rect -2800 18805 -2795 18835
rect -2765 18805 -2760 18835
rect -2800 18800 -2760 18805
rect -2720 18835 -2680 18840
rect -2720 18805 -2715 18835
rect -2685 18805 -2680 18835
rect -2720 18800 -2680 18805
rect -2640 18835 -2600 18840
rect -2640 18805 -2635 18835
rect -2605 18805 -2600 18835
rect -2640 18800 -2600 18805
rect -2560 18835 -2520 18840
rect -2560 18805 -2555 18835
rect -2525 18805 -2520 18835
rect -2560 18800 -2520 18805
rect -2480 18835 -2440 18840
rect -2480 18805 -2475 18835
rect -2445 18805 -2440 18835
rect -2480 18800 -2440 18805
rect -2400 18835 -2360 18840
rect -2400 18805 -2395 18835
rect -2365 18805 -2360 18835
rect -2400 18800 -2360 18805
rect -2320 18835 -2280 18840
rect -2320 18805 -2315 18835
rect -2285 18805 -2280 18835
rect -2320 18800 -2280 18805
rect -2240 18835 -2200 18840
rect -2240 18805 -2235 18835
rect -2205 18805 -2200 18835
rect -2240 18800 -2200 18805
rect -2160 18835 -2120 18840
rect -2160 18805 -2155 18835
rect -2125 18805 -2120 18835
rect -2160 18800 -2120 18805
rect -2080 18835 -2040 18840
rect -2080 18805 -2075 18835
rect -2045 18805 -2040 18835
rect -2080 18800 -2040 18805
rect -2000 18835 -1960 18840
rect -2000 18805 -1995 18835
rect -1965 18805 -1960 18835
rect -2000 18800 -1960 18805
rect -1920 18835 -1880 18840
rect -1920 18805 -1915 18835
rect -1885 18805 -1880 18835
rect -1920 18800 -1880 18805
rect -1840 18835 -1800 18840
rect -1840 18805 -1835 18835
rect -1805 18805 -1800 18835
rect -1840 18800 -1800 18805
rect -1760 18835 -1720 18840
rect -1760 18805 -1755 18835
rect -1725 18805 -1720 18835
rect -1760 18800 -1720 18805
rect -1680 18835 -1640 18840
rect -1680 18805 -1675 18835
rect -1645 18805 -1640 18835
rect -1680 18800 -1640 18805
rect -1600 18835 -1560 18840
rect -1600 18805 -1595 18835
rect -1565 18805 -1560 18835
rect -1600 18800 -1560 18805
rect -1520 18835 -1480 18840
rect -1520 18805 -1515 18835
rect -1485 18805 -1480 18835
rect -1520 18800 -1480 18805
rect -1440 18835 -1400 18840
rect -1440 18805 -1435 18835
rect -1405 18805 -1400 18835
rect -1440 18800 -1400 18805
rect -1360 18835 -1320 18840
rect -1360 18805 -1355 18835
rect -1325 18805 -1320 18835
rect -1360 18800 -1320 18805
rect -1280 18835 -1240 18840
rect -1280 18805 -1275 18835
rect -1245 18805 -1240 18835
rect -1280 18800 -1240 18805
rect -1200 18835 -1160 18840
rect -1200 18805 -1195 18835
rect -1165 18805 -1160 18835
rect -1200 18800 -1160 18805
rect -1120 18835 -1080 18840
rect -1120 18805 -1115 18835
rect -1085 18805 -1080 18835
rect -1120 18800 -1080 18805
rect -1040 18835 -1000 18840
rect -1040 18805 -1035 18835
rect -1005 18805 -1000 18835
rect -1040 18800 -1000 18805
rect -960 18835 -920 18840
rect -960 18805 -955 18835
rect -925 18805 -920 18835
rect -960 18800 -920 18805
rect -880 18835 -840 18840
rect -880 18805 -875 18835
rect -845 18805 -840 18835
rect -880 18800 -840 18805
rect -800 18835 -760 18840
rect -800 18805 -795 18835
rect -765 18805 -760 18835
rect -800 18800 -760 18805
rect -720 18835 -680 18840
rect -720 18805 -715 18835
rect -685 18805 -680 18835
rect -720 18800 -680 18805
rect -640 18835 -600 18840
rect -640 18805 -635 18835
rect -605 18805 -600 18835
rect -640 18800 -600 18805
rect -560 18835 -520 18840
rect -560 18805 -555 18835
rect -525 18805 -520 18835
rect -560 18800 -520 18805
rect -480 18835 -440 18840
rect -480 18805 -475 18835
rect -445 18805 -440 18835
rect -480 18800 -440 18805
rect -400 18835 -360 18840
rect -400 18805 -395 18835
rect -365 18805 -360 18835
rect -400 18800 -360 18805
rect -320 18835 -280 18840
rect -320 18805 -315 18835
rect -285 18805 -280 18835
rect -320 18800 -280 18805
rect -240 18835 -200 18840
rect -240 18805 -235 18835
rect -205 18805 -200 18835
rect -240 18800 -200 18805
rect -160 18835 -120 18840
rect -160 18805 -155 18835
rect -125 18805 -120 18835
rect -160 18800 -120 18805
rect -80 18835 -40 18840
rect -80 18805 -75 18835
rect -45 18805 -40 18835
rect -80 18800 -40 18805
rect 0 18835 40 18840
rect 0 18805 5 18835
rect 35 18805 40 18835
rect 0 18800 40 18805
rect 38360 18315 38400 18320
rect 38360 18285 38365 18315
rect 38395 18285 38400 18315
rect 38360 18280 38400 18285
rect 38440 18315 38480 18320
rect 38440 18285 38445 18315
rect 38475 18285 38480 18315
rect 38440 18280 38480 18285
rect 38360 18155 38400 18160
rect 38360 18125 38365 18155
rect 38395 18125 38400 18155
rect 38360 18120 38400 18125
rect 38440 18155 38480 18160
rect 38440 18125 38445 18155
rect 38475 18125 38480 18155
rect 38440 18120 38480 18125
rect -1280 17635 -1240 17640
rect -1280 17605 -1275 17635
rect -1245 17605 -1240 17635
rect -1280 17600 -1240 17605
rect -1200 17635 -1160 17640
rect -1200 17605 -1195 17635
rect -1165 17605 -1160 17635
rect -1200 17600 -1160 17605
rect -1120 17635 -1080 17640
rect -1120 17605 -1115 17635
rect -1085 17605 -1080 17635
rect -1120 17600 -1080 17605
rect -1040 17635 -1000 17640
rect -1040 17605 -1035 17635
rect -1005 17605 -1000 17635
rect -1040 17600 -1000 17605
rect -960 17635 -920 17640
rect -960 17605 -955 17635
rect -925 17605 -920 17635
rect -960 17600 -920 17605
rect -880 17635 -840 17640
rect -880 17605 -875 17635
rect -845 17605 -840 17635
rect -880 17600 -840 17605
rect -800 17635 -760 17640
rect -800 17605 -795 17635
rect -765 17605 -760 17635
rect -800 17600 -760 17605
rect -720 17635 -680 17640
rect -720 17605 -715 17635
rect -685 17605 -680 17635
rect -720 17600 -680 17605
rect -640 17635 -600 17640
rect -640 17605 -635 17635
rect -605 17605 -600 17635
rect -640 17600 -600 17605
rect -560 17635 -520 17640
rect -560 17605 -555 17635
rect -525 17605 -520 17635
rect -560 17600 -520 17605
rect -480 17635 -440 17640
rect -480 17605 -475 17635
rect -445 17605 -440 17635
rect -480 17600 -440 17605
rect -400 17635 -360 17640
rect -400 17605 -395 17635
rect -365 17605 -360 17635
rect -400 17600 -360 17605
rect -320 17635 -280 17640
rect -320 17605 -315 17635
rect -285 17605 -280 17635
rect -320 17600 -280 17605
rect -240 17635 -200 17640
rect -240 17605 -235 17635
rect -205 17605 -200 17635
rect -240 17600 -200 17605
rect -160 17635 -120 17640
rect -160 17605 -155 17635
rect -125 17605 -120 17635
rect -160 17600 -120 17605
rect -80 17635 -40 17640
rect -80 17605 -75 17635
rect -45 17605 -40 17635
rect -80 17600 -40 17605
rect 0 17635 40 17640
rect 0 17605 5 17635
rect 35 17605 40 17635
rect 0 17600 40 17605
rect -1280 17475 -1240 17480
rect -1280 17445 -1275 17475
rect -1245 17445 -1240 17475
rect -1280 17440 -1240 17445
rect -1200 17475 -1160 17480
rect -1200 17445 -1195 17475
rect -1165 17445 -1160 17475
rect -1200 17440 -1160 17445
rect -1120 17475 -1080 17480
rect -1120 17445 -1115 17475
rect -1085 17445 -1080 17475
rect -1120 17440 -1080 17445
rect -1040 17475 -1000 17480
rect -1040 17445 -1035 17475
rect -1005 17445 -1000 17475
rect -1040 17440 -1000 17445
rect -960 17475 -920 17480
rect -960 17445 -955 17475
rect -925 17445 -920 17475
rect -960 17440 -920 17445
rect -880 17475 -840 17480
rect -880 17445 -875 17475
rect -845 17445 -840 17475
rect -880 17440 -840 17445
rect -800 17475 -760 17480
rect -800 17445 -795 17475
rect -765 17445 -760 17475
rect -800 17440 -760 17445
rect -720 17475 -680 17480
rect -720 17445 -715 17475
rect -685 17445 -680 17475
rect -720 17440 -680 17445
rect -640 17475 -600 17480
rect -640 17445 -635 17475
rect -605 17445 -600 17475
rect -640 17440 -600 17445
rect -560 17475 -520 17480
rect -560 17445 -555 17475
rect -525 17445 -520 17475
rect -560 17440 -520 17445
rect -480 17475 -440 17480
rect -480 17445 -475 17475
rect -445 17445 -440 17475
rect -480 17440 -440 17445
rect -400 17475 -360 17480
rect -400 17445 -395 17475
rect -365 17445 -360 17475
rect -400 17440 -360 17445
rect -320 17475 -280 17480
rect -320 17445 -315 17475
rect -285 17445 -280 17475
rect -320 17440 -280 17445
rect -240 17475 -200 17480
rect -240 17445 -235 17475
rect -205 17445 -200 17475
rect -240 17440 -200 17445
rect -160 17475 -120 17480
rect -160 17445 -155 17475
rect -125 17445 -120 17475
rect -160 17440 -120 17445
rect -80 17475 -40 17480
rect -80 17445 -75 17475
rect -45 17445 -40 17475
rect -80 17440 -40 17445
rect 0 17475 40 17480
rect 0 17445 5 17475
rect 35 17445 40 17475
rect 0 17440 40 17445
<< via1 >>
rect -475 20950 -445 20955
rect -475 20930 -470 20950
rect -470 20930 -450 20950
rect -450 20930 -445 20950
rect -475 20925 -445 20930
rect -395 20950 -365 20955
rect -395 20930 -390 20950
rect -390 20930 -370 20950
rect -370 20930 -365 20950
rect -395 20925 -365 20930
rect -315 20950 -285 20955
rect -315 20930 -310 20950
rect -310 20930 -290 20950
rect -290 20930 -285 20950
rect -315 20925 -285 20930
rect -235 20950 -205 20955
rect -235 20930 -230 20950
rect -230 20930 -210 20950
rect -210 20930 -205 20950
rect -235 20925 -205 20930
rect -155 20950 -125 20955
rect -155 20930 -150 20950
rect -150 20930 -130 20950
rect -130 20930 -125 20950
rect -155 20925 -125 20930
rect -75 20950 -45 20955
rect -75 20930 -70 20950
rect -70 20930 -50 20950
rect -50 20930 -45 20950
rect -75 20925 -45 20930
rect 5 20950 35 20955
rect 5 20930 10 20950
rect 10 20930 30 20950
rect 30 20930 35 20950
rect 5 20925 35 20930
rect -475 20790 -445 20795
rect -475 20770 -470 20790
rect -470 20770 -450 20790
rect -450 20770 -445 20790
rect -475 20765 -445 20770
rect -395 20790 -365 20795
rect -395 20770 -390 20790
rect -390 20770 -370 20790
rect -370 20770 -365 20790
rect -395 20765 -365 20770
rect -315 20790 -285 20795
rect -315 20770 -310 20790
rect -310 20770 -290 20790
rect -290 20770 -285 20790
rect -315 20765 -285 20770
rect -235 20790 -205 20795
rect -235 20770 -230 20790
rect -230 20770 -210 20790
rect -210 20770 -205 20790
rect -235 20765 -205 20770
rect -155 20790 -125 20795
rect -155 20770 -150 20790
rect -150 20770 -130 20790
rect -130 20770 -125 20790
rect -155 20765 -125 20770
rect -75 20790 -45 20795
rect -75 20770 -70 20790
rect -70 20770 -50 20790
rect -50 20770 -45 20790
rect -75 20765 -45 20770
rect 5 20790 35 20795
rect 5 20770 10 20790
rect 10 20770 30 20790
rect 30 20770 35 20790
rect 5 20765 35 20770
rect 38365 20310 38395 20315
rect 38365 20290 38370 20310
rect 38370 20290 38390 20310
rect 38390 20290 38395 20310
rect 38365 20285 38395 20290
rect 38445 20310 38475 20315
rect 38445 20290 38450 20310
rect 38450 20290 38470 20310
rect 38470 20290 38475 20310
rect 38445 20285 38475 20290
rect 38365 20150 38395 20155
rect 38365 20130 38370 20150
rect 38370 20130 38390 20150
rect 38390 20130 38395 20150
rect 38365 20125 38395 20130
rect 38445 20150 38475 20155
rect 38445 20130 38450 20150
rect 38450 20130 38470 20150
rect 38470 20130 38475 20150
rect 38445 20125 38475 20130
rect -3515 19150 -3485 19155
rect -3515 19130 -3510 19150
rect -3510 19130 -3490 19150
rect -3490 19130 -3485 19150
rect -3515 19125 -3485 19130
rect -3435 19150 -3405 19155
rect -3435 19130 -3430 19150
rect -3430 19130 -3410 19150
rect -3410 19130 -3405 19150
rect -3435 19125 -3405 19130
rect -3355 19150 -3325 19155
rect -3355 19130 -3350 19150
rect -3350 19130 -3330 19150
rect -3330 19130 -3325 19150
rect -3355 19125 -3325 19130
rect -3275 19150 -3245 19155
rect -3275 19130 -3270 19150
rect -3270 19130 -3250 19150
rect -3250 19130 -3245 19150
rect -3275 19125 -3245 19130
rect -3195 19150 -3165 19155
rect -3195 19130 -3190 19150
rect -3190 19130 -3170 19150
rect -3170 19130 -3165 19150
rect -3195 19125 -3165 19130
rect -3115 19150 -3085 19155
rect -3115 19130 -3110 19150
rect -3110 19130 -3090 19150
rect -3090 19130 -3085 19150
rect -3115 19125 -3085 19130
rect -3035 19150 -3005 19155
rect -3035 19130 -3030 19150
rect -3030 19130 -3010 19150
rect -3010 19130 -3005 19150
rect -3035 19125 -3005 19130
rect -2955 19150 -2925 19155
rect -2955 19130 -2950 19150
rect -2950 19130 -2930 19150
rect -2930 19130 -2925 19150
rect -2955 19125 -2925 19130
rect -2875 19150 -2845 19155
rect -2875 19130 -2870 19150
rect -2870 19130 -2850 19150
rect -2850 19130 -2845 19150
rect -2875 19125 -2845 19130
rect -2795 19150 -2765 19155
rect -2795 19130 -2790 19150
rect -2790 19130 -2770 19150
rect -2770 19130 -2765 19150
rect -2795 19125 -2765 19130
rect -2715 19150 -2685 19155
rect -2715 19130 -2710 19150
rect -2710 19130 -2690 19150
rect -2690 19130 -2685 19150
rect -2715 19125 -2685 19130
rect -2635 19150 -2605 19155
rect -2635 19130 -2630 19150
rect -2630 19130 -2610 19150
rect -2610 19130 -2605 19150
rect -2635 19125 -2605 19130
rect -2555 19150 -2525 19155
rect -2555 19130 -2550 19150
rect -2550 19130 -2530 19150
rect -2530 19130 -2525 19150
rect -2555 19125 -2525 19130
rect -2475 19150 -2445 19155
rect -2475 19130 -2470 19150
rect -2470 19130 -2450 19150
rect -2450 19130 -2445 19150
rect -2475 19125 -2445 19130
rect -2395 19150 -2365 19155
rect -2395 19130 -2390 19150
rect -2390 19130 -2370 19150
rect -2370 19130 -2365 19150
rect -2395 19125 -2365 19130
rect -2315 19150 -2285 19155
rect -2315 19130 -2310 19150
rect -2310 19130 -2290 19150
rect -2290 19130 -2285 19150
rect -2315 19125 -2285 19130
rect -2235 19150 -2205 19155
rect -2235 19130 -2230 19150
rect -2230 19130 -2210 19150
rect -2210 19130 -2205 19150
rect -2235 19125 -2205 19130
rect -2155 19150 -2125 19155
rect -2155 19130 -2150 19150
rect -2150 19130 -2130 19150
rect -2130 19130 -2125 19150
rect -2155 19125 -2125 19130
rect -2075 19150 -2045 19155
rect -2075 19130 -2070 19150
rect -2070 19130 -2050 19150
rect -2050 19130 -2045 19150
rect -2075 19125 -2045 19130
rect -1995 19150 -1965 19155
rect -1995 19130 -1990 19150
rect -1990 19130 -1970 19150
rect -1970 19130 -1965 19150
rect -1995 19125 -1965 19130
rect -1915 19150 -1885 19155
rect -1915 19130 -1910 19150
rect -1910 19130 -1890 19150
rect -1890 19130 -1885 19150
rect -1915 19125 -1885 19130
rect -1835 19150 -1805 19155
rect -1835 19130 -1830 19150
rect -1830 19130 -1810 19150
rect -1810 19130 -1805 19150
rect -1835 19125 -1805 19130
rect -1755 19150 -1725 19155
rect -1755 19130 -1750 19150
rect -1750 19130 -1730 19150
rect -1730 19130 -1725 19150
rect -1755 19125 -1725 19130
rect -1675 19150 -1645 19155
rect -1675 19130 -1670 19150
rect -1670 19130 -1650 19150
rect -1650 19130 -1645 19150
rect -1675 19125 -1645 19130
rect -1595 19150 -1565 19155
rect -1595 19130 -1590 19150
rect -1590 19130 -1570 19150
rect -1570 19130 -1565 19150
rect -1595 19125 -1565 19130
rect -1515 19150 -1485 19155
rect -1515 19130 -1510 19150
rect -1510 19130 -1490 19150
rect -1490 19130 -1485 19150
rect -1515 19125 -1485 19130
rect -1435 19150 -1405 19155
rect -1435 19130 -1430 19150
rect -1430 19130 -1410 19150
rect -1410 19130 -1405 19150
rect -1435 19125 -1405 19130
rect -1355 19150 -1325 19155
rect -1355 19130 -1350 19150
rect -1350 19130 -1330 19150
rect -1330 19130 -1325 19150
rect -1355 19125 -1325 19130
rect -1275 19150 -1245 19155
rect -1275 19130 -1270 19150
rect -1270 19130 -1250 19150
rect -1250 19130 -1245 19150
rect -1275 19125 -1245 19130
rect -1195 19150 -1165 19155
rect -1195 19130 -1190 19150
rect -1190 19130 -1170 19150
rect -1170 19130 -1165 19150
rect -1195 19125 -1165 19130
rect -1115 19150 -1085 19155
rect -1115 19130 -1110 19150
rect -1110 19130 -1090 19150
rect -1090 19130 -1085 19150
rect -1115 19125 -1085 19130
rect -1035 19150 -1005 19155
rect -1035 19130 -1030 19150
rect -1030 19130 -1010 19150
rect -1010 19130 -1005 19150
rect -1035 19125 -1005 19130
rect -955 19150 -925 19155
rect -955 19130 -950 19150
rect -950 19130 -930 19150
rect -930 19130 -925 19150
rect -955 19125 -925 19130
rect -875 19150 -845 19155
rect -875 19130 -870 19150
rect -870 19130 -850 19150
rect -850 19130 -845 19150
rect -875 19125 -845 19130
rect -795 19150 -765 19155
rect -795 19130 -790 19150
rect -790 19130 -770 19150
rect -770 19130 -765 19150
rect -795 19125 -765 19130
rect -715 19150 -685 19155
rect -715 19130 -710 19150
rect -710 19130 -690 19150
rect -690 19130 -685 19150
rect -715 19125 -685 19130
rect -635 19150 -605 19155
rect -635 19130 -630 19150
rect -630 19130 -610 19150
rect -610 19130 -605 19150
rect -635 19125 -605 19130
rect -555 19150 -525 19155
rect -555 19130 -550 19150
rect -550 19130 -530 19150
rect -530 19130 -525 19150
rect -555 19125 -525 19130
rect -475 19150 -445 19155
rect -475 19130 -470 19150
rect -470 19130 -450 19150
rect -450 19130 -445 19150
rect -475 19125 -445 19130
rect -395 19150 -365 19155
rect -395 19130 -390 19150
rect -390 19130 -370 19150
rect -370 19130 -365 19150
rect -395 19125 -365 19130
rect -315 19150 -285 19155
rect -315 19130 -310 19150
rect -310 19130 -290 19150
rect -290 19130 -285 19150
rect -315 19125 -285 19130
rect -235 19150 -205 19155
rect -235 19130 -230 19150
rect -230 19130 -210 19150
rect -210 19130 -205 19150
rect -235 19125 -205 19130
rect -155 19150 -125 19155
rect -155 19130 -150 19150
rect -150 19130 -130 19150
rect -130 19130 -125 19150
rect -155 19125 -125 19130
rect -75 19150 -45 19155
rect -75 19130 -70 19150
rect -70 19130 -50 19150
rect -50 19130 -45 19150
rect -75 19125 -45 19130
rect 5 19150 35 19155
rect 5 19130 10 19150
rect 10 19130 30 19150
rect 30 19130 35 19150
rect 5 19125 35 19130
rect -3515 18990 -3485 18995
rect -3515 18970 -3510 18990
rect -3510 18970 -3490 18990
rect -3490 18970 -3485 18990
rect -3515 18965 -3485 18970
rect -3435 18990 -3405 18995
rect -3435 18970 -3430 18990
rect -3430 18970 -3410 18990
rect -3410 18970 -3405 18990
rect -3435 18965 -3405 18970
rect -3355 18990 -3325 18995
rect -3355 18970 -3350 18990
rect -3350 18970 -3330 18990
rect -3330 18970 -3325 18990
rect -3355 18965 -3325 18970
rect -3275 18990 -3245 18995
rect -3275 18970 -3270 18990
rect -3270 18970 -3250 18990
rect -3250 18970 -3245 18990
rect -3275 18965 -3245 18970
rect -3195 18990 -3165 18995
rect -3195 18970 -3190 18990
rect -3190 18970 -3170 18990
rect -3170 18970 -3165 18990
rect -3195 18965 -3165 18970
rect -3115 18990 -3085 18995
rect -3115 18970 -3110 18990
rect -3110 18970 -3090 18990
rect -3090 18970 -3085 18990
rect -3115 18965 -3085 18970
rect -3035 18990 -3005 18995
rect -3035 18970 -3030 18990
rect -3030 18970 -3010 18990
rect -3010 18970 -3005 18990
rect -3035 18965 -3005 18970
rect -2955 18990 -2925 18995
rect -2955 18970 -2950 18990
rect -2950 18970 -2930 18990
rect -2930 18970 -2925 18990
rect -2955 18965 -2925 18970
rect -2875 18990 -2845 18995
rect -2875 18970 -2870 18990
rect -2870 18970 -2850 18990
rect -2850 18970 -2845 18990
rect -2875 18965 -2845 18970
rect -2795 18990 -2765 18995
rect -2795 18970 -2790 18990
rect -2790 18970 -2770 18990
rect -2770 18970 -2765 18990
rect -2795 18965 -2765 18970
rect -2715 18990 -2685 18995
rect -2715 18970 -2710 18990
rect -2710 18970 -2690 18990
rect -2690 18970 -2685 18990
rect -2715 18965 -2685 18970
rect -2635 18990 -2605 18995
rect -2635 18970 -2630 18990
rect -2630 18970 -2610 18990
rect -2610 18970 -2605 18990
rect -2635 18965 -2605 18970
rect -2555 18990 -2525 18995
rect -2555 18970 -2550 18990
rect -2550 18970 -2530 18990
rect -2530 18970 -2525 18990
rect -2555 18965 -2525 18970
rect -2475 18990 -2445 18995
rect -2475 18970 -2470 18990
rect -2470 18970 -2450 18990
rect -2450 18970 -2445 18990
rect -2475 18965 -2445 18970
rect -2395 18990 -2365 18995
rect -2395 18970 -2390 18990
rect -2390 18970 -2370 18990
rect -2370 18970 -2365 18990
rect -2395 18965 -2365 18970
rect -2315 18990 -2285 18995
rect -2315 18970 -2310 18990
rect -2310 18970 -2290 18990
rect -2290 18970 -2285 18990
rect -2315 18965 -2285 18970
rect -2235 18990 -2205 18995
rect -2235 18970 -2230 18990
rect -2230 18970 -2210 18990
rect -2210 18970 -2205 18990
rect -2235 18965 -2205 18970
rect -2155 18990 -2125 18995
rect -2155 18970 -2150 18990
rect -2150 18970 -2130 18990
rect -2130 18970 -2125 18990
rect -2155 18965 -2125 18970
rect -2075 18990 -2045 18995
rect -2075 18970 -2070 18990
rect -2070 18970 -2050 18990
rect -2050 18970 -2045 18990
rect -2075 18965 -2045 18970
rect -1995 18990 -1965 18995
rect -1995 18970 -1990 18990
rect -1990 18970 -1970 18990
rect -1970 18970 -1965 18990
rect -1995 18965 -1965 18970
rect -1915 18990 -1885 18995
rect -1915 18970 -1910 18990
rect -1910 18970 -1890 18990
rect -1890 18970 -1885 18990
rect -1915 18965 -1885 18970
rect -1835 18990 -1805 18995
rect -1835 18970 -1830 18990
rect -1830 18970 -1810 18990
rect -1810 18970 -1805 18990
rect -1835 18965 -1805 18970
rect -1755 18990 -1725 18995
rect -1755 18970 -1750 18990
rect -1750 18970 -1730 18990
rect -1730 18970 -1725 18990
rect -1755 18965 -1725 18970
rect -1675 18990 -1645 18995
rect -1675 18970 -1670 18990
rect -1670 18970 -1650 18990
rect -1650 18970 -1645 18990
rect -1675 18965 -1645 18970
rect -1595 18990 -1565 18995
rect -1595 18970 -1590 18990
rect -1590 18970 -1570 18990
rect -1570 18970 -1565 18990
rect -1595 18965 -1565 18970
rect -1515 18990 -1485 18995
rect -1515 18970 -1510 18990
rect -1510 18970 -1490 18990
rect -1490 18970 -1485 18990
rect -1515 18965 -1485 18970
rect -1435 18990 -1405 18995
rect -1435 18970 -1430 18990
rect -1430 18970 -1410 18990
rect -1410 18970 -1405 18990
rect -1435 18965 -1405 18970
rect -1355 18990 -1325 18995
rect -1355 18970 -1350 18990
rect -1350 18970 -1330 18990
rect -1330 18970 -1325 18990
rect -1355 18965 -1325 18970
rect -1275 18990 -1245 18995
rect -1275 18970 -1270 18990
rect -1270 18970 -1250 18990
rect -1250 18970 -1245 18990
rect -1275 18965 -1245 18970
rect -1195 18990 -1165 18995
rect -1195 18970 -1190 18990
rect -1190 18970 -1170 18990
rect -1170 18970 -1165 18990
rect -1195 18965 -1165 18970
rect -1115 18990 -1085 18995
rect -1115 18970 -1110 18990
rect -1110 18970 -1090 18990
rect -1090 18970 -1085 18990
rect -1115 18965 -1085 18970
rect -1035 18990 -1005 18995
rect -1035 18970 -1030 18990
rect -1030 18970 -1010 18990
rect -1010 18970 -1005 18990
rect -1035 18965 -1005 18970
rect -955 18990 -925 18995
rect -955 18970 -950 18990
rect -950 18970 -930 18990
rect -930 18970 -925 18990
rect -955 18965 -925 18970
rect -875 18990 -845 18995
rect -875 18970 -870 18990
rect -870 18970 -850 18990
rect -850 18970 -845 18990
rect -875 18965 -845 18970
rect -795 18990 -765 18995
rect -795 18970 -790 18990
rect -790 18970 -770 18990
rect -770 18970 -765 18990
rect -795 18965 -765 18970
rect -715 18990 -685 18995
rect -715 18970 -710 18990
rect -710 18970 -690 18990
rect -690 18970 -685 18990
rect -715 18965 -685 18970
rect -635 18990 -605 18995
rect -635 18970 -630 18990
rect -630 18970 -610 18990
rect -610 18970 -605 18990
rect -635 18965 -605 18970
rect -555 18990 -525 18995
rect -555 18970 -550 18990
rect -550 18970 -530 18990
rect -530 18970 -525 18990
rect -555 18965 -525 18970
rect -475 18990 -445 18995
rect -475 18970 -470 18990
rect -470 18970 -450 18990
rect -450 18970 -445 18990
rect -475 18965 -445 18970
rect -395 18990 -365 18995
rect -395 18970 -390 18990
rect -390 18970 -370 18990
rect -370 18970 -365 18990
rect -395 18965 -365 18970
rect -315 18990 -285 18995
rect -315 18970 -310 18990
rect -310 18970 -290 18990
rect -290 18970 -285 18990
rect -315 18965 -285 18970
rect -235 18990 -205 18995
rect -235 18970 -230 18990
rect -230 18970 -210 18990
rect -210 18970 -205 18990
rect -235 18965 -205 18970
rect -155 18990 -125 18995
rect -155 18970 -150 18990
rect -150 18970 -130 18990
rect -130 18970 -125 18990
rect -155 18965 -125 18970
rect -75 18990 -45 18995
rect -75 18970 -70 18990
rect -70 18970 -50 18990
rect -50 18970 -45 18990
rect -75 18965 -45 18970
rect 5 18990 35 18995
rect 5 18970 10 18990
rect 10 18970 30 18990
rect 30 18970 35 18990
rect 5 18965 35 18970
rect -3515 18830 -3485 18835
rect -3515 18810 -3510 18830
rect -3510 18810 -3490 18830
rect -3490 18810 -3485 18830
rect -3515 18805 -3485 18810
rect -3435 18830 -3405 18835
rect -3435 18810 -3430 18830
rect -3430 18810 -3410 18830
rect -3410 18810 -3405 18830
rect -3435 18805 -3405 18810
rect -3355 18830 -3325 18835
rect -3355 18810 -3350 18830
rect -3350 18810 -3330 18830
rect -3330 18810 -3325 18830
rect -3355 18805 -3325 18810
rect -3275 18830 -3245 18835
rect -3275 18810 -3270 18830
rect -3270 18810 -3250 18830
rect -3250 18810 -3245 18830
rect -3275 18805 -3245 18810
rect -3195 18830 -3165 18835
rect -3195 18810 -3190 18830
rect -3190 18810 -3170 18830
rect -3170 18810 -3165 18830
rect -3195 18805 -3165 18810
rect -3115 18830 -3085 18835
rect -3115 18810 -3110 18830
rect -3110 18810 -3090 18830
rect -3090 18810 -3085 18830
rect -3115 18805 -3085 18810
rect -3035 18830 -3005 18835
rect -3035 18810 -3030 18830
rect -3030 18810 -3010 18830
rect -3010 18810 -3005 18830
rect -3035 18805 -3005 18810
rect -2955 18830 -2925 18835
rect -2955 18810 -2950 18830
rect -2950 18810 -2930 18830
rect -2930 18810 -2925 18830
rect -2955 18805 -2925 18810
rect -2875 18830 -2845 18835
rect -2875 18810 -2870 18830
rect -2870 18810 -2850 18830
rect -2850 18810 -2845 18830
rect -2875 18805 -2845 18810
rect -2795 18830 -2765 18835
rect -2795 18810 -2790 18830
rect -2790 18810 -2770 18830
rect -2770 18810 -2765 18830
rect -2795 18805 -2765 18810
rect -2715 18830 -2685 18835
rect -2715 18810 -2710 18830
rect -2710 18810 -2690 18830
rect -2690 18810 -2685 18830
rect -2715 18805 -2685 18810
rect -2635 18830 -2605 18835
rect -2635 18810 -2630 18830
rect -2630 18810 -2610 18830
rect -2610 18810 -2605 18830
rect -2635 18805 -2605 18810
rect -2555 18830 -2525 18835
rect -2555 18810 -2550 18830
rect -2550 18810 -2530 18830
rect -2530 18810 -2525 18830
rect -2555 18805 -2525 18810
rect -2475 18830 -2445 18835
rect -2475 18810 -2470 18830
rect -2470 18810 -2450 18830
rect -2450 18810 -2445 18830
rect -2475 18805 -2445 18810
rect -2395 18830 -2365 18835
rect -2395 18810 -2390 18830
rect -2390 18810 -2370 18830
rect -2370 18810 -2365 18830
rect -2395 18805 -2365 18810
rect -2315 18830 -2285 18835
rect -2315 18810 -2310 18830
rect -2310 18810 -2290 18830
rect -2290 18810 -2285 18830
rect -2315 18805 -2285 18810
rect -2235 18830 -2205 18835
rect -2235 18810 -2230 18830
rect -2230 18810 -2210 18830
rect -2210 18810 -2205 18830
rect -2235 18805 -2205 18810
rect -2155 18830 -2125 18835
rect -2155 18810 -2150 18830
rect -2150 18810 -2130 18830
rect -2130 18810 -2125 18830
rect -2155 18805 -2125 18810
rect -2075 18830 -2045 18835
rect -2075 18810 -2070 18830
rect -2070 18810 -2050 18830
rect -2050 18810 -2045 18830
rect -2075 18805 -2045 18810
rect -1995 18830 -1965 18835
rect -1995 18810 -1990 18830
rect -1990 18810 -1970 18830
rect -1970 18810 -1965 18830
rect -1995 18805 -1965 18810
rect -1915 18830 -1885 18835
rect -1915 18810 -1910 18830
rect -1910 18810 -1890 18830
rect -1890 18810 -1885 18830
rect -1915 18805 -1885 18810
rect -1835 18830 -1805 18835
rect -1835 18810 -1830 18830
rect -1830 18810 -1810 18830
rect -1810 18810 -1805 18830
rect -1835 18805 -1805 18810
rect -1755 18830 -1725 18835
rect -1755 18810 -1750 18830
rect -1750 18810 -1730 18830
rect -1730 18810 -1725 18830
rect -1755 18805 -1725 18810
rect -1675 18830 -1645 18835
rect -1675 18810 -1670 18830
rect -1670 18810 -1650 18830
rect -1650 18810 -1645 18830
rect -1675 18805 -1645 18810
rect -1595 18830 -1565 18835
rect -1595 18810 -1590 18830
rect -1590 18810 -1570 18830
rect -1570 18810 -1565 18830
rect -1595 18805 -1565 18810
rect -1515 18830 -1485 18835
rect -1515 18810 -1510 18830
rect -1510 18810 -1490 18830
rect -1490 18810 -1485 18830
rect -1515 18805 -1485 18810
rect -1435 18830 -1405 18835
rect -1435 18810 -1430 18830
rect -1430 18810 -1410 18830
rect -1410 18810 -1405 18830
rect -1435 18805 -1405 18810
rect -1355 18830 -1325 18835
rect -1355 18810 -1350 18830
rect -1350 18810 -1330 18830
rect -1330 18810 -1325 18830
rect -1355 18805 -1325 18810
rect -1275 18830 -1245 18835
rect -1275 18810 -1270 18830
rect -1270 18810 -1250 18830
rect -1250 18810 -1245 18830
rect -1275 18805 -1245 18810
rect -1195 18830 -1165 18835
rect -1195 18810 -1190 18830
rect -1190 18810 -1170 18830
rect -1170 18810 -1165 18830
rect -1195 18805 -1165 18810
rect -1115 18830 -1085 18835
rect -1115 18810 -1110 18830
rect -1110 18810 -1090 18830
rect -1090 18810 -1085 18830
rect -1115 18805 -1085 18810
rect -1035 18830 -1005 18835
rect -1035 18810 -1030 18830
rect -1030 18810 -1010 18830
rect -1010 18810 -1005 18830
rect -1035 18805 -1005 18810
rect -955 18830 -925 18835
rect -955 18810 -950 18830
rect -950 18810 -930 18830
rect -930 18810 -925 18830
rect -955 18805 -925 18810
rect -875 18830 -845 18835
rect -875 18810 -870 18830
rect -870 18810 -850 18830
rect -850 18810 -845 18830
rect -875 18805 -845 18810
rect -795 18830 -765 18835
rect -795 18810 -790 18830
rect -790 18810 -770 18830
rect -770 18810 -765 18830
rect -795 18805 -765 18810
rect -715 18830 -685 18835
rect -715 18810 -710 18830
rect -710 18810 -690 18830
rect -690 18810 -685 18830
rect -715 18805 -685 18810
rect -635 18830 -605 18835
rect -635 18810 -630 18830
rect -630 18810 -610 18830
rect -610 18810 -605 18830
rect -635 18805 -605 18810
rect -555 18830 -525 18835
rect -555 18810 -550 18830
rect -550 18810 -530 18830
rect -530 18810 -525 18830
rect -555 18805 -525 18810
rect -475 18830 -445 18835
rect -475 18810 -470 18830
rect -470 18810 -450 18830
rect -450 18810 -445 18830
rect -475 18805 -445 18810
rect -395 18830 -365 18835
rect -395 18810 -390 18830
rect -390 18810 -370 18830
rect -370 18810 -365 18830
rect -395 18805 -365 18810
rect -315 18830 -285 18835
rect -315 18810 -310 18830
rect -310 18810 -290 18830
rect -290 18810 -285 18830
rect -315 18805 -285 18810
rect -235 18830 -205 18835
rect -235 18810 -230 18830
rect -230 18810 -210 18830
rect -210 18810 -205 18830
rect -235 18805 -205 18810
rect -155 18830 -125 18835
rect -155 18810 -150 18830
rect -150 18810 -130 18830
rect -130 18810 -125 18830
rect -155 18805 -125 18810
rect -75 18830 -45 18835
rect -75 18810 -70 18830
rect -70 18810 -50 18830
rect -50 18810 -45 18830
rect -75 18805 -45 18810
rect 5 18830 35 18835
rect 5 18810 10 18830
rect 10 18810 30 18830
rect 30 18810 35 18830
rect 5 18805 35 18810
rect 38365 18310 38395 18315
rect 38365 18290 38370 18310
rect 38370 18290 38390 18310
rect 38390 18290 38395 18310
rect 38365 18285 38395 18290
rect 38445 18310 38475 18315
rect 38445 18290 38450 18310
rect 38450 18290 38470 18310
rect 38470 18290 38475 18310
rect 38445 18285 38475 18290
rect 38365 18150 38395 18155
rect 38365 18130 38370 18150
rect 38370 18130 38390 18150
rect 38390 18130 38395 18150
rect 38365 18125 38395 18130
rect 38445 18150 38475 18155
rect 38445 18130 38450 18150
rect 38450 18130 38470 18150
rect 38470 18130 38475 18150
rect 38445 18125 38475 18130
rect -1275 17630 -1245 17635
rect -1275 17610 -1270 17630
rect -1270 17610 -1250 17630
rect -1250 17610 -1245 17630
rect -1275 17605 -1245 17610
rect -1195 17630 -1165 17635
rect -1195 17610 -1190 17630
rect -1190 17610 -1170 17630
rect -1170 17610 -1165 17630
rect -1195 17605 -1165 17610
rect -1115 17630 -1085 17635
rect -1115 17610 -1110 17630
rect -1110 17610 -1090 17630
rect -1090 17610 -1085 17630
rect -1115 17605 -1085 17610
rect -1035 17630 -1005 17635
rect -1035 17610 -1030 17630
rect -1030 17610 -1010 17630
rect -1010 17610 -1005 17630
rect -1035 17605 -1005 17610
rect -955 17630 -925 17635
rect -955 17610 -950 17630
rect -950 17610 -930 17630
rect -930 17610 -925 17630
rect -955 17605 -925 17610
rect -875 17630 -845 17635
rect -875 17610 -870 17630
rect -870 17610 -850 17630
rect -850 17610 -845 17630
rect -875 17605 -845 17610
rect -795 17630 -765 17635
rect -795 17610 -790 17630
rect -790 17610 -770 17630
rect -770 17610 -765 17630
rect -795 17605 -765 17610
rect -715 17630 -685 17635
rect -715 17610 -710 17630
rect -710 17610 -690 17630
rect -690 17610 -685 17630
rect -715 17605 -685 17610
rect -635 17630 -605 17635
rect -635 17610 -630 17630
rect -630 17610 -610 17630
rect -610 17610 -605 17630
rect -635 17605 -605 17610
rect -555 17630 -525 17635
rect -555 17610 -550 17630
rect -550 17610 -530 17630
rect -530 17610 -525 17630
rect -555 17605 -525 17610
rect -475 17630 -445 17635
rect -475 17610 -470 17630
rect -470 17610 -450 17630
rect -450 17610 -445 17630
rect -475 17605 -445 17610
rect -395 17630 -365 17635
rect -395 17610 -390 17630
rect -390 17610 -370 17630
rect -370 17610 -365 17630
rect -395 17605 -365 17610
rect -315 17630 -285 17635
rect -315 17610 -310 17630
rect -310 17610 -290 17630
rect -290 17610 -285 17630
rect -315 17605 -285 17610
rect -235 17630 -205 17635
rect -235 17610 -230 17630
rect -230 17610 -210 17630
rect -210 17610 -205 17630
rect -235 17605 -205 17610
rect -155 17630 -125 17635
rect -155 17610 -150 17630
rect -150 17610 -130 17630
rect -130 17610 -125 17630
rect -155 17605 -125 17610
rect -75 17630 -45 17635
rect -75 17610 -70 17630
rect -70 17610 -50 17630
rect -50 17610 -45 17630
rect -75 17605 -45 17610
rect 5 17630 35 17635
rect 5 17610 10 17630
rect 10 17610 30 17630
rect 30 17610 35 17630
rect 5 17605 35 17610
rect -1275 17470 -1245 17475
rect -1275 17450 -1270 17470
rect -1270 17450 -1250 17470
rect -1250 17450 -1245 17470
rect -1275 17445 -1245 17450
rect -1195 17470 -1165 17475
rect -1195 17450 -1190 17470
rect -1190 17450 -1170 17470
rect -1170 17450 -1165 17470
rect -1195 17445 -1165 17450
rect -1115 17470 -1085 17475
rect -1115 17450 -1110 17470
rect -1110 17450 -1090 17470
rect -1090 17450 -1085 17470
rect -1115 17445 -1085 17450
rect -1035 17470 -1005 17475
rect -1035 17450 -1030 17470
rect -1030 17450 -1010 17470
rect -1010 17450 -1005 17470
rect -1035 17445 -1005 17450
rect -955 17470 -925 17475
rect -955 17450 -950 17470
rect -950 17450 -930 17470
rect -930 17450 -925 17470
rect -955 17445 -925 17450
rect -875 17470 -845 17475
rect -875 17450 -870 17470
rect -870 17450 -850 17470
rect -850 17450 -845 17470
rect -875 17445 -845 17450
rect -795 17470 -765 17475
rect -795 17450 -790 17470
rect -790 17450 -770 17470
rect -770 17450 -765 17470
rect -795 17445 -765 17450
rect -715 17470 -685 17475
rect -715 17450 -710 17470
rect -710 17450 -690 17470
rect -690 17450 -685 17470
rect -715 17445 -685 17450
rect -635 17470 -605 17475
rect -635 17450 -630 17470
rect -630 17450 -610 17470
rect -610 17450 -605 17470
rect -635 17445 -605 17450
rect -555 17470 -525 17475
rect -555 17450 -550 17470
rect -550 17450 -530 17470
rect -530 17450 -525 17470
rect -555 17445 -525 17450
rect -475 17470 -445 17475
rect -475 17450 -470 17470
rect -470 17450 -450 17470
rect -450 17450 -445 17470
rect -475 17445 -445 17450
rect -395 17470 -365 17475
rect -395 17450 -390 17470
rect -390 17450 -370 17470
rect -370 17450 -365 17470
rect -395 17445 -365 17450
rect -315 17470 -285 17475
rect -315 17450 -310 17470
rect -310 17450 -290 17470
rect -290 17450 -285 17470
rect -315 17445 -285 17450
rect -235 17470 -205 17475
rect -235 17450 -230 17470
rect -230 17450 -210 17470
rect -210 17450 -205 17470
rect -235 17445 -205 17450
rect -155 17470 -125 17475
rect -155 17450 -150 17470
rect -150 17450 -130 17470
rect -130 17450 -125 17470
rect -155 17445 -125 17450
rect -75 17470 -45 17475
rect -75 17450 -70 17470
rect -70 17450 -50 17470
rect -50 17450 -45 17470
rect -75 17445 -45 17450
rect 5 17470 35 17475
rect 5 17450 10 17470
rect 10 17450 30 17470
rect 30 17450 35 17470
rect 5 17445 35 17450
<< metal2 >>
rect 38440 22235 38720 22240
rect 38440 22205 38445 22235
rect 38475 22205 38720 22235
rect 38440 22200 38720 22205
rect 38520 21835 38720 21840
rect 38520 21805 38525 21835
rect 38555 21805 38685 21835
rect 38715 21805 38720 21835
rect 38520 21800 38720 21805
rect 38600 21755 38720 21760
rect 38600 21725 38605 21755
rect 38635 21725 38720 21755
rect 38600 21720 38720 21725
rect 38520 21675 38720 21680
rect 38520 21645 38525 21675
rect 38555 21645 38685 21675
rect 38715 21645 38720 21675
rect 38520 21640 38720 21645
rect 38520 21595 38720 21600
rect 38520 21565 38525 21595
rect 38555 21565 38685 21595
rect 38715 21565 38720 21595
rect 38520 21560 38720 21565
rect 38520 21515 38720 21520
rect 38520 21485 38525 21515
rect 38555 21485 38685 21515
rect 38715 21485 38720 21515
rect 38520 21480 38720 21485
rect 38520 21435 38720 21440
rect 38520 21405 38525 21435
rect 38555 21405 38685 21435
rect 38715 21405 38720 21435
rect 38520 21400 38720 21405
rect 38520 21355 38720 21360
rect 38520 21325 38525 21355
rect 38555 21325 38685 21355
rect 38715 21325 38720 21355
rect 38520 21320 38720 21325
rect 63320 21320 63520 21360
rect 38600 21275 38720 21280
rect 38600 21245 38605 21275
rect 38635 21245 38720 21275
rect 38600 21240 38720 21245
rect 63320 21200 63360 21320
rect 63480 21200 63520 21320
rect 38520 21195 38720 21200
rect 38520 21165 38525 21195
rect 38555 21165 38685 21195
rect 38715 21165 38720 21195
rect 38520 21160 38720 21165
rect 63320 21160 63520 21200
rect -720 20920 -520 20960
rect -480 20955 80 20960
rect -480 20925 -475 20955
rect -445 20925 -395 20955
rect -365 20925 -315 20955
rect -285 20925 -235 20955
rect -205 20925 -155 20955
rect -125 20925 -75 20955
rect -45 20925 5 20955
rect 35 20925 80 20955
rect -480 20920 80 20925
rect -720 20800 -680 20920
rect -560 20880 -520 20920
rect -560 20840 40 20880
rect 38320 20875 38480 20880
rect 38320 20845 38445 20875
rect 38475 20845 38480 20875
rect 38320 20840 38480 20845
rect 38520 20875 38720 20880
rect 38520 20845 38525 20875
rect 38555 20845 38685 20875
rect 38715 20845 38720 20875
rect 38520 20840 38720 20845
rect -560 20800 -520 20840
rect -720 20760 -520 20800
rect -480 20795 80 20800
rect -480 20765 -475 20795
rect -445 20765 -395 20795
rect -365 20765 -315 20795
rect -285 20765 -235 20795
rect -205 20765 -155 20795
rect -125 20765 -75 20795
rect -45 20765 5 20795
rect 35 20765 80 20795
rect -480 20760 80 20765
rect 38600 20795 38720 20800
rect 38600 20765 38605 20795
rect 38635 20765 38720 20795
rect 38600 20760 38720 20765
rect 38520 20715 38720 20720
rect 38520 20685 38525 20715
rect 38555 20685 38685 20715
rect 38715 20685 38720 20715
rect 38520 20680 38720 20685
rect 38520 20635 38720 20640
rect 38520 20605 38525 20635
rect 38555 20605 38685 20635
rect 38715 20605 38720 20635
rect 38520 20600 38720 20605
rect 38520 20555 38720 20560
rect 38520 20525 38525 20555
rect 38555 20525 38685 20555
rect 38715 20525 38720 20555
rect 38520 20520 38720 20525
rect 38520 20475 38720 20480
rect 38520 20445 38525 20475
rect 38555 20445 38685 20475
rect 38715 20445 38720 20475
rect 38520 20440 38720 20445
rect 38520 20395 38720 20400
rect 38520 20365 38525 20395
rect 38555 20365 38685 20395
rect 38715 20365 38720 20395
rect 38520 20360 38720 20365
rect 38240 20315 38720 20320
rect 38240 20285 38365 20315
rect 38395 20285 38445 20315
rect 38475 20285 38525 20315
rect 38555 20285 38685 20315
rect 38715 20285 38720 20315
rect 38240 20280 38720 20285
rect 38320 20235 38720 20240
rect 38320 20205 38605 20235
rect 38635 20205 38720 20235
rect 38320 20200 38720 20205
rect 38240 20155 38720 20160
rect 38240 20125 38365 20155
rect 38395 20125 38445 20155
rect 38475 20125 38525 20155
rect 38555 20125 38685 20155
rect 38715 20125 38720 20155
rect 38240 20120 38720 20125
rect -3520 19155 80 19160
rect -3520 19125 -3515 19155
rect -3485 19125 -3435 19155
rect -3405 19125 -3355 19155
rect -3325 19125 -3275 19155
rect -3245 19125 -3195 19155
rect -3165 19125 -3115 19155
rect -3085 19125 -3035 19155
rect -3005 19125 -2955 19155
rect -2925 19125 -2875 19155
rect -2845 19125 -2795 19155
rect -2765 19125 -2715 19155
rect -2685 19125 -2635 19155
rect -2605 19125 -2555 19155
rect -2525 19125 -2475 19155
rect -2445 19125 -2395 19155
rect -2365 19125 -2315 19155
rect -2285 19125 -2235 19155
rect -2205 19125 -2155 19155
rect -2125 19125 -2075 19155
rect -2045 19125 -1995 19155
rect -1965 19125 -1915 19155
rect -1885 19125 -1835 19155
rect -1805 19125 -1755 19155
rect -1725 19125 -1675 19155
rect -1645 19125 -1595 19155
rect -1565 19125 -1515 19155
rect -1485 19125 -1435 19155
rect -1405 19125 -1355 19155
rect -1325 19125 -1275 19155
rect -1245 19125 -1195 19155
rect -1165 19125 -1115 19155
rect -1085 19125 -1035 19155
rect -1005 19125 -955 19155
rect -925 19125 -875 19155
rect -845 19125 -795 19155
rect -765 19125 -715 19155
rect -685 19125 -635 19155
rect -605 19125 -555 19155
rect -525 19125 -475 19155
rect -445 19125 -395 19155
rect -365 19125 -315 19155
rect -285 19125 -235 19155
rect -205 19125 -155 19155
rect -125 19125 -75 19155
rect -45 19125 5 19155
rect 35 19125 80 19155
rect -3520 19120 80 19125
rect -3520 19075 40 19080
rect -3520 19045 -3035 19075
rect -3005 19045 40 19075
rect -3520 19040 40 19045
rect -3520 18995 80 19000
rect -3520 18965 -3515 18995
rect -3485 18965 -3435 18995
rect -3405 18965 -3355 18995
rect -3325 18965 -3275 18995
rect -3245 18965 -3195 18995
rect -3165 18965 -3115 18995
rect -3085 18965 -3035 18995
rect -3005 18965 -2955 18995
rect -2925 18965 -2875 18995
rect -2845 18965 -2795 18995
rect -2765 18965 -2715 18995
rect -2685 18965 -2635 18995
rect -2605 18965 -2555 18995
rect -2525 18965 -2475 18995
rect -2445 18965 -2395 18995
rect -2365 18965 -2315 18995
rect -2285 18965 -2235 18995
rect -2205 18965 -2155 18995
rect -2125 18965 -2075 18995
rect -2045 18965 -1995 18995
rect -1965 18965 -1915 18995
rect -1885 18965 -1835 18995
rect -1805 18965 -1755 18995
rect -1725 18965 -1675 18995
rect -1645 18965 -1595 18995
rect -1565 18965 -1515 18995
rect -1485 18965 -1435 18995
rect -1405 18965 -1355 18995
rect -1325 18965 -1275 18995
rect -1245 18965 -1195 18995
rect -1165 18965 -1115 18995
rect -1085 18965 -1035 18995
rect -1005 18965 -955 18995
rect -925 18965 -875 18995
rect -845 18965 -795 18995
rect -765 18965 -715 18995
rect -685 18965 -635 18995
rect -605 18965 -555 18995
rect -525 18965 -475 18995
rect -445 18965 -395 18995
rect -365 18965 -315 18995
rect -285 18965 -235 18995
rect -205 18965 -155 18995
rect -125 18965 -75 18995
rect -45 18965 5 18995
rect 35 18965 80 18995
rect -3520 18960 80 18965
rect -3520 18915 40 18920
rect -3520 18885 -2235 18915
rect -2205 18885 40 18915
rect -3520 18880 40 18885
rect -3520 18835 80 18840
rect -3520 18805 -3515 18835
rect -3485 18805 -3435 18835
rect -3405 18805 -3355 18835
rect -3325 18805 -3275 18835
rect -3245 18805 -3195 18835
rect -3165 18805 -3115 18835
rect -3085 18805 -3035 18835
rect -3005 18805 -2955 18835
rect -2925 18805 -2875 18835
rect -2845 18805 -2795 18835
rect -2765 18805 -2715 18835
rect -2685 18805 -2635 18835
rect -2605 18805 -2555 18835
rect -2525 18805 -2475 18835
rect -2445 18805 -2395 18835
rect -2365 18805 -2315 18835
rect -2285 18805 -2235 18835
rect -2205 18805 -2155 18835
rect -2125 18805 -2075 18835
rect -2045 18805 -1995 18835
rect -1965 18805 -1915 18835
rect -1885 18805 -1835 18835
rect -1805 18805 -1755 18835
rect -1725 18805 -1675 18835
rect -1645 18805 -1595 18835
rect -1565 18805 -1515 18835
rect -1485 18805 -1435 18835
rect -1405 18805 -1355 18835
rect -1325 18805 -1275 18835
rect -1245 18805 -1195 18835
rect -1165 18805 -1115 18835
rect -1085 18805 -1035 18835
rect -1005 18805 -955 18835
rect -925 18805 -875 18835
rect -845 18805 -795 18835
rect -765 18805 -715 18835
rect -685 18805 -635 18835
rect -605 18805 -555 18835
rect -525 18805 -475 18835
rect -445 18805 -395 18835
rect -365 18805 -315 18835
rect -285 18805 -235 18835
rect -205 18805 -155 18835
rect -125 18805 -75 18835
rect -45 18805 5 18835
rect 35 18805 80 18835
rect -3520 18800 80 18805
rect 38520 18475 38720 18480
rect 38520 18445 38525 18475
rect 38555 18445 38685 18475
rect 38715 18445 38720 18475
rect 38520 18440 38720 18445
rect 38600 18395 38720 18400
rect 38600 18365 38605 18395
rect 38635 18365 38720 18395
rect 38600 18360 38720 18365
rect 38240 18315 38720 18320
rect 38240 18285 38365 18315
rect 38395 18285 38445 18315
rect 38475 18285 38525 18315
rect 38555 18285 38685 18315
rect 38715 18285 38720 18315
rect 38240 18280 38720 18285
rect 38320 18235 38640 18240
rect 38320 18205 38605 18235
rect 38635 18205 38640 18235
rect 38320 18200 38640 18205
rect 38240 18155 38720 18160
rect 38240 18125 38365 18155
rect 38395 18125 38445 18155
rect 38475 18125 38525 18155
rect 38555 18125 38685 18155
rect 38715 18125 38720 18155
rect 38240 18120 38720 18125
rect 38520 17995 38720 18000
rect 38520 17965 38525 17995
rect 38555 17965 38685 17995
rect 38715 17965 38720 17995
rect 38520 17960 38720 17965
rect 63320 17960 63520 18000
rect 38600 17915 38720 17920
rect 38600 17885 38605 17915
rect 38635 17885 38720 17915
rect 38600 17880 38720 17885
rect 63320 17840 63360 17960
rect 63480 17840 63520 17960
rect 38520 17835 38720 17840
rect 38520 17805 38525 17835
rect 38555 17805 38685 17835
rect 38715 17805 38720 17835
rect 38520 17800 38720 17805
rect 63320 17800 63520 17840
rect 38520 17755 38720 17760
rect 38520 17725 38525 17755
rect 38555 17725 38685 17755
rect 38715 17725 38720 17755
rect 38520 17720 38720 17725
rect 38520 17675 38720 17680
rect 38520 17645 38525 17675
rect 38555 17645 38685 17675
rect 38715 17645 38720 17675
rect 38520 17640 38720 17645
rect -1520 17600 -1320 17640
rect -1280 17635 80 17640
rect -1280 17605 -1275 17635
rect -1245 17605 -1195 17635
rect -1165 17605 -1115 17635
rect -1085 17605 -1035 17635
rect -1005 17605 -955 17635
rect -925 17605 -875 17635
rect -845 17605 -795 17635
rect -765 17605 -715 17635
rect -685 17605 -635 17635
rect -605 17605 -555 17635
rect -525 17605 -475 17635
rect -445 17605 -395 17635
rect -365 17605 -315 17635
rect -285 17605 -235 17635
rect -205 17605 -155 17635
rect -125 17605 -75 17635
rect -45 17605 5 17635
rect 35 17605 80 17635
rect -1280 17600 80 17605
rect -1520 17480 -1480 17600
rect -1360 17560 -1320 17600
rect 38520 17595 38720 17600
rect 38520 17565 38525 17595
rect 38555 17565 38685 17595
rect 38715 17565 38720 17595
rect 38520 17560 38720 17565
rect -1360 17520 40 17560
rect -1360 17480 -1320 17520
rect 38520 17515 38720 17520
rect 38520 17485 38525 17515
rect 38555 17485 38685 17515
rect 38715 17485 38720 17515
rect 38520 17480 38720 17485
rect -1520 17440 -1320 17480
rect -1280 17475 80 17480
rect -1280 17445 -1275 17475
rect -1245 17445 -1195 17475
rect -1165 17445 -1115 17475
rect -1085 17445 -1035 17475
rect -1005 17445 -955 17475
rect -925 17445 -875 17475
rect -845 17445 -795 17475
rect -765 17445 -715 17475
rect -685 17445 -635 17475
rect -605 17445 -555 17475
rect -525 17445 -475 17475
rect -445 17445 -395 17475
rect -365 17445 -315 17475
rect -285 17445 -235 17475
rect -205 17445 -155 17475
rect -125 17445 -75 17475
rect -45 17445 5 17475
rect 35 17445 80 17475
rect -1280 17440 80 17445
rect 38600 17435 38720 17440
rect 38600 17405 38605 17435
rect 38635 17405 38720 17435
rect 38600 17400 38720 17405
rect 38520 17355 38720 17360
rect 38520 17325 38525 17355
rect 38555 17325 38685 17355
rect 38715 17325 38720 17355
rect 38520 17320 38720 17325
<< via2 >>
rect 38445 22205 38475 22235
rect 38525 21805 38555 21835
rect 38685 21805 38715 21835
rect 38605 21725 38635 21755
rect 38525 21645 38555 21675
rect 38685 21645 38715 21675
rect 38525 21565 38555 21595
rect 38685 21565 38715 21595
rect 38525 21485 38555 21515
rect 38685 21485 38715 21515
rect 38525 21405 38555 21435
rect 38685 21405 38715 21435
rect 38525 21325 38555 21355
rect 38685 21325 38715 21355
rect 38605 21245 38635 21275
rect 63360 21200 63480 21320
rect 38525 21165 38555 21195
rect 38685 21165 38715 21195
rect -475 20925 -445 20955
rect -395 20925 -365 20955
rect -315 20925 -285 20955
rect -235 20925 -205 20955
rect -155 20925 -125 20955
rect -75 20925 -45 20955
rect 5 20925 35 20955
rect -680 20800 -560 20920
rect 38445 20845 38475 20875
rect 38525 20845 38555 20875
rect 38685 20845 38715 20875
rect -475 20765 -445 20795
rect -395 20765 -365 20795
rect -315 20765 -285 20795
rect -235 20765 -205 20795
rect -155 20765 -125 20795
rect -75 20765 -45 20795
rect 5 20765 35 20795
rect 38605 20765 38635 20795
rect 38525 20685 38555 20715
rect 38685 20685 38715 20715
rect 38525 20605 38555 20635
rect 38685 20605 38715 20635
rect 38525 20525 38555 20555
rect 38685 20525 38715 20555
rect 38525 20445 38555 20475
rect 38685 20445 38715 20475
rect 38525 20365 38555 20395
rect 38685 20365 38715 20395
rect 38365 20285 38395 20315
rect 38445 20285 38475 20315
rect 38525 20285 38555 20315
rect 38685 20285 38715 20315
rect 38605 20205 38635 20235
rect 38365 20125 38395 20155
rect 38445 20125 38475 20155
rect 38525 20125 38555 20155
rect 38685 20125 38715 20155
rect -3515 19125 -3485 19155
rect -3435 19125 -3405 19155
rect -3355 19125 -3325 19155
rect -3275 19125 -3245 19155
rect -3195 19125 -3165 19155
rect -2875 19125 -2845 19155
rect -2795 19125 -2765 19155
rect -2715 19125 -2685 19155
rect -2635 19125 -2605 19155
rect -2555 19125 -2525 19155
rect -2475 19125 -2445 19155
rect -2395 19125 -2365 19155
rect -2075 19125 -2045 19155
rect -1995 19125 -1965 19155
rect -1915 19125 -1885 19155
rect -1835 19125 -1805 19155
rect -1755 19125 -1725 19155
rect -1675 19125 -1645 19155
rect -1595 19125 -1565 19155
rect -1515 19125 -1485 19155
rect -1435 19125 -1405 19155
rect -1355 19125 -1325 19155
rect -1275 19125 -1245 19155
rect -1195 19125 -1165 19155
rect -1115 19125 -1085 19155
rect -1035 19125 -1005 19155
rect -955 19125 -925 19155
rect -875 19125 -845 19155
rect -795 19125 -765 19155
rect -715 19125 -685 19155
rect -635 19125 -605 19155
rect -555 19125 -525 19155
rect -475 19125 -445 19155
rect -395 19125 -365 19155
rect -315 19125 -285 19155
rect -235 19125 -205 19155
rect -155 19125 -125 19155
rect -75 19125 -45 19155
rect 5 19125 35 19155
rect -3035 19045 -3005 19075
rect -3515 18965 -3485 18995
rect -3435 18965 -3405 18995
rect -3355 18965 -3325 18995
rect -3275 18965 -3245 18995
rect -3195 18965 -3165 18995
rect -2875 18965 -2845 18995
rect -2795 18965 -2765 18995
rect -2715 18965 -2685 18995
rect -2635 18965 -2605 18995
rect -2555 18965 -2525 18995
rect -2475 18965 -2445 18995
rect -2395 18965 -2365 18995
rect -2075 18965 -2045 18995
rect -1995 18965 -1965 18995
rect -1915 18965 -1885 18995
rect -1835 18965 -1805 18995
rect -1755 18965 -1725 18995
rect -1675 18965 -1645 18995
rect -1595 18965 -1565 18995
rect -1515 18965 -1485 18995
rect -1435 18965 -1405 18995
rect -1355 18965 -1325 18995
rect -1275 18965 -1245 18995
rect -1195 18965 -1165 18995
rect -1115 18965 -1085 18995
rect -1035 18965 -1005 18995
rect -955 18965 -925 18995
rect -875 18965 -845 18995
rect -795 18965 -765 18995
rect -715 18965 -685 18995
rect -635 18965 -605 18995
rect -555 18965 -525 18995
rect -475 18965 -445 18995
rect -395 18965 -365 18995
rect -315 18965 -285 18995
rect -235 18965 -205 18995
rect -155 18965 -125 18995
rect -75 18965 -45 18995
rect 5 18965 35 18995
rect -2235 18885 -2205 18915
rect -3515 18805 -3485 18835
rect -3435 18805 -3405 18835
rect -3355 18805 -3325 18835
rect -3275 18805 -3245 18835
rect -3195 18805 -3165 18835
rect -2875 18805 -2845 18835
rect -2795 18805 -2765 18835
rect -2715 18805 -2685 18835
rect -2635 18805 -2605 18835
rect -2555 18805 -2525 18835
rect -2475 18805 -2445 18835
rect -2395 18805 -2365 18835
rect -2075 18805 -2045 18835
rect -1995 18805 -1965 18835
rect -1915 18805 -1885 18835
rect -1835 18805 -1805 18835
rect -1755 18805 -1725 18835
rect -1675 18805 -1645 18835
rect -1595 18805 -1565 18835
rect -1515 18805 -1485 18835
rect -1435 18805 -1405 18835
rect -1355 18805 -1325 18835
rect -1275 18805 -1245 18835
rect -1195 18805 -1165 18835
rect -1115 18805 -1085 18835
rect -1035 18805 -1005 18835
rect -955 18805 -925 18835
rect -875 18805 -845 18835
rect -795 18805 -765 18835
rect -715 18805 -685 18835
rect -635 18805 -605 18835
rect -555 18805 -525 18835
rect -475 18805 -445 18835
rect -395 18805 -365 18835
rect -315 18805 -285 18835
rect -235 18805 -205 18835
rect -155 18805 -125 18835
rect -75 18805 -45 18835
rect 5 18805 35 18835
rect 38525 18445 38555 18475
rect 38685 18445 38715 18475
rect 38605 18365 38635 18395
rect 38365 18285 38395 18315
rect 38445 18285 38475 18315
rect 38525 18285 38555 18315
rect 38685 18285 38715 18315
rect 38605 18205 38635 18235
rect 38365 18125 38395 18155
rect 38445 18125 38475 18155
rect 38525 18125 38555 18155
rect 38685 18125 38715 18155
rect 38525 17965 38555 17995
rect 38685 17965 38715 17995
rect 38605 17885 38635 17915
rect 63360 17840 63480 17960
rect 38525 17805 38555 17835
rect 38685 17805 38715 17835
rect 38525 17725 38555 17755
rect 38685 17725 38715 17755
rect 38525 17645 38555 17675
rect 38685 17645 38715 17675
rect -1275 17605 -1245 17635
rect -1195 17605 -1165 17635
rect -1115 17605 -1085 17635
rect -1035 17605 -1005 17635
rect -955 17605 -925 17635
rect -875 17605 -845 17635
rect -795 17605 -765 17635
rect -715 17605 -685 17635
rect -635 17605 -605 17635
rect -555 17605 -525 17635
rect -475 17605 -445 17635
rect -395 17605 -365 17635
rect -315 17605 -285 17635
rect -235 17605 -205 17635
rect -155 17605 -125 17635
rect -75 17605 -45 17635
rect 5 17605 35 17635
rect -1480 17480 -1360 17600
rect 38525 17565 38555 17595
rect 38685 17565 38715 17595
rect 38525 17485 38555 17515
rect 38685 17485 38715 17515
rect -1275 17445 -1245 17475
rect -1195 17445 -1165 17475
rect -1115 17445 -1085 17475
rect -1035 17445 -1005 17475
rect -955 17445 -925 17475
rect -875 17445 -845 17475
rect -795 17445 -765 17475
rect -715 17445 -685 17475
rect -635 17445 -605 17475
rect -555 17445 -525 17475
rect -475 17445 -445 17475
rect -395 17445 -365 17475
rect -315 17445 -285 17475
rect -235 17445 -205 17475
rect -155 17445 -125 17475
rect -75 17445 -45 17475
rect 5 17445 35 17475
rect 38605 17405 38635 17435
rect 38525 17325 38555 17355
rect 38685 17325 38715 17355
<< metal3 >>
rect 38440 22235 38480 22240
rect 38440 22205 38445 22235
rect 38475 22205 38480 22235
rect -720 20920 -520 20960
rect -720 20800 -680 20920
rect -560 20800 -520 20920
rect -720 20760 -520 20800
rect -480 20955 -440 20960
rect -480 20925 -475 20955
rect -445 20925 -440 20955
rect -480 20795 -440 20925
rect -480 20765 -475 20795
rect -445 20765 -440 20795
rect -480 20760 -440 20765
rect -400 20955 -360 20960
rect -400 20925 -395 20955
rect -365 20925 -360 20955
rect -400 20795 -360 20925
rect -400 20765 -395 20795
rect -365 20765 -360 20795
rect -400 20760 -360 20765
rect -320 20955 -280 20960
rect -320 20925 -315 20955
rect -285 20925 -280 20955
rect -320 20795 -280 20925
rect -320 20765 -315 20795
rect -285 20765 -280 20795
rect -320 20760 -280 20765
rect -240 20955 -200 20960
rect -240 20925 -235 20955
rect -205 20925 -200 20955
rect -240 20795 -200 20925
rect -240 20765 -235 20795
rect -205 20765 -200 20795
rect -240 20760 -200 20765
rect -160 20955 -120 20960
rect -160 20925 -155 20955
rect -125 20925 -120 20955
rect -160 20795 -120 20925
rect -160 20765 -155 20795
rect -125 20765 -120 20795
rect -160 20760 -120 20765
rect -80 20955 -40 20960
rect -80 20925 -75 20955
rect -45 20925 -40 20955
rect -80 20795 -40 20925
rect -80 20765 -75 20795
rect -45 20765 -40 20795
rect -80 20760 -40 20765
rect 0 20955 40 20960
rect 0 20925 5 20955
rect 35 20925 40 20955
rect 0 20795 40 20925
rect 38440 20875 38480 22205
rect 38520 21836 38560 21840
rect 38520 21804 38524 21836
rect 38556 21804 38560 21836
rect 38520 21676 38560 21804
rect 38680 21836 38720 21840
rect 38680 21804 38684 21836
rect 38716 21804 38720 21836
rect 38520 21644 38524 21676
rect 38556 21644 38560 21676
rect 38520 21596 38560 21644
rect 38520 21564 38524 21596
rect 38556 21564 38560 21596
rect 38520 21516 38560 21564
rect 38520 21484 38524 21516
rect 38556 21484 38560 21516
rect 38520 21436 38560 21484
rect 38520 21404 38524 21436
rect 38556 21404 38560 21436
rect 38520 21356 38560 21404
rect 38520 21324 38524 21356
rect 38556 21324 38560 21356
rect 38520 21196 38560 21324
rect 38600 21755 38640 21760
rect 38600 21725 38605 21755
rect 38635 21725 38640 21755
rect 38600 21275 38640 21725
rect 38600 21245 38605 21275
rect 38635 21245 38640 21275
rect 38600 21240 38640 21245
rect 38680 21676 38720 21804
rect 38680 21644 38684 21676
rect 38716 21644 38720 21676
rect 38680 21596 38720 21644
rect 38680 21564 38684 21596
rect 38716 21564 38720 21596
rect 38680 21516 38720 21564
rect 38680 21484 38684 21516
rect 38716 21484 38720 21516
rect 38680 21436 38720 21484
rect 38680 21404 38684 21436
rect 38716 21404 38720 21436
rect 38680 21356 38720 21404
rect 38680 21324 38684 21356
rect 38716 21324 38720 21356
rect 38520 21164 38524 21196
rect 38556 21164 38560 21196
rect 38520 21160 38560 21164
rect 38680 21196 38720 21324
rect 38680 21164 38684 21196
rect 38716 21164 38720 21196
rect 38680 21160 38720 21164
rect 63320 21320 63520 21360
rect 63320 21200 63360 21320
rect 63480 21200 63520 21320
rect 38440 20845 38445 20875
rect 38475 20845 38480 20875
rect 38440 20840 38480 20845
rect 38520 20876 38560 20880
rect 38520 20844 38524 20876
rect 38556 20844 38560 20876
rect 0 20765 5 20795
rect 35 20765 40 20795
rect 0 20760 40 20765
rect 38520 20716 38560 20844
rect 38520 20684 38524 20716
rect 38556 20684 38560 20716
rect 38520 20636 38560 20684
rect 38520 20604 38524 20636
rect 38556 20604 38560 20636
rect 38520 20556 38560 20604
rect 38520 20524 38524 20556
rect 38556 20524 38560 20556
rect 38520 20476 38560 20524
rect 38520 20444 38524 20476
rect 38556 20444 38560 20476
rect 38520 20396 38560 20444
rect 38520 20364 38524 20396
rect 38556 20364 38560 20396
rect 38360 20315 38400 20320
rect 38360 20285 38365 20315
rect 38395 20285 38400 20315
rect 38360 20155 38400 20285
rect 38360 20125 38365 20155
rect 38395 20125 38400 20155
rect 38360 20120 38400 20125
rect 38440 20315 38480 20320
rect 38440 20285 38445 20315
rect 38475 20285 38480 20315
rect 38440 20155 38480 20285
rect 38440 20125 38445 20155
rect 38475 20125 38480 20155
rect 38440 20120 38480 20125
rect 38520 20316 38560 20364
rect 38520 20284 38524 20316
rect 38556 20284 38560 20316
rect 38520 20156 38560 20284
rect 38520 20124 38524 20156
rect 38556 20124 38560 20156
rect 38520 20120 38560 20124
rect 38600 20795 38640 20880
rect 38600 20765 38605 20795
rect 38635 20765 38640 20795
rect 38600 20235 38640 20765
rect 38600 20205 38605 20235
rect 38635 20205 38640 20235
rect 38600 20120 38640 20205
rect 38680 20876 38720 20880
rect 38680 20844 38684 20876
rect 38716 20844 38720 20876
rect 38680 20716 38720 20844
rect 38680 20684 38684 20716
rect 38716 20684 38720 20716
rect 38680 20636 38720 20684
rect 38680 20604 38684 20636
rect 38716 20604 38720 20636
rect 38680 20556 38720 20604
rect 38680 20524 38684 20556
rect 38716 20524 38720 20556
rect 38680 20476 38720 20524
rect 38680 20444 38684 20476
rect 38716 20444 38720 20476
rect 38680 20396 38720 20444
rect 38680 20364 38684 20396
rect 38716 20364 38720 20396
rect 38680 20316 38720 20364
rect 38680 20284 38684 20316
rect 38716 20284 38720 20316
rect 38680 20156 38720 20284
rect 38680 20124 38684 20156
rect 38716 20124 38720 20156
rect 38680 20120 38720 20124
rect 63320 20040 63520 21200
rect 63320 19920 63360 20040
rect 63480 19920 63520 20040
rect 63320 19880 63520 19920
rect 63320 19240 63520 19280
rect -3520 19155 -3480 19160
rect -3520 19125 -3515 19155
rect -3485 19125 -3480 19155
rect -3520 18995 -3480 19125
rect -3520 18965 -3515 18995
rect -3485 18965 -3480 18995
rect -3520 18835 -3480 18965
rect -3520 18805 -3515 18835
rect -3485 18805 -3480 18835
rect -3520 18800 -3480 18805
rect -3440 19155 -3400 19160
rect -3440 19125 -3435 19155
rect -3405 19125 -3400 19155
rect -3440 18995 -3400 19125
rect -3440 18965 -3435 18995
rect -3405 18965 -3400 18995
rect -3440 18835 -3400 18965
rect -3440 18805 -3435 18835
rect -3405 18805 -3400 18835
rect -3440 18800 -3400 18805
rect -3360 19155 -3320 19160
rect -3360 19125 -3355 19155
rect -3325 19125 -3320 19155
rect -3360 18995 -3320 19125
rect -3360 18965 -3355 18995
rect -3325 18965 -3320 18995
rect -3360 18835 -3320 18965
rect -3360 18805 -3355 18835
rect -3325 18805 -3320 18835
rect -3360 18800 -3320 18805
rect -3280 19155 -3240 19160
rect -3280 19125 -3275 19155
rect -3245 19125 -3240 19155
rect -3280 18995 -3240 19125
rect -3280 18965 -3275 18995
rect -3245 18965 -3240 18995
rect -3280 18835 -3240 18965
rect -3280 18805 -3275 18835
rect -3245 18805 -3240 18835
rect -3280 18800 -3240 18805
rect -3200 19155 -3160 19160
rect -3200 19125 -3195 19155
rect -3165 19125 -3160 19155
rect -3200 18995 -3160 19125
rect -3200 18965 -3195 18995
rect -3165 18965 -3160 18995
rect -3200 18835 -3160 18965
rect -3120 19120 -2920 19160
rect -3120 19000 -3080 19120
rect -2960 19000 -2920 19120
rect -3120 18960 -2920 19000
rect -2880 19155 -2840 19160
rect -2880 19125 -2875 19155
rect -2845 19125 -2840 19155
rect -2880 18995 -2840 19125
rect -2880 18965 -2875 18995
rect -2845 18965 -2840 18995
rect -3200 18805 -3195 18835
rect -3165 18805 -3160 18835
rect -3200 18800 -3160 18805
rect -2880 18835 -2840 18965
rect -2880 18805 -2875 18835
rect -2845 18805 -2840 18835
rect -2880 18800 -2840 18805
rect -2800 19155 -2760 19160
rect -2800 19125 -2795 19155
rect -2765 19125 -2760 19155
rect -2800 18995 -2760 19125
rect -2800 18965 -2795 18995
rect -2765 18965 -2760 18995
rect -2800 18835 -2760 18965
rect -2800 18805 -2795 18835
rect -2765 18805 -2760 18835
rect -2800 18800 -2760 18805
rect -2720 19155 -2680 19160
rect -2720 19125 -2715 19155
rect -2685 19125 -2680 19155
rect -2720 18995 -2680 19125
rect -2720 18965 -2715 18995
rect -2685 18965 -2680 18995
rect -2720 18835 -2680 18965
rect -2720 18805 -2715 18835
rect -2685 18805 -2680 18835
rect -2720 18800 -2680 18805
rect -2640 19155 -2600 19160
rect -2640 19125 -2635 19155
rect -2605 19125 -2600 19155
rect -2640 18995 -2600 19125
rect -2640 18965 -2635 18995
rect -2605 18965 -2600 18995
rect -2640 18835 -2600 18965
rect -2640 18805 -2635 18835
rect -2605 18805 -2600 18835
rect -2640 18800 -2600 18805
rect -2560 19155 -2520 19160
rect -2560 19125 -2555 19155
rect -2525 19125 -2520 19155
rect -2560 18995 -2520 19125
rect -2560 18965 -2555 18995
rect -2525 18965 -2520 18995
rect -2560 18835 -2520 18965
rect -2560 18805 -2555 18835
rect -2525 18805 -2520 18835
rect -2560 18800 -2520 18805
rect -2480 19155 -2440 19160
rect -2480 19125 -2475 19155
rect -2445 19125 -2440 19155
rect -2480 18995 -2440 19125
rect -2480 18965 -2475 18995
rect -2445 18965 -2440 18995
rect -2480 18835 -2440 18965
rect -2480 18805 -2475 18835
rect -2445 18805 -2440 18835
rect -2480 18800 -2440 18805
rect -2400 19155 -2360 19160
rect -2400 19125 -2395 19155
rect -2365 19125 -2360 19155
rect -2400 18995 -2360 19125
rect -2080 19155 -2040 19160
rect -2080 19125 -2075 19155
rect -2045 19125 -2040 19155
rect -2400 18965 -2395 18995
rect -2365 18965 -2360 18995
rect -2400 18835 -2360 18965
rect -2400 18805 -2395 18835
rect -2365 18805 -2360 18835
rect -2400 18800 -2360 18805
rect -2320 18960 -2120 19000
rect -2320 18840 -2280 18960
rect -2160 18840 -2120 18960
rect -2320 18800 -2120 18840
rect -2080 18995 -2040 19125
rect -2080 18965 -2075 18995
rect -2045 18965 -2040 18995
rect -2080 18835 -2040 18965
rect -2080 18805 -2075 18835
rect -2045 18805 -2040 18835
rect -2080 18800 -2040 18805
rect -2000 19155 -1960 19160
rect -2000 19125 -1995 19155
rect -1965 19125 -1960 19155
rect -2000 18995 -1960 19125
rect -2000 18965 -1995 18995
rect -1965 18965 -1960 18995
rect -2000 18835 -1960 18965
rect -2000 18805 -1995 18835
rect -1965 18805 -1960 18835
rect -2000 18800 -1960 18805
rect -1920 19155 -1880 19160
rect -1920 19125 -1915 19155
rect -1885 19125 -1880 19155
rect -1920 18995 -1880 19125
rect -1920 18965 -1915 18995
rect -1885 18965 -1880 18995
rect -1920 18835 -1880 18965
rect -1920 18805 -1915 18835
rect -1885 18805 -1880 18835
rect -1920 18800 -1880 18805
rect -1840 19155 -1800 19160
rect -1840 19125 -1835 19155
rect -1805 19125 -1800 19155
rect -1840 18995 -1800 19125
rect -1840 18965 -1835 18995
rect -1805 18965 -1800 18995
rect -1840 18835 -1800 18965
rect -1840 18805 -1835 18835
rect -1805 18805 -1800 18835
rect -1840 18800 -1800 18805
rect -1760 19155 -1720 19160
rect -1760 19125 -1755 19155
rect -1725 19125 -1720 19155
rect -1760 18995 -1720 19125
rect -1760 18965 -1755 18995
rect -1725 18965 -1720 18995
rect -1760 18835 -1720 18965
rect -1760 18805 -1755 18835
rect -1725 18805 -1720 18835
rect -1760 18800 -1720 18805
rect -1680 19155 -1640 19160
rect -1680 19125 -1675 19155
rect -1645 19125 -1640 19155
rect -1680 18995 -1640 19125
rect -1680 18965 -1675 18995
rect -1645 18965 -1640 18995
rect -1680 18835 -1640 18965
rect -1680 18805 -1675 18835
rect -1645 18805 -1640 18835
rect -1680 18800 -1640 18805
rect -1600 19155 -1560 19160
rect -1600 19125 -1595 19155
rect -1565 19125 -1560 19155
rect -1600 18995 -1560 19125
rect -1600 18965 -1595 18995
rect -1565 18965 -1560 18995
rect -1600 18835 -1560 18965
rect -1600 18805 -1595 18835
rect -1565 18805 -1560 18835
rect -1600 18800 -1560 18805
rect -1520 19155 -1480 19160
rect -1520 19125 -1515 19155
rect -1485 19125 -1480 19155
rect -1520 18995 -1480 19125
rect -1520 18965 -1515 18995
rect -1485 18965 -1480 18995
rect -1520 18835 -1480 18965
rect -1520 18805 -1515 18835
rect -1485 18805 -1480 18835
rect -1520 18800 -1480 18805
rect -1440 19155 -1400 19160
rect -1440 19125 -1435 19155
rect -1405 19125 -1400 19155
rect -1440 18995 -1400 19125
rect -1440 18965 -1435 18995
rect -1405 18965 -1400 18995
rect -1440 18835 -1400 18965
rect -1440 18805 -1435 18835
rect -1405 18805 -1400 18835
rect -1440 18800 -1400 18805
rect -1360 19155 -1320 19160
rect -1360 19125 -1355 19155
rect -1325 19125 -1320 19155
rect -1360 18995 -1320 19125
rect -1360 18965 -1355 18995
rect -1325 18965 -1320 18995
rect -1360 18835 -1320 18965
rect -1360 18805 -1355 18835
rect -1325 18805 -1320 18835
rect -1360 18800 -1320 18805
rect -1280 19155 -1240 19160
rect -1280 19125 -1275 19155
rect -1245 19125 -1240 19155
rect -1280 18995 -1240 19125
rect -1280 18965 -1275 18995
rect -1245 18965 -1240 18995
rect -1280 18835 -1240 18965
rect -1280 18805 -1275 18835
rect -1245 18805 -1240 18835
rect -1280 18800 -1240 18805
rect -1200 19155 -1160 19160
rect -1200 19125 -1195 19155
rect -1165 19125 -1160 19155
rect -1200 18995 -1160 19125
rect -1200 18965 -1195 18995
rect -1165 18965 -1160 18995
rect -1200 18835 -1160 18965
rect -1200 18805 -1195 18835
rect -1165 18805 -1160 18835
rect -1200 18800 -1160 18805
rect -1120 19155 -1080 19160
rect -1120 19125 -1115 19155
rect -1085 19125 -1080 19155
rect -1120 18995 -1080 19125
rect -1120 18965 -1115 18995
rect -1085 18965 -1080 18995
rect -1120 18835 -1080 18965
rect -1120 18805 -1115 18835
rect -1085 18805 -1080 18835
rect -1120 18800 -1080 18805
rect -1040 19155 -1000 19160
rect -1040 19125 -1035 19155
rect -1005 19125 -1000 19155
rect -1040 18995 -1000 19125
rect -1040 18965 -1035 18995
rect -1005 18965 -1000 18995
rect -1040 18835 -1000 18965
rect -1040 18805 -1035 18835
rect -1005 18805 -1000 18835
rect -1040 18800 -1000 18805
rect -960 19155 -920 19160
rect -960 19125 -955 19155
rect -925 19125 -920 19155
rect -960 18995 -920 19125
rect -960 18965 -955 18995
rect -925 18965 -920 18995
rect -960 18835 -920 18965
rect -960 18805 -955 18835
rect -925 18805 -920 18835
rect -960 18800 -920 18805
rect -880 19155 -840 19160
rect -880 19125 -875 19155
rect -845 19125 -840 19155
rect -880 18995 -840 19125
rect -880 18965 -875 18995
rect -845 18965 -840 18995
rect -880 18835 -840 18965
rect -880 18805 -875 18835
rect -845 18805 -840 18835
rect -880 18800 -840 18805
rect -800 19155 -760 19160
rect -800 19125 -795 19155
rect -765 19125 -760 19155
rect -800 18995 -760 19125
rect -800 18965 -795 18995
rect -765 18965 -760 18995
rect -800 18835 -760 18965
rect -800 18805 -795 18835
rect -765 18805 -760 18835
rect -800 18800 -760 18805
rect -720 19155 -680 19160
rect -720 19125 -715 19155
rect -685 19125 -680 19155
rect -720 18995 -680 19125
rect -720 18965 -715 18995
rect -685 18965 -680 18995
rect -720 18835 -680 18965
rect -720 18805 -715 18835
rect -685 18805 -680 18835
rect -720 18800 -680 18805
rect -640 19155 -600 19160
rect -640 19125 -635 19155
rect -605 19125 -600 19155
rect -640 18995 -600 19125
rect -640 18965 -635 18995
rect -605 18965 -600 18995
rect -640 18835 -600 18965
rect -640 18805 -635 18835
rect -605 18805 -600 18835
rect -640 18800 -600 18805
rect -560 19155 -520 19160
rect -560 19125 -555 19155
rect -525 19125 -520 19155
rect -560 18995 -520 19125
rect -560 18965 -555 18995
rect -525 18965 -520 18995
rect -560 18835 -520 18965
rect -560 18805 -555 18835
rect -525 18805 -520 18835
rect -560 18800 -520 18805
rect -480 19155 -440 19160
rect -480 19125 -475 19155
rect -445 19125 -440 19155
rect -480 18995 -440 19125
rect -480 18965 -475 18995
rect -445 18965 -440 18995
rect -480 18835 -440 18965
rect -480 18805 -475 18835
rect -445 18805 -440 18835
rect -480 18800 -440 18805
rect -400 19155 -360 19160
rect -400 19125 -395 19155
rect -365 19125 -360 19155
rect -400 18995 -360 19125
rect -400 18965 -395 18995
rect -365 18965 -360 18995
rect -400 18835 -360 18965
rect -400 18805 -395 18835
rect -365 18805 -360 18835
rect -400 18800 -360 18805
rect -320 19155 -280 19160
rect -320 19125 -315 19155
rect -285 19125 -280 19155
rect -320 18995 -280 19125
rect -320 18965 -315 18995
rect -285 18965 -280 18995
rect -320 18835 -280 18965
rect -320 18805 -315 18835
rect -285 18805 -280 18835
rect -320 18800 -280 18805
rect -240 19155 -200 19160
rect -240 19125 -235 19155
rect -205 19125 -200 19155
rect -240 18995 -200 19125
rect -240 18965 -235 18995
rect -205 18965 -200 18995
rect -240 18835 -200 18965
rect -240 18805 -235 18835
rect -205 18805 -200 18835
rect -240 18800 -200 18805
rect -160 19155 -120 19160
rect -160 19125 -155 19155
rect -125 19125 -120 19155
rect -160 18995 -120 19125
rect -160 18965 -155 18995
rect -125 18965 -120 18995
rect -160 18835 -120 18965
rect -160 18805 -155 18835
rect -125 18805 -120 18835
rect -160 18800 -120 18805
rect -80 19155 -40 19160
rect -80 19125 -75 19155
rect -45 19125 -40 19155
rect -80 18995 -40 19125
rect -80 18965 -75 18995
rect -45 18965 -40 18995
rect -80 18835 -40 18965
rect -80 18805 -75 18835
rect -45 18805 -40 18835
rect -80 18800 -40 18805
rect 0 19155 40 19160
rect 0 19125 5 19155
rect 35 19125 40 19155
rect 0 18995 40 19125
rect 0 18965 5 18995
rect 35 18965 40 18995
rect 0 18835 40 18965
rect 0 18805 5 18835
rect 35 18805 40 18835
rect 0 18800 40 18805
rect 63320 19120 63360 19240
rect 63480 19120 63520 19240
rect 38520 18476 38560 18480
rect 38520 18444 38524 18476
rect 38556 18444 38560 18476
rect 38360 18315 38400 18320
rect 38360 18285 38365 18315
rect 38395 18285 38400 18315
rect 38360 18155 38400 18285
rect 38360 18125 38365 18155
rect 38395 18125 38400 18155
rect 38360 18120 38400 18125
rect 38440 18315 38480 18320
rect 38440 18285 38445 18315
rect 38475 18285 38480 18315
rect 38440 18155 38480 18285
rect 38440 18125 38445 18155
rect 38475 18125 38480 18155
rect 38440 18120 38480 18125
rect 38520 18316 38560 18444
rect 38520 18284 38524 18316
rect 38556 18284 38560 18316
rect 38520 18156 38560 18284
rect 38520 18124 38524 18156
rect 38556 18124 38560 18156
rect 38520 18120 38560 18124
rect 38600 18395 38640 18480
rect 38600 18365 38605 18395
rect 38635 18365 38640 18395
rect 38600 18235 38640 18365
rect 38600 18205 38605 18235
rect 38635 18205 38640 18235
rect 38600 18120 38640 18205
rect 38680 18476 38720 18480
rect 38680 18444 38684 18476
rect 38716 18444 38720 18476
rect 38680 18316 38720 18444
rect 38680 18284 38684 18316
rect 38716 18284 38720 18316
rect 38680 18156 38720 18284
rect 38680 18124 38684 18156
rect 38716 18124 38720 18156
rect 38680 18120 38720 18124
rect 38520 17996 38560 18000
rect 38520 17964 38524 17996
rect 38556 17964 38560 17996
rect 38520 17836 38560 17964
rect 38680 17996 38720 18000
rect 38680 17964 38684 17996
rect 38716 17964 38720 17996
rect 38520 17804 38524 17836
rect 38556 17804 38560 17836
rect 38520 17756 38560 17804
rect 38520 17724 38524 17756
rect 38556 17724 38560 17756
rect 38520 17676 38560 17724
rect 38520 17644 38524 17676
rect 38556 17644 38560 17676
rect -1520 17600 -1320 17640
rect -1520 17480 -1480 17600
rect -1360 17480 -1320 17600
rect -1520 17440 -1320 17480
rect -1280 17635 -1240 17640
rect -1280 17605 -1275 17635
rect -1245 17605 -1240 17635
rect -1280 17475 -1240 17605
rect -1280 17445 -1275 17475
rect -1245 17445 -1240 17475
rect -1280 17440 -1240 17445
rect -1200 17635 -1160 17640
rect -1200 17605 -1195 17635
rect -1165 17605 -1160 17635
rect -1200 17475 -1160 17605
rect -1200 17445 -1195 17475
rect -1165 17445 -1160 17475
rect -1200 17440 -1160 17445
rect -1120 17635 -1080 17640
rect -1120 17605 -1115 17635
rect -1085 17605 -1080 17635
rect -1120 17475 -1080 17605
rect -1120 17445 -1115 17475
rect -1085 17445 -1080 17475
rect -1120 17440 -1080 17445
rect -1040 17635 -1000 17640
rect -1040 17605 -1035 17635
rect -1005 17605 -1000 17635
rect -1040 17475 -1000 17605
rect -1040 17445 -1035 17475
rect -1005 17445 -1000 17475
rect -1040 17440 -1000 17445
rect -960 17635 -920 17640
rect -960 17605 -955 17635
rect -925 17605 -920 17635
rect -960 17475 -920 17605
rect -960 17445 -955 17475
rect -925 17445 -920 17475
rect -960 17440 -920 17445
rect -880 17635 -840 17640
rect -880 17605 -875 17635
rect -845 17605 -840 17635
rect -880 17475 -840 17605
rect -880 17445 -875 17475
rect -845 17445 -840 17475
rect -880 17440 -840 17445
rect -800 17635 -760 17640
rect -800 17605 -795 17635
rect -765 17605 -760 17635
rect -800 17475 -760 17605
rect -800 17445 -795 17475
rect -765 17445 -760 17475
rect -800 17440 -760 17445
rect -720 17635 -680 17640
rect -720 17605 -715 17635
rect -685 17605 -680 17635
rect -720 17475 -680 17605
rect -720 17445 -715 17475
rect -685 17445 -680 17475
rect -720 17440 -680 17445
rect -640 17635 -600 17640
rect -640 17605 -635 17635
rect -605 17605 -600 17635
rect -640 17475 -600 17605
rect -640 17445 -635 17475
rect -605 17445 -600 17475
rect -640 17440 -600 17445
rect -560 17635 -520 17640
rect -560 17605 -555 17635
rect -525 17605 -520 17635
rect -560 17475 -520 17605
rect -560 17445 -555 17475
rect -525 17445 -520 17475
rect -560 17440 -520 17445
rect -480 17635 -440 17640
rect -480 17605 -475 17635
rect -445 17605 -440 17635
rect -480 17475 -440 17605
rect -480 17445 -475 17475
rect -445 17445 -440 17475
rect -480 17440 -440 17445
rect -400 17635 -360 17640
rect -400 17605 -395 17635
rect -365 17605 -360 17635
rect -400 17475 -360 17605
rect -400 17445 -395 17475
rect -365 17445 -360 17475
rect -400 17440 -360 17445
rect -320 17635 -280 17640
rect -320 17605 -315 17635
rect -285 17605 -280 17635
rect -320 17475 -280 17605
rect -320 17445 -315 17475
rect -285 17445 -280 17475
rect -320 17440 -280 17445
rect -240 17635 -200 17640
rect -240 17605 -235 17635
rect -205 17605 -200 17635
rect -240 17475 -200 17605
rect -240 17445 -235 17475
rect -205 17445 -200 17475
rect -240 17440 -200 17445
rect -160 17635 -120 17640
rect -160 17605 -155 17635
rect -125 17605 -120 17635
rect -160 17475 -120 17605
rect -160 17445 -155 17475
rect -125 17445 -120 17475
rect -160 17440 -120 17445
rect -80 17635 -40 17640
rect -80 17605 -75 17635
rect -45 17605 -40 17635
rect -80 17475 -40 17605
rect -80 17445 -75 17475
rect -45 17445 -40 17475
rect -80 17440 -40 17445
rect 0 17635 40 17640
rect 0 17605 5 17635
rect 35 17605 40 17635
rect 0 17475 40 17605
rect 0 17445 5 17475
rect 35 17445 40 17475
rect 0 17440 40 17445
rect 38520 17596 38560 17644
rect 38520 17564 38524 17596
rect 38556 17564 38560 17596
rect 38520 17516 38560 17564
rect 38520 17484 38524 17516
rect 38556 17484 38560 17516
rect 38520 17356 38560 17484
rect 38520 17324 38524 17356
rect 38556 17324 38560 17356
rect 38520 17320 38560 17324
rect 38600 17915 38640 17920
rect 38600 17885 38605 17915
rect 38635 17885 38640 17915
rect 38600 17435 38640 17885
rect 38600 17405 38605 17435
rect 38635 17405 38640 17435
rect 38600 17320 38640 17405
rect 38680 17836 38720 17964
rect 38680 17804 38684 17836
rect 38716 17804 38720 17836
rect 38680 17756 38720 17804
rect 63320 17960 63520 19120
rect 63320 17840 63360 17960
rect 63480 17840 63520 17960
rect 63320 17800 63520 17840
rect 38680 17724 38684 17756
rect 38716 17724 38720 17756
rect 38680 17676 38720 17724
rect 38680 17644 38684 17676
rect 38716 17644 38720 17676
rect 38680 17596 38720 17644
rect 38680 17564 38684 17596
rect 38716 17564 38720 17596
rect 38680 17516 38720 17564
rect 38680 17484 38684 17516
rect 38716 17484 38720 17516
rect 38680 17356 38720 17484
rect 38680 17324 38684 17356
rect 38716 17324 38720 17356
rect 38680 17320 38720 17324
<< via3 >>
rect -680 20800 -560 20920
rect 38524 21835 38556 21836
rect 38524 21805 38525 21835
rect 38525 21805 38555 21835
rect 38555 21805 38556 21835
rect 38524 21804 38556 21805
rect 38684 21835 38716 21836
rect 38684 21805 38685 21835
rect 38685 21805 38715 21835
rect 38715 21805 38716 21835
rect 38684 21804 38716 21805
rect 38524 21675 38556 21676
rect 38524 21645 38525 21675
rect 38525 21645 38555 21675
rect 38555 21645 38556 21675
rect 38524 21644 38556 21645
rect 38524 21595 38556 21596
rect 38524 21565 38525 21595
rect 38525 21565 38555 21595
rect 38555 21565 38556 21595
rect 38524 21564 38556 21565
rect 38524 21515 38556 21516
rect 38524 21485 38525 21515
rect 38525 21485 38555 21515
rect 38555 21485 38556 21515
rect 38524 21484 38556 21485
rect 38524 21435 38556 21436
rect 38524 21405 38525 21435
rect 38525 21405 38555 21435
rect 38555 21405 38556 21435
rect 38524 21404 38556 21405
rect 38524 21355 38556 21356
rect 38524 21325 38525 21355
rect 38525 21325 38555 21355
rect 38555 21325 38556 21355
rect 38524 21324 38556 21325
rect 38684 21675 38716 21676
rect 38684 21645 38685 21675
rect 38685 21645 38715 21675
rect 38715 21645 38716 21675
rect 38684 21644 38716 21645
rect 38684 21595 38716 21596
rect 38684 21565 38685 21595
rect 38685 21565 38715 21595
rect 38715 21565 38716 21595
rect 38684 21564 38716 21565
rect 38684 21515 38716 21516
rect 38684 21485 38685 21515
rect 38685 21485 38715 21515
rect 38715 21485 38716 21515
rect 38684 21484 38716 21485
rect 38684 21435 38716 21436
rect 38684 21405 38685 21435
rect 38685 21405 38715 21435
rect 38715 21405 38716 21435
rect 38684 21404 38716 21405
rect 38684 21355 38716 21356
rect 38684 21325 38685 21355
rect 38685 21325 38715 21355
rect 38715 21325 38716 21355
rect 38684 21324 38716 21325
rect 38524 21195 38556 21196
rect 38524 21165 38525 21195
rect 38525 21165 38555 21195
rect 38555 21165 38556 21195
rect 38524 21164 38556 21165
rect 38684 21195 38716 21196
rect 38684 21165 38685 21195
rect 38685 21165 38715 21195
rect 38715 21165 38716 21195
rect 38684 21164 38716 21165
rect 38524 20875 38556 20876
rect 38524 20845 38525 20875
rect 38525 20845 38555 20875
rect 38555 20845 38556 20875
rect 38524 20844 38556 20845
rect 38524 20715 38556 20716
rect 38524 20685 38525 20715
rect 38525 20685 38555 20715
rect 38555 20685 38556 20715
rect 38524 20684 38556 20685
rect 38524 20635 38556 20636
rect 38524 20605 38525 20635
rect 38525 20605 38555 20635
rect 38555 20605 38556 20635
rect 38524 20604 38556 20605
rect 38524 20555 38556 20556
rect 38524 20525 38525 20555
rect 38525 20525 38555 20555
rect 38555 20525 38556 20555
rect 38524 20524 38556 20525
rect 38524 20475 38556 20476
rect 38524 20445 38525 20475
rect 38525 20445 38555 20475
rect 38555 20445 38556 20475
rect 38524 20444 38556 20445
rect 38524 20395 38556 20396
rect 38524 20365 38525 20395
rect 38525 20365 38555 20395
rect 38555 20365 38556 20395
rect 38524 20364 38556 20365
rect 38524 20315 38556 20316
rect 38524 20285 38525 20315
rect 38525 20285 38555 20315
rect 38555 20285 38556 20315
rect 38524 20284 38556 20285
rect 38524 20155 38556 20156
rect 38524 20125 38525 20155
rect 38525 20125 38555 20155
rect 38555 20125 38556 20155
rect 38524 20124 38556 20125
rect 38684 20875 38716 20876
rect 38684 20845 38685 20875
rect 38685 20845 38715 20875
rect 38715 20845 38716 20875
rect 38684 20844 38716 20845
rect 38684 20715 38716 20716
rect 38684 20685 38685 20715
rect 38685 20685 38715 20715
rect 38715 20685 38716 20715
rect 38684 20684 38716 20685
rect 38684 20635 38716 20636
rect 38684 20605 38685 20635
rect 38685 20605 38715 20635
rect 38715 20605 38716 20635
rect 38684 20604 38716 20605
rect 38684 20555 38716 20556
rect 38684 20525 38685 20555
rect 38685 20525 38715 20555
rect 38715 20525 38716 20555
rect 38684 20524 38716 20525
rect 38684 20475 38716 20476
rect 38684 20445 38685 20475
rect 38685 20445 38715 20475
rect 38715 20445 38716 20475
rect 38684 20444 38716 20445
rect 38684 20395 38716 20396
rect 38684 20365 38685 20395
rect 38685 20365 38715 20395
rect 38715 20365 38716 20395
rect 38684 20364 38716 20365
rect 38684 20315 38716 20316
rect 38684 20285 38685 20315
rect 38685 20285 38715 20315
rect 38715 20285 38716 20315
rect 38684 20284 38716 20285
rect 38684 20155 38716 20156
rect 38684 20125 38685 20155
rect 38685 20125 38715 20155
rect 38715 20125 38716 20155
rect 38684 20124 38716 20125
rect 63360 19920 63480 20040
rect -3080 19075 -2960 19120
rect -3080 19045 -3035 19075
rect -3035 19045 -3005 19075
rect -3005 19045 -2960 19075
rect -3080 19000 -2960 19045
rect -2280 18915 -2160 18960
rect -2280 18885 -2235 18915
rect -2235 18885 -2205 18915
rect -2205 18885 -2160 18915
rect -2280 18840 -2160 18885
rect 63360 19120 63480 19240
rect 38524 18475 38556 18476
rect 38524 18445 38525 18475
rect 38525 18445 38555 18475
rect 38555 18445 38556 18475
rect 38524 18444 38556 18445
rect 38524 18315 38556 18316
rect 38524 18285 38525 18315
rect 38525 18285 38555 18315
rect 38555 18285 38556 18315
rect 38524 18284 38556 18285
rect 38524 18155 38556 18156
rect 38524 18125 38525 18155
rect 38525 18125 38555 18155
rect 38555 18125 38556 18155
rect 38524 18124 38556 18125
rect 38684 18475 38716 18476
rect 38684 18445 38685 18475
rect 38685 18445 38715 18475
rect 38715 18445 38716 18475
rect 38684 18444 38716 18445
rect 38684 18315 38716 18316
rect 38684 18285 38685 18315
rect 38685 18285 38715 18315
rect 38715 18285 38716 18315
rect 38684 18284 38716 18285
rect 38684 18155 38716 18156
rect 38684 18125 38685 18155
rect 38685 18125 38715 18155
rect 38715 18125 38716 18155
rect 38684 18124 38716 18125
rect 38524 17995 38556 17996
rect 38524 17965 38525 17995
rect 38525 17965 38555 17995
rect 38555 17965 38556 17995
rect 38524 17964 38556 17965
rect 38684 17995 38716 17996
rect 38684 17965 38685 17995
rect 38685 17965 38715 17995
rect 38715 17965 38716 17995
rect 38684 17964 38716 17965
rect 38524 17835 38556 17836
rect 38524 17805 38525 17835
rect 38525 17805 38555 17835
rect 38555 17805 38556 17835
rect 38524 17804 38556 17805
rect 38524 17755 38556 17756
rect 38524 17725 38525 17755
rect 38525 17725 38555 17755
rect 38555 17725 38556 17755
rect 38524 17724 38556 17725
rect 38524 17675 38556 17676
rect 38524 17645 38525 17675
rect 38525 17645 38555 17675
rect 38555 17645 38556 17675
rect 38524 17644 38556 17645
rect -1480 17480 -1360 17600
rect 38524 17595 38556 17596
rect 38524 17565 38525 17595
rect 38525 17565 38555 17595
rect 38555 17565 38556 17595
rect 38524 17564 38556 17565
rect 38524 17515 38556 17516
rect 38524 17485 38525 17515
rect 38525 17485 38555 17515
rect 38555 17485 38556 17515
rect 38524 17484 38556 17485
rect 38524 17355 38556 17356
rect 38524 17325 38525 17355
rect 38525 17325 38555 17355
rect 38555 17325 38556 17355
rect 38524 17324 38556 17325
rect 38684 17835 38716 17836
rect 38684 17805 38685 17835
rect 38685 17805 38715 17835
rect 38715 17805 38716 17835
rect 38684 17804 38716 17805
rect 38684 17755 38716 17756
rect 38684 17725 38685 17755
rect 38685 17725 38715 17755
rect 38715 17725 38716 17755
rect 38684 17724 38716 17725
rect 38684 17675 38716 17676
rect 38684 17645 38685 17675
rect 38685 17645 38715 17675
rect 38715 17645 38716 17675
rect 38684 17644 38716 17645
rect 38684 17595 38716 17596
rect 38684 17565 38685 17595
rect 38685 17565 38715 17595
rect 38715 17565 38716 17595
rect 38684 17564 38716 17565
rect 38684 17515 38716 17516
rect 38684 17485 38685 17515
rect 38685 17485 38715 17515
rect 38715 17485 38716 17515
rect 38684 17484 38716 17485
rect 38684 17355 38716 17356
rect 38684 17325 38685 17355
rect 38685 17325 38715 17355
rect 38715 17325 38716 17355
rect 38684 17324 38716 17325
<< metal4 >>
rect 38240 39760 40160 39800
rect 38240 39640 38800 39760
rect 38920 39640 40160 39760
rect 38240 39600 40160 39640
rect 38240 39520 40160 39560
rect 38240 39400 39600 39520
rect 39720 39400 40160 39520
rect 38240 39360 40160 39400
rect 38240 39280 40160 39320
rect 38240 39160 40000 39280
rect 40120 39160 40160 39280
rect 38240 39120 40160 39160
rect 38520 21836 38720 21840
rect 38520 21804 38524 21836
rect 38556 21804 38684 21836
rect 38716 21804 38720 21836
rect 38520 21800 38720 21804
rect 38520 21676 38720 21680
rect 38520 21644 38524 21676
rect 38556 21644 38684 21676
rect 38716 21644 38720 21676
rect 38520 21640 38720 21644
rect 38520 21596 38720 21600
rect 38520 21564 38524 21596
rect 38556 21564 38684 21596
rect 38716 21564 38720 21596
rect 38520 21560 38720 21564
rect 38520 21516 38720 21520
rect 38520 21484 38524 21516
rect 38556 21484 38684 21516
rect 38716 21484 38720 21516
rect 38520 21480 38720 21484
rect 38520 21436 38720 21440
rect 38520 21404 38524 21436
rect 38556 21404 38684 21436
rect 38716 21404 38720 21436
rect 38520 21400 38720 21404
rect 38520 21356 38720 21360
rect 38520 21324 38524 21356
rect 38556 21324 38684 21356
rect 38716 21324 38720 21356
rect 38520 21320 38720 21324
rect 38520 21196 38720 21200
rect 38520 21164 38524 21196
rect 38556 21164 38684 21196
rect 38716 21164 38720 21196
rect 38520 21160 38720 21164
rect -720 20920 -520 20960
rect -720 20800 -680 20920
rect -560 20800 -520 20920
rect 38520 20876 38720 20880
rect 38520 20844 38524 20876
rect 38556 20844 38684 20876
rect 38716 20844 38720 20876
rect 38520 20840 38720 20844
rect -720 20760 -520 20800
rect 38520 20716 38720 20720
rect 38520 20684 38524 20716
rect 38556 20684 38684 20716
rect 38716 20684 38720 20716
rect 38520 20680 38720 20684
rect 38520 20636 38720 20640
rect 38520 20604 38524 20636
rect 38556 20604 38684 20636
rect 38716 20604 38720 20636
rect 38520 20600 38720 20604
rect 38520 20556 38720 20560
rect 38520 20524 38524 20556
rect 38556 20524 38684 20556
rect 38716 20524 38720 20556
rect 38520 20520 38720 20524
rect 38520 20476 38720 20480
rect 38520 20444 38524 20476
rect 38556 20444 38684 20476
rect 38716 20444 38720 20476
rect 38520 20440 38720 20444
rect 62200 20440 63720 20480
rect 38520 20396 38720 20400
rect 38520 20364 38524 20396
rect 38556 20364 38684 20396
rect 38716 20364 38720 20396
rect 38520 20360 38720 20364
rect 62200 20320 62240 20440
rect 62360 20320 63720 20440
rect 38520 20316 38720 20320
rect 38520 20284 38524 20316
rect 38556 20284 38684 20316
rect 38716 20284 38720 20316
rect 38520 20280 38720 20284
rect 62200 20280 63720 20320
rect 38520 20156 38720 20160
rect 38520 20124 38524 20156
rect 38556 20124 38684 20156
rect 38716 20124 38720 20156
rect 38520 20120 38720 20124
rect 63320 20040 63720 20080
rect 63320 19920 63360 20040
rect 63480 19920 63720 20040
rect 63320 19880 63720 19920
rect 62200 19640 63720 19680
rect 62200 19520 62240 19640
rect 62360 19520 63720 19640
rect 62200 19480 63720 19520
rect 63320 19240 63720 19280
rect -3120 19120 -2920 19160
rect -3120 19000 -3080 19120
rect -2960 19000 -2920 19120
rect 63320 19120 63360 19240
rect 63480 19120 63720 19240
rect 63320 19080 63720 19120
rect -3120 18960 -2920 19000
rect -2320 18960 -2120 19000
rect -2320 18840 -2280 18960
rect -2160 18840 -2120 18960
rect -2320 18800 -2120 18840
rect 62200 18840 63720 18880
rect 62200 18720 62240 18840
rect 62360 18720 63720 18840
rect 62200 18680 63720 18720
rect 38520 18476 38720 18480
rect 38520 18444 38524 18476
rect 38556 18444 38684 18476
rect 38716 18444 38720 18476
rect 38520 18440 38720 18444
rect 38520 18316 38720 18320
rect 38520 18284 38524 18316
rect 38556 18284 38684 18316
rect 38716 18284 38720 18316
rect 38520 18280 38720 18284
rect 38520 18156 38720 18160
rect 38520 18124 38524 18156
rect 38556 18124 38684 18156
rect 38716 18124 38720 18156
rect 38520 18120 38720 18124
rect 38520 17996 38720 18000
rect 38520 17964 38524 17996
rect 38556 17964 38684 17996
rect 38716 17964 38720 17996
rect 38520 17960 38720 17964
rect 38520 17836 38720 17840
rect 38520 17804 38524 17836
rect 38556 17804 38684 17836
rect 38716 17804 38720 17836
rect 38520 17800 38720 17804
rect 38520 17756 38720 17760
rect 38520 17724 38524 17756
rect 38556 17724 38684 17756
rect 38716 17724 38720 17756
rect 38520 17720 38720 17724
rect 38520 17676 38720 17680
rect 38520 17644 38524 17676
rect 38556 17644 38684 17676
rect 38716 17644 38720 17676
rect 38520 17640 38720 17644
rect -1520 17600 -1320 17640
rect -1520 17480 -1480 17600
rect -1360 17480 -1320 17600
rect 38520 17596 38720 17600
rect 38520 17564 38524 17596
rect 38556 17564 38684 17596
rect 38716 17564 38720 17596
rect 38520 17560 38720 17564
rect 38520 17516 38720 17520
rect 38520 17484 38524 17516
rect 38556 17484 38684 17516
rect 38716 17484 38720 17516
rect 38520 17480 38720 17484
rect -1520 17440 -1320 17480
rect 38520 17356 38720 17360
rect 38520 17324 38524 17356
rect 38556 17324 38684 17356
rect 38716 17324 38720 17356
rect 38520 17320 38720 17324
<< via4 >>
rect 38800 39640 38920 39760
rect 39600 39400 39720 39520
rect 40000 39160 40120 39280
rect -680 20800 -560 20920
rect 62240 20320 62360 20440
rect 62240 19520 62360 19640
rect -3080 19000 -2960 19120
rect -2280 18840 -2160 18960
rect 62240 18720 62360 18840
rect -1480 17480 -1360 17600
<< metal5 >>
rect -3520 18800 -3320 39880
rect -3120 19120 -2920 39880
rect -3120 19000 -3080 19120
rect -2960 19000 -2920 19120
rect -3120 18800 -2920 19000
rect -2720 18800 -2520 39880
rect -2320 18960 -2120 39880
rect -2320 18840 -2280 18960
rect -2160 18840 -2120 18960
rect -2320 18800 -2120 18840
rect -1920 17440 -1720 39880
rect -1520 17600 -1320 39880
rect -1520 17480 -1480 17600
rect -1360 17480 -1320 17600
rect -1520 17440 -1320 17480
rect -1120 17440 -920 39880
rect -720 20920 -520 39880
rect -720 20800 -680 20920
rect -560 20800 -520 20920
rect -720 20760 -520 20800
rect -320 19480 -120 39880
rect 80 39840 280 39880
rect 480 39840 680 39880
rect 880 39840 1080 39880
rect 38760 39760 38960 39800
rect 38760 39640 38800 39760
rect 38920 39640 38960 39760
rect 38760 39360 38960 39640
rect 39560 39520 39760 39800
rect 39560 39400 39600 39520
rect 39720 39400 39760 39520
rect 39560 39360 39760 39400
rect 39960 39360 40160 39800
rect 62200 20440 62400 20480
rect 62200 20320 62240 20440
rect 62360 20320 62400 20440
rect 62200 20280 62400 20320
rect 62600 20280 62800 20480
rect 63000 20280 63200 20480
rect 62200 18840 62400 18880
rect 62200 18720 62240 18840
rect 62360 18720 62400 18840
rect 62200 18680 62400 18720
rect 62600 18680 62800 18880
rect 63000 18680 63200 18880
use opamp_pair  buffer ../../opamp/mag
timestamp 1638409325
transform 1 0 40360 0 1 22360
box -1640 -23720 22960 17000
use lna  lna ../../lna/mag
timestamp 1638398216
transform 1 0 16640 0 1 280
box -16640 -2120 21680 39560
<< labels >>
rlabel metal2 38320 20200 38360 20240 1 xp
rlabel metal2 38320 18200 38360 18240 1 xm
rlabel metal2 -40 19040 0 19080 0 ip
port 1 nsew
rlabel metal2 -40 18880 0 18920 0 im
port 2 nsew
rlabel metal5 -3120 39840 -2920 39880 0 ip
port 3 nsew
rlabel metal5 -2320 39840 -2120 39880 0 im
port 4 nsew
rlabel metal5 -1520 39840 -1320 39880 0 fsb
port 7 nsew
rlabel metal5 -720 39840 -520 39880 0 ib
port 8 nsew
rlabel metal5 80 39840 280 39880 0 vdda
port 9 nsew
rlabel metal5 480 39840 680 39880 0 gnda
port 10 nsew
rlabel metal5 880 39840 1080 39880 0 vssa
port 11 nsew
rlabel metal4 63680 19880 63720 20080 0 op
port 6 nsew
rlabel metal4 63680 19080 63720 19280 0 om
port 5 nsew
<< end >>
