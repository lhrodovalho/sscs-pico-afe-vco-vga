magic
tech sky130A
timestamp 1634766937
<< nwell >>
rect 6860 40 6920 60
rect 6860 10 6950 40
rect 6860 -2720 6920 10
rect 7790 0 7840 50
rect 22920 0 22970 50
rect 23840 40 23900 60
rect 23770 10 23900 40
rect 6860 -2750 6950 -2720
rect 6860 -2770 6920 -2750
rect 7790 -2760 7840 -2710
rect 22920 -2760 22970 -2710
rect 23840 -2720 23900 10
rect 23770 -2750 23900 -2720
rect 23840 -2770 23900 -2750
rect 6860 -3290 6920 -3270
rect 6860 -3320 6950 -3290
rect 6860 -6050 6920 -3320
rect 7790 -3330 7840 -3280
rect 22920 -3330 22970 -3280
rect 23840 -3290 23900 -3270
rect 23770 -3320 23900 -3290
rect 6860 -6080 6950 -6050
rect 6860 -6100 6920 -6080
rect 7790 -6090 7840 -6040
rect 22920 -6090 22970 -6040
rect 23840 -6050 23900 -3320
rect 23770 -6080 23900 -6050
rect 23840 -6100 23900 -6080
rect 6860 -6550 6920 -6530
rect 6860 -6580 6950 -6550
rect 6860 -9310 6920 -6580
rect 7790 -6590 7840 -6540
rect 22920 -6590 22970 -6540
rect 6860 -9340 6950 -9310
rect 6860 -9360 6920 -9340
rect 22920 -9350 22970 -9300
rect 23840 -9310 23900 -6530
rect 23820 -9340 23900 -9310
rect 23840 -9360 23900 -9340
<< pwell >>
rect 10620 80 10740 130
rect 12500 80 12620 130
rect 14380 80 14500 130
rect 16260 80 16380 130
rect 18140 80 18260 130
rect 20020 80 20140 130
rect 21900 80 22020 130
rect 6940 -11180 6990 -11130
rect 23770 -11180 23820 -11130
<< psubdiff >>
rect 6810 80 6920 110
rect 10620 80 10740 110
rect 12500 80 12620 110
rect 14380 80 14500 110
rect 16260 80 16380 110
rect 18140 80 18260 110
rect 20020 80 20140 110
rect 21900 80 22020 110
rect 23840 80 23950 110
rect 6810 -2820 6860 -2790
rect 23900 -2820 23950 -2790
rect 6810 -3220 6840 -2820
rect 23920 -3220 23950 -2820
rect 6810 -3250 6920 -3220
rect 23840 -3250 23950 -3220
rect 6810 -6150 6860 -6120
rect 23900 -6150 23950 -6120
rect 6810 -6480 6840 -6150
rect 23920 -6480 23950 -6150
rect 6810 -6510 6920 -6480
rect 23840 -6510 23950 -6480
rect 6810 -9410 6860 -9380
rect 23900 -9410 23950 -9380
rect 6810 -9980 6840 -9410
rect 23920 -9980 23950 -9410
rect 6810 -10010 6920 -9980
rect 23840 -10010 23950 -9980
rect 6810 -11170 6920 -11140
rect 6940 -11170 6990 -11140
rect 23770 -11170 23820 -11140
rect 23840 -11170 23950 -11140
<< nsubdiff >>
rect 6880 10 6950 40
rect 7790 10 7840 40
rect 22920 10 22970 40
rect 23770 10 23880 40
rect 6880 -2750 6950 -2720
rect 7790 -2750 7840 -2720
rect 22920 -2750 22970 -2720
rect 23770 -2750 23880 -2720
rect 6880 -3320 6950 -3290
rect 7790 -3320 7840 -3290
rect 22920 -3320 22970 -3290
rect 23770 -3320 23880 -3290
rect 6880 -6080 6950 -6050
rect 7790 -6080 7840 -6050
rect 22920 -6080 22970 -6050
rect 23770 -6080 23880 -6050
rect 6880 -6580 6950 -6550
rect 7790 -6580 7840 -6550
rect 22920 -6580 22970 -6550
rect 23820 -6580 23880 -6550
rect 6880 -9340 6950 -9310
rect 22920 -9340 22970 -9310
rect 23820 -9340 23880 -9310
<< psubdiffcont >>
rect 6810 -2790 6840 80
rect 23920 -2790 23950 80
rect 6860 -2820 23900 -2790
rect 6810 -6120 6840 -3250
rect 23920 -6120 23950 -3250
rect 6860 -6150 23900 -6120
rect 6810 -9380 6840 -6510
rect 23920 -9380 23950 -6510
rect 6860 -9410 23900 -9380
rect 6810 -11140 6840 -10010
rect 23920 -11140 23950 -10010
<< nsubdiffcont >>
rect 6880 -2720 6910 10
rect 23850 -2720 23880 10
rect 6880 -6050 6910 -3320
rect 23850 -6050 23880 -3320
rect 6880 -9310 6910 -6580
rect 23850 -9310 23880 -6580
<< locali >>
rect 5130 -2880 5300 940
rect 5330 -2880 5500 940
rect 5530 -2880 5700 940
rect 5730 -2880 5900 940
rect 6810 80 6920 110
rect 10620 80 10740 110
rect 12500 80 12620 110
rect 14380 80 14500 110
rect 16260 80 16380 110
rect 18140 80 18260 110
rect 20020 80 20140 110
rect 21900 80 22020 110
rect 23840 80 23950 110
rect 7790 40 7840 50
rect 6880 10 6950 40
rect 7790 10 7800 40
rect 7830 10 7840 40
rect 7790 0 7840 10
rect 22920 40 22970 50
rect 22920 10 22930 40
rect 22960 10 22970 40
rect 23770 10 23880 40
rect 22920 0 22970 10
rect 7790 -2720 7840 -2710
rect 6880 -2750 6950 -2720
rect 7790 -2750 7800 -2720
rect 7830 -2750 7840 -2720
rect 7790 -2760 7840 -2750
rect 22920 -2720 22970 -2710
rect 22920 -2750 22930 -2720
rect 22960 -2750 22970 -2720
rect 23770 -2750 23880 -2720
rect 22920 -2760 22970 -2750
rect 6810 -2820 6860 -2790
rect 23900 -2820 23950 -2790
rect 5130 -2970 23840 -2880
rect 5130 -6210 5300 -2970
rect 5330 -6210 5500 -2970
rect 5530 -6210 5700 -2970
rect 5730 -6210 5900 -2970
rect 23920 -3220 23950 -2820
rect 6810 -3250 6920 -3220
rect 23840 -3250 23950 -3220
rect 7790 -3290 7840 -3280
rect 6880 -3320 6950 -3290
rect 7790 -3320 7800 -3290
rect 7830 -3320 7840 -3290
rect 7790 -3330 7840 -3320
rect 22920 -3290 22970 -3280
rect 22920 -3320 22930 -3290
rect 22960 -3320 22970 -3290
rect 23770 -3320 23880 -3290
rect 22920 -3330 22970 -3320
rect 7790 -6050 7840 -6040
rect 6880 -6080 6950 -6050
rect 7790 -6080 7800 -6050
rect 7830 -6080 7840 -6050
rect 7790 -6090 7840 -6080
rect 22920 -6050 22970 -6040
rect 22920 -6080 22930 -6050
rect 22960 -6080 22970 -6050
rect 23770 -6080 23880 -6050
rect 22920 -6090 22970 -6080
rect 6810 -6150 6860 -6120
rect 23900 -6150 23950 -6120
rect 5100 -6300 23840 -6210
rect 5130 -6330 5300 -6300
rect 5330 -6330 5500 -6300
rect 5530 -6330 5700 -6300
rect 5730 -6330 5900 -6300
rect 5100 -6420 23840 -6330
rect 5130 -9470 5300 -6420
rect 5330 -9470 5500 -6420
rect 5530 -9470 5700 -6420
rect 5730 -9470 5900 -6420
rect 23920 -6480 23950 -6150
rect 6810 -6510 6920 -6480
rect 23840 -6510 23950 -6480
rect 7790 -6550 7840 -6540
rect 6880 -6580 6950 -6550
rect 7790 -6580 7800 -6550
rect 7830 -6580 7840 -6550
rect 7790 -6590 7840 -6580
rect 22920 -6550 22970 -6540
rect 22920 -6580 22930 -6550
rect 22960 -6580 22970 -6550
rect 23840 -6580 23880 -6550
rect 22920 -6590 22970 -6580
rect 7790 -9310 7840 -9300
rect 6880 -9340 6950 -9310
rect 7790 -9340 7800 -9310
rect 7830 -9340 7840 -9310
rect 7790 -9350 7840 -9340
rect 22920 -9310 22970 -9300
rect 22920 -9340 22930 -9310
rect 22960 -9340 22970 -9310
rect 23820 -9340 23880 -9310
rect 22920 -9350 22970 -9340
rect 6810 -9410 6860 -9380
rect 23900 -9410 23950 -9380
rect 5100 -9560 23840 -9470
rect 5130 -9590 5300 -9560
rect 5330 -9590 5500 -9560
rect 5530 -9590 5700 -9560
rect 5730 -9590 5900 -9560
rect 5100 -9680 23840 -9590
rect 5130 -9710 5300 -9680
rect 5330 -9710 5500 -9680
rect 5530 -9710 5700 -9680
rect 5730 -9710 5900 -9680
rect 5100 -9800 23840 -9710
rect 5130 -9830 5300 -9800
rect 5330 -9830 5500 -9800
rect 5530 -9830 5700 -9800
rect 5730 -9830 5900 -9800
rect 5100 -9920 23840 -9830
rect 5130 -12000 5300 -9920
rect 5330 -12000 5500 -9920
rect 5530 -12000 5700 -9920
rect 5730 -12000 5900 -9920
rect 23770 -9980 23820 -9970
rect 23920 -9980 23950 -9410
rect 6810 -10010 6920 -9980
rect 23770 -10010 23780 -9980
rect 23810 -10010 23820 -9980
rect 23840 -10010 23950 -9980
rect 23770 -10020 23820 -10010
rect 23770 -11140 23820 -11130
rect 6810 -11170 6920 -11140
rect 6940 -11170 6950 -11140
rect 6980 -11170 6990 -11140
rect 23770 -11170 23780 -11140
rect 23810 -11170 23820 -11140
rect 23830 -11170 23950 -11140
rect 23770 -11180 23820 -11170
<< viali >>
rect 7800 10 7830 40
rect 22930 10 22960 40
rect 7800 -2750 7830 -2720
rect 22930 -2750 22960 -2720
rect 7800 -3320 7830 -3290
rect 22930 -3320 22960 -3290
rect 7800 -6080 7830 -6050
rect 22930 -6080 22960 -6050
rect 7800 -6580 7830 -6550
rect 22930 -6580 22960 -6550
rect 7800 -9340 7830 -9310
rect 22930 -9340 22960 -9310
rect 6950 -10010 6980 -9980
rect 23780 -10010 23810 -9980
rect 6950 -11170 6980 -11140
rect 23780 -11170 23810 -11140
<< metal1 >>
rect 5100 -2840 5130 940
rect 5300 -2840 5330 940
rect 5500 -2840 5530 940
rect 5700 -2840 5730 940
rect 5900 -2840 5930 940
rect 7800 50 7830 130
rect 8740 110 8770 130
rect 8830 110 8860 130
rect 10620 110 10650 130
rect 10710 110 10740 130
rect 12500 110 12530 130
rect 12590 110 12620 130
rect 14380 110 14410 130
rect 14470 110 14500 130
rect 16260 110 16290 130
rect 16350 110 16380 130
rect 18140 110 18170 130
rect 18230 110 18260 130
rect 20020 110 20050 130
rect 20110 110 20140 130
rect 21900 110 21930 130
rect 21990 110 22020 130
rect 22930 50 22960 130
rect 7790 40 7840 50
rect 7790 10 7800 40
rect 7830 10 7840 40
rect 7790 0 7840 10
rect 22920 40 22970 50
rect 22920 10 22930 40
rect 22960 10 22970 40
rect 22920 0 22970 10
rect 7800 -2710 7830 0
rect 22930 -2710 22960 0
rect 7790 -2720 7840 -2710
rect 7790 -2750 7800 -2720
rect 7830 -2750 7840 -2720
rect 7790 -2760 7840 -2750
rect 22920 -2720 22970 -2710
rect 22920 -2750 22930 -2720
rect 22960 -2750 22970 -2720
rect 22920 -2760 22970 -2750
rect 5090 -2850 5140 -2840
rect 5090 -2880 5100 -2850
rect 5130 -2880 5140 -2850
rect 5090 -2890 5140 -2880
rect 5290 -2850 5340 -2840
rect 5290 -2880 5300 -2850
rect 5330 -2880 5340 -2850
rect 5290 -2890 5340 -2880
rect 5490 -2850 5540 -2840
rect 5490 -2880 5500 -2850
rect 5530 -2880 5540 -2850
rect 5490 -2890 5540 -2880
rect 5690 -2850 5740 -2840
rect 5690 -2880 5700 -2850
rect 5730 -2880 5740 -2850
rect 5690 -2890 5740 -2880
rect 5890 -2850 5940 -2840
rect 5890 -2880 5900 -2850
rect 5930 -2880 5940 -2850
rect 5890 -2890 5940 -2880
rect 5100 -2960 5130 -2890
rect 5300 -2960 5330 -2890
rect 5500 -2960 5530 -2890
rect 5700 -2960 5730 -2890
rect 5790 -2950 5840 -2900
rect 5900 -2960 5930 -2890
rect 7070 -2910 7100 -2840
rect 7070 -2950 7100 -2940
rect 5090 -2970 5140 -2960
rect 5090 -3000 5100 -2970
rect 5130 -3000 5140 -2970
rect 5090 -3010 5140 -3000
rect 5290 -2970 5340 -2960
rect 5290 -3000 5300 -2970
rect 5330 -3000 5340 -2970
rect 5290 -3010 5340 -3000
rect 5490 -2970 5540 -2960
rect 5490 -3000 5500 -2970
rect 5530 -3000 5540 -2970
rect 5490 -3010 5540 -3000
rect 5690 -2970 5740 -2960
rect 5690 -3000 5700 -2970
rect 5730 -3000 5740 -2970
rect 5690 -3010 5740 -3000
rect 5890 -2970 5940 -2960
rect 5890 -3000 5900 -2970
rect 5930 -3000 5940 -2970
rect 5890 -3010 5940 -3000
rect 5100 -6170 5130 -3010
rect 5300 -6170 5330 -3010
rect 5500 -6170 5530 -3010
rect 5700 -6170 5730 -3010
rect 5900 -6170 5930 -3010
rect 7800 -3040 7830 -2760
rect 8010 -2910 8040 -2840
rect 8010 -2950 8040 -2940
rect 8740 -2910 8770 -2840
rect 8740 -2950 8770 -2940
rect 7800 -3280 7830 -3180
rect 8740 -3040 8770 -3030
rect 8740 -3200 8770 -3180
rect 8830 -3040 8860 -2840
rect 9560 -2910 9590 -2840
rect 9560 -2950 9590 -2940
rect 9890 -2910 9920 -2840
rect 9890 -2950 9920 -2940
rect 8830 -3200 8860 -3180
rect 10620 -3040 10650 -2840
rect 10710 -2910 10740 -2840
rect 10710 -2950 10740 -2940
rect 11440 -2910 11470 -2840
rect 11440 -2950 11470 -2940
rect 11770 -2910 11800 -2840
rect 11770 -2950 11800 -2940
rect 12500 -2910 12530 -2840
rect 12500 -2950 12530 -2940
rect 10620 -3200 10650 -3180
rect 10710 -3040 10740 -3030
rect 10710 -3200 10740 -3180
rect 12500 -3040 12530 -3030
rect 12500 -3200 12530 -3180
rect 12590 -3040 12620 -2840
rect 13320 -2910 13350 -2840
rect 13320 -2950 13350 -2940
rect 13650 -2910 13680 -2840
rect 13650 -2950 13680 -2940
rect 12590 -3200 12620 -3180
rect 14380 -3040 14410 -2840
rect 14470 -2910 14500 -2840
rect 14470 -2950 14500 -2940
rect 15200 -2910 15230 -2840
rect 15200 -2950 15230 -2940
rect 15530 -2910 15560 -2840
rect 15530 -2950 15560 -2940
rect 16260 -2910 16290 -2840
rect 16260 -2950 16290 -2940
rect 14380 -3200 14410 -3180
rect 14470 -3040 14500 -3030
rect 14470 -3200 14500 -3180
rect 16260 -3040 16290 -3030
rect 16260 -3200 16290 -3180
rect 16350 -3040 16380 -2840
rect 17080 -2910 17110 -2840
rect 17080 -2950 17110 -2940
rect 17410 -2910 17440 -2840
rect 17410 -2950 17440 -2940
rect 16350 -3200 16380 -3180
rect 18140 -3040 18170 -2840
rect 18230 -2910 18260 -2840
rect 18230 -2950 18260 -2940
rect 18960 -2910 18990 -2840
rect 18960 -2950 18990 -2940
rect 19290 -2910 19320 -2840
rect 19290 -2950 19320 -2940
rect 20020 -2910 20050 -2840
rect 20020 -2950 20050 -2940
rect 18140 -3200 18170 -3180
rect 18230 -3040 18260 -3030
rect 18230 -3200 18260 -3180
rect 20020 -3040 20050 -3030
rect 20020 -3200 20050 -3180
rect 20110 -3040 20140 -2840
rect 20840 -2910 20870 -2840
rect 20840 -2950 20870 -2940
rect 21170 -2910 21200 -2840
rect 21170 -2950 21200 -2940
rect 20110 -3200 20140 -3180
rect 21900 -3040 21930 -2840
rect 21990 -2910 22020 -2840
rect 21990 -2950 22020 -2940
rect 22720 -2910 22750 -2840
rect 22720 -2950 22750 -2940
rect 21900 -3200 21930 -3180
rect 21990 -3040 22020 -3030
rect 21990 -3200 22020 -3180
rect 22930 -3280 22960 -2760
rect 23660 -2910 23690 -2840
rect 23660 -2950 23690 -2940
rect 7790 -3290 7840 -3280
rect 7790 -3320 7800 -3290
rect 7830 -3320 7840 -3290
rect 7790 -3330 7840 -3320
rect 22920 -3290 22970 -3280
rect 22920 -3320 22930 -3290
rect 22960 -3320 22970 -3290
rect 22920 -3330 22970 -3320
rect 5090 -6180 5140 -6170
rect 5090 -6210 5100 -6180
rect 5130 -6210 5140 -6180
rect 5090 -6220 5140 -6210
rect 5290 -6180 5340 -6170
rect 5290 -6210 5300 -6180
rect 5330 -6210 5340 -6180
rect 5290 -6220 5340 -6210
rect 5490 -6180 5540 -6170
rect 5490 -6210 5500 -6180
rect 5530 -6210 5540 -6180
rect 5490 -6220 5540 -6210
rect 5690 -6180 5740 -6170
rect 5690 -6210 5700 -6180
rect 5730 -6210 5740 -6180
rect 5690 -6220 5740 -6210
rect 5890 -6180 5940 -6170
rect 5890 -6210 5900 -6180
rect 5930 -6210 5940 -6180
rect 5890 -6220 5940 -6210
rect 5100 -6290 5130 -6220
rect 5300 -6290 5330 -6220
rect 5500 -6290 5530 -6220
rect 5700 -6290 5730 -6220
rect 5900 -6290 5930 -6220
rect 7070 -6240 7100 -6030
rect 7800 -6040 7830 -3330
rect 22930 -6040 22960 -3330
rect 7790 -6050 7840 -6040
rect 7790 -6080 7800 -6050
rect 7830 -6080 7840 -6050
rect 7790 -6090 7840 -6080
rect 22920 -6050 22970 -6040
rect 22920 -6080 22930 -6050
rect 22960 -6080 22970 -6050
rect 22920 -6090 22970 -6080
rect 7070 -6280 7100 -6270
rect 5090 -6300 5140 -6290
rect 5090 -6330 5100 -6300
rect 5130 -6330 5140 -6300
rect 5090 -6340 5140 -6330
rect 5290 -6300 5340 -6290
rect 5290 -6330 5300 -6300
rect 5330 -6330 5340 -6300
rect 5290 -6340 5340 -6330
rect 5490 -6300 5540 -6290
rect 5490 -6330 5500 -6300
rect 5530 -6330 5540 -6300
rect 5490 -6340 5540 -6330
rect 5690 -6300 5740 -6290
rect 5690 -6330 5700 -6300
rect 5730 -6330 5740 -6300
rect 5690 -6340 5740 -6330
rect 5890 -6300 5940 -6290
rect 5890 -6330 5900 -6300
rect 5930 -6330 5940 -6300
rect 5890 -6340 5940 -6330
rect 5100 -6410 5130 -6340
rect 5300 -6410 5330 -6340
rect 5500 -6410 5530 -6340
rect 5700 -6410 5730 -6340
rect 5900 -6410 5930 -6340
rect 5090 -6420 5140 -6410
rect 5090 -6450 5100 -6420
rect 5130 -6450 5140 -6420
rect 5090 -6460 5140 -6450
rect 5290 -6420 5340 -6410
rect 5290 -6450 5300 -6420
rect 5330 -6450 5340 -6420
rect 5290 -6460 5340 -6450
rect 5490 -6420 5540 -6410
rect 5490 -6450 5500 -6420
rect 5530 -6450 5540 -6420
rect 5490 -6460 5540 -6450
rect 5690 -6420 5740 -6410
rect 5690 -6450 5700 -6420
rect 5730 -6450 5740 -6420
rect 5690 -6460 5740 -6450
rect 5890 -6420 5940 -6410
rect 5890 -6450 5900 -6420
rect 5930 -6450 5940 -6420
rect 5890 -6460 5940 -6450
rect 5100 -9430 5130 -6460
rect 5300 -9430 5330 -6460
rect 5500 -9430 5530 -6460
rect 5700 -9430 5730 -6460
rect 5900 -9430 5930 -6460
rect 7800 -6540 7830 -6090
rect 8010 -6240 8040 -6170
rect 8010 -6280 8040 -6270
rect 8740 -6360 8770 -6170
rect 8740 -6460 8770 -6390
rect 8830 -6360 8860 -6170
rect 9560 -6240 9590 -6170
rect 9560 -6280 9590 -6270
rect 9890 -6240 9920 -6170
rect 9890 -6280 9920 -6270
rect 8830 -6460 8860 -6390
rect 10620 -6360 10650 -6170
rect 10620 -6460 10650 -6390
rect 10710 -6360 10740 -6170
rect 11440 -6240 11470 -6170
rect 11440 -6280 11470 -6270
rect 11770 -6240 11800 -6170
rect 11770 -6280 11800 -6270
rect 10710 -6460 10740 -6390
rect 12500 -6360 12530 -6170
rect 12500 -6460 12530 -6390
rect 12590 -6360 12620 -6170
rect 13320 -6240 13350 -6170
rect 13320 -6280 13350 -6270
rect 13650 -6240 13680 -6170
rect 13650 -6280 13680 -6270
rect 12590 -6460 12620 -6390
rect 14380 -6360 14410 -6170
rect 14380 -6460 14410 -6390
rect 14470 -6360 14500 -6170
rect 15200 -6240 15230 -6170
rect 15200 -6280 15230 -6270
rect 15530 -6240 15560 -6170
rect 15530 -6280 15560 -6270
rect 14470 -6460 14500 -6390
rect 16260 -6360 16290 -6170
rect 16260 -6460 16290 -6390
rect 16350 -6360 16380 -6170
rect 17080 -6240 17110 -6170
rect 17080 -6280 17110 -6270
rect 17410 -6240 17440 -6170
rect 17410 -6280 17440 -6270
rect 16350 -6460 16380 -6390
rect 18140 -6360 18170 -6170
rect 18140 -6460 18170 -6390
rect 18230 -6360 18260 -6170
rect 18960 -6240 18990 -6170
rect 18960 -6280 18990 -6270
rect 19290 -6240 19320 -6170
rect 19290 -6280 19320 -6270
rect 18230 -6460 18260 -6390
rect 20020 -6360 20050 -6170
rect 20020 -6460 20050 -6390
rect 20110 -6360 20140 -6170
rect 20840 -6240 20870 -6170
rect 20840 -6280 20870 -6270
rect 21170 -6240 21200 -6170
rect 21170 -6280 21200 -6270
rect 20110 -6460 20140 -6390
rect 21900 -6360 21930 -6170
rect 21900 -6460 21930 -6390
rect 21990 -6360 22020 -6170
rect 22720 -6240 22750 -6170
rect 22720 -6280 22750 -6270
rect 21990 -6460 22020 -6390
rect 22930 -6540 22960 -6090
rect 23660 -6240 23690 -6170
rect 23660 -6280 23690 -6270
rect 7790 -6550 7840 -6540
rect 7790 -6580 7800 -6550
rect 7830 -6580 7840 -6550
rect 7790 -6590 7840 -6580
rect 22920 -6550 22970 -6540
rect 22920 -6580 22930 -6550
rect 22960 -6580 22970 -6550
rect 22920 -6590 22970 -6580
rect 7800 -9300 7830 -6590
rect 22930 -9300 22960 -6590
rect 7790 -9310 7840 -9300
rect 7790 -9340 7800 -9310
rect 7830 -9340 7840 -9310
rect 7790 -9350 7840 -9340
rect 22920 -9310 22970 -9300
rect 22920 -9340 22930 -9310
rect 22960 -9340 22970 -9310
rect 22920 -9350 22970 -9340
rect 7800 -9430 7830 -9350
rect 22930 -9430 22960 -9350
rect 5090 -9440 5140 -9430
rect 5090 -9470 5100 -9440
rect 5130 -9470 5140 -9440
rect 5090 -9480 5140 -9470
rect 5290 -9440 5340 -9430
rect 5290 -9470 5300 -9440
rect 5330 -9470 5340 -9440
rect 5290 -9480 5340 -9470
rect 5490 -9440 5540 -9430
rect 5490 -9470 5500 -9440
rect 5530 -9470 5540 -9440
rect 5490 -9480 5540 -9470
rect 5690 -9440 5740 -9430
rect 5690 -9470 5700 -9440
rect 5730 -9470 5740 -9440
rect 5690 -9480 5740 -9470
rect 5890 -9440 5940 -9430
rect 5890 -9470 5900 -9440
rect 5930 -9470 5940 -9440
rect 5890 -9480 5940 -9470
rect 5100 -9550 5130 -9480
rect 5300 -9550 5330 -9480
rect 5500 -9550 5530 -9480
rect 5700 -9550 5730 -9480
rect 5900 -9550 5930 -9480
rect 5090 -9560 5140 -9550
rect 5090 -9590 5100 -9560
rect 5130 -9590 5140 -9560
rect 5090 -9600 5140 -9590
rect 5290 -9560 5340 -9550
rect 5290 -9590 5300 -9560
rect 5330 -9590 5340 -9560
rect 5290 -9600 5340 -9590
rect 5490 -9560 5540 -9550
rect 5490 -9590 5500 -9560
rect 5530 -9590 5540 -9560
rect 5490 -9600 5540 -9590
rect 5690 -9560 5740 -9550
rect 5690 -9590 5700 -9560
rect 5730 -9590 5740 -9560
rect 5690 -9600 5740 -9590
rect 5890 -9560 5940 -9550
rect 5890 -9590 5900 -9560
rect 5930 -9590 5940 -9560
rect 5890 -9600 5940 -9590
rect 5100 -9670 5130 -9600
rect 5300 -9670 5330 -9600
rect 5500 -9670 5530 -9600
rect 5700 -9670 5730 -9600
rect 5900 -9670 5930 -9600
rect 5090 -9680 5140 -9670
rect 5090 -9710 5100 -9680
rect 5130 -9710 5140 -9680
rect 5090 -9720 5140 -9710
rect 5290 -9680 5340 -9670
rect 5290 -9710 5300 -9680
rect 5330 -9710 5340 -9680
rect 5290 -9720 5340 -9710
rect 5490 -9680 5540 -9670
rect 5490 -9710 5500 -9680
rect 5530 -9710 5540 -9680
rect 5490 -9720 5540 -9710
rect 5690 -9680 5740 -9670
rect 5690 -9710 5700 -9680
rect 5730 -9710 5740 -9680
rect 5690 -9720 5740 -9710
rect 5890 -9680 5940 -9670
rect 5890 -9710 5900 -9680
rect 5930 -9710 5940 -9680
rect 5890 -9720 5940 -9710
rect 5100 -9790 5130 -9720
rect 5300 -9790 5330 -9720
rect 5500 -9790 5530 -9720
rect 5700 -9790 5730 -9720
rect 5900 -9790 5930 -9720
rect 7070 -9740 7100 -9430
rect 8010 -9500 8040 -9430
rect 8010 -9540 8040 -9530
rect 7070 -9780 7100 -9770
rect 7680 -9740 7710 -9730
rect 5090 -9800 5140 -9790
rect 5090 -9830 5100 -9800
rect 5130 -9830 5140 -9800
rect 5090 -9840 5140 -9830
rect 5290 -9800 5340 -9790
rect 5290 -9830 5300 -9800
rect 5330 -9830 5340 -9800
rect 5290 -9840 5340 -9830
rect 5490 -9800 5540 -9790
rect 5490 -9830 5500 -9800
rect 5530 -9830 5540 -9800
rect 5490 -9840 5540 -9830
rect 5690 -9800 5740 -9790
rect 5690 -9830 5700 -9800
rect 5730 -9830 5740 -9800
rect 5690 -9840 5740 -9830
rect 5890 -9800 5940 -9790
rect 5890 -9830 5900 -9800
rect 5930 -9830 5940 -9800
rect 5890 -9840 5940 -9830
rect 5100 -9910 5130 -9840
rect 5300 -9910 5330 -9840
rect 5500 -9910 5530 -9840
rect 5700 -9910 5730 -9840
rect 5900 -9910 5930 -9840
rect 5090 -9920 5140 -9910
rect 5090 -9950 5100 -9920
rect 5130 -9950 5140 -9920
rect 5090 -9960 5140 -9950
rect 5290 -9920 5340 -9910
rect 5290 -9950 5300 -9920
rect 5330 -9950 5340 -9920
rect 5290 -9960 5340 -9950
rect 5490 -9920 5540 -9910
rect 5490 -9950 5500 -9920
rect 5530 -9950 5540 -9920
rect 5490 -9960 5540 -9950
rect 5690 -9920 5740 -9910
rect 5690 -9950 5700 -9920
rect 5730 -9950 5740 -9920
rect 5690 -9960 5740 -9950
rect 5890 -9920 5940 -9910
rect 5890 -9950 5900 -9920
rect 5930 -9950 5940 -9920
rect 5890 -9960 5940 -9950
rect 7680 -9960 7710 -9770
rect 7890 -9740 7920 -9730
rect 7890 -9960 7920 -9770
rect 8620 -9740 8650 -9730
rect 8620 -9960 8650 -9770
rect 8740 -9740 8770 -9430
rect 8740 -9780 8770 -9770
rect 8830 -9860 8860 -9430
rect 9560 -9620 9590 -9430
rect 9560 -9660 9590 -9650
rect 9890 -9620 9920 -9430
rect 9890 -9660 9920 -9650
rect 8830 -9900 8860 -9890
rect 8950 -9740 8980 -9730
rect 8950 -9960 8980 -9770
rect 10500 -9740 10530 -9730
rect 9680 -9860 9710 -9850
rect 9680 -9960 9710 -9890
rect 9770 -9860 9800 -9850
rect 9770 -9960 9800 -9890
rect 10500 -9960 10530 -9770
rect 10620 -9860 10650 -9430
rect 10710 -9740 10740 -9430
rect 11440 -9500 11470 -9430
rect 11440 -9540 11470 -9530
rect 11770 -9500 11800 -9430
rect 11770 -9540 11800 -9530
rect 10710 -9780 10740 -9770
rect 10830 -9740 10860 -9730
rect 10620 -9900 10650 -9890
rect 10830 -9960 10860 -9770
rect 11560 -9740 11590 -9730
rect 11560 -9960 11590 -9770
rect 11650 -9740 11680 -9730
rect 11650 -9960 11680 -9770
rect 12380 -9740 12410 -9730
rect 12380 -9960 12410 -9770
rect 12500 -9740 12530 -9430
rect 12500 -9780 12530 -9770
rect 12590 -9860 12620 -9430
rect 13320 -9620 13350 -9430
rect 13320 -9660 13350 -9650
rect 13650 -9620 13680 -9430
rect 13650 -9660 13680 -9650
rect 12590 -9900 12620 -9890
rect 12710 -9740 12740 -9730
rect 12710 -9960 12740 -9770
rect 14260 -9740 14290 -9730
rect 13440 -9860 13470 -9850
rect 13440 -9960 13470 -9890
rect 13530 -9860 13560 -9850
rect 13530 -9960 13560 -9890
rect 14260 -9960 14290 -9770
rect 14380 -9860 14410 -9430
rect 14470 -9740 14500 -9430
rect 15200 -9500 15230 -9430
rect 15200 -9540 15230 -9530
rect 15530 -9500 15560 -9430
rect 15530 -9540 15560 -9530
rect 14470 -9780 14500 -9770
rect 14590 -9740 14620 -9730
rect 14380 -9900 14410 -9890
rect 14590 -9960 14620 -9770
rect 15320 -9740 15350 -9730
rect 15320 -9960 15350 -9770
rect 15410 -9740 15440 -9730
rect 15410 -9960 15440 -9770
rect 16140 -9740 16170 -9730
rect 16140 -9960 16170 -9770
rect 16260 -9740 16290 -9430
rect 16260 -9780 16290 -9770
rect 16350 -9860 16380 -9430
rect 17080 -9620 17110 -9430
rect 17080 -9660 17110 -9650
rect 17410 -9620 17440 -9430
rect 17410 -9660 17440 -9650
rect 16350 -9900 16380 -9890
rect 16470 -9740 16500 -9730
rect 16470 -9960 16500 -9770
rect 18020 -9740 18050 -9730
rect 17200 -9860 17230 -9850
rect 17200 -9960 17230 -9890
rect 17290 -9860 17320 -9850
rect 17290 -9960 17320 -9890
rect 18020 -9960 18050 -9770
rect 18140 -9860 18170 -9430
rect 18230 -9740 18260 -9430
rect 18960 -9500 18990 -9430
rect 18960 -9540 18990 -9530
rect 19290 -9500 19320 -9430
rect 19290 -9540 19320 -9530
rect 18230 -9780 18260 -9770
rect 18350 -9740 18380 -9730
rect 18140 -9900 18170 -9890
rect 18350 -9960 18380 -9770
rect 19080 -9740 19110 -9730
rect 19080 -9960 19110 -9770
rect 19170 -9740 19200 -9730
rect 19170 -9960 19200 -9770
rect 19900 -9740 19930 -9730
rect 19900 -9960 19930 -9770
rect 20020 -9740 20050 -9430
rect 20020 -9780 20050 -9770
rect 20110 -9860 20140 -9430
rect 20840 -9620 20870 -9430
rect 20840 -9660 20870 -9650
rect 21170 -9620 21200 -9430
rect 21170 -9660 21200 -9650
rect 20110 -9900 20140 -9890
rect 20230 -9740 20260 -9730
rect 20230 -9960 20260 -9770
rect 21780 -9740 21810 -9730
rect 20960 -9860 20990 -9850
rect 20960 -9960 20990 -9890
rect 21050 -9860 21080 -9850
rect 21050 -9960 21080 -9890
rect 21780 -9960 21810 -9770
rect 21900 -9860 21930 -9430
rect 21990 -9740 22020 -9430
rect 22720 -9500 22750 -9430
rect 22720 -9540 22750 -9530
rect 21990 -9780 22020 -9770
rect 22110 -9740 22140 -9730
rect 21900 -9900 21930 -9890
rect 22110 -9960 22140 -9770
rect 22840 -9740 22870 -9730
rect 22840 -9960 22870 -9770
rect 23050 -9740 23080 -9730
rect 23050 -9960 23080 -9770
rect 23660 -9740 23690 -9430
rect 23660 -9780 23690 -9770
rect 5100 -12000 5130 -9960
rect 5300 -12000 5330 -9960
rect 5500 -12000 5530 -9960
rect 5700 -12000 5730 -9960
rect 5900 -12000 5930 -9960
rect 6950 -9970 6980 -9960
rect 23780 -9970 23810 -9960
rect 6940 -9980 6990 -9970
rect 6940 -10010 6950 -9980
rect 6980 -10010 6990 -9980
rect 6940 -10020 6990 -10010
rect 23770 -9980 23820 -9970
rect 23770 -10010 23780 -9980
rect 23810 -10010 23820 -9980
rect 23770 -10020 23820 -10010
rect 6950 -11130 6980 -10020
rect 23780 -11130 23810 -10020
rect 6940 -11140 6990 -11130
rect 6940 -11170 6950 -11140
rect 6980 -11170 6990 -11140
rect 6940 -11180 6990 -11170
rect 23770 -11140 23820 -11130
rect 23770 -11170 23780 -11140
rect 23810 -11170 23820 -11140
rect 23770 -11180 23820 -11170
rect 6950 -11210 6980 -11180
rect 6950 -11360 6980 -11350
rect 7890 -11210 7920 -11190
rect 7890 -11360 7920 -11350
rect 9680 -11210 9710 -11190
rect 9680 -11360 9710 -11350
rect 9770 -11210 9800 -11190
rect 9770 -11360 9800 -11350
rect 11560 -11210 11590 -11190
rect 11560 -11360 11590 -11350
rect 11650 -11210 11680 -11190
rect 11650 -11360 11680 -11350
rect 13440 -11210 13470 -11190
rect 13440 -11360 13470 -11350
rect 13530 -11210 13560 -11190
rect 13530 -11360 13560 -11350
rect 15320 -11210 15350 -11190
rect 15320 -11360 15350 -11350
rect 15410 -11210 15440 -11190
rect 15410 -11360 15440 -11350
rect 17200 -11210 17230 -11190
rect 17200 -11360 17230 -11350
rect 17290 -11210 17320 -11190
rect 17290 -11360 17320 -11350
rect 19080 -11210 19110 -11190
rect 19080 -11360 19110 -11350
rect 19170 -11210 19200 -11190
rect 19170 -11360 19200 -11350
rect 20960 -11210 20990 -11190
rect 20960 -11360 20990 -11350
rect 21050 -11210 21080 -11190
rect 21050 -11360 21080 -11350
rect 22840 -11210 22870 -11190
rect 22840 -11360 22870 -11350
rect 23780 -11210 23810 -11180
rect 23780 -11360 23810 -11350
<< via1 >>
rect 8740 80 8770 110
rect 8830 80 8860 110
rect 10620 80 10650 110
rect 10710 80 10740 110
rect 12500 80 12530 110
rect 12590 80 12620 110
rect 14380 80 14410 110
rect 14470 80 14500 110
rect 16260 80 16290 110
rect 16350 80 16380 110
rect 18140 80 18170 110
rect 18230 80 18260 110
rect 20020 80 20050 110
rect 20110 80 20140 110
rect 21900 80 21930 110
rect 21990 80 22020 110
rect 5100 -2880 5130 -2850
rect 5300 -2880 5330 -2850
rect 5500 -2880 5530 -2850
rect 5700 -2880 5730 -2850
rect 5900 -2880 5930 -2850
rect 7070 -2940 7100 -2910
rect 5100 -3000 5130 -2970
rect 5300 -3000 5330 -2970
rect 5500 -3000 5530 -2970
rect 5700 -3000 5730 -2970
rect 5900 -3000 5930 -2970
rect 8010 -2940 8040 -2910
rect 8740 -2940 8770 -2910
rect 7800 -3180 7830 -3040
rect 8740 -3180 8770 -3040
rect 9560 -2940 9590 -2910
rect 9890 -2940 9920 -2910
rect 8830 -3180 8860 -3040
rect 10710 -2940 10740 -2910
rect 11440 -2940 11470 -2910
rect 11770 -2940 11800 -2910
rect 12500 -2940 12530 -2910
rect 10620 -3180 10650 -3040
rect 10710 -3180 10740 -3040
rect 12500 -3180 12530 -3040
rect 13320 -2940 13350 -2910
rect 13650 -2940 13680 -2910
rect 12590 -3180 12620 -3040
rect 14470 -2940 14500 -2910
rect 15200 -2940 15230 -2910
rect 15530 -2940 15560 -2910
rect 16260 -2940 16290 -2910
rect 14380 -3180 14410 -3040
rect 14470 -3180 14500 -3040
rect 16260 -3180 16290 -3040
rect 17080 -2940 17110 -2910
rect 17410 -2940 17440 -2910
rect 16350 -3180 16380 -3040
rect 18230 -2940 18260 -2910
rect 18960 -2940 18990 -2910
rect 19290 -2940 19320 -2910
rect 20020 -2940 20050 -2910
rect 18140 -3180 18170 -3040
rect 18230 -3180 18260 -3040
rect 20020 -3180 20050 -3040
rect 20840 -2940 20870 -2910
rect 21170 -2940 21200 -2910
rect 20110 -3180 20140 -3040
rect 21990 -2940 22020 -2910
rect 22720 -2940 22750 -2910
rect 21900 -3180 21930 -3040
rect 21990 -3180 22020 -3040
rect 23660 -2940 23690 -2910
rect 5100 -6210 5130 -6180
rect 5300 -6210 5330 -6180
rect 5500 -6210 5530 -6180
rect 5700 -6210 5730 -6180
rect 5900 -6210 5930 -6180
rect 7070 -6270 7100 -6240
rect 5100 -6330 5130 -6300
rect 5300 -6330 5330 -6300
rect 5500 -6330 5530 -6300
rect 5700 -6330 5730 -6300
rect 5900 -6330 5930 -6300
rect 5100 -6450 5130 -6420
rect 5300 -6450 5330 -6420
rect 5500 -6450 5530 -6420
rect 5700 -6450 5730 -6420
rect 5900 -6450 5930 -6420
rect 8010 -6270 8040 -6240
rect 8740 -6390 8770 -6360
rect 9560 -6270 9590 -6240
rect 9890 -6270 9920 -6240
rect 8830 -6390 8860 -6360
rect 10620 -6390 10650 -6360
rect 11440 -6270 11470 -6240
rect 11770 -6270 11800 -6240
rect 10710 -6390 10740 -6360
rect 12500 -6390 12530 -6360
rect 13320 -6270 13350 -6240
rect 13650 -6270 13680 -6240
rect 12590 -6390 12620 -6360
rect 14380 -6390 14410 -6360
rect 15200 -6270 15230 -6240
rect 15530 -6270 15560 -6240
rect 14470 -6390 14500 -6360
rect 16260 -6390 16290 -6360
rect 17080 -6270 17110 -6240
rect 17410 -6270 17440 -6240
rect 16350 -6390 16380 -6360
rect 18140 -6390 18170 -6360
rect 18960 -6270 18990 -6240
rect 19290 -6270 19320 -6240
rect 18230 -6390 18260 -6360
rect 20020 -6390 20050 -6360
rect 20840 -6270 20870 -6240
rect 21170 -6270 21200 -6240
rect 20110 -6390 20140 -6360
rect 21900 -6390 21930 -6360
rect 22720 -6270 22750 -6240
rect 21990 -6390 22020 -6360
rect 23660 -6270 23690 -6240
rect 5100 -9470 5130 -9440
rect 5300 -9470 5330 -9440
rect 5500 -9470 5530 -9440
rect 5700 -9470 5730 -9440
rect 5900 -9470 5930 -9440
rect 5100 -9590 5130 -9560
rect 5300 -9590 5330 -9560
rect 5500 -9590 5530 -9560
rect 5700 -9590 5730 -9560
rect 5900 -9590 5930 -9560
rect 5100 -9710 5130 -9680
rect 5300 -9710 5330 -9680
rect 5500 -9710 5530 -9680
rect 5700 -9710 5730 -9680
rect 5900 -9710 5930 -9680
rect 8010 -9530 8040 -9500
rect 7070 -9770 7100 -9740
rect 7680 -9770 7710 -9740
rect 5100 -9830 5130 -9800
rect 5300 -9830 5330 -9800
rect 5500 -9830 5530 -9800
rect 5700 -9830 5730 -9800
rect 5900 -9830 5930 -9800
rect 5100 -9950 5130 -9920
rect 5300 -9950 5330 -9920
rect 5500 -9950 5530 -9920
rect 5700 -9950 5730 -9920
rect 5900 -9950 5930 -9920
rect 7890 -9770 7920 -9740
rect 8620 -9770 8650 -9740
rect 8740 -9770 8770 -9740
rect 9560 -9650 9590 -9620
rect 9890 -9650 9920 -9620
rect 8830 -9890 8860 -9860
rect 8950 -9770 8980 -9740
rect 10500 -9770 10530 -9740
rect 9680 -9890 9710 -9860
rect 9770 -9890 9800 -9860
rect 11440 -9530 11470 -9500
rect 11770 -9530 11800 -9500
rect 10710 -9770 10740 -9740
rect 10830 -9770 10860 -9740
rect 10620 -9890 10650 -9860
rect 11560 -9770 11590 -9740
rect 11650 -9770 11680 -9740
rect 12380 -9770 12410 -9740
rect 12500 -9770 12530 -9740
rect 13320 -9650 13350 -9620
rect 13650 -9650 13680 -9620
rect 12590 -9890 12620 -9860
rect 12710 -9770 12740 -9740
rect 14260 -9770 14290 -9740
rect 13440 -9890 13470 -9860
rect 13530 -9890 13560 -9860
rect 15200 -9530 15230 -9500
rect 15530 -9530 15560 -9500
rect 14470 -9770 14500 -9740
rect 14590 -9770 14620 -9740
rect 14380 -9890 14410 -9860
rect 15320 -9770 15350 -9740
rect 15410 -9770 15440 -9740
rect 16140 -9770 16170 -9740
rect 16260 -9770 16290 -9740
rect 17080 -9650 17110 -9620
rect 17410 -9650 17440 -9620
rect 16350 -9890 16380 -9860
rect 16470 -9770 16500 -9740
rect 18020 -9770 18050 -9740
rect 17200 -9890 17230 -9860
rect 17290 -9890 17320 -9860
rect 18960 -9530 18990 -9500
rect 19290 -9530 19320 -9500
rect 18230 -9770 18260 -9740
rect 18350 -9770 18380 -9740
rect 18140 -9890 18170 -9860
rect 19080 -9770 19110 -9740
rect 19170 -9770 19200 -9740
rect 19900 -9770 19930 -9740
rect 20020 -9770 20050 -9740
rect 20840 -9650 20870 -9620
rect 21170 -9650 21200 -9620
rect 20110 -9890 20140 -9860
rect 20230 -9770 20260 -9740
rect 21780 -9770 21810 -9740
rect 20960 -9890 20990 -9860
rect 21050 -9890 21080 -9860
rect 22720 -9530 22750 -9500
rect 21990 -9770 22020 -9740
rect 22110 -9770 22140 -9740
rect 21900 -9890 21930 -9860
rect 22840 -9770 22870 -9740
rect 23050 -9770 23080 -9740
rect 23660 -9770 23690 -9740
rect 6950 -11350 6980 -11210
rect 7890 -11350 7920 -11210
rect 9680 -11350 9710 -11210
rect 9770 -11350 9800 -11210
rect 11560 -11350 11590 -11210
rect 11650 -11350 11680 -11210
rect 13440 -11350 13470 -11210
rect 13530 -11350 13560 -11210
rect 15320 -11350 15350 -11210
rect 15410 -11350 15440 -11210
rect 17200 -11350 17230 -11210
rect 17290 -11350 17320 -11210
rect 19080 -11350 19110 -11210
rect 19170 -11350 19200 -11210
rect 20960 -11350 20990 -11210
rect 21050 -11350 21080 -11210
rect 22840 -11350 22870 -11210
rect 23780 -11350 23810 -11210
<< metal2 >>
rect 8730 80 8740 110
rect 8770 80 8830 110
rect 8860 80 10620 110
rect 10650 80 10710 110
rect 10740 80 12500 110
rect 12530 80 12590 110
rect 12620 80 14380 110
rect 14410 80 14470 110
rect 14500 80 16260 110
rect 16290 80 16350 110
rect 16380 80 18140 110
rect 18170 80 18230 110
rect 18260 80 20020 110
rect 20050 80 20110 110
rect 20140 80 21900 110
rect 21930 80 21990 110
rect 22020 80 22030 110
rect 5090 -2850 5140 -2840
rect 5290 -2850 5340 -2840
rect 5490 -2850 5540 -2840
rect 5690 -2850 5740 -2840
rect 5890 -2850 5940 -2840
rect 6290 -2850 6470 -2840
rect 5090 -2880 5100 -2850
rect 5130 -2880 5300 -2850
rect 5330 -2880 5500 -2850
rect 5530 -2880 5700 -2850
rect 5730 -2880 5900 -2850
rect 5930 -2880 6300 -2850
rect 6460 -2880 23840 -2850
rect 5090 -2890 5140 -2880
rect 5290 -2890 5340 -2880
rect 5490 -2890 5540 -2880
rect 5690 -2890 5740 -2880
rect 5890 -2890 5940 -2880
rect 6290 -2890 6470 -2880
rect 5790 -2910 5840 -2900
rect 5130 -2940 5800 -2910
rect 5830 -2940 7070 -2910
rect 7100 -2940 8010 -2910
rect 8040 -2940 8740 -2910
rect 8770 -2940 9560 -2910
rect 9590 -2940 9890 -2910
rect 9920 -2940 10710 -2910
rect 10740 -2940 11440 -2910
rect 11470 -2940 11770 -2910
rect 11800 -2940 12500 -2910
rect 12530 -2940 13320 -2910
rect 13350 -2940 13650 -2910
rect 13680 -2940 14470 -2910
rect 14500 -2940 15200 -2910
rect 15230 -2940 15530 -2910
rect 15560 -2940 16260 -2910
rect 16290 -2940 17080 -2910
rect 17110 -2940 17410 -2910
rect 17440 -2940 18230 -2910
rect 18260 -2940 18960 -2910
rect 18990 -2940 19290 -2910
rect 19320 -2940 20020 -2910
rect 20050 -2940 20840 -2910
rect 20870 -2940 21170 -2910
rect 21200 -2940 21990 -2910
rect 22020 -2940 22720 -2910
rect 22750 -2940 23660 -2910
rect 23690 -2940 23840 -2910
rect 5790 -2950 5840 -2940
rect 5090 -2970 5140 -2960
rect 5290 -2970 5340 -2960
rect 5490 -2970 5540 -2960
rect 5690 -2970 5740 -2960
rect 5890 -2970 5940 -2960
rect 6290 -2970 6470 -2960
rect 5090 -3000 5100 -2970
rect 5130 -3000 5300 -2970
rect 5330 -3000 5500 -2970
rect 5530 -3000 5700 -2970
rect 5730 -3000 5900 -2970
rect 5930 -3000 6300 -2970
rect 6460 -3000 23840 -2970
rect 5090 -3010 5140 -3000
rect 5290 -3010 5340 -3000
rect 5490 -3010 5540 -3000
rect 5690 -3010 5740 -3000
rect 5890 -3010 5940 -3000
rect 6290 -3010 6470 -3000
rect 5100 -3040 23840 -3030
rect 5100 -3180 5990 -3040
rect 6130 -3180 7800 -3040
rect 7830 -3180 8740 -3040
rect 8770 -3180 8830 -3040
rect 8860 -3180 10620 -3040
rect 10650 -3180 10710 -3040
rect 10740 -3180 12500 -3040
rect 12530 -3180 12590 -3040
rect 12620 -3180 14380 -3040
rect 14410 -3180 14470 -3040
rect 14500 -3180 16260 -3040
rect 16290 -3180 16350 -3040
rect 16380 -3180 18140 -3040
rect 18170 -3180 18230 -3040
rect 18260 -3180 20020 -3040
rect 20050 -3180 20110 -3040
rect 20140 -3180 21900 -3040
rect 21930 -3180 21990 -3040
rect 22020 -3180 23840 -3040
rect 5100 -3190 23840 -3180
rect 5090 -6180 5140 -6170
rect 5290 -6180 5340 -6170
rect 5490 -6180 5540 -6170
rect 5690 -6180 5740 -6170
rect 5890 -6180 5940 -6170
rect 6290 -6180 6470 -6170
rect 5090 -6210 5100 -6180
rect 5130 -6210 5300 -6180
rect 5330 -6210 5500 -6180
rect 5530 -6210 5700 -6180
rect 5730 -6210 5900 -6180
rect 5930 -6210 6300 -6180
rect 6460 -6210 23840 -6180
rect 5090 -6220 5140 -6210
rect 5290 -6220 5340 -6210
rect 5490 -6220 5540 -6210
rect 5690 -6220 5740 -6210
rect 5890 -6220 5940 -6210
rect 6290 -6220 6470 -6210
rect 5790 -6240 5840 -6230
rect 5100 -6270 5800 -6240
rect 5830 -6270 7070 -6240
rect 7100 -6270 8010 -6240
rect 8040 -6270 9560 -6240
rect 9590 -6270 9890 -6240
rect 9920 -6270 11440 -6240
rect 11470 -6270 11770 -6240
rect 11800 -6270 13320 -6240
rect 13350 -6270 13650 -6240
rect 13680 -6270 15200 -6240
rect 15230 -6270 15530 -6240
rect 15560 -6270 17080 -6240
rect 17110 -6270 17410 -6240
rect 17440 -6270 18960 -6240
rect 18990 -6270 19290 -6240
rect 19320 -6270 20840 -6240
rect 20870 -6270 21170 -6240
rect 21200 -6270 22720 -6240
rect 22750 -6270 23660 -6240
rect 23690 -6270 23840 -6240
rect 5790 -6280 5840 -6270
rect 5090 -6300 5140 -6290
rect 5290 -6300 5340 -6290
rect 5490 -6300 5540 -6290
rect 5690 -6300 5740 -6290
rect 5890 -6300 5940 -6290
rect 6290 -6300 6470 -6290
rect 5090 -6330 5100 -6300
rect 5130 -6330 5300 -6300
rect 5330 -6330 5500 -6300
rect 5530 -6330 5700 -6300
rect 5730 -6330 5900 -6300
rect 5930 -6330 6300 -6300
rect 6460 -6330 23840 -6300
rect 5090 -6340 5140 -6330
rect 5290 -6340 5340 -6330
rect 5490 -6340 5540 -6330
rect 5690 -6340 5740 -6330
rect 5890 -6340 5940 -6330
rect 6290 -6340 6470 -6330
rect 5100 -6390 5930 -6360
rect 6810 -6390 8740 -6360
rect 8770 -6390 8830 -6360
rect 8860 -6390 10620 -6360
rect 10650 -6390 10710 -6360
rect 10740 -6390 12500 -6360
rect 12530 -6390 12590 -6360
rect 12620 -6390 14380 -6360
rect 14410 -6390 14470 -6360
rect 14500 -6390 16260 -6360
rect 16290 -6390 16350 -6360
rect 16380 -6390 18140 -6360
rect 18170 -6390 18230 -6360
rect 18260 -6390 20020 -6360
rect 20050 -6390 20110 -6360
rect 20140 -6390 21900 -6360
rect 21930 -6390 21990 -6360
rect 22020 -6390 23840 -6360
rect 5090 -6420 5140 -6410
rect 5290 -6420 5340 -6410
rect 5490 -6420 5540 -6410
rect 5690 -6420 5740 -6410
rect 5890 -6420 5940 -6410
rect 5090 -6450 5100 -6420
rect 5130 -6450 5300 -6420
rect 5330 -6450 5500 -6420
rect 5530 -6450 5700 -6420
rect 5730 -6450 5900 -6420
rect 5930 -6430 23840 -6420
rect 5930 -6450 6300 -6430
rect 5090 -6460 5140 -6450
rect 5290 -6460 5340 -6450
rect 5490 -6460 5540 -6450
rect 5690 -6460 5740 -6450
rect 5890 -6460 5940 -6450
rect 6290 -6460 6300 -6450
rect 6460 -6450 23840 -6430
rect 6460 -6460 6470 -6450
rect 6290 -6470 6470 -6460
rect 5090 -9440 5140 -9430
rect 5290 -9440 5340 -9430
rect 5490 -9440 5540 -9430
rect 5690 -9440 5740 -9430
rect 5890 -9440 5940 -9430
rect 6290 -9440 6470 -9430
rect 5090 -9470 5100 -9440
rect 5130 -9470 5300 -9440
rect 5330 -9470 5500 -9440
rect 5530 -9470 5700 -9440
rect 5730 -9470 5900 -9440
rect 5930 -9470 6300 -9440
rect 6460 -9470 23840 -9440
rect 5090 -9480 5140 -9470
rect 5290 -9480 5340 -9470
rect 5490 -9480 5540 -9470
rect 5690 -9480 5740 -9470
rect 5890 -9480 5940 -9470
rect 6290 -9480 6470 -9470
rect 5390 -9500 5440 -9490
rect 5100 -9530 5400 -9500
rect 5430 -9530 8010 -9500
rect 8040 -9530 11440 -9500
rect 11470 -9530 11770 -9500
rect 11800 -9530 15200 -9500
rect 15230 -9530 15530 -9500
rect 15560 -9530 18960 -9500
rect 18990 -9530 19290 -9500
rect 19320 -9530 22720 -9500
rect 22750 -9530 23840 -9500
rect 5390 -9540 5440 -9530
rect 5090 -9560 5140 -9550
rect 5290 -9560 5340 -9550
rect 5490 -9560 5540 -9550
rect 5690 -9560 5740 -9550
rect 5890 -9560 5940 -9550
rect 6290 -9560 6470 -9550
rect 5090 -9590 5100 -9560
rect 5130 -9590 5300 -9560
rect 5330 -9590 5500 -9560
rect 5530 -9590 5700 -9560
rect 5730 -9590 5900 -9560
rect 5930 -9590 6300 -9560
rect 6460 -9590 23840 -9560
rect 5090 -9600 5140 -9590
rect 5290 -9600 5340 -9590
rect 5490 -9600 5540 -9590
rect 5690 -9600 5740 -9590
rect 5890 -9600 5940 -9590
rect 6290 -9600 6470 -9590
rect 5190 -9620 5240 -9610
rect 5100 -9650 5200 -9620
rect 5230 -9650 9560 -9620
rect 9590 -9650 9890 -9620
rect 9920 -9650 13320 -9620
rect 13350 -9650 13650 -9620
rect 13680 -9650 17080 -9620
rect 17110 -9650 17410 -9620
rect 17440 -9650 20840 -9620
rect 20870 -9650 21170 -9620
rect 21200 -9650 23840 -9620
rect 5190 -9660 5240 -9650
rect 5090 -9680 5140 -9670
rect 5290 -9680 5340 -9670
rect 5490 -9680 5540 -9670
rect 5690 -9680 5740 -9670
rect 5890 -9680 5940 -9670
rect 6290 -9680 6470 -9670
rect 5090 -9710 5100 -9680
rect 5130 -9710 5300 -9680
rect 5330 -9710 5500 -9680
rect 5530 -9710 5700 -9680
rect 5730 -9710 5900 -9680
rect 5930 -9710 6300 -9680
rect 6460 -9710 23840 -9680
rect 5090 -9720 5140 -9710
rect 5290 -9720 5340 -9710
rect 5490 -9720 5540 -9710
rect 5690 -9720 5740 -9710
rect 5890 -9720 5940 -9710
rect 6290 -9720 6470 -9710
rect 5100 -9770 5930 -9740
rect 6840 -9770 7070 -9740
rect 7100 -9770 7680 -9740
rect 7710 -9770 7890 -9740
rect 7920 -9770 8620 -9740
rect 8650 -9770 8740 -9740
rect 8770 -9770 8950 -9740
rect 8980 -9770 10500 -9740
rect 10530 -9770 10710 -9740
rect 10740 -9770 10830 -9740
rect 10860 -9770 11560 -9740
rect 11590 -9770 11650 -9740
rect 11680 -9770 12380 -9740
rect 12410 -9770 12500 -9740
rect 12530 -9770 12710 -9740
rect 12740 -9770 14260 -9740
rect 14290 -9770 14470 -9740
rect 14500 -9770 14590 -9740
rect 14620 -9770 15320 -9740
rect 15350 -9770 15410 -9740
rect 15440 -9770 16140 -9740
rect 16170 -9770 16260 -9740
rect 16290 -9770 16470 -9740
rect 16500 -9770 18020 -9740
rect 18050 -9770 18230 -9740
rect 18260 -9770 18350 -9740
rect 18380 -9770 19080 -9740
rect 19110 -9770 19170 -9740
rect 19200 -9770 19900 -9740
rect 19930 -9770 20020 -9740
rect 20050 -9770 20230 -9740
rect 20260 -9770 21780 -9740
rect 21810 -9770 21990 -9740
rect 22020 -9770 22110 -9740
rect 22140 -9770 22840 -9740
rect 22870 -9770 23050 -9740
rect 23080 -9770 23660 -9740
rect 23690 -9770 23840 -9740
rect 5090 -9800 5140 -9790
rect 5290 -9800 5340 -9790
rect 5490 -9800 5540 -9790
rect 5690 -9800 5740 -9790
rect 5890 -9800 5940 -9790
rect 6290 -9800 6470 -9790
rect 5090 -9830 5100 -9800
rect 5130 -9830 5300 -9800
rect 5330 -9830 5500 -9800
rect 5530 -9830 5700 -9800
rect 5730 -9830 5900 -9800
rect 5930 -9830 6300 -9800
rect 6460 -9830 23840 -9800
rect 5090 -9840 5140 -9830
rect 5290 -9840 5340 -9830
rect 5490 -9840 5540 -9830
rect 5690 -9840 5740 -9830
rect 5890 -9840 5940 -9830
rect 6290 -9840 6470 -9830
rect 5590 -9860 5640 -9850
rect 5100 -9890 5600 -9860
rect 5630 -9890 8830 -9860
rect 8860 -9890 9680 -9860
rect 9710 -9890 9770 -9860
rect 9800 -9890 10620 -9860
rect 10650 -9890 12590 -9860
rect 12620 -9890 13440 -9860
rect 13470 -9890 13530 -9860
rect 13560 -9890 14380 -9860
rect 14410 -9890 16350 -9860
rect 16380 -9890 17200 -9860
rect 17230 -9890 17290 -9860
rect 17320 -9890 18140 -9860
rect 18170 -9890 20110 -9860
rect 20140 -9890 20960 -9860
rect 20990 -9890 21050 -9860
rect 21080 -9890 21900 -9860
rect 21930 -9890 23840 -9860
rect 5590 -9900 5640 -9890
rect 5090 -9920 5140 -9910
rect 5290 -9920 5340 -9910
rect 5490 -9920 5540 -9910
rect 5690 -9920 5740 -9910
rect 5890 -9920 5940 -9910
rect 6290 -9920 6470 -9910
rect 5090 -9950 5100 -9920
rect 5130 -9950 5300 -9920
rect 5330 -9950 5500 -9920
rect 5530 -9950 5700 -9920
rect 5730 -9950 5900 -9920
rect 5930 -9950 6300 -9920
rect 6460 -9950 23840 -9920
rect 5090 -9960 5140 -9950
rect 5290 -9960 5340 -9950
rect 5490 -9960 5540 -9950
rect 5690 -9960 5740 -9950
rect 5890 -9960 5940 -9950
rect 6290 -9960 6470 -9950
rect 6620 -11210 24140 -11200
rect 6620 -11350 6630 -11210
rect 6770 -11350 6950 -11210
rect 6980 -11350 7890 -11210
rect 7920 -11350 9680 -11210
rect 9710 -11350 9770 -11210
rect 9800 -11350 11560 -11210
rect 11590 -11350 11650 -11210
rect 11680 -11350 13440 -11210
rect 13470 -11350 13530 -11210
rect 13560 -11350 15320 -11210
rect 15350 -11350 15410 -11210
rect 15440 -11350 17200 -11210
rect 17230 -11350 17290 -11210
rect 17320 -11350 19080 -11210
rect 19110 -11350 19170 -11210
rect 19200 -11350 20960 -11210
rect 20990 -11350 21050 -11210
rect 21080 -11350 22840 -11210
rect 22870 -11350 23780 -11210
rect 23810 -11350 23990 -11210
rect 24130 -11350 24140 -11210
rect 6620 -11360 24140 -11350
<< via2 >>
rect 5100 -2880 5130 -2850
rect 5300 -2880 5330 -2850
rect 5500 -2880 5530 -2850
rect 5700 -2880 5730 -2850
rect 5900 -2880 5930 -2850
rect 6300 -2880 6460 -2850
rect 5800 -2940 5830 -2910
rect 5100 -3000 5130 -2970
rect 5300 -3000 5330 -2970
rect 5500 -3000 5530 -2970
rect 5700 -3000 5730 -2970
rect 5900 -3000 5930 -2970
rect 6300 -3000 6460 -2970
rect 5990 -3180 6130 -3040
rect 5100 -6210 5130 -6180
rect 5300 -6210 5330 -6180
rect 5500 -6210 5530 -6180
rect 5700 -6210 5730 -6180
rect 5900 -6210 5930 -6180
rect 6300 -6210 6460 -6180
rect 5800 -6270 5830 -6240
rect 5100 -6330 5130 -6300
rect 5300 -6330 5330 -6300
rect 5500 -6330 5530 -6300
rect 5700 -6330 5730 -6300
rect 5900 -6330 5930 -6300
rect 6300 -6330 6460 -6300
rect 5100 -6450 5130 -6420
rect 5300 -6450 5330 -6420
rect 5500 -6450 5530 -6420
rect 5700 -6450 5730 -6420
rect 5900 -6450 5930 -6420
rect 6300 -6460 6460 -6430
rect 5100 -9470 5130 -9440
rect 5300 -9470 5330 -9440
rect 5500 -9470 5530 -9440
rect 5700 -9470 5730 -9440
rect 5900 -9470 5930 -9440
rect 6300 -9470 6460 -9440
rect 5400 -9530 5430 -9500
rect 5100 -9590 5130 -9560
rect 5300 -9590 5330 -9560
rect 5500 -9590 5530 -9560
rect 5700 -9590 5730 -9560
rect 5900 -9590 5930 -9560
rect 6300 -9590 6460 -9560
rect 5200 -9650 5230 -9620
rect 5100 -9710 5130 -9680
rect 5300 -9710 5330 -9680
rect 5500 -9710 5530 -9680
rect 5700 -9710 5730 -9680
rect 5900 -9710 5930 -9680
rect 6300 -9710 6460 -9680
rect 5100 -9830 5130 -9800
rect 5300 -9830 5330 -9800
rect 5500 -9830 5530 -9800
rect 5700 -9830 5730 -9800
rect 5900 -9830 5930 -9800
rect 6300 -9830 6460 -9800
rect 5600 -9890 5630 -9860
rect 5100 -9950 5130 -9920
rect 5300 -9950 5330 -9920
rect 5500 -9950 5530 -9920
rect 5700 -9950 5730 -9920
rect 5900 -9950 5930 -9920
rect 6300 -9950 6460 -9920
rect 6630 -11350 6770 -11210
rect 23990 -11350 24130 -11210
<< metal3 >>
rect 5100 -2840 5130 940
rect 5090 -2850 5140 -2840
rect 5090 -2880 5100 -2850
rect 5130 -2880 5140 -2850
rect 5090 -2890 5140 -2880
rect 5100 -2960 5130 -2890
rect 5090 -2970 5140 -2960
rect 5090 -3000 5100 -2970
rect 5130 -3000 5140 -2970
rect 5090 -3010 5140 -3000
rect 5100 -6170 5130 -3010
rect 5090 -6180 5140 -6170
rect 5090 -6210 5100 -6180
rect 5130 -6210 5140 -6180
rect 5090 -6220 5140 -6210
rect 5100 -6290 5130 -6220
rect 5090 -6300 5140 -6290
rect 5090 -6330 5100 -6300
rect 5130 -6330 5140 -6300
rect 5090 -6340 5140 -6330
rect 5100 -6410 5130 -6340
rect 5090 -6420 5140 -6410
rect 5090 -6450 5100 -6420
rect 5130 -6450 5140 -6420
rect 5090 -6460 5140 -6450
rect 5100 -9430 5130 -6460
rect 5090 -9440 5140 -9430
rect 5090 -9470 5100 -9440
rect 5130 -9470 5140 -9440
rect 5090 -9480 5140 -9470
rect 5100 -9550 5130 -9480
rect 5090 -9560 5140 -9550
rect 5090 -9590 5100 -9560
rect 5130 -9590 5140 -9560
rect 5090 -9600 5140 -9590
rect 5100 -9670 5130 -9600
rect 5200 -9610 5230 970
rect 5300 -2840 5330 940
rect 5290 -2850 5340 -2840
rect 5290 -2880 5300 -2850
rect 5330 -2880 5340 -2850
rect 5290 -2890 5340 -2880
rect 5300 -2960 5330 -2890
rect 5290 -2970 5340 -2960
rect 5290 -3000 5300 -2970
rect 5330 -3000 5340 -2970
rect 5290 -3010 5340 -3000
rect 5300 -6170 5330 -3010
rect 5290 -6180 5340 -6170
rect 5290 -6210 5300 -6180
rect 5330 -6210 5340 -6180
rect 5290 -6220 5340 -6210
rect 5300 -6290 5330 -6220
rect 5290 -6300 5340 -6290
rect 5290 -6330 5300 -6300
rect 5330 -6330 5340 -6300
rect 5290 -6340 5340 -6330
rect 5300 -6410 5330 -6340
rect 5290 -6420 5340 -6410
rect 5290 -6450 5300 -6420
rect 5330 -6450 5340 -6420
rect 5290 -6460 5340 -6450
rect 5300 -9430 5330 -6460
rect 5290 -9440 5340 -9430
rect 5290 -9470 5300 -9440
rect 5330 -9470 5340 -9440
rect 5290 -9480 5340 -9470
rect 5300 -9550 5330 -9480
rect 5400 -9490 5430 970
rect 5500 -2840 5530 940
rect 5490 -2850 5540 -2840
rect 5490 -2880 5500 -2850
rect 5530 -2880 5540 -2850
rect 5490 -2890 5540 -2880
rect 5500 -2960 5530 -2890
rect 5490 -2970 5540 -2960
rect 5490 -3000 5500 -2970
rect 5530 -3000 5540 -2970
rect 5490 -3010 5540 -3000
rect 5500 -6170 5530 -3010
rect 5490 -6180 5540 -6170
rect 5490 -6210 5500 -6180
rect 5530 -6210 5540 -6180
rect 5490 -6220 5540 -6210
rect 5500 -6290 5530 -6220
rect 5490 -6300 5540 -6290
rect 5490 -6330 5500 -6300
rect 5530 -6330 5540 -6300
rect 5490 -6340 5540 -6330
rect 5500 -6410 5530 -6340
rect 5490 -6420 5540 -6410
rect 5490 -6450 5500 -6420
rect 5530 -6450 5540 -6420
rect 5490 -6460 5540 -6450
rect 5500 -9430 5530 -6460
rect 5490 -9440 5540 -9430
rect 5490 -9470 5500 -9440
rect 5530 -9470 5540 -9440
rect 5490 -9480 5540 -9470
rect 5390 -9500 5440 -9490
rect 5390 -9530 5400 -9500
rect 5430 -9530 5440 -9500
rect 5390 -9540 5440 -9530
rect 5290 -9560 5340 -9550
rect 5290 -9590 5300 -9560
rect 5330 -9590 5340 -9560
rect 5290 -9600 5340 -9590
rect 5190 -9620 5240 -9610
rect 5190 -9650 5200 -9620
rect 5230 -9650 5240 -9620
rect 5190 -9660 5240 -9650
rect 5090 -9680 5140 -9670
rect 5090 -9710 5100 -9680
rect 5130 -9710 5140 -9680
rect 5090 -9720 5140 -9710
rect 5100 -9790 5130 -9720
rect 5090 -9800 5140 -9790
rect 5090 -9830 5100 -9800
rect 5130 -9830 5140 -9800
rect 5090 -9840 5140 -9830
rect 5100 -9910 5130 -9840
rect 5090 -9920 5140 -9910
rect 5090 -9950 5100 -9920
rect 5130 -9950 5140 -9920
rect 5090 -9960 5140 -9950
rect 5100 -12000 5130 -9960
rect 5200 -12000 5230 -9660
rect 5300 -9670 5330 -9600
rect 5290 -9680 5340 -9670
rect 5290 -9710 5300 -9680
rect 5330 -9710 5340 -9680
rect 5290 -9720 5340 -9710
rect 5300 -9790 5330 -9720
rect 5290 -9800 5340 -9790
rect 5290 -9830 5300 -9800
rect 5330 -9830 5340 -9800
rect 5290 -9840 5340 -9830
rect 5300 -9910 5330 -9840
rect 5290 -9920 5340 -9910
rect 5290 -9950 5300 -9920
rect 5330 -9950 5340 -9920
rect 5290 -9960 5340 -9950
rect 5300 -12000 5330 -9960
rect 5400 -12000 5430 -9540
rect 5500 -9550 5530 -9480
rect 5490 -9560 5540 -9550
rect 5490 -9590 5500 -9560
rect 5530 -9590 5540 -9560
rect 5490 -9600 5540 -9590
rect 5500 -9670 5530 -9600
rect 5490 -9680 5540 -9670
rect 5490 -9710 5500 -9680
rect 5530 -9710 5540 -9680
rect 5490 -9720 5540 -9710
rect 5500 -9790 5530 -9720
rect 5490 -9800 5540 -9790
rect 5490 -9830 5500 -9800
rect 5530 -9830 5540 -9800
rect 5490 -9840 5540 -9830
rect 5500 -9910 5530 -9840
rect 5600 -9850 5630 970
rect 5700 -2840 5730 940
rect 5690 -2850 5740 -2840
rect 5690 -2880 5700 -2850
rect 5730 -2880 5740 -2850
rect 5690 -2890 5740 -2880
rect 5700 -2960 5730 -2890
rect 5800 -2900 5830 970
rect 5900 -2840 5930 940
rect 5980 930 6140 970
rect 5980 790 5990 930
rect 6130 790 6140 930
rect 5890 -2850 5940 -2840
rect 5890 -2880 5900 -2850
rect 5930 -2880 5940 -2850
rect 5890 -2890 5940 -2880
rect 5790 -2910 5840 -2900
rect 5790 -2940 5800 -2910
rect 5830 -2940 5840 -2910
rect 5790 -2950 5840 -2940
rect 5690 -2970 5740 -2960
rect 5690 -3000 5700 -2970
rect 5730 -3000 5740 -2970
rect 5690 -3010 5740 -3000
rect 5700 -6170 5730 -3010
rect 5690 -6180 5740 -6170
rect 5690 -6210 5700 -6180
rect 5730 -6210 5740 -6180
rect 5690 -6220 5740 -6210
rect 5700 -6290 5730 -6220
rect 5800 -6230 5830 -2950
rect 5900 -2960 5930 -2890
rect 5890 -2970 5940 -2960
rect 5890 -3000 5900 -2970
rect 5930 -3000 5940 -2970
rect 5890 -3010 5940 -3000
rect 5900 -6170 5930 -3010
rect 5980 -3040 6140 790
rect 6300 610 6460 970
rect 6300 470 6310 610
rect 6450 470 6460 610
rect 6300 -2840 6460 470
rect 6620 290 6780 970
rect 24620 930 24780 940
rect 24620 790 24630 930
rect 24770 790 24780 930
rect 24300 610 24460 620
rect 24300 470 24310 610
rect 24450 470 24460 610
rect 6620 150 6630 290
rect 6770 150 6780 290
rect 6290 -2850 6470 -2840
rect 6290 -2880 6300 -2850
rect 6460 -2880 6470 -2850
rect 6290 -2890 6470 -2880
rect 6300 -2960 6460 -2890
rect 6290 -2970 6470 -2960
rect 6290 -3000 6300 -2970
rect 6460 -3000 6470 -2970
rect 6290 -3010 6470 -3000
rect 5980 -3180 5990 -3040
rect 6130 -3180 6140 -3040
rect 5890 -6180 5940 -6170
rect 5890 -6210 5900 -6180
rect 5930 -6210 5940 -6180
rect 5890 -6220 5940 -6210
rect 5790 -6240 5840 -6230
rect 5790 -6270 5800 -6240
rect 5830 -6270 5840 -6240
rect 5790 -6280 5840 -6270
rect 5690 -6300 5740 -6290
rect 5690 -6330 5700 -6300
rect 5730 -6330 5740 -6300
rect 5690 -6340 5740 -6330
rect 5700 -6410 5730 -6340
rect 5690 -6420 5740 -6410
rect 5690 -6450 5700 -6420
rect 5730 -6450 5740 -6420
rect 5690 -6460 5740 -6450
rect 5700 -9430 5730 -6460
rect 5690 -9440 5740 -9430
rect 5690 -9470 5700 -9440
rect 5730 -9470 5740 -9440
rect 5690 -9480 5740 -9470
rect 5700 -9550 5730 -9480
rect 5690 -9560 5740 -9550
rect 5690 -9590 5700 -9560
rect 5730 -9590 5740 -9560
rect 5690 -9600 5740 -9590
rect 5700 -9670 5730 -9600
rect 5690 -9680 5740 -9670
rect 5690 -9710 5700 -9680
rect 5730 -9710 5740 -9680
rect 5690 -9720 5740 -9710
rect 5700 -9790 5730 -9720
rect 5690 -9800 5740 -9790
rect 5690 -9830 5700 -9800
rect 5730 -9830 5740 -9800
rect 5690 -9840 5740 -9830
rect 5590 -9860 5640 -9850
rect 5590 -9890 5600 -9860
rect 5630 -9890 5640 -9860
rect 5590 -9900 5640 -9890
rect 5490 -9920 5540 -9910
rect 5490 -9950 5500 -9920
rect 5530 -9950 5540 -9920
rect 5490 -9960 5540 -9950
rect 5500 -12000 5530 -9960
rect 5600 -12000 5630 -9900
rect 5700 -9910 5730 -9840
rect 5690 -9920 5740 -9910
rect 5690 -9950 5700 -9920
rect 5730 -9950 5740 -9920
rect 5690 -9960 5740 -9950
rect 5700 -12000 5730 -9960
rect 5800 -12000 5830 -6280
rect 5900 -6290 5930 -6220
rect 5890 -6300 5940 -6290
rect 5890 -6330 5900 -6300
rect 5930 -6330 5940 -6300
rect 5890 -6340 5940 -6330
rect 5900 -6410 5930 -6340
rect 5890 -6420 5940 -6410
rect 5890 -6450 5900 -6420
rect 5930 -6450 5940 -6420
rect 5890 -6460 5940 -6450
rect 5900 -9430 5930 -6460
rect 5890 -9440 5940 -9430
rect 5890 -9470 5900 -9440
rect 5930 -9470 5940 -9440
rect 5890 -9480 5940 -9470
rect 5900 -9550 5930 -9480
rect 5890 -9560 5940 -9550
rect 5890 -9590 5900 -9560
rect 5930 -9590 5940 -9560
rect 5890 -9600 5940 -9590
rect 5900 -9670 5930 -9600
rect 5890 -9680 5940 -9670
rect 5890 -9710 5900 -9680
rect 5930 -9710 5940 -9680
rect 5890 -9720 5940 -9710
rect 5900 -9790 5930 -9720
rect 5890 -9800 5940 -9790
rect 5890 -9830 5900 -9800
rect 5930 -9830 5940 -9800
rect 5890 -9840 5940 -9830
rect 5900 -9910 5930 -9840
rect 5890 -9920 5940 -9910
rect 5890 -9950 5900 -9920
rect 5930 -9950 5940 -9920
rect 5890 -9960 5940 -9950
rect 5900 -12000 5930 -9960
rect 5980 -11850 6140 -3180
rect 6300 -6170 6460 -3010
rect 6290 -6180 6470 -6170
rect 6290 -6210 6300 -6180
rect 6460 -6210 6470 -6180
rect 6290 -6220 6470 -6210
rect 6300 -6290 6460 -6220
rect 6290 -6300 6470 -6290
rect 6290 -6330 6300 -6300
rect 6460 -6330 6470 -6300
rect 6290 -6340 6470 -6330
rect 6300 -6420 6460 -6340
rect 6290 -6430 6470 -6420
rect 6290 -6460 6300 -6430
rect 6460 -6460 6470 -6430
rect 6290 -6470 6470 -6460
rect 6300 -9430 6460 -6470
rect 6290 -9440 6470 -9430
rect 6290 -9470 6300 -9440
rect 6460 -9470 6470 -9440
rect 6290 -9480 6470 -9470
rect 6300 -9550 6460 -9480
rect 6290 -9560 6470 -9550
rect 6290 -9590 6300 -9560
rect 6460 -9590 6470 -9560
rect 6290 -9600 6470 -9590
rect 6300 -9670 6460 -9600
rect 6290 -9680 6470 -9670
rect 6290 -9710 6300 -9680
rect 6460 -9710 6470 -9680
rect 6290 -9720 6470 -9710
rect 6300 -9790 6460 -9720
rect 6290 -9800 6470 -9790
rect 6290 -9830 6300 -9800
rect 6460 -9830 6470 -9800
rect 6290 -9840 6470 -9830
rect 6300 -9910 6460 -9840
rect 6290 -9920 6470 -9910
rect 6290 -9950 6300 -9920
rect 6460 -9950 6470 -9920
rect 6290 -9960 6470 -9950
rect 6300 -11530 6460 -9960
rect 6620 -11210 6780 150
rect 6620 -11350 6630 -11210
rect 6770 -11350 6780 -11210
rect 6620 -11360 6780 -11350
rect 23980 290 24140 300
rect 23980 150 23990 290
rect 24130 150 24140 290
rect 23980 -11210 24140 150
rect 23980 -11350 23990 -11210
rect 24130 -11350 24140 -11210
rect 23980 -11360 24140 -11350
rect 6300 -11670 6310 -11530
rect 6450 -11670 6460 -11530
rect 6300 -11680 6460 -11670
rect 24300 -11530 24460 470
rect 24300 -11670 24310 -11530
rect 24450 -11670 24460 -11530
rect 24300 -11680 24460 -11670
rect 5980 -11990 5990 -11850
rect 6130 -11990 6140 -11850
rect 5980 -12000 6140 -11990
rect 24620 -11850 24780 790
rect 24620 -11990 24630 -11850
rect 24770 -11990 24780 -11850
rect 24620 -12000 24780 -11990
<< via3 >>
rect 5990 790 6130 930
rect 6310 470 6450 610
rect 24630 790 24770 930
rect 24310 470 24450 610
rect 6630 150 6770 290
rect 23990 150 24130 290
rect 6310 -11670 6450 -11530
rect 24310 -11670 24450 -11530
rect 5990 -11990 6130 -11850
rect 24630 -11990 24770 -11850
<< metal4 >>
rect 5980 930 24780 940
rect 5980 790 5990 930
rect 6130 790 24630 930
rect 24770 790 24780 930
rect 5980 780 24780 790
rect 6300 610 24460 620
rect 6300 470 6310 610
rect 6450 470 24310 610
rect 24450 470 24460 610
rect 6300 460 24460 470
rect 6620 290 24140 300
rect 6620 150 6630 290
rect 6770 150 23990 290
rect 24130 150 24140 290
rect 6620 140 24140 150
rect 5130 -3000 23840 -2850
rect 5100 -6390 23840 -6240
rect 5100 -9650 23840 -9500
rect 5100 -9890 23840 -9740
rect 6300 -11530 24460 -11520
rect 6300 -11670 6310 -11530
rect 6450 -11670 24310 -11530
rect 24450 -11670 24460 -11530
rect 6300 -11680 24460 -11670
rect 5980 -11850 24780 -11840
rect 5980 -11990 5990 -11850
rect 6130 -11990 24630 -11850
rect 24770 -11990 24780 -11850
rect 5980 -12000 24780 -11990
<< metal5 >>
rect 5200 -12000 5430 940
rect 5600 -12000 5830 940
use n1_8  n1_8_0
timestamp 1634337365
transform 1 0 7860 0 1 -11190
box 0 0 940 1230
use p1_8  p1_8_5
timestamp 1634440922
transform 1 0 7860 0 1 -9430
box 0 0 940 2970
use n1_8  n1_8_16
timestamp 1634337365
transform 1 0 6920 0 1 -11190
box 0 0 940 1230
use p1_8  p1_8_48
timestamp 1634440922
transform 1 0 6920 0 1 -9430
box 0 0 940 2970
use p1_8  p1_8_4
timestamp 1634440922
transform -1 0 9740 0 1 -9430
box 0 0 940 2970
use n1_8  n1_8_1
timestamp 1634337365
transform -1 0 9740 0 1 -11190
box 0 0 940 1230
use n1_8  n1_8_3
timestamp 1634337365
transform 1 0 9740 0 1 -11190
box 0 0 940 1230
use p1_8  p1_8_11
timestamp 1634440922
transform 1 0 9740 0 1 -9430
box 0 0 940 2970
use n1_8  n1_8_2
timestamp 1634337365
transform -1 0 11620 0 1 -11190
box 0 0 940 1230
use p1_8  p1_8_10
timestamp 1634440922
transform -1 0 11620 0 1 -9430
box 0 0 940 2970
use p1_8  p1_8_13
timestamp 1634440922
transform 1 0 11620 0 1 -9430
box 0 0 940 2970
use n1_8  n1_8_5
timestamp 1634337365
transform 1 0 11620 0 1 -11190
box 0 0 940 1230
use p1_8  p1_8_12
timestamp 1634440922
transform -1 0 13500 0 1 -9430
box 0 0 940 2970
use n1_8  n1_8_4
timestamp 1634337365
transform -1 0 13500 0 1 -11190
box 0 0 940 1230
use n1_8  n1_8_6
timestamp 1634337365
transform 1 0 13500 0 1 -11190
box 0 0 940 1230
use p1_8  p1_8_14
timestamp 1634440922
transform 1 0 13500 0 1 -9430
box 0 0 940 2970
use n1_8  n1_8_7
timestamp 1634337365
transform -1 0 15380 0 1 -11190
box 0 0 940 1230
use p1_8  p1_8_15
timestamp 1634440922
transform -1 0 15380 0 1 -9430
box 0 0 940 2970
use p1_8  p1_8_25
timestamp 1634440922
transform 1 0 15380 0 1 -9430
box 0 0 940 2970
use n1_8  n1_8_9
timestamp 1634337365
transform 1 0 15380 0 1 -11190
box 0 0 940 1230
use p1_8  p1_8_26
timestamp 1634440922
transform -1 0 17260 0 1 -9430
box 0 0 940 2970
use n1_8  n1_8_10
timestamp 1634337365
transform -1 0 17260 0 1 -11190
box 0 0 940 1230
use p1_8  p1_8_24
timestamp 1634440922
transform 1 0 17260 0 1 -9430
box 0 0 940 2970
use n1_8  n1_8_8
timestamp 1634337365
transform 1 0 17260 0 1 -11190
box 0 0 940 1230
use p1_8  p1_8_29
timestamp 1634440922
transform -1 0 19140 0 1 -9430
box 0 0 940 2970
use n1_8  n1_8_13
timestamp 1634337365
transform -1 0 19140 0 1 -11190
box 0 0 940 1230
use p1_8  p1_8_30
timestamp 1634440922
transform 1 0 19140 0 1 -9430
box 0 0 940 2970
use n1_8  n1_8_14
timestamp 1634337365
transform 1 0 19140 0 1 -11190
box 0 0 940 1230
use p1_8  p1_8_28
timestamp 1634440922
transform -1 0 21020 0 1 -9430
box 0 0 940 2970
use n1_8  n1_8_12
timestamp 1634337365
transform -1 0 21020 0 1 -11190
box 0 0 940 1230
use p1_8  p1_8_27
timestamp 1634440922
transform 1 0 21020 0 1 -9430
box 0 0 940 2970
use n1_8  n1_8_11
timestamp 1634337365
transform 1 0 21020 0 1 -11190
box 0 0 940 1230
use n1_8  n1_8_15
timestamp 1634337365
transform -1 0 22900 0 1 -11190
box 0 0 940 1230
use p1_8  p1_8_31
timestamp 1634440922
transform -1 0 22900 0 1 -9430
box 0 0 940 2970
use n1_8  n1_8_17
timestamp 1634337365
transform -1 0 23840 0 1 -11190
box 0 0 940 1230
use p1_8  p1_8_51
timestamp 1634440922
transform -1 0 23840 0 1 -9430
box 0 0 940 2970
use p1_8  p1_8_2
timestamp 1634440922
transform 1 0 7860 0 1 -6170
box 0 0 940 2970
use p1_8  p1_8_49
timestamp 1634440922
transform 1 0 6920 0 1 -6170
box 0 0 940 2970
use p1_8  p1_8_3
timestamp 1634440922
transform -1 0 9740 0 1 -6170
box 0 0 940 2970
use p1_8  p1_8_9
timestamp 1634440922
transform 1 0 9740 0 1 -6170
box 0 0 940 2970
use p1_8  p1_8_8
timestamp 1634440922
transform -1 0 11620 0 1 -6170
box 0 0 940 2970
use p1_8  p1_8_17
timestamp 1634440922
transform 1 0 11620 0 1 -6170
box 0 0 940 2970
use p1_8  p1_8_16
timestamp 1634440922
transform -1 0 13500 0 1 -6170
box 0 0 940 2970
use p1_8  p1_8_18
timestamp 1634440922
transform 1 0 13500 0 1 -6170
box 0 0 940 2970
use p1_8  p1_8_19
timestamp 1634440922
transform -1 0 15380 0 1 -6170
box 0 0 940 2970
use p1_8  p1_8_33
timestamp 1634440922
transform 1 0 15380 0 1 -6170
box 0 0 940 2970
use p1_8  p1_8_34
timestamp 1634440922
transform -1 0 17260 0 1 -6170
box 0 0 940 2970
use p1_8  p1_8_32
timestamp 1634440922
transform 1 0 17260 0 1 -6170
box 0 0 940 2970
use p1_8  p1_8_37
timestamp 1634440922
transform -1 0 19140 0 1 -6170
box 0 0 940 2970
use p1_8  p1_8_38
timestamp 1634440922
transform 1 0 19140 0 1 -6170
box 0 0 940 2970
use p1_8  p1_8_35
timestamp 1634440922
transform -1 0 21020 0 1 -6170
box 0 0 940 2970
use p1_8  p1_8_36
timestamp 1634440922
transform 1 0 21020 0 1 -6170
box 0 0 940 2970
use p1_8  p1_8_39
timestamp 1634440922
transform -1 0 22900 0 1 -6170
box 0 0 940 2970
use p1_8  p1_8_52
timestamp 1634440922
transform -1 0 23840 0 1 -6170
box 0 0 940 2970
use p1_8  p1_8_0
timestamp 1634440922
transform 1 0 7860 0 1 -2840
box 0 0 940 2970
use p1_8  p1_8_50
timestamp 1634440922
transform 1 0 6920 0 1 -2840
box 0 0 940 2970
use p1_8  p1_8_1
timestamp 1634440922
transform -1 0 9740 0 1 -2840
box 0 0 940 2970
use p1_8  p1_8_6
timestamp 1634440922
transform 1 0 9740 0 1 -2840
box 0 0 940 2970
use p1_8  p1_8_7
timestamp 1634440922
transform -1 0 11620 0 1 -2840
box 0 0 940 2970
use p1_8  p1_8_20
timestamp 1634440922
transform 1 0 11620 0 1 -2840
box 0 0 940 2970
use p1_8  p1_8_21
timestamp 1634440922
transform -1 0 13500 0 1 -2840
box 0 0 940 2970
use p1_8  p1_8_22
timestamp 1634440922
transform 1 0 13500 0 1 -2840
box 0 0 940 2970
use p1_8  p1_8_23
timestamp 1634440922
transform -1 0 15380 0 1 -2840
box 0 0 940 2970
use p1_8  p1_8_42
timestamp 1634440922
transform 1 0 15380 0 1 -2840
box 0 0 940 2970
use p1_8  p1_8_41
timestamp 1634440922
transform -1 0 17260 0 1 -2840
box 0 0 940 2970
use p1_8  p1_8_40
timestamp 1634440922
transform 1 0 17260 0 1 -2840
box 0 0 940 2970
use p1_8  p1_8_45
timestamp 1634440922
transform -1 0 19140 0 1 -2840
box 0 0 940 2970
use p1_8  p1_8_46
timestamp 1634440922
transform 1 0 19140 0 1 -2840
box 0 0 940 2970
use p1_8  p1_8_44
timestamp 1634440922
transform -1 0 21020 0 1 -2840
box 0 0 940 2970
use p1_8  p1_8_43
timestamp 1634440922
transform 1 0 21020 0 1 -2840
box 0 0 940 2970
use p1_8  p1_8_47
timestamp 1634440922
transform -1 0 22900 0 1 -2840
box 0 0 940 2970
use p1_8  p1_8_53
timestamp 1634440922
transform -1 0 23840 0 1 -2840
box 0 0 940 2970
<< labels >>
rlabel metal3 5200 940 5230 970 1 inm
port 1 n
rlabel metal3 5400 940 5430 970 1 inp
port 2 n
rlabel metal3 5600 940 5630 970 1 out
port 3 n
rlabel metal3 5800 940 5830 970 1 ib
port 4 n
rlabel metal3 5980 940 6140 970 1 vdda
port 5 n
rlabel metal3 6300 940 6460 970 1 gnda
port 6 n
rlabel metal3 6620 940 6780 970 1 vssa
port 7 n
rlabel metal2 8780 80 8810 110 1 z
rlabel metal2 6840 -6390 6870 -6360 0 x
rlabel metal2 6840 -9770 6870 -9740 0 y
<< end >>
